magic
tech EFS8A
magscale 1 2
timestamp 1602530518
<< locali >>
rect 9631 23137 9758 23171
rect 10885 22049 11046 22083
rect 16439 22049 16474 22083
rect 10885 21947 10919 22049
rect 19349 21471 19383 21641
rect 19349 21335 19383 21437
rect 10149 20383 10183 20485
rect 11799 20009 11805 20043
rect 13547 20009 13553 20043
rect 11799 19941 11833 20009
rect 13547 19941 13581 20009
rect 2881 19873 3042 19907
rect 9631 19873 9758 19907
rect 15243 19873 15370 19907
rect 20855 19873 20982 19907
rect 2881 19703 2915 19873
rect 23995 19465 24133 19499
rect 5819 18921 5825 18955
rect 5819 18853 5853 18921
rect 2881 18785 3042 18819
rect 22879 18785 22914 18819
rect 25455 18785 25490 18819
rect 2881 18751 2915 18785
rect 20821 18139 20855 18309
rect 6187 17833 6193 17867
rect 6187 17765 6221 17833
rect 15703 17697 15738 17731
rect 11891 16745 11897 16779
rect 11891 16677 11925 16745
rect 24035 15657 24041 15691
rect 24035 15589 24069 15657
rect 25455 15521 25490 15555
rect 16589 15351 16623 15521
rect 12259 13481 12265 13515
rect 12259 13413 12293 13481
rect 8027 12393 8033 12427
rect 8027 12325 8061 12393
rect 19435 11305 19441 11339
rect 22287 11305 22293 11339
rect 19435 11237 19469 11305
rect 22287 11237 22321 11305
rect 15335 11169 15462 11203
rect 20855 11169 20982 11203
rect 13645 10455 13679 10625
rect 15427 10081 15554 10115
rect 3433 9571 3467 9673
rect 3893 8993 4110 9027
rect 3893 8959 3927 8993
rect 4364 7973 4432 8007
rect 5181 7803 5215 7973
rect 17963 6953 17969 6987
rect 2455 6885 2500 6919
rect 17963 6885 17997 6953
rect 19475 6817 19602 6851
rect 25375 6409 25513 6443
rect 1443 5729 1478 5763
rect 21315 5729 21350 5763
rect 7383 4777 7389 4811
rect 19435 4777 19441 4811
rect 7383 4709 7417 4777
rect 19435 4709 19469 4777
rect 1903 4641 2030 4675
rect 3007 4641 3042 4675
rect 13587 4233 13771 4267
rect 15847 3689 15853 3723
rect 15847 3621 15881 3689
rect 17693 3451 17727 3553
rect 20913 3043 20947 3145
rect 5089 2363 5123 2465
<< viali >>
rect 25145 24905 25179 24939
rect 24660 24701 24694 24735
rect 12449 24565 12483 24599
rect 24731 24565 24765 24599
rect 24777 24361 24811 24395
rect 12700 24225 12734 24259
rect 13712 24225 13746 24259
rect 24593 24225 24627 24259
rect 12771 24021 12805 24055
rect 13783 24021 13817 24055
rect 5365 23817 5399 23851
rect 7021 23817 7055 23851
rect 7481 23817 7515 23851
rect 12633 23817 12667 23851
rect 13369 23817 13403 23851
rect 15945 23817 15979 23851
rect 24777 23817 24811 23851
rect 14703 23749 14737 23783
rect 1460 23613 1494 23647
rect 1869 23613 1903 23647
rect 4972 23613 5006 23647
rect 6837 23613 6871 23647
rect 12449 23613 12483 23647
rect 13001 23613 13035 23647
rect 13588 23613 13622 23647
rect 14632 23613 14666 23647
rect 15117 23613 15151 23647
rect 15761 23613 15795 23647
rect 16313 23613 16347 23647
rect 18061 23613 18095 23647
rect 24593 23613 24627 23647
rect 1547 23545 1581 23579
rect 14473 23545 14507 23579
rect 18613 23545 18647 23579
rect 5043 23477 5077 23511
rect 13691 23477 13725 23511
rect 14105 23477 14139 23511
rect 18245 23477 18279 23511
rect 24409 23477 24443 23511
rect 25237 23477 25271 23511
rect 24777 23273 24811 23307
rect 1476 23137 1510 23171
rect 9597 23137 9631 23171
rect 11228 23137 11262 23171
rect 13252 23137 13286 23171
rect 15368 23137 15402 23171
rect 16380 23137 16414 23171
rect 24593 23137 24627 23171
rect 12173 23069 12207 23103
rect 14197 23069 14231 23103
rect 9827 23001 9861 23035
rect 1547 22933 1581 22967
rect 11299 22933 11333 22967
rect 13323 22933 13357 22967
rect 15439 22933 15473 22967
rect 16451 22933 16485 22967
rect 1593 22729 1627 22763
rect 7665 22729 7699 22763
rect 10885 22729 10919 22763
rect 15669 22729 15703 22763
rect 24685 22729 24719 22763
rect 10149 22661 10183 22695
rect 10609 22661 10643 22695
rect 15347 22593 15381 22627
rect 16359 22593 16393 22627
rect 7481 22525 7515 22559
rect 8033 22525 8067 22559
rect 8712 22525 8746 22559
rect 9137 22525 9171 22559
rect 9756 22525 9790 22559
rect 10701 22525 10735 22559
rect 12884 22525 12918 22559
rect 13737 22525 13771 22559
rect 14264 22525 14298 22559
rect 15260 22525 15294 22559
rect 16256 22525 16290 22559
rect 8815 22457 8849 22491
rect 16681 22457 16715 22491
rect 9827 22389 9861 22423
rect 11345 22389 11379 22423
rect 12955 22389 12989 22423
rect 13369 22389 13403 22423
rect 14335 22389 14369 22423
rect 14749 22389 14783 22423
rect 16129 22389 16163 22423
rect 17049 22389 17083 22423
rect 6883 22185 6917 22219
rect 14013 22185 14047 22219
rect 13093 22117 13127 22151
rect 13185 22117 13219 22151
rect 17555 22117 17589 22151
rect 6812 22049 6846 22083
rect 8008 22049 8042 22083
rect 9724 22049 9758 22083
rect 10793 22049 10827 22083
rect 12056 22049 12090 22083
rect 15393 22049 15427 22083
rect 16405 22049 16439 22083
rect 17452 22049 17486 22083
rect 18496 22049 18530 22083
rect 20964 22049 20998 22083
rect 21051 21981 21085 22015
rect 10885 21913 10919 21947
rect 13645 21913 13679 21947
rect 18567 21913 18601 21947
rect 8079 21845 8113 21879
rect 8677 21845 8711 21879
rect 9045 21845 9079 21879
rect 9827 21845 9861 21879
rect 11115 21845 11149 21879
rect 12127 21845 12161 21879
rect 15577 21845 15611 21879
rect 16543 21845 16577 21879
rect 10287 21641 10321 21675
rect 14381 21641 14415 21675
rect 16773 21641 16807 21675
rect 19349 21641 19383 21675
rect 20913 21641 20947 21675
rect 21281 21641 21315 21675
rect 8493 21573 8527 21607
rect 9689 21573 9723 21607
rect 11069 21573 11103 21607
rect 15071 21573 15105 21607
rect 16405 21573 16439 21607
rect 19211 21573 19245 21607
rect 8677 21505 8711 21539
rect 13461 21505 13495 21539
rect 15761 21505 15795 21539
rect 17877 21505 17911 21539
rect 18613 21505 18647 21539
rect 7640 21437 7674 21471
rect 10216 21437 10250 21471
rect 10609 21437 10643 21471
rect 11228 21437 11262 21471
rect 14968 21437 15002 21471
rect 15485 21437 15519 21471
rect 16012 21437 16046 21471
rect 17008 21437 17042 21471
rect 18061 21437 18095 21471
rect 19140 21437 19174 21471
rect 19349 21437 19383 21471
rect 20504 21437 20538 21471
rect 20591 21437 20625 21471
rect 8769 21369 8803 21403
rect 9321 21369 9355 21403
rect 13553 21369 13587 21403
rect 14105 21369 14139 21403
rect 17095 21369 17129 21403
rect 5733 21301 5767 21335
rect 7113 21301 7147 21335
rect 7711 21301 7745 21335
rect 8125 21301 8159 21335
rect 11299 21301 11333 21335
rect 11713 21301 11747 21335
rect 12081 21301 12115 21335
rect 12909 21301 12943 21335
rect 13185 21301 13219 21335
rect 16083 21301 16117 21335
rect 17417 21301 17451 21335
rect 18245 21301 18279 21335
rect 18889 21301 18923 21335
rect 19349 21301 19383 21335
rect 19625 21301 19659 21335
rect 8125 21029 8159 21063
rect 8217 21029 8251 21063
rect 9873 21029 9907 21063
rect 11713 21029 11747 21063
rect 12265 21029 12299 21063
rect 13185 21029 13219 21063
rect 13277 21029 13311 21063
rect 1568 20961 1602 20995
rect 4848 20961 4882 20995
rect 5917 20961 5951 20995
rect 6285 20961 6319 20995
rect 15393 20961 15427 20995
rect 15853 20961 15887 20995
rect 17024 20961 17058 20995
rect 18036 20961 18070 20995
rect 19016 20961 19050 20995
rect 20948 20961 20982 20995
rect 5733 20893 5767 20927
rect 6561 20893 6595 20927
rect 6837 20893 6871 20927
rect 8401 20893 8435 20927
rect 9781 20893 9815 20927
rect 10057 20893 10091 20927
rect 11437 20893 11471 20927
rect 11621 20893 11655 20927
rect 15945 20893 15979 20927
rect 13737 20825 13771 20859
rect 16773 20825 16807 20859
rect 21051 20825 21085 20859
rect 1639 20757 1673 20791
rect 4951 20757 4985 20791
rect 16497 20757 16531 20791
rect 17095 20757 17129 20791
rect 18107 20757 18141 20791
rect 19119 20757 19153 20791
rect 1593 20553 1627 20587
rect 4721 20553 4755 20587
rect 8125 20553 8159 20587
rect 8769 20553 8803 20587
rect 11437 20553 11471 20587
rect 12909 20553 12943 20587
rect 15669 20553 15703 20587
rect 17325 20553 17359 20587
rect 21649 20553 21683 20587
rect 4077 20485 4111 20519
rect 10149 20485 10183 20519
rect 10241 20485 10275 20519
rect 14105 20485 14139 20519
rect 14473 20485 14507 20519
rect 16129 20485 16163 20519
rect 6837 20417 6871 20451
rect 8953 20417 8987 20451
rect 11897 20417 11931 20451
rect 12173 20417 12207 20451
rect 13185 20417 13219 20451
rect 14749 20417 14783 20451
rect 15025 20417 15059 20451
rect 21373 20417 21407 20451
rect 1409 20349 1443 20383
rect 1961 20349 1995 20383
rect 3893 20349 3927 20383
rect 4905 20349 4939 20383
rect 5457 20349 5491 20383
rect 10149 20349 10183 20383
rect 10425 20349 10459 20383
rect 10885 20349 10919 20383
rect 18061 20349 18095 20383
rect 18613 20349 18647 20383
rect 19876 20349 19910 20383
rect 20856 20349 20890 20383
rect 21884 20349 21918 20383
rect 22293 20349 22327 20383
rect 5641 20281 5675 20315
rect 6653 20281 6687 20315
rect 7199 20281 7233 20315
rect 9045 20281 9079 20315
rect 9597 20281 9631 20315
rect 11161 20281 11195 20315
rect 13277 20281 13311 20315
rect 13829 20281 13863 20315
rect 14841 20281 14875 20315
rect 16405 20281 16439 20315
rect 16497 20281 16531 20315
rect 17049 20281 17083 20315
rect 18797 20281 18831 20315
rect 21971 20281 22005 20315
rect 2421 20213 2455 20247
rect 3709 20213 3743 20247
rect 4445 20213 4479 20247
rect 6009 20213 6043 20247
rect 7757 20213 7791 20247
rect 9965 20213 9999 20247
rect 17877 20213 17911 20247
rect 19073 20213 19107 20247
rect 19947 20213 19981 20247
rect 20361 20213 20395 20247
rect 20959 20213 20993 20247
rect 5181 20009 5215 20043
rect 7205 20009 7239 20043
rect 8401 20009 8435 20043
rect 8953 20009 8987 20043
rect 9505 20009 9539 20043
rect 9827 20009 9861 20043
rect 11805 20009 11839 20043
rect 12357 20009 12391 20043
rect 13093 20009 13127 20043
rect 13553 20009 13587 20043
rect 14105 20009 14139 20043
rect 14749 20009 14783 20043
rect 16313 20009 16347 20043
rect 18061 20009 18095 20043
rect 1547 19941 1581 19975
rect 6003 19941 6037 19975
rect 7481 19941 7515 19975
rect 7573 19941 7607 19975
rect 16589 19941 16623 19975
rect 1444 19873 1478 19907
rect 4629 19873 4663 19907
rect 5641 19873 5675 19907
rect 9597 19873 9631 19907
rect 11437 19873 11471 19907
rect 15209 19873 15243 19907
rect 18797 19873 18831 19907
rect 19073 19873 19107 19907
rect 20821 19873 20855 19907
rect 5549 19805 5583 19839
rect 8125 19805 8159 19839
rect 13185 19805 13219 19839
rect 15439 19805 15473 19839
rect 16497 19805 16531 19839
rect 19349 19805 19383 19839
rect 22661 19805 22695 19839
rect 23673 19805 23707 19839
rect 24685 19805 24719 19839
rect 6561 19737 6595 19771
rect 17049 19737 17083 19771
rect 2881 19669 2915 19703
rect 3111 19669 3145 19703
rect 4813 19669 4847 19703
rect 10517 19669 10551 19703
rect 12633 19669 12667 19703
rect 18521 19669 18555 19703
rect 19625 19669 19659 19703
rect 21051 19669 21085 19703
rect 2237 19465 2271 19499
rect 5089 19465 5123 19499
rect 8125 19465 8159 19499
rect 8493 19465 8527 19499
rect 11805 19465 11839 19499
rect 12265 19465 12299 19499
rect 13645 19465 13679 19499
rect 15945 19465 15979 19499
rect 16313 19465 16347 19499
rect 19073 19465 19107 19499
rect 24133 19465 24167 19499
rect 5825 19397 5859 19431
rect 7757 19397 7791 19431
rect 11529 19397 11563 19431
rect 22385 19397 22419 19431
rect 5273 19329 5307 19363
rect 6653 19329 6687 19363
rect 7205 19329 7239 19363
rect 8769 19329 8803 19363
rect 9413 19329 9447 19363
rect 11161 19329 11195 19363
rect 14013 19329 14047 19363
rect 14657 19329 14691 19363
rect 16497 19329 16531 19363
rect 18429 19329 18463 19363
rect 1476 19261 1510 19295
rect 1869 19261 1903 19295
rect 3208 19261 3242 19295
rect 3295 19261 3329 19295
rect 6193 19261 6227 19295
rect 10425 19261 10459 19295
rect 10977 19261 11011 19295
rect 12449 19261 12483 19295
rect 17141 19261 17175 19295
rect 19625 19261 19659 19295
rect 20085 19261 20119 19295
rect 21256 19261 21290 19295
rect 22201 19261 22235 19295
rect 22661 19261 22695 19295
rect 23924 19261 23958 19295
rect 5365 19193 5399 19227
rect 7297 19193 7331 19227
rect 8861 19193 8895 19227
rect 12811 19193 12845 19227
rect 14289 19193 14323 19227
rect 14381 19193 14415 19227
rect 16589 19193 16623 19227
rect 18153 19193 18187 19227
rect 18245 19193 18279 19227
rect 19441 19193 19475 19227
rect 24409 19193 24443 19227
rect 1547 19125 1581 19159
rect 2973 19125 3007 19159
rect 3617 19125 3651 19159
rect 4169 19125 4203 19159
rect 4721 19125 4755 19159
rect 9689 19125 9723 19159
rect 10241 19125 10275 19159
rect 13369 19125 13403 19159
rect 15301 19125 15335 19159
rect 17417 19125 17451 19159
rect 17877 19125 17911 19159
rect 19717 19125 19751 19159
rect 20913 19125 20947 19159
rect 21327 19125 21361 19159
rect 21741 19125 21775 19159
rect 24869 19125 24903 19159
rect 1593 18921 1627 18955
rect 5825 18921 5859 18955
rect 7481 18921 7515 18955
rect 7941 18921 7975 18955
rect 14381 18921 14415 18955
rect 16681 18921 16715 18955
rect 16957 18921 16991 18955
rect 18705 18921 18739 18955
rect 19165 18921 19199 18955
rect 8125 18853 8159 18887
rect 8217 18853 8251 18887
rect 9873 18853 9907 18887
rect 11897 18853 11931 18887
rect 13461 18853 13495 18887
rect 14657 18853 14691 18887
rect 16082 18853 16116 18887
rect 17693 18853 17727 18887
rect 1409 18785 1443 18819
rect 4512 18785 4546 18819
rect 5365 18785 5399 18819
rect 6377 18785 6411 18819
rect 19073 18785 19107 18819
rect 19533 18785 19567 18819
rect 21557 18785 21591 18819
rect 21741 18785 21775 18819
rect 22845 18785 22879 18819
rect 24476 18785 24510 18819
rect 25421 18785 25455 18819
rect 2881 18717 2915 18751
rect 5457 18717 5491 18751
rect 8769 18717 8803 18751
rect 9781 18717 9815 18751
rect 10057 18717 10091 18751
rect 11805 18717 11839 18751
rect 13369 18717 13403 18751
rect 13737 18717 13771 18751
rect 15761 18717 15795 18751
rect 17601 18717 17635 18751
rect 17877 18717 17911 18751
rect 21833 18717 21867 18751
rect 4583 18649 4617 18683
rect 12357 18649 12391 18683
rect 3111 18581 3145 18615
rect 4997 18581 5031 18615
rect 9137 18581 9171 18615
rect 10885 18581 10919 18615
rect 12725 18581 12759 18615
rect 15669 18581 15703 18615
rect 20085 18581 20119 18615
rect 21189 18581 21223 18615
rect 22983 18581 23017 18615
rect 24547 18581 24581 18615
rect 25559 18581 25593 18615
rect 1593 18377 1627 18411
rect 2053 18377 2087 18411
rect 8585 18377 8619 18411
rect 8953 18377 8987 18411
rect 10609 18377 10643 18411
rect 11897 18377 11931 18411
rect 13645 18377 13679 18411
rect 16957 18377 16991 18411
rect 17509 18377 17543 18411
rect 18199 18377 18233 18411
rect 18613 18377 18647 18411
rect 20913 18377 20947 18411
rect 24777 18377 24811 18411
rect 3065 18309 3099 18343
rect 4537 18309 4571 18343
rect 9781 18309 9815 18343
rect 20821 18309 20855 18343
rect 5549 18241 5583 18275
rect 6193 18241 6227 18275
rect 10149 18241 10183 18275
rect 11529 18241 11563 18275
rect 14933 18241 14967 18275
rect 20269 18241 20303 18275
rect 1409 18173 1443 18207
rect 3249 18173 3283 18207
rect 3801 18173 3835 18207
rect 4997 18173 5031 18207
rect 5273 18173 5307 18207
rect 7385 18173 7419 18207
rect 8309 18173 8343 18207
rect 10793 18173 10827 18207
rect 11253 18173 11287 18207
rect 12449 18173 12483 18207
rect 13369 18173 13403 18207
rect 14013 18173 14047 18207
rect 16037 18173 16071 18207
rect 18128 18173 18162 18207
rect 20637 18173 20671 18207
rect 21465 18241 21499 18275
rect 24133 18173 24167 18207
rect 24593 18173 24627 18207
rect 3985 18105 4019 18139
rect 7710 18105 7744 18139
rect 9229 18105 9263 18139
rect 9321 18105 9355 18139
rect 12770 18105 12804 18139
rect 14289 18105 14323 18139
rect 14381 18105 14415 18139
rect 16358 18105 16392 18139
rect 19625 18105 19659 18139
rect 19717 18105 19751 18139
rect 20821 18105 20855 18139
rect 21189 18105 21223 18139
rect 21281 18105 21315 18139
rect 2605 18037 2639 18071
rect 5917 18037 5951 18071
rect 7205 18037 7239 18071
rect 12265 18037 12299 18071
rect 15485 18037 15519 18071
rect 15853 18037 15887 18071
rect 19073 18037 19107 18071
rect 22109 18037 22143 18071
rect 22845 18037 22879 18071
rect 24501 18037 24535 18071
rect 25513 18037 25547 18071
rect 3893 17833 3927 17867
rect 5273 17833 5307 17867
rect 6193 17833 6227 17867
rect 6745 17833 6779 17867
rect 7389 17833 7423 17867
rect 8493 17833 8527 17867
rect 9229 17833 9263 17867
rect 9873 17833 9907 17867
rect 11805 17833 11839 17867
rect 13369 17833 13403 17867
rect 13829 17833 13863 17867
rect 14381 17833 14415 17867
rect 15807 17833 15841 17867
rect 17693 17833 17727 17867
rect 18981 17833 19015 17867
rect 19993 17833 20027 17867
rect 20269 17833 20303 17867
rect 21005 17833 21039 17867
rect 21925 17833 21959 17867
rect 3525 17765 3559 17799
rect 7935 17765 7969 17799
rect 11345 17765 11379 17799
rect 12494 17765 12528 17799
rect 16865 17765 16899 17799
rect 19394 17765 19428 17799
rect 2973 17697 3007 17731
rect 4537 17697 4571 17731
rect 4721 17697 4755 17731
rect 4997 17697 5031 17731
rect 7573 17697 7607 17731
rect 10609 17697 10643 17731
rect 11161 17697 11195 17731
rect 13988 17697 14022 17731
rect 15669 17697 15703 17731
rect 19073 17697 19107 17731
rect 20913 17697 20947 17731
rect 21465 17697 21499 17731
rect 23029 17697 23063 17731
rect 23213 17697 23247 17731
rect 24593 17697 24627 17731
rect 1961 17629 1995 17663
rect 5825 17629 5859 17663
rect 12173 17629 12207 17663
rect 16773 17629 16807 17663
rect 17417 17629 17451 17663
rect 23489 17629 23523 17663
rect 16589 17561 16623 17595
rect 1593 17493 1627 17527
rect 3157 17493 3191 17527
rect 8861 17493 8895 17527
rect 13093 17493 13127 17527
rect 14059 17493 14093 17527
rect 16221 17493 16255 17527
rect 22661 17493 22695 17527
rect 24777 17493 24811 17527
rect 1593 17289 1627 17323
rect 2053 17289 2087 17323
rect 2973 17289 3007 17323
rect 8677 17289 8711 17323
rect 10609 17289 10643 17323
rect 11897 17289 11931 17323
rect 13369 17289 13403 17323
rect 17417 17289 17451 17323
rect 18613 17289 18647 17323
rect 19993 17289 20027 17323
rect 23029 17289 23063 17323
rect 25421 17289 25455 17323
rect 14197 17221 14231 17255
rect 15531 17221 15565 17255
rect 17049 17221 17083 17255
rect 20361 17221 20395 17255
rect 22707 17221 22741 17255
rect 24685 17221 24719 17255
rect 5825 17153 5859 17187
rect 6469 17153 6503 17187
rect 9505 17153 9539 17187
rect 11529 17153 11563 17187
rect 13645 17153 13679 17187
rect 16497 17153 16531 17187
rect 17785 17153 17819 17187
rect 18199 17153 18233 17187
rect 19073 17153 19107 17187
rect 20637 17153 20671 17187
rect 20913 17153 20947 17187
rect 1409 17085 1443 17119
rect 3065 17085 3099 17119
rect 3893 17085 3927 17119
rect 4077 17085 4111 17119
rect 4997 17085 5031 17119
rect 5181 17085 5215 17119
rect 5549 17085 5583 17119
rect 7113 17085 7147 17119
rect 7481 17085 7515 17119
rect 7665 17085 7699 17119
rect 10793 17085 10827 17119
rect 11253 17085 11287 17119
rect 12500 17085 12534 17119
rect 15428 17085 15462 17119
rect 15853 17085 15887 17119
rect 18112 17085 18146 17119
rect 22636 17085 22670 17119
rect 23489 17085 23523 17119
rect 23673 17085 23707 17119
rect 24133 17085 24167 17119
rect 25237 17085 25271 17119
rect 25789 17085 25823 17119
rect 7941 17017 7975 17051
rect 8861 17017 8895 17051
rect 8953 17017 8987 17051
rect 12587 17017 12621 17051
rect 13737 17017 13771 17051
rect 16221 17017 16255 17051
rect 16589 17017 16623 17051
rect 19394 17017 19428 17051
rect 21005 17017 21039 17051
rect 21557 17017 21591 17051
rect 22477 17017 22511 17051
rect 3249 16949 3283 16983
rect 3617 16949 3651 16983
rect 4261 16949 4295 16983
rect 4629 16949 4663 16983
rect 6101 16949 6135 16983
rect 8309 16949 8343 16983
rect 9965 16949 9999 16983
rect 10241 16949 10275 16983
rect 12173 16949 12207 16983
rect 13001 16949 13035 16983
rect 14657 16949 14691 16983
rect 18889 16949 18923 16983
rect 21833 16949 21867 16983
rect 23765 16949 23799 16983
rect 1593 16745 1627 16779
rect 2329 16745 2363 16779
rect 4261 16745 4295 16779
rect 5273 16745 5307 16779
rect 7573 16745 7607 16779
rect 10793 16745 10827 16779
rect 11897 16745 11931 16779
rect 12449 16745 12483 16779
rect 17049 16745 17083 16779
rect 20729 16745 20763 16779
rect 5549 16677 5583 16711
rect 5825 16677 5859 16711
rect 5917 16677 5951 16711
rect 7297 16677 7331 16711
rect 9873 16677 9907 16711
rect 12725 16677 12759 16711
rect 13369 16677 13403 16711
rect 13645 16677 13679 16711
rect 16450 16677 16484 16711
rect 17325 16677 17359 16711
rect 18061 16677 18095 16711
rect 19579 16677 19613 16711
rect 21097 16677 21131 16711
rect 21649 16677 21683 16711
rect 24317 16677 24351 16711
rect 24409 16677 24443 16711
rect 1409 16609 1443 16643
rect 3040 16609 3074 16643
rect 4721 16609 4755 16643
rect 8033 16609 8067 16643
rect 8493 16609 8527 16643
rect 19492 16609 19526 16643
rect 22845 16609 22879 16643
rect 23121 16609 23155 16643
rect 6469 16541 6503 16575
rect 8769 16541 8803 16575
rect 9505 16541 9539 16575
rect 9781 16541 9815 16575
rect 11529 16541 11563 16575
rect 13553 16541 13587 16575
rect 13829 16541 13863 16575
rect 16129 16541 16163 16575
rect 17969 16541 18003 16575
rect 18429 16541 18463 16575
rect 21005 16541 21039 16575
rect 23397 16541 23431 16575
rect 24961 16541 24995 16575
rect 3111 16473 3145 16507
rect 4905 16473 4939 16507
rect 10333 16473 10367 16507
rect 19901 16473 19935 16507
rect 1961 16405 1995 16439
rect 3709 16405 3743 16439
rect 19073 16405 19107 16439
rect 23673 16405 23707 16439
rect 24041 16405 24075 16439
rect 2421 16201 2455 16235
rect 6193 16201 6227 16235
rect 9965 16201 9999 16235
rect 15025 16201 15059 16235
rect 16957 16201 16991 16235
rect 17785 16201 17819 16235
rect 22293 16201 22327 16235
rect 22753 16201 22787 16235
rect 24593 16201 24627 16235
rect 25237 16201 25271 16235
rect 25605 16201 25639 16235
rect 3893 16133 3927 16167
rect 15485 16133 15519 16167
rect 15853 16133 15887 16167
rect 24869 16133 24903 16167
rect 3764 16065 3798 16099
rect 3985 16065 4019 16099
rect 11253 16065 11287 16099
rect 12541 16065 12575 16099
rect 16037 16065 16071 16099
rect 17233 16065 17267 16099
rect 19441 16065 19475 16099
rect 21281 16065 21315 16099
rect 23673 16065 23707 16099
rect 1409 15997 1443 16031
rect 2656 15997 2690 16031
rect 3617 15997 3651 16031
rect 4629 15997 4663 16031
rect 5089 15997 5123 16031
rect 5365 15997 5399 16031
rect 5733 15997 5767 16031
rect 7205 15997 7239 16031
rect 7389 15997 7423 16031
rect 7665 15997 7699 16031
rect 8493 15997 8527 16031
rect 10333 15997 10367 16031
rect 10517 15997 10551 16031
rect 10977 15997 11011 16031
rect 13921 15997 13955 16031
rect 14197 15997 14231 16031
rect 14473 15997 14507 16031
rect 18061 15997 18095 16031
rect 18521 15997 18555 16031
rect 25421 15997 25455 16031
rect 25973 15997 26007 16031
rect 2743 15929 2777 15963
rect 4353 15929 4387 15963
rect 6653 15929 6687 15963
rect 8814 15929 8848 15963
rect 12633 15929 12667 15963
rect 13185 15929 13219 15963
rect 13553 15929 13587 15963
rect 16358 15929 16392 15963
rect 19762 15929 19796 15963
rect 21373 15929 21407 15963
rect 21925 15929 21959 15963
rect 24035 15929 24069 15963
rect 1593 15861 1627 15895
rect 2053 15861 2087 15895
rect 3065 15861 3099 15895
rect 3525 15861 3559 15895
rect 5273 15861 5307 15895
rect 7941 15861 7975 15895
rect 8309 15861 8343 15895
rect 9413 15861 9447 15895
rect 11621 15861 11655 15895
rect 12265 15861 12299 15895
rect 14105 15861 14139 15895
rect 18245 15861 18279 15895
rect 18889 15861 18923 15895
rect 19349 15861 19383 15895
rect 20361 15861 20395 15895
rect 21005 15861 21039 15895
rect 23029 15861 23063 15895
rect 23397 15861 23431 15895
rect 5273 15657 5307 15691
rect 6285 15657 6319 15691
rect 7021 15657 7055 15691
rect 8677 15657 8711 15691
rect 9505 15657 9539 15691
rect 11529 15657 11563 15691
rect 12633 15657 12667 15691
rect 14473 15657 14507 15691
rect 16037 15657 16071 15691
rect 16773 15657 16807 15691
rect 19717 15657 19751 15691
rect 21281 15657 21315 15691
rect 21557 15657 21591 15691
rect 24041 15657 24075 15691
rect 3709 15589 3743 15623
rect 5727 15589 5761 15623
rect 7434 15589 7468 15623
rect 10286 15589 10320 15623
rect 12034 15589 12068 15623
rect 13277 15589 13311 15623
rect 13553 15589 13587 15623
rect 13645 15589 13679 15623
rect 18842 15589 18876 15623
rect 22062 15589 22096 15623
rect 1961 15521 1995 15555
rect 2973 15521 3007 15555
rect 4420 15521 4454 15555
rect 5365 15521 5399 15555
rect 9965 15521 9999 15555
rect 10885 15521 10919 15555
rect 15761 15521 15795 15555
rect 16313 15521 16347 15555
rect 16589 15521 16623 15555
rect 17325 15521 17359 15555
rect 19441 15521 19475 15555
rect 21741 15521 21775 15555
rect 23673 15521 23707 15555
rect 25421 15521 25455 15555
rect 2881 15453 2915 15487
rect 7113 15453 7147 15487
rect 11713 15453 11747 15487
rect 13829 15453 13863 15487
rect 4491 15385 4525 15419
rect 8401 15385 8435 15419
rect 18521 15453 18555 15487
rect 17877 15385 17911 15419
rect 1869 15317 1903 15351
rect 2421 15317 2455 15351
rect 3157 15317 3191 15351
rect 4813 15317 4847 15351
rect 6561 15317 6595 15351
rect 8033 15317 8067 15351
rect 16589 15317 16623 15351
rect 17509 15317 17543 15351
rect 22661 15317 22695 15351
rect 24593 15317 24627 15351
rect 24961 15317 24995 15351
rect 25559 15317 25593 15351
rect 2126 15113 2160 15147
rect 4537 15113 4571 15147
rect 9413 15113 9447 15147
rect 10057 15113 10091 15147
rect 13001 15113 13035 15147
rect 13461 15113 13495 15147
rect 16681 15113 16715 15147
rect 17325 15113 17359 15147
rect 19625 15113 19659 15147
rect 23397 15113 23431 15147
rect 24409 15113 24443 15147
rect 2237 15045 2271 15079
rect 2973 15045 3007 15079
rect 6561 15045 6595 15079
rect 12265 15045 12299 15079
rect 22661 15045 22695 15079
rect 23857 15045 23891 15079
rect 2329 14977 2363 15011
rect 4261 14977 4295 15011
rect 5825 14977 5859 15011
rect 7389 14977 7423 15011
rect 8493 14977 8527 15011
rect 13737 14977 13771 15011
rect 14841 14977 14875 15011
rect 16221 14977 16255 15011
rect 19349 14977 19383 15011
rect 20545 14977 20579 15011
rect 20821 14977 20855 15011
rect 22109 14977 22143 15011
rect 23029 14977 23063 15011
rect 24593 14977 24627 15011
rect 25237 14977 25271 15011
rect 1961 14909 1995 14943
rect 3433 14909 3467 14943
rect 3801 14909 3835 14943
rect 3985 14909 4019 14943
rect 5181 14909 5215 14943
rect 5549 14909 5583 14943
rect 10701 14909 10735 14943
rect 11069 14909 11103 14943
rect 11253 14909 11287 14943
rect 12516 14909 12550 14943
rect 15945 14909 15979 14943
rect 16129 14909 16163 14943
rect 18613 14909 18647 14943
rect 19165 14909 19199 14943
rect 2697 14841 2731 14875
rect 6929 14841 6963 14875
rect 7021 14841 7055 14875
rect 8814 14841 8848 14875
rect 11529 14841 11563 14875
rect 13829 14841 13863 14875
rect 14381 14841 14415 14875
rect 15209 14841 15243 14875
rect 15577 14841 15611 14875
rect 20637 14841 20671 14875
rect 22201 14841 22235 14875
rect 24685 14841 24719 14875
rect 1685 14773 1719 14807
rect 4997 14773 5031 14807
rect 6193 14773 6227 14807
rect 7849 14773 7883 14807
rect 8309 14773 8343 14807
rect 11897 14773 11931 14807
rect 12587 14773 12621 14807
rect 17785 14773 17819 14807
rect 18429 14773 18463 14807
rect 20361 14773 20395 14807
rect 21741 14773 21775 14807
rect 25513 14773 25547 14807
rect 1777 14569 1811 14603
rect 2973 14569 3007 14603
rect 3617 14569 3651 14603
rect 5457 14569 5491 14603
rect 6929 14569 6963 14603
rect 7205 14569 7239 14603
rect 8493 14569 8527 14603
rect 9505 14569 9539 14603
rect 10793 14569 10827 14603
rect 14197 14569 14231 14603
rect 14657 14569 14691 14603
rect 16957 14569 16991 14603
rect 18981 14569 19015 14603
rect 20545 14569 20579 14603
rect 22109 14569 22143 14603
rect 23673 14569 23707 14603
rect 2053 14501 2087 14535
rect 4169 14501 4203 14535
rect 4261 14501 4295 14535
rect 7665 14501 7699 14535
rect 9873 14501 9907 14535
rect 10425 14501 10459 14535
rect 11805 14501 11839 14535
rect 13369 14501 13403 14535
rect 13921 14501 13955 14535
rect 15485 14501 15519 14535
rect 18705 14501 18739 14535
rect 19441 14501 19475 14535
rect 21097 14501 21131 14535
rect 21649 14501 21683 14535
rect 22385 14501 22419 14535
rect 23305 14501 23339 14535
rect 24225 14501 24259 14535
rect 24317 14501 24351 14535
rect 5641 14433 5675 14467
rect 6101 14433 6135 14467
rect 17141 14433 17175 14467
rect 17325 14433 17359 14467
rect 22845 14433 22879 14467
rect 23121 14433 23155 14467
rect 1961 14365 1995 14399
rect 2605 14365 2639 14399
rect 5181 14365 5215 14399
rect 6377 14365 6411 14399
rect 7573 14365 7607 14399
rect 9781 14365 9815 14399
rect 11713 14365 11747 14399
rect 12357 14365 12391 14399
rect 13277 14365 13311 14399
rect 15393 14365 15427 14399
rect 15669 14365 15703 14399
rect 19349 14365 19383 14399
rect 19993 14365 20027 14399
rect 21005 14365 21039 14399
rect 24869 14365 24903 14399
rect 4721 14297 4755 14331
rect 8125 14297 8159 14331
rect 8861 14229 8895 14263
rect 2697 14025 2731 14059
rect 2973 14025 3007 14059
rect 4445 14025 4479 14059
rect 9689 14025 9723 14059
rect 9965 14025 9999 14059
rect 11805 14025 11839 14059
rect 13369 14025 13403 14059
rect 15393 14025 15427 14059
rect 17233 14025 17267 14059
rect 17601 14025 17635 14059
rect 19533 14025 19567 14059
rect 19901 14025 19935 14059
rect 20821 14025 20855 14059
rect 21925 14025 21959 14059
rect 22937 14025 22971 14059
rect 24593 14025 24627 14059
rect 24869 14025 24903 14059
rect 25559 14025 25593 14059
rect 4721 13957 4755 13991
rect 5457 13957 5491 13991
rect 9229 13957 9263 13991
rect 22385 13957 22419 13991
rect 1777 13889 1811 13923
rect 5089 13889 5123 13923
rect 6837 13889 6871 13923
rect 8033 13889 8067 13923
rect 8677 13889 8711 13923
rect 10241 13889 10275 13923
rect 12449 13889 12483 13923
rect 14289 13889 14323 13923
rect 14933 13889 14967 13923
rect 16221 13889 16255 13923
rect 16497 13889 16531 13923
rect 18613 13889 18647 13923
rect 21005 13889 21039 13923
rect 23673 13889 23707 13923
rect 3525 13821 3559 13855
rect 5265 13821 5299 13855
rect 5825 13821 5859 13855
rect 11529 13821 11563 13855
rect 21649 13821 21683 13855
rect 22477 13821 22511 13855
rect 25456 13821 25490 13855
rect 25881 13821 25915 13855
rect 1685 13753 1719 13787
rect 2098 13753 2132 13787
rect 3341 13753 3375 13787
rect 3846 13753 3880 13787
rect 6561 13753 6595 13787
rect 7158 13753 7192 13787
rect 8769 13753 8803 13787
rect 10333 13753 10367 13787
rect 10885 13753 10919 13787
rect 12770 13753 12804 13787
rect 14381 13753 14415 13787
rect 16037 13753 16071 13787
rect 16313 13753 16347 13787
rect 18934 13753 18968 13787
rect 20453 13753 20487 13787
rect 21097 13753 21131 13787
rect 23994 13753 24028 13787
rect 6193 13685 6227 13719
rect 7757 13685 7791 13719
rect 8401 13685 8435 13719
rect 12173 13685 12207 13719
rect 13645 13685 13679 13719
rect 14013 13685 14047 13719
rect 18429 13685 18463 13719
rect 22661 13685 22695 13719
rect 23397 13685 23431 13719
rect 1777 13481 1811 13515
rect 3065 13481 3099 13515
rect 3709 13481 3743 13515
rect 5181 13481 5215 13515
rect 5641 13481 5675 13515
rect 7297 13481 7331 13515
rect 7665 13481 7699 13515
rect 8309 13481 8343 13515
rect 8953 13481 8987 13515
rect 9505 13481 9539 13515
rect 10701 13481 10735 13515
rect 11713 13481 11747 13515
rect 12265 13481 12299 13515
rect 12817 13481 12851 13515
rect 13461 13481 13495 13515
rect 15025 13481 15059 13515
rect 16221 13481 16255 13515
rect 19349 13481 19383 13515
rect 21833 13481 21867 13515
rect 24685 13481 24719 13515
rect 25145 13481 25179 13515
rect 6698 13413 6732 13447
rect 9873 13413 9907 13447
rect 10425 13413 10459 13447
rect 13829 13413 13863 13447
rect 16773 13413 16807 13447
rect 16865 13413 16899 13447
rect 18337 13413 18371 13447
rect 18429 13413 18463 13447
rect 21275 13413 21309 13447
rect 23851 13413 23885 13447
rect 1961 13345 1995 13379
rect 2513 13345 2547 13379
rect 4353 13345 4387 13379
rect 4537 13345 4571 13379
rect 4813 13345 4847 13379
rect 7941 13345 7975 13379
rect 8125 13345 8159 13379
rect 15301 13345 15335 13379
rect 19809 13345 19843 13379
rect 23489 13345 23523 13379
rect 25237 13345 25271 13379
rect 2329 13277 2363 13311
rect 6377 13277 6411 13311
rect 8585 13277 8619 13311
rect 9781 13277 9815 13311
rect 11897 13277 11931 13311
rect 13737 13277 13771 13311
rect 14013 13277 14047 13311
rect 17049 13277 17083 13311
rect 20913 13277 20947 13311
rect 15485 13209 15519 13243
rect 18889 13209 18923 13243
rect 19993 13209 20027 13243
rect 3341 13141 3375 13175
rect 6193 13141 6227 13175
rect 13093 13141 13127 13175
rect 15853 13141 15887 13175
rect 20729 13141 20763 13175
rect 22477 13141 22511 13175
rect 24409 13141 24443 13175
rect 25421 13141 25455 13175
rect 1961 12937 1995 12971
rect 2329 12937 2363 12971
rect 2789 12937 2823 12971
rect 4353 12937 4387 12971
rect 6469 12937 6503 12971
rect 7021 12937 7055 12971
rect 10885 12937 10919 12971
rect 13645 12937 13679 12971
rect 17233 12937 17267 12971
rect 17877 12937 17911 12971
rect 18337 12937 18371 12971
rect 20177 12937 20211 12971
rect 21741 12937 21775 12971
rect 23489 12937 23523 12971
rect 23857 12937 23891 12971
rect 25421 12937 25455 12971
rect 4629 12869 4663 12903
rect 10517 12869 10551 12903
rect 15485 12869 15519 12903
rect 16589 12869 16623 12903
rect 22109 12869 22143 12903
rect 24961 12869 24995 12903
rect 1832 12801 1866 12835
rect 2053 12801 2087 12835
rect 3065 12801 3099 12835
rect 5917 12801 5951 12835
rect 7941 12801 7975 12835
rect 8125 12801 8159 12835
rect 9965 12801 9999 12835
rect 12541 12801 12575 12835
rect 15117 12801 15151 12835
rect 20821 12801 20855 12835
rect 21097 12801 21131 12835
rect 24409 12801 24443 12835
rect 1685 12733 1719 12767
rect 3249 12733 3283 12767
rect 3709 12733 3743 12767
rect 5089 12733 5123 12767
rect 5365 12733 5399 12767
rect 5733 12733 5767 12767
rect 6837 12733 6871 12767
rect 9045 12733 9079 12767
rect 14105 12733 14139 12767
rect 14565 12733 14599 12767
rect 15669 12733 15703 12767
rect 18981 12733 19015 12767
rect 22360 12733 22394 12767
rect 8447 12665 8481 12699
rect 9413 12665 9447 12699
rect 10057 12665 10091 12699
rect 12633 12665 12667 12699
rect 13185 12665 13219 12699
rect 13921 12665 13955 12699
rect 14841 12665 14875 12699
rect 15990 12665 16024 12699
rect 18797 12665 18831 12699
rect 19302 12665 19336 12699
rect 20545 12665 20579 12699
rect 20913 12665 20947 12699
rect 24501 12665 24535 12699
rect 3341 12597 3375 12631
rect 7573 12597 7607 12631
rect 9781 12597 9815 12631
rect 11529 12597 11563 12631
rect 11897 12597 11931 12631
rect 16865 12597 16899 12631
rect 19901 12597 19935 12631
rect 22431 12597 22465 12631
rect 22845 12597 22879 12631
rect 3249 12393 3283 12427
rect 4721 12393 4755 12427
rect 7021 12393 7055 12427
rect 8033 12393 8067 12427
rect 9413 12393 9447 12427
rect 10793 12393 10827 12427
rect 11529 12393 11563 12427
rect 14473 12393 14507 12427
rect 17693 12393 17727 12427
rect 21051 12393 21085 12427
rect 21373 12393 21407 12427
rect 24409 12393 24443 12427
rect 2145 12325 2179 12359
rect 2237 12325 2271 12359
rect 4077 12325 4111 12359
rect 5733 12325 5767 12359
rect 7481 12325 7515 12359
rect 9781 12325 9815 12359
rect 9873 12325 9907 12359
rect 13001 12325 13035 12359
rect 14197 12325 14231 12359
rect 16174 12325 16208 12359
rect 19441 12325 19475 12359
rect 19993 12325 20027 12359
rect 22477 12325 22511 12359
rect 24685 12325 24719 12359
rect 25237 12325 25271 12359
rect 2329 12257 2363 12291
rect 5365 12257 5399 12291
rect 6009 12257 6043 12291
rect 6469 12257 6503 12291
rect 8861 12257 8895 12291
rect 11529 12257 11563 12291
rect 11805 12257 11839 12291
rect 17601 12257 17635 12291
rect 18153 12257 18187 12291
rect 20980 12257 21014 12291
rect 4224 12189 4258 12223
rect 4445 12189 4479 12223
rect 6653 12189 6687 12223
rect 7665 12189 7699 12223
rect 10149 12189 10183 12223
rect 12909 12189 12943 12223
rect 15853 12189 15887 12223
rect 19349 12189 19383 12223
rect 22385 12189 22419 12223
rect 22661 12189 22695 12223
rect 24593 12189 24627 12223
rect 8585 12121 8619 12155
rect 13461 12121 13495 12155
rect 19073 12121 19107 12155
rect 1777 12053 1811 12087
rect 3893 12053 3927 12087
rect 4353 12053 4387 12087
rect 12541 12053 12575 12087
rect 15669 12053 15703 12087
rect 16773 12053 16807 12087
rect 17049 12053 17083 12087
rect 18613 12053 18647 12087
rect 21925 12053 21959 12087
rect 2053 11849 2087 11883
rect 2513 11849 2547 11883
rect 2881 11849 2915 11883
rect 4077 11849 4111 11883
rect 4445 11849 4479 11883
rect 5641 11849 5675 11883
rect 6561 11849 6595 11883
rect 10241 11849 10275 11883
rect 12173 11849 12207 11883
rect 14105 11849 14139 11883
rect 19533 11849 19567 11883
rect 22937 11849 22971 11883
rect 24225 11849 24259 11883
rect 25421 11849 25455 11883
rect 3249 11781 3283 11815
rect 3709 11781 3743 11815
rect 4905 11781 4939 11815
rect 8769 11781 8803 11815
rect 17325 11781 17359 11815
rect 23305 11781 23339 11815
rect 25053 11781 25087 11815
rect 2384 11713 2418 11747
rect 2605 11713 2639 11747
rect 4169 11713 4203 11747
rect 7757 11713 7791 11747
rect 9321 11713 9355 11747
rect 9965 11713 9999 11747
rect 12725 11713 12759 11747
rect 15301 11713 15335 11747
rect 15853 11713 15887 11747
rect 16221 11713 16255 11747
rect 16497 11713 16531 11747
rect 17601 11713 17635 11747
rect 20453 11713 20487 11747
rect 20729 11713 20763 11747
rect 22661 11713 22695 11747
rect 24501 11713 24535 11747
rect 1777 11645 1811 11679
rect 2237 11645 2271 11679
rect 3948 11645 3982 11679
rect 5365 11645 5399 11679
rect 5549 11645 5583 11679
rect 6193 11645 6227 11679
rect 8401 11645 8435 11679
rect 10793 11645 10827 11679
rect 11253 11645 11287 11679
rect 14473 11645 14507 11679
rect 14749 11645 14783 11679
rect 15117 11645 15151 11679
rect 18521 11645 18555 11679
rect 18981 11645 19015 11679
rect 3801 11577 3835 11611
rect 5181 11577 5215 11611
rect 7849 11577 7883 11611
rect 9413 11577 9447 11611
rect 11529 11577 11563 11611
rect 12817 11577 12851 11611
rect 13369 11577 13403 11611
rect 16313 11577 16347 11611
rect 20545 11577 20579 11611
rect 22017 11577 22051 11611
rect 22109 11577 22143 11611
rect 24593 11577 24627 11611
rect 7205 11509 7239 11543
rect 7573 11509 7607 11543
rect 9045 11509 9079 11543
rect 10609 11509 10643 11543
rect 11897 11509 11931 11543
rect 13645 11509 13679 11543
rect 18337 11509 18371 11543
rect 18797 11509 18831 11543
rect 20269 11509 20303 11543
rect 21465 11509 21499 11543
rect 21741 11509 21775 11543
rect 23949 11509 23983 11543
rect 3801 11305 3835 11339
rect 5457 11305 5491 11339
rect 5825 11305 5859 11339
rect 6101 11305 6135 11339
rect 7573 11305 7607 11339
rect 8585 11305 8619 11339
rect 9321 11305 9355 11339
rect 14013 11305 14047 11339
rect 14657 11305 14691 11339
rect 15531 11305 15565 11339
rect 16221 11305 16255 11339
rect 18153 11305 18187 11339
rect 18889 11305 18923 11339
rect 19441 11305 19475 11339
rect 20361 11305 20395 11339
rect 22293 11305 22327 11339
rect 22845 11305 22879 11339
rect 24869 11305 24903 11339
rect 3433 11237 3467 11271
rect 4813 11237 4847 11271
rect 6469 11237 6503 11271
rect 7015 11237 7049 11271
rect 9873 11237 9907 11271
rect 11615 11237 11649 11271
rect 13185 11237 13219 11271
rect 13737 11237 13771 11271
rect 16589 11237 16623 11271
rect 18521 11237 18555 11271
rect 23994 11237 24028 11271
rect 1409 11169 1443 11203
rect 2421 11169 2455 11203
rect 2881 11169 2915 11203
rect 4077 11169 4111 11203
rect 5641 11169 5675 11203
rect 6653 11169 6687 11203
rect 8217 11169 8251 11203
rect 8401 11169 8435 11203
rect 15301 11169 15335 11203
rect 17969 11169 18003 11203
rect 19073 11169 19107 11203
rect 20821 11169 20855 11203
rect 24593 11169 24627 11203
rect 25456 11169 25490 11203
rect 1961 11101 1995 11135
rect 3157 11101 3191 11135
rect 4224 11101 4258 11135
rect 4445 11101 4479 11135
rect 5089 11101 5123 11135
rect 9781 11101 9815 11135
rect 10057 11101 10091 11135
rect 11253 11101 11287 11135
rect 13093 11101 13127 11135
rect 16497 11101 16531 11135
rect 16957 11101 16991 11135
rect 21925 11101 21959 11135
rect 23673 11101 23707 11135
rect 1593 11033 1627 11067
rect 2329 11033 2363 11067
rect 10793 11033 10827 11067
rect 12173 11033 12207 11067
rect 19993 11033 20027 11067
rect 25559 11033 25593 11067
rect 4353 10965 4387 10999
rect 7849 10965 7883 10999
rect 8861 10965 8895 10999
rect 12633 10965 12667 10999
rect 17509 10965 17543 10999
rect 21051 10965 21085 10999
rect 21373 10965 21407 10999
rect 1685 10761 1719 10795
rect 4261 10761 4295 10795
rect 4813 10761 4847 10795
rect 5273 10761 5307 10795
rect 6653 10761 6687 10795
rect 14105 10761 14139 10795
rect 15945 10761 15979 10795
rect 17877 10761 17911 10795
rect 21649 10761 21683 10795
rect 23489 10761 23523 10795
rect 24593 10761 24627 10795
rect 25237 10761 25271 10795
rect 25605 10761 25639 10795
rect 3617 10693 3651 10727
rect 3939 10693 3973 10727
rect 4077 10693 4111 10727
rect 22615 10693 22649 10727
rect 3249 10625 3283 10659
rect 4169 10625 4203 10659
rect 6193 10625 6227 10659
rect 7113 10625 7147 10659
rect 9229 10625 9263 10659
rect 12817 10625 12851 10659
rect 13645 10625 13679 10659
rect 14381 10625 14415 10659
rect 14657 10625 14691 10659
rect 16129 10625 16163 10659
rect 19901 10625 19935 10659
rect 20729 10625 20763 10659
rect 2053 10557 2087 10591
rect 2329 10557 2363 10591
rect 3801 10557 3835 10591
rect 5549 10557 5583 10591
rect 8033 10557 8067 10591
rect 10149 10557 10183 10591
rect 10609 10557 10643 10591
rect 11529 10557 11563 10591
rect 12173 10557 12207 10591
rect 5365 10489 5399 10523
rect 7434 10489 7468 10523
rect 8953 10489 8987 10523
rect 9045 10489 9079 10523
rect 10517 10489 10551 10523
rect 10930 10489 10964 10523
rect 11805 10489 11839 10523
rect 12909 10489 12943 10523
rect 13461 10489 13495 10523
rect 15485 10557 15519 10591
rect 18188 10557 18222 10591
rect 18613 10557 18647 10591
rect 19257 10557 19291 10591
rect 19625 10557 19659 10591
rect 22544 10557 22578 10591
rect 22937 10557 22971 10591
rect 23673 10557 23707 10591
rect 24869 10557 24903 10591
rect 25421 10557 25455 10591
rect 25973 10557 26007 10591
rect 13737 10489 13771 10523
rect 14473 10489 14507 10523
rect 16450 10489 16484 10523
rect 18981 10489 19015 10523
rect 20177 10489 20211 10523
rect 21050 10489 21084 10523
rect 21925 10489 21959 10523
rect 23994 10489 24028 10523
rect 2513 10421 2547 10455
rect 5641 10421 5675 10455
rect 8401 10421 8435 10455
rect 13645 10421 13679 10455
rect 17049 10421 17083 10455
rect 17325 10421 17359 10455
rect 18291 10421 18325 10455
rect 20637 10421 20671 10455
rect 22293 10421 22327 10455
rect 4721 10217 4755 10251
rect 5733 10217 5767 10251
rect 7389 10217 7423 10251
rect 9873 10217 9907 10251
rect 10241 10217 10275 10251
rect 11161 10217 11195 10251
rect 11529 10217 11563 10251
rect 12357 10217 12391 10251
rect 14013 10217 14047 10251
rect 15623 10217 15657 10251
rect 18245 10217 18279 10251
rect 19809 10217 19843 10251
rect 23765 10217 23799 10251
rect 24593 10217 24627 10251
rect 7113 10149 7147 10183
rect 12633 10149 12667 10183
rect 13093 10149 13127 10183
rect 14381 10149 14415 10183
rect 16129 10149 16163 10183
rect 16681 10149 16715 10183
rect 18521 10149 18555 10183
rect 18613 10149 18647 10183
rect 21097 10149 21131 10183
rect 23489 10149 23523 10183
rect 24133 10149 24167 10183
rect 1409 10081 1443 10115
rect 3065 10081 3099 10115
rect 4077 10081 4111 10115
rect 6101 10081 6135 10115
rect 6377 10081 6411 10115
rect 6837 10081 6871 10115
rect 7757 10081 7791 10115
rect 7941 10081 7975 10115
rect 8217 10081 8251 10115
rect 10149 10081 10183 10115
rect 10701 10081 10735 10115
rect 11713 10081 11747 10115
rect 15393 10081 15427 10115
rect 22753 10081 22787 10115
rect 23213 10081 23247 10115
rect 24317 10081 24351 10115
rect 24777 10081 24811 10115
rect 3157 10013 3191 10047
rect 4445 10013 4479 10047
rect 8401 10013 8435 10047
rect 13001 10013 13035 10047
rect 16589 10013 16623 10047
rect 18889 10013 18923 10047
rect 21005 10013 21039 10047
rect 21281 10013 21315 10047
rect 1593 9945 1627 9979
rect 4353 9945 4387 9979
rect 5365 9945 5399 9979
rect 8033 9945 8067 9979
rect 9321 9945 9355 9979
rect 11897 9945 11931 9979
rect 13553 9945 13587 9979
rect 17141 9945 17175 9979
rect 2145 9877 2179 9911
rect 3433 9877 3467 9911
rect 3893 9877 3927 9911
rect 4242 9877 4276 9911
rect 8953 9877 8987 9911
rect 19441 9877 19475 9911
rect 2053 9673 2087 9707
rect 3433 9673 3467 9707
rect 3847 9673 3881 9707
rect 4721 9673 4755 9707
rect 10149 9673 10183 9707
rect 12173 9673 12207 9707
rect 13645 9673 13679 9707
rect 21005 9673 21039 9707
rect 22753 9673 22787 9707
rect 25053 9673 25087 9707
rect 25421 9673 25455 9707
rect 2283 9605 2317 9639
rect 2421 9605 2455 9639
rect 3985 9605 4019 9639
rect 5089 9605 5123 9639
rect 9873 9605 9907 9639
rect 11805 9605 11839 9639
rect 2513 9537 2547 9571
rect 3433 9537 3467 9571
rect 4077 9537 4111 9571
rect 4445 9537 4479 9571
rect 7389 9537 7423 9571
rect 8861 9537 8895 9571
rect 12725 9537 12759 9571
rect 13001 9537 13035 9571
rect 14289 9537 14323 9571
rect 14749 9537 14783 9571
rect 15945 9537 15979 9571
rect 18337 9537 18371 9571
rect 20085 9537 20119 9571
rect 20361 9537 20395 9571
rect 22293 9537 22327 9571
rect 24225 9537 24259 9571
rect 1685 9469 1719 9503
rect 2145 9469 2179 9503
rect 3249 9469 3283 9503
rect 5273 9469 5307 9503
rect 5825 9469 5859 9503
rect 6837 9469 6871 9503
rect 7297 9469 7331 9503
rect 8401 9469 8435 9503
rect 8493 9469 8527 9503
rect 8677 9469 8711 9503
rect 10793 9469 10827 9503
rect 11253 9469 11287 9503
rect 16313 9469 16347 9503
rect 16405 9469 16439 9503
rect 16865 9469 16899 9503
rect 21557 9469 21591 9503
rect 22109 9469 22143 9503
rect 23397 9469 23431 9503
rect 23673 9469 23707 9503
rect 24133 9469 24167 9503
rect 25237 9469 25271 9503
rect 25789 9469 25823 9503
rect 3709 9401 3743 9435
rect 9413 9401 9447 9435
rect 11529 9401 11563 9435
rect 12817 9401 12851 9435
rect 14381 9401 14415 9435
rect 15577 9401 15611 9435
rect 17141 9401 17175 9435
rect 17877 9401 17911 9435
rect 18429 9401 18463 9435
rect 18981 9401 19015 9435
rect 19901 9401 19935 9435
rect 20177 9401 20211 9435
rect 24685 9401 24719 9435
rect 2789 9333 2823 9367
rect 3525 9333 3559 9367
rect 5457 9333 5491 9367
rect 6469 9333 6503 9367
rect 8033 9333 8067 9367
rect 10701 9333 10735 9367
rect 14013 9333 14047 9367
rect 19257 9333 19291 9367
rect 21373 9333 21407 9367
rect 2237 9129 2271 9163
rect 5917 9129 5951 9163
rect 6377 9129 6411 9163
rect 7481 9129 7515 9163
rect 10333 9129 10367 9163
rect 12173 9129 12207 9163
rect 13645 9129 13679 9163
rect 14565 9129 14599 9163
rect 16589 9129 16623 9163
rect 17969 9129 18003 9163
rect 18613 9129 18647 9163
rect 21097 9129 21131 9163
rect 22753 9129 22787 9163
rect 23121 9129 23155 9163
rect 24133 9129 24167 9163
rect 3157 9061 3191 9095
rect 10701 9061 10735 9095
rect 11247 9061 11281 9095
rect 12449 9061 12483 9095
rect 13046 9061 13080 9095
rect 14197 9061 14231 9095
rect 17370 9061 17404 9095
rect 19118 9061 19152 9095
rect 20085 9061 20119 9095
rect 20729 9061 20763 9095
rect 21649 9061 21683 9095
rect 24731 9061 24765 9095
rect 1409 8993 1443 9027
rect 2421 8993 2455 9027
rect 2697 8993 2731 9027
rect 6469 8993 6503 9027
rect 6745 8993 6779 9027
rect 8033 8993 8067 9027
rect 8309 8993 8343 9027
rect 9873 8993 9907 9027
rect 10885 8993 10919 9027
rect 15669 8993 15703 9027
rect 15945 8993 15979 9027
rect 18797 8993 18831 9027
rect 19717 8993 19751 9027
rect 23029 8993 23063 9027
rect 23489 8993 23523 9027
rect 24644 8993 24678 9027
rect 3893 8925 3927 8959
rect 4445 8925 4479 8959
rect 5089 8925 5123 8959
rect 5457 8925 5491 8959
rect 6929 8925 6963 8959
rect 8769 8925 8803 8959
rect 12725 8925 12759 8959
rect 16221 8925 16255 8959
rect 17049 8925 17083 8959
rect 21557 8925 21591 8959
rect 21833 8925 21867 8959
rect 2513 8857 2547 8891
rect 4215 8857 4249 8891
rect 6561 8857 6595 8891
rect 8125 8857 8159 8891
rect 10057 8857 10091 8891
rect 16957 8857 16991 8891
rect 1593 8789 1627 8823
rect 3709 8789 3743 8823
rect 4353 8789 4387 8823
rect 4537 8789 4571 8823
rect 7849 8789 7883 8823
rect 9045 8789 9079 8823
rect 11805 8789 11839 8823
rect 18337 8789 18371 8823
rect 2421 8585 2455 8619
rect 3157 8585 3191 8619
rect 4077 8585 4111 8619
rect 5549 8585 5583 8619
rect 8033 8585 8067 8619
rect 10701 8585 10735 8619
rect 12265 8585 12299 8619
rect 17233 8585 17267 8619
rect 19165 8585 19199 8619
rect 19625 8585 19659 8619
rect 20913 8585 20947 8619
rect 22293 8585 22327 8619
rect 22661 8585 22695 8619
rect 25421 8585 25455 8619
rect 5181 8517 5215 8551
rect 5917 8517 5951 8551
rect 11437 8517 11471 8551
rect 16129 8517 16163 8551
rect 20361 8517 20395 8551
rect 23397 8517 23431 8551
rect 4261 8449 4295 8483
rect 9965 8449 9999 8483
rect 12449 8449 12483 8483
rect 13645 8449 13679 8483
rect 14289 8449 14323 8483
rect 14565 8449 14599 8483
rect 16957 8449 16991 8483
rect 17601 8449 17635 8483
rect 18889 8449 18923 8483
rect 19809 8449 19843 8483
rect 21373 8449 21407 8483
rect 24041 8449 24075 8483
rect 1501 8381 1535 8415
rect 2973 8381 3007 8415
rect 5733 8381 5767 8415
rect 7389 8381 7423 8415
rect 8401 8381 8435 8415
rect 9229 8381 9263 8415
rect 9689 8381 9723 8415
rect 13369 8381 13403 8415
rect 14013 8381 14047 8415
rect 16497 8381 16531 8415
rect 16681 8381 16715 8415
rect 25237 8381 25271 8415
rect 25789 8381 25823 8415
rect 4353 8313 4387 8347
rect 4905 8313 4939 8347
rect 6837 8313 6871 8347
rect 10333 8313 10367 8347
rect 10885 8313 10919 8347
rect 10977 8313 11011 8347
rect 11805 8313 11839 8347
rect 12770 8313 12804 8347
rect 14381 8313 14415 8347
rect 18245 8313 18279 8347
rect 18337 8313 18371 8347
rect 19901 8313 19935 8347
rect 21694 8313 21728 8347
rect 23765 8313 23799 8347
rect 23857 8313 23891 8347
rect 1869 8245 1903 8279
rect 2881 8245 2915 8279
rect 3617 8245 3651 8279
rect 6561 8245 6595 8279
rect 9137 8245 9171 8279
rect 15577 8245 15611 8279
rect 21189 8245 21223 8279
rect 23029 8245 23063 8279
rect 24777 8245 24811 8279
rect 1593 8041 1627 8075
rect 2237 8041 2271 8075
rect 3525 8041 3559 8075
rect 5733 8041 5767 8075
rect 6929 8041 6963 8075
rect 7941 8041 7975 8075
rect 9321 8041 9355 8075
rect 13553 8041 13587 8075
rect 15577 8041 15611 8075
rect 17325 8041 17359 8075
rect 18337 8041 18371 8075
rect 20637 8041 20671 8075
rect 24639 8041 24673 8075
rect 4330 7973 4364 8007
rect 5181 7973 5215 8007
rect 5365 7973 5399 8007
rect 8769 7973 8803 8007
rect 12678 7973 12712 8007
rect 13921 7973 13955 8007
rect 17738 7973 17772 8007
rect 18797 7973 18831 8007
rect 19349 7973 19383 8007
rect 21097 7973 21131 8007
rect 21649 7973 21683 8007
rect 23074 7973 23108 8007
rect 1409 7905 1443 7939
rect 2697 7905 2731 7939
rect 2973 7905 3007 7939
rect 3157 7837 3191 7871
rect 4077 7837 4111 7871
rect 6285 7905 6319 7939
rect 6469 7905 6503 7939
rect 6745 7905 6779 7939
rect 8033 7905 8067 7939
rect 8309 7905 8343 7939
rect 9689 7905 9723 7939
rect 10793 7905 10827 7939
rect 11253 7905 11287 7939
rect 14105 7905 14139 7939
rect 15577 7905 15611 7939
rect 15853 7905 15887 7939
rect 23673 7905 23707 7939
rect 24317 7905 24351 7939
rect 24568 7905 24602 7939
rect 11529 7837 11563 7871
rect 12357 7837 12391 7871
rect 17417 7837 17451 7871
rect 19257 7837 19291 7871
rect 19533 7837 19567 7871
rect 21005 7837 21039 7871
rect 22753 7837 22787 7871
rect 1869 7769 1903 7803
rect 5181 7769 5215 7803
rect 6561 7769 6595 7803
rect 7481 7769 7515 7803
rect 8125 7769 8159 7803
rect 10609 7769 10643 7803
rect 15025 7769 15059 7803
rect 3893 7701 3927 7735
rect 4997 7701 5031 7735
rect 9873 7701 9907 7735
rect 13277 7701 13311 7735
rect 14289 7701 14323 7735
rect 16405 7701 16439 7735
rect 20177 7701 20211 7735
rect 22017 7701 22051 7735
rect 22661 7701 22695 7735
rect 24041 7701 24075 7735
rect 1593 7497 1627 7531
rect 1961 7497 1995 7531
rect 5917 7497 5951 7531
rect 7205 7497 7239 7531
rect 7481 7497 7515 7531
rect 9689 7497 9723 7531
rect 12173 7497 12207 7531
rect 12633 7497 12667 7531
rect 13277 7497 13311 7531
rect 14381 7497 14415 7531
rect 16037 7497 16071 7531
rect 16405 7497 16439 7531
rect 19441 7497 19475 7531
rect 21465 7497 21499 7531
rect 23029 7497 23063 7531
rect 2513 7429 2547 7463
rect 5641 7429 5675 7463
rect 19165 7429 19199 7463
rect 25375 7429 25409 7463
rect 9321 7361 9355 7395
rect 10609 7361 10643 7395
rect 13461 7361 13495 7395
rect 17509 7361 17543 7395
rect 18797 7361 18831 7395
rect 20545 7361 20579 7395
rect 23397 7361 23431 7395
rect 1409 7293 1443 7327
rect 2881 7293 2915 7327
rect 3157 7293 3191 7327
rect 4261 7293 4295 7327
rect 4721 7293 4755 7327
rect 5733 7293 5767 7327
rect 7297 7293 7331 7327
rect 8125 7293 8159 7327
rect 8309 7293 8343 7327
rect 8401 7293 8435 7327
rect 8585 7293 8619 7327
rect 10793 7293 10827 7327
rect 11253 7293 11287 7327
rect 11805 7293 11839 7327
rect 14841 7293 14875 7327
rect 15209 7293 15243 7327
rect 15393 7293 15427 7327
rect 16716 7293 16750 7327
rect 17141 7293 17175 7327
rect 22017 7293 22051 7327
rect 22477 7293 22511 7327
rect 23673 7293 23707 7327
rect 24133 7293 24167 7327
rect 25272 7293 25306 7327
rect 25697 7293 25731 7327
rect 3709 7225 3743 7259
rect 9045 7225 9079 7259
rect 11529 7225 11563 7259
rect 13553 7225 13587 7259
rect 14105 7225 14139 7259
rect 15669 7225 15703 7259
rect 16819 7225 16853 7259
rect 18153 7225 18187 7259
rect 18245 7225 18279 7259
rect 20637 7225 20671 7259
rect 21189 7225 21223 7259
rect 22753 7225 22787 7259
rect 2697 7157 2731 7191
rect 4077 7157 4111 7191
rect 4445 7157 4479 7191
rect 5181 7157 5215 7191
rect 6469 7157 6503 7191
rect 10241 7157 10275 7191
rect 19809 7157 19843 7191
rect 20361 7157 20395 7191
rect 21833 7157 21867 7191
rect 23765 7157 23799 7191
rect 24685 7157 24719 7191
rect 1685 6953 1719 6987
rect 3709 6953 3743 6987
rect 4261 6953 4295 6987
rect 6101 6953 6135 6987
rect 8309 6953 8343 6987
rect 11437 6953 11471 6987
rect 12633 6953 12667 6987
rect 15025 6953 15059 6987
rect 17969 6953 18003 6987
rect 18797 6953 18831 6987
rect 19671 6953 19705 6987
rect 21833 6953 21867 6987
rect 23581 6953 23615 6987
rect 2421 6885 2455 6919
rect 5181 6885 5215 6919
rect 6377 6885 6411 6919
rect 7573 6885 7607 6919
rect 8953 6885 8987 6919
rect 13369 6885 13403 6919
rect 19165 6885 19199 6919
rect 20269 6885 20303 6919
rect 21234 6885 21268 6919
rect 22982 6885 23016 6919
rect 24501 6885 24535 6919
rect 24593 6885 24627 6919
rect 2145 6817 2179 6851
rect 6561 6817 6595 6851
rect 7021 6817 7055 6851
rect 7941 6817 7975 6851
rect 8125 6817 8159 6851
rect 10057 6817 10091 6851
rect 10609 6817 10643 6851
rect 11897 6817 11931 6851
rect 12173 6817 12207 6851
rect 15577 6817 15611 6851
rect 15761 6817 15795 6851
rect 17601 6817 17635 6851
rect 18521 6817 18555 6851
rect 19441 6817 19475 6851
rect 2053 6749 2087 6783
rect 5089 6749 5123 6783
rect 7113 6749 7147 6783
rect 10793 6749 10827 6783
rect 12357 6749 12391 6783
rect 13277 6749 13311 6783
rect 13553 6749 13587 6783
rect 15853 6749 15887 6783
rect 20913 6749 20947 6783
rect 22661 6749 22695 6783
rect 24777 6749 24811 6783
rect 5641 6681 5675 6715
rect 17417 6681 17451 6715
rect 3065 6613 3099 6647
rect 3433 6613 3467 6647
rect 4721 6613 4755 6647
rect 8677 6613 8711 6647
rect 11069 6613 11103 6647
rect 20637 6613 20671 6647
rect 23857 6613 23891 6647
rect 1593 6409 1627 6443
rect 3433 6409 3467 6443
rect 5273 6409 5307 6443
rect 6285 6409 6319 6443
rect 11897 6409 11931 6443
rect 12265 6409 12299 6443
rect 13645 6409 13679 6443
rect 16681 6409 16715 6443
rect 18291 6409 18325 6443
rect 21005 6409 21039 6443
rect 23029 6409 23063 6443
rect 24685 6409 24719 6443
rect 25053 6409 25087 6443
rect 25513 6409 25547 6443
rect 11529 6341 11563 6375
rect 15301 6341 15335 6375
rect 17601 6341 17635 6375
rect 22753 6341 22787 6375
rect 23489 6341 23523 6375
rect 2789 6273 2823 6307
rect 3893 6273 3927 6307
rect 4353 6273 4387 6307
rect 5917 6273 5951 6307
rect 7021 6273 7055 6307
rect 8861 6273 8895 6307
rect 9137 6273 9171 6307
rect 12449 6273 12483 6307
rect 15393 6273 15427 6307
rect 16957 6273 16991 6307
rect 19073 6273 19107 6307
rect 1409 6205 1443 6239
rect 8217 6205 8251 6239
rect 10701 6205 10735 6239
rect 10885 6205 10919 6239
rect 14232 6205 14266 6239
rect 14657 6205 14691 6239
rect 18220 6205 18254 6239
rect 18705 6205 18739 6239
rect 19349 6205 19383 6239
rect 19625 6205 19659 6239
rect 21465 6205 21499 6239
rect 21833 6205 21867 6239
rect 22017 6205 22051 6239
rect 23673 6205 23707 6239
rect 24225 6205 24259 6239
rect 25272 6205 25306 6239
rect 25697 6205 25731 6239
rect 2513 6137 2547 6171
rect 2605 6137 2639 6171
rect 4674 6137 4708 6171
rect 6561 6137 6595 6171
rect 7342 6137 7376 6171
rect 8585 6137 8619 6171
rect 8953 6137 8987 6171
rect 11161 6137 11195 6171
rect 12770 6137 12804 6171
rect 14013 6137 14047 6171
rect 15714 6137 15748 6171
rect 19901 6137 19935 6171
rect 20637 6137 20671 6171
rect 2237 6069 2271 6103
rect 4169 6069 4203 6103
rect 7941 6069 7975 6103
rect 10057 6069 10091 6103
rect 13369 6069 13403 6103
rect 14335 6069 14369 6103
rect 16313 6069 16347 6103
rect 20177 6069 20211 6103
rect 21833 6069 21867 6103
rect 23765 6069 23799 6103
rect 1547 5865 1581 5899
rect 2145 5865 2179 5899
rect 2881 5865 2915 5899
rect 3525 5865 3559 5899
rect 3893 5865 3927 5899
rect 5365 5865 5399 5899
rect 5733 5865 5767 5899
rect 7113 5865 7147 5899
rect 9045 5865 9079 5899
rect 11713 5865 11747 5899
rect 12725 5865 12759 5899
rect 15577 5865 15611 5899
rect 17509 5865 17543 5899
rect 18429 5865 18463 5899
rect 19257 5865 19291 5899
rect 20177 5865 20211 5899
rect 24133 5865 24167 5899
rect 4490 5797 4524 5831
rect 6101 5797 6135 5831
rect 8217 5797 8251 5831
rect 10425 5797 10459 5831
rect 12167 5797 12201 5831
rect 13737 5797 13771 5831
rect 15990 5797 16024 5831
rect 22655 5797 22689 5831
rect 23765 5797 23799 5831
rect 1409 5729 1443 5763
rect 3065 5729 3099 5763
rect 5089 5729 5123 5763
rect 14289 5729 14323 5763
rect 15669 5729 15703 5763
rect 17417 5729 17451 5763
rect 17969 5729 18003 5763
rect 19165 5729 19199 5763
rect 19717 5729 19751 5763
rect 21281 5729 21315 5763
rect 22293 5729 22327 5763
rect 24225 5729 24259 5763
rect 24593 5729 24627 5763
rect 4169 5661 4203 5695
rect 6009 5661 6043 5695
rect 6469 5661 6503 5695
rect 7941 5661 7975 5695
rect 8125 5661 8159 5695
rect 10333 5661 10367 5695
rect 11805 5661 11839 5695
rect 13645 5661 13679 5695
rect 21741 5661 21775 5695
rect 7573 5593 7607 5627
rect 8677 5593 8711 5627
rect 10885 5593 10919 5627
rect 13369 5593 13403 5627
rect 21419 5593 21453 5627
rect 10149 5525 10183 5559
rect 14565 5525 14599 5559
rect 16589 5525 16623 5559
rect 23213 5525 23247 5559
rect 1593 5321 1627 5355
rect 2513 5321 2547 5355
rect 4629 5321 4663 5355
rect 6009 5321 6043 5355
rect 7849 5321 7883 5355
rect 10885 5321 10919 5355
rect 11897 5321 11931 5355
rect 12173 5321 12207 5355
rect 13737 5321 13771 5355
rect 15393 5321 15427 5355
rect 17417 5321 17451 5355
rect 17877 5321 17911 5355
rect 18337 5321 18371 5355
rect 18567 5321 18601 5355
rect 23029 5321 23063 5355
rect 23397 5321 23431 5355
rect 24685 5321 24719 5355
rect 5365 5253 5399 5287
rect 7481 5253 7515 5287
rect 11253 5253 11287 5287
rect 20729 5253 20763 5287
rect 3893 5185 3927 5219
rect 4813 5185 4847 5219
rect 6285 5185 6319 5219
rect 7067 5185 7101 5219
rect 8953 5185 8987 5219
rect 9597 5185 9631 5219
rect 9873 5185 9907 5219
rect 12449 5185 12483 5219
rect 14289 5185 14323 5219
rect 14933 5185 14967 5219
rect 15669 5185 15703 5219
rect 16313 5185 16347 5219
rect 19533 5185 19567 5219
rect 21833 5185 21867 5219
rect 24041 5185 24075 5219
rect 25237 5185 25271 5219
rect 1409 5117 1443 5151
rect 1961 5117 1995 5151
rect 3065 5117 3099 5151
rect 3433 5117 3467 5151
rect 3709 5117 3743 5151
rect 6964 5117 6998 5151
rect 11069 5117 11103 5151
rect 13369 5117 13403 5151
rect 14013 5117 14047 5151
rect 18464 5117 18498 5151
rect 18889 5117 18923 5151
rect 19441 5117 19475 5151
rect 21649 5117 21683 5151
rect 4905 5049 4939 5083
rect 8033 5049 8067 5083
rect 8125 5049 8159 5083
rect 8677 5049 8711 5083
rect 9413 5049 9447 5083
rect 9689 5049 9723 5083
rect 12770 5049 12804 5083
rect 14381 5049 14415 5083
rect 16129 5049 16163 5083
rect 16405 5049 16439 5083
rect 16957 5049 16991 5083
rect 19854 5049 19888 5083
rect 22154 5049 22188 5083
rect 23765 5049 23799 5083
rect 23857 5049 23891 5083
rect 4169 4981 4203 5015
rect 10609 4981 10643 5015
rect 20453 4981 20487 5015
rect 21281 4981 21315 5015
rect 22753 4981 22787 5015
rect 1593 4777 1627 4811
rect 2099 4777 2133 4811
rect 2513 4777 2547 4811
rect 3525 4777 3559 4811
rect 3893 4777 3927 4811
rect 7389 4777 7423 4811
rect 7941 4777 7975 4811
rect 8309 4777 8343 4811
rect 13001 4777 13035 4811
rect 15669 4777 15703 4811
rect 16773 4777 16807 4811
rect 19441 4777 19475 4811
rect 19993 4777 20027 4811
rect 21925 4777 21959 4811
rect 22293 4777 22327 4811
rect 24409 4777 24443 4811
rect 24777 4777 24811 4811
rect 3111 4709 3145 4743
rect 4905 4709 4939 4743
rect 5457 4709 5491 4743
rect 6009 4709 6043 4743
rect 11799 4709 11833 4743
rect 13461 4709 13495 4743
rect 13553 4709 13587 4743
rect 14105 4709 14139 4743
rect 15945 4709 15979 4743
rect 17646 4709 17680 4743
rect 21097 4709 21131 4743
rect 23029 4709 23063 4743
rect 1869 4641 1903 4675
rect 2973 4641 3007 4675
rect 9873 4641 9907 4675
rect 10333 4641 10367 4675
rect 10609 4641 10643 4675
rect 12633 4641 12667 4675
rect 17325 4641 17359 4675
rect 19073 4641 19107 4675
rect 24593 4641 24627 4675
rect 4813 4573 4847 4607
rect 7021 4573 7055 4607
rect 11437 4573 11471 4607
rect 15853 4573 15887 4607
rect 16221 4573 16255 4607
rect 21005 4573 21039 4607
rect 21281 4573 21315 4607
rect 22937 4573 22971 4607
rect 23213 4573 23247 4607
rect 10977 4505 11011 4539
rect 4261 4437 4295 4471
rect 8861 4437 8895 4471
rect 12357 4437 12391 4471
rect 14473 4437 14507 4471
rect 18245 4437 18279 4471
rect 18613 4437 18647 4471
rect 24133 4437 24167 4471
rect 1593 4233 1627 4267
rect 1961 4233 1995 4267
rect 2283 4233 2317 4267
rect 5089 4233 5123 4267
rect 5365 4233 5399 4267
rect 12173 4233 12207 4267
rect 13553 4233 13587 4267
rect 15393 4233 15427 4267
rect 17049 4233 17083 4267
rect 17877 4233 17911 4267
rect 19717 4233 19751 4267
rect 20913 4233 20947 4267
rect 23305 4233 23339 4267
rect 24823 4233 24857 4267
rect 25237 4233 25271 4267
rect 2973 4165 3007 4199
rect 9873 4165 9907 4199
rect 13369 4165 13403 4199
rect 19349 4165 19383 4199
rect 21603 4165 21637 4199
rect 24225 4165 24259 4199
rect 24593 4165 24627 4199
rect 2697 4097 2731 4131
rect 4169 4097 4203 4131
rect 8861 4097 8895 4131
rect 9137 4097 9171 4131
rect 10701 4097 10735 4131
rect 11529 4097 11563 4131
rect 12817 4097 12851 4131
rect 14381 4097 14415 4131
rect 15025 4097 15059 4131
rect 17325 4097 17359 4131
rect 18429 4097 18463 4131
rect 20637 4097 20671 4131
rect 22385 4097 22419 4131
rect 2212 4029 2246 4063
rect 3157 4029 3191 4063
rect 3617 4029 3651 4063
rect 7021 4029 7055 4063
rect 21532 4029 21566 4063
rect 21925 4029 21959 4063
rect 22512 4029 22546 4063
rect 22937 4029 22971 4063
rect 23740 4029 23774 4063
rect 24720 4029 24754 4063
rect 3985 3961 4019 3995
rect 4490 3961 4524 3995
rect 6285 3961 6319 3995
rect 7342 3961 7376 3995
rect 8953 3961 8987 3995
rect 10885 3961 10919 3995
rect 10977 3961 11011 3995
rect 12909 3961 12943 3995
rect 14197 3961 14231 3995
rect 14473 3961 14507 3995
rect 15945 3961 15979 3995
rect 16037 3961 16071 3995
rect 16589 3961 16623 3995
rect 18521 3961 18555 3995
rect 19073 3961 19107 3995
rect 19993 3961 20027 3995
rect 20085 3961 20119 3995
rect 21281 3961 21315 3995
rect 3341 3893 3375 3927
rect 6561 3893 6595 3927
rect 7941 3893 7975 3927
rect 8585 3893 8619 3927
rect 10241 3893 10275 3927
rect 11805 3893 11839 3927
rect 15761 3893 15795 3927
rect 22615 3893 22649 3927
rect 23811 3893 23845 3927
rect 4353 3689 4387 3723
rect 7205 3689 7239 3723
rect 12173 3689 12207 3723
rect 12817 3689 12851 3723
rect 14381 3689 14415 3723
rect 15853 3689 15887 3723
rect 16681 3689 16715 3723
rect 19487 3689 19521 3723
rect 19993 3689 20027 3723
rect 20269 3689 20303 3723
rect 24087 3689 24121 3723
rect 25145 3689 25179 3723
rect 6929 3621 6963 3655
rect 7573 3621 7607 3655
rect 8125 3621 8159 3655
rect 8677 3621 8711 3655
rect 11615 3621 11649 3655
rect 13185 3621 13219 3655
rect 17969 3621 18003 3655
rect 1961 3553 1995 3587
rect 2973 3553 3007 3587
rect 4169 3553 4203 3587
rect 4537 3553 4571 3587
rect 6193 3553 6227 3587
rect 6653 3553 6687 3587
rect 9689 3553 9723 3587
rect 10149 3553 10183 3587
rect 17693 3553 17727 3587
rect 19416 3553 19450 3587
rect 20980 3553 21014 3587
rect 21992 3553 22026 3587
rect 23004 3553 23038 3587
rect 24016 3553 24050 3587
rect 24961 3553 24995 3587
rect 8033 3485 8067 3519
rect 10425 3485 10459 3519
rect 11253 3485 11287 3519
rect 13093 3485 13127 3519
rect 15485 3485 15519 3519
rect 17877 3485 17911 3519
rect 3157 3417 3191 3451
rect 13645 3417 13679 3451
rect 14657 3417 14691 3451
rect 17693 3417 17727 3451
rect 18429 3417 18463 3451
rect 22063 3417 22097 3451
rect 23075 3417 23109 3451
rect 2145 3349 2179 3383
rect 5089 3349 5123 3383
rect 10701 3349 10735 3383
rect 11069 3349 11103 3383
rect 16405 3349 16439 3383
rect 21051 3349 21085 3383
rect 22477 3349 22511 3383
rect 1961 3145 1995 3179
rect 3065 3145 3099 3179
rect 4169 3145 4203 3179
rect 4491 3145 4525 3179
rect 6561 3145 6595 3179
rect 7941 3145 7975 3179
rect 8217 3145 8251 3179
rect 10057 3145 10091 3179
rect 12173 3145 12207 3179
rect 12725 3145 12759 3179
rect 14013 3145 14047 3179
rect 15117 3145 15151 3179
rect 16865 3145 16899 3179
rect 17877 3145 17911 3179
rect 18245 3145 18279 3179
rect 18889 3145 18923 3179
rect 20913 3145 20947 3179
rect 22017 3145 22051 3179
rect 23811 3145 23845 3179
rect 25145 3145 25179 3179
rect 3479 3077 3513 3111
rect 17233 3077 17267 3111
rect 19625 3077 19659 3111
rect 20269 3077 20303 3111
rect 23029 3077 23063 3111
rect 24225 3077 24259 3111
rect 3893 3009 3927 3043
rect 9781 3009 9815 3043
rect 10609 3009 10643 3043
rect 13001 3009 13035 3043
rect 13645 3009 13679 3043
rect 15945 3009 15979 3043
rect 16589 3009 16623 3043
rect 20913 3009 20947 3043
rect 25513 3009 25547 3043
rect 3408 2941 3442 2975
rect 4420 2941 4454 2975
rect 5549 2941 5583 2975
rect 5768 2941 5802 2975
rect 6193 2941 6227 2975
rect 6837 2941 6871 2975
rect 7389 2941 7423 2975
rect 8861 2941 8895 2975
rect 9045 2941 9079 2975
rect 9505 2941 9539 2975
rect 14473 2941 14507 2975
rect 18981 2941 19015 2975
rect 20085 2941 20119 2975
rect 21224 2941 21258 2975
rect 22268 2941 22302 2975
rect 23740 2941 23774 2975
rect 24501 2941 24535 2975
rect 24720 2941 24754 2975
rect 2329 2873 2363 2907
rect 10517 2873 10551 2907
rect 10971 2873 11005 2907
rect 13093 2873 13127 2907
rect 15485 2873 15519 2907
rect 16037 2873 16071 2907
rect 20729 2873 20763 2907
rect 24823 2873 24857 2907
rect 4905 2805 4939 2839
rect 5871 2805 5905 2839
rect 6929 2805 6963 2839
rect 11529 2805 11563 2839
rect 11897 2805 11931 2839
rect 14657 2805 14691 2839
rect 19165 2805 19199 2839
rect 21005 2805 21039 2839
rect 21327 2805 21361 2839
rect 22339 2805 22373 2839
rect 2099 2601 2133 2635
rect 3525 2601 3559 2635
rect 4353 2601 4387 2635
rect 4951 2601 4985 2635
rect 7849 2601 7883 2635
rect 9919 2601 9953 2635
rect 11989 2601 12023 2635
rect 13001 2601 13035 2635
rect 18061 2601 18095 2635
rect 21005 2601 21039 2635
rect 6377 2533 6411 2567
rect 6745 2533 6779 2567
rect 10885 2533 10919 2567
rect 11161 2533 11195 2567
rect 13277 2533 13311 2567
rect 13645 2533 13679 2567
rect 15945 2533 15979 2567
rect 16405 2533 16439 2567
rect 17233 2533 17267 2567
rect 18521 2533 18555 2567
rect 19441 2533 19475 2567
rect 2028 2465 2062 2499
rect 3024 2465 3058 2499
rect 4880 2465 4914 2499
rect 5089 2465 5123 2499
rect 5825 2465 5859 2499
rect 6929 2465 6963 2499
rect 8033 2465 8067 2499
rect 9848 2465 9882 2499
rect 10241 2465 10275 2499
rect 11713 2465 11747 2499
rect 17601 2465 17635 2499
rect 19901 2465 19935 2499
rect 20453 2465 20487 2499
rect 22109 2465 22143 2499
rect 24593 2465 24627 2499
rect 25145 2465 25179 2499
rect 3111 2397 3145 2431
rect 7481 2397 7515 2431
rect 11069 2397 11103 2431
rect 13553 2397 13587 2431
rect 16313 2397 16347 2431
rect 18429 2397 18463 2431
rect 18889 2397 18923 2431
rect 22661 2397 22695 2431
rect 5089 2329 5123 2363
rect 5365 2329 5399 2363
rect 8677 2329 8711 2363
rect 14105 2329 14139 2363
rect 16865 2329 16899 2363
rect 20085 2329 20119 2363
rect 22293 2329 22327 2363
rect 24777 2329 24811 2363
rect 2513 2261 2547 2295
rect 6009 2261 6043 2295
rect 7113 2261 7147 2295
rect 8217 2261 8251 2295
rect 9045 2261 9079 2295
rect 9505 2261 9539 2295
rect 12449 2261 12483 2295
rect 14565 2261 14599 2295
<< metal1 >>
rect 14 27480 20 27532
rect 72 27520 78 27532
rect 750 27520 756 27532
rect 72 27492 756 27520
rect 72 27480 78 27492
rect 750 27480 756 27492
rect 808 27480 814 27532
rect 2866 27480 2872 27532
rect 2924 27520 2930 27532
rect 3694 27520 3700 27532
rect 2924 27492 3700 27520
rect 2924 27480 2930 27492
rect 3694 27480 3700 27492
rect 3752 27480 3758 27532
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 25130 24936 25136 24948
rect 25091 24908 25136 24936
rect 25130 24896 25136 24908
rect 25188 24896 25194 24948
rect 24648 24735 24706 24741
rect 24648 24701 24660 24735
rect 24694 24732 24706 24735
rect 25130 24732 25136 24744
rect 24694 24704 25136 24732
rect 24694 24701 24706 24704
rect 24648 24695 24706 24701
rect 25130 24692 25136 24704
rect 25188 24692 25194 24744
rect 11422 24556 11428 24608
rect 11480 24596 11486 24608
rect 12437 24599 12495 24605
rect 12437 24596 12449 24599
rect 11480 24568 12449 24596
rect 11480 24556 11486 24568
rect 12437 24565 12449 24568
rect 12483 24565 12495 24599
rect 12437 24559 12495 24565
rect 21266 24556 21272 24608
rect 21324 24596 21330 24608
rect 24719 24599 24777 24605
rect 24719 24596 24731 24599
rect 21324 24568 24731 24596
rect 21324 24556 21330 24568
rect 24719 24565 24731 24568
rect 24765 24565 24777 24599
rect 24719 24559 24777 24565
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 24765 24395 24823 24401
rect 24765 24361 24777 24395
rect 24811 24392 24823 24395
rect 25774 24392 25780 24404
rect 24811 24364 25780 24392
rect 24811 24361 24823 24364
rect 24765 24355 24823 24361
rect 25774 24352 25780 24364
rect 25832 24352 25838 24404
rect 12688 24259 12746 24265
rect 12688 24225 12700 24259
rect 12734 24256 12746 24259
rect 13354 24256 13360 24268
rect 12734 24228 13360 24256
rect 12734 24225 12746 24228
rect 12688 24219 12746 24225
rect 13354 24216 13360 24228
rect 13412 24216 13418 24268
rect 13700 24259 13758 24265
rect 13700 24225 13712 24259
rect 13746 24256 13758 24259
rect 14090 24256 14096 24268
rect 13746 24228 14096 24256
rect 13746 24225 13758 24228
rect 13700 24219 13758 24225
rect 14090 24216 14096 24228
rect 14148 24216 14154 24268
rect 24026 24216 24032 24268
rect 24084 24256 24090 24268
rect 24581 24259 24639 24265
rect 24581 24256 24593 24259
rect 24084 24228 24593 24256
rect 24084 24216 24090 24228
rect 24581 24225 24593 24228
rect 24627 24225 24639 24259
rect 24581 24219 24639 24225
rect 11698 24148 11704 24200
rect 11756 24188 11762 24200
rect 13998 24188 14004 24200
rect 11756 24160 14004 24188
rect 11756 24148 11762 24160
rect 13998 24148 14004 24160
rect 14056 24148 14062 24200
rect 12759 24055 12817 24061
rect 12759 24021 12771 24055
rect 12805 24052 12817 24055
rect 13078 24052 13084 24064
rect 12805 24024 13084 24052
rect 12805 24021 12817 24024
rect 12759 24015 12817 24021
rect 13078 24012 13084 24024
rect 13136 24012 13142 24064
rect 13771 24055 13829 24061
rect 13771 24021 13783 24055
rect 13817 24052 13829 24055
rect 13998 24052 14004 24064
rect 13817 24024 14004 24052
rect 13817 24021 13829 24024
rect 13771 24015 13829 24021
rect 13998 24012 14004 24024
rect 14056 24012 14062 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 5350 23848 5356 23860
rect 5311 23820 5356 23848
rect 5350 23808 5356 23820
rect 5408 23808 5414 23860
rect 6638 23808 6644 23860
rect 6696 23848 6702 23860
rect 7009 23851 7067 23857
rect 7009 23848 7021 23851
rect 6696 23820 7021 23848
rect 6696 23808 6702 23820
rect 7009 23817 7021 23820
rect 7055 23817 7067 23851
rect 7009 23811 7067 23817
rect 7469 23851 7527 23857
rect 7469 23817 7481 23851
rect 7515 23848 7527 23851
rect 9582 23848 9588 23860
rect 7515 23820 9588 23848
rect 7515 23817 7527 23820
rect 7469 23811 7527 23817
rect 1448 23647 1506 23653
rect 1448 23613 1460 23647
rect 1494 23644 1506 23647
rect 1854 23644 1860 23656
rect 1494 23616 1860 23644
rect 1494 23613 1506 23616
rect 1448 23607 1506 23613
rect 1854 23604 1860 23616
rect 1912 23604 1918 23656
rect 4960 23647 5018 23653
rect 4960 23613 4972 23647
rect 5006 23644 5018 23647
rect 5350 23644 5356 23656
rect 5006 23616 5356 23644
rect 5006 23613 5018 23616
rect 4960 23607 5018 23613
rect 5350 23604 5356 23616
rect 5408 23604 5414 23656
rect 6178 23604 6184 23656
rect 6236 23644 6242 23656
rect 6825 23647 6883 23653
rect 6825 23644 6837 23647
rect 6236 23616 6837 23644
rect 6236 23604 6242 23616
rect 6825 23613 6837 23616
rect 6871 23644 6883 23647
rect 7484 23644 7512 23811
rect 9582 23808 9588 23820
rect 9640 23808 9646 23860
rect 12618 23848 12624 23860
rect 12579 23820 12624 23848
rect 12618 23808 12624 23820
rect 12676 23808 12682 23860
rect 13354 23848 13360 23860
rect 13315 23820 13360 23848
rect 13354 23808 13360 23820
rect 13412 23808 13418 23860
rect 15933 23851 15991 23857
rect 15933 23817 15945 23851
rect 15979 23848 15991 23851
rect 16942 23848 16948 23860
rect 15979 23820 16948 23848
rect 15979 23817 15991 23820
rect 15933 23811 15991 23817
rect 16942 23808 16948 23820
rect 17000 23808 17006 23860
rect 24762 23848 24768 23860
rect 24723 23820 24768 23848
rect 24762 23808 24768 23820
rect 24820 23808 24826 23860
rect 13538 23740 13544 23792
rect 13596 23780 13602 23792
rect 14691 23783 14749 23789
rect 14691 23780 14703 23783
rect 13596 23752 14703 23780
rect 13596 23740 13602 23752
rect 14691 23749 14703 23752
rect 14737 23749 14749 23783
rect 14691 23743 14749 23749
rect 12066 23672 12072 23724
rect 12124 23712 12130 23724
rect 12124 23684 15792 23712
rect 12124 23672 12130 23684
rect 6871 23616 7512 23644
rect 12437 23647 12495 23653
rect 6871 23613 6883 23616
rect 6825 23607 6883 23613
rect 12437 23613 12449 23647
rect 12483 23644 12495 23647
rect 12986 23644 12992 23656
rect 12483 23616 12992 23644
rect 12483 23613 12495 23616
rect 12437 23607 12495 23613
rect 12986 23604 12992 23616
rect 13044 23604 13050 23656
rect 13170 23604 13176 23656
rect 13228 23644 13234 23656
rect 13576 23647 13634 23653
rect 13576 23644 13588 23647
rect 13228 23616 13588 23644
rect 13228 23604 13234 23616
rect 13576 23613 13588 23616
rect 13622 23644 13634 23647
rect 13622 23616 13814 23644
rect 13622 23613 13634 23616
rect 13576 23607 13634 23613
rect 1535 23579 1593 23585
rect 1535 23545 1547 23579
rect 1581 23576 1593 23579
rect 2774 23576 2780 23588
rect 1581 23548 2780 23576
rect 1581 23545 1593 23548
rect 1535 23539 1593 23545
rect 2774 23536 2780 23548
rect 2832 23536 2838 23588
rect 13786 23576 13814 23616
rect 13906 23604 13912 23656
rect 13964 23644 13970 23656
rect 14620 23647 14678 23653
rect 14620 23644 14632 23647
rect 13964 23616 14632 23644
rect 13964 23604 13970 23616
rect 14620 23613 14632 23616
rect 14666 23644 14678 23647
rect 15105 23647 15163 23653
rect 15105 23644 15117 23647
rect 14666 23616 15117 23644
rect 14666 23613 14678 23616
rect 14620 23607 14678 23613
rect 15105 23613 15117 23616
rect 15151 23644 15163 23647
rect 15654 23644 15660 23656
rect 15151 23616 15660 23644
rect 15151 23613 15163 23616
rect 15105 23607 15163 23613
rect 15654 23604 15660 23616
rect 15712 23604 15718 23656
rect 15764 23653 15792 23684
rect 15749 23647 15807 23653
rect 15749 23613 15761 23647
rect 15795 23644 15807 23647
rect 16301 23647 16359 23653
rect 16301 23644 16313 23647
rect 15795 23616 16313 23644
rect 15795 23613 15807 23616
rect 15749 23607 15807 23613
rect 16301 23613 16313 23616
rect 16347 23644 16359 23647
rect 16390 23644 16396 23656
rect 16347 23616 16396 23644
rect 16347 23613 16359 23616
rect 16301 23607 16359 23613
rect 16390 23604 16396 23616
rect 16448 23604 16454 23656
rect 18049 23647 18107 23653
rect 18049 23613 18061 23647
rect 18095 23613 18107 23647
rect 18049 23607 18107 23613
rect 24581 23647 24639 23653
rect 24581 23613 24593 23647
rect 24627 23644 24639 23647
rect 24627 23616 25268 23644
rect 24627 23613 24639 23616
rect 24581 23607 24639 23613
rect 14461 23579 14519 23585
rect 14461 23576 14473 23579
rect 13786 23548 14473 23576
rect 14461 23545 14473 23548
rect 14507 23576 14519 23579
rect 16482 23576 16488 23588
rect 14507 23548 16488 23576
rect 14507 23545 14519 23548
rect 14461 23539 14519 23545
rect 16482 23536 16488 23548
rect 16540 23536 16546 23588
rect 18064 23576 18092 23607
rect 18506 23576 18512 23588
rect 18064 23548 18512 23576
rect 5031 23511 5089 23517
rect 5031 23477 5043 23511
rect 5077 23508 5089 23511
rect 7190 23508 7196 23520
rect 5077 23480 7196 23508
rect 5077 23477 5089 23480
rect 5031 23471 5089 23477
rect 7190 23468 7196 23480
rect 7248 23468 7254 23520
rect 13446 23468 13452 23520
rect 13504 23508 13510 23520
rect 13679 23511 13737 23517
rect 13679 23508 13691 23511
rect 13504 23480 13691 23508
rect 13504 23468 13510 23480
rect 13679 23477 13691 23480
rect 13725 23477 13737 23511
rect 14090 23508 14096 23520
rect 14003 23480 14096 23508
rect 13679 23471 13737 23477
rect 14090 23468 14096 23480
rect 14148 23508 14154 23520
rect 18064 23508 18092 23548
rect 18506 23536 18512 23548
rect 18564 23576 18570 23588
rect 18601 23579 18659 23585
rect 18601 23576 18613 23579
rect 18564 23548 18613 23576
rect 18564 23536 18570 23548
rect 18601 23545 18613 23548
rect 18647 23545 18659 23579
rect 18601 23539 18659 23545
rect 18230 23508 18236 23520
rect 14148 23480 18092 23508
rect 18191 23480 18236 23508
rect 14148 23468 14154 23480
rect 18230 23468 18236 23480
rect 18288 23468 18294 23520
rect 24026 23468 24032 23520
rect 24084 23508 24090 23520
rect 25240 23517 25268 23616
rect 24397 23511 24455 23517
rect 24397 23508 24409 23511
rect 24084 23480 24409 23508
rect 24084 23468 24090 23480
rect 24397 23477 24409 23480
rect 24443 23477 24455 23511
rect 24397 23471 24455 23477
rect 25225 23511 25283 23517
rect 25225 23477 25237 23511
rect 25271 23508 25283 23511
rect 25314 23508 25320 23520
rect 25271 23480 25320 23508
rect 25271 23477 25283 23480
rect 25225 23471 25283 23477
rect 25314 23468 25320 23480
rect 25372 23468 25378 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 9582 23264 9588 23316
rect 9640 23304 9646 23316
rect 13170 23304 13176 23316
rect 9640 23276 13176 23304
rect 9640 23264 9646 23276
rect 13170 23264 13176 23276
rect 13228 23264 13234 23316
rect 16482 23264 16488 23316
rect 16540 23304 16546 23316
rect 18046 23304 18052 23316
rect 16540 23276 18052 23304
rect 16540 23264 16546 23276
rect 18046 23264 18052 23276
rect 18104 23264 18110 23316
rect 24765 23307 24823 23313
rect 24765 23273 24777 23307
rect 24811 23304 24823 23307
rect 27246 23304 27252 23316
rect 24811 23276 27252 23304
rect 24811 23273 24823 23276
rect 24765 23267 24823 23273
rect 27246 23264 27252 23276
rect 27304 23264 27310 23316
rect 1464 23171 1522 23177
rect 1464 23137 1476 23171
rect 1510 23168 1522 23171
rect 1578 23168 1584 23180
rect 1510 23140 1584 23168
rect 1510 23137 1522 23140
rect 1464 23131 1522 23137
rect 1578 23128 1584 23140
rect 1636 23128 1642 23180
rect 9585 23171 9643 23177
rect 9585 23137 9597 23171
rect 9631 23168 9643 23171
rect 9674 23168 9680 23180
rect 9631 23140 9680 23168
rect 9631 23137 9643 23140
rect 9585 23131 9643 23137
rect 9674 23128 9680 23140
rect 9732 23128 9738 23180
rect 11216 23171 11274 23177
rect 11216 23137 11228 23171
rect 11262 23168 11274 23171
rect 11330 23168 11336 23180
rect 11262 23140 11336 23168
rect 11262 23137 11274 23140
rect 11216 23131 11274 23137
rect 11330 23128 11336 23140
rect 11388 23128 11394 23180
rect 13240 23171 13298 23177
rect 13240 23137 13252 23171
rect 13286 23168 13298 23171
rect 13906 23168 13912 23180
rect 13286 23140 13912 23168
rect 13286 23137 13298 23140
rect 13240 23131 13298 23137
rect 13906 23128 13912 23140
rect 13964 23128 13970 23180
rect 15356 23171 15414 23177
rect 15356 23137 15368 23171
rect 15402 23168 15414 23171
rect 15470 23168 15476 23180
rect 15402 23140 15476 23168
rect 15402 23137 15414 23140
rect 15356 23131 15414 23137
rect 15470 23128 15476 23140
rect 15528 23128 15534 23180
rect 16368 23171 16426 23177
rect 16368 23137 16380 23171
rect 16414 23168 16426 23171
rect 16758 23168 16764 23180
rect 16414 23140 16764 23168
rect 16414 23137 16426 23140
rect 16368 23131 16426 23137
rect 16758 23128 16764 23140
rect 16816 23128 16822 23180
rect 24581 23171 24639 23177
rect 24581 23137 24593 23171
rect 24627 23168 24639 23171
rect 24670 23168 24676 23180
rect 24627 23140 24676 23168
rect 24627 23137 24639 23140
rect 24581 23131 24639 23137
rect 24670 23128 24676 23140
rect 24728 23128 24734 23180
rect 12158 23100 12164 23112
rect 12119 23072 12164 23100
rect 12158 23060 12164 23072
rect 12216 23060 12222 23112
rect 12710 23060 12716 23112
rect 12768 23100 12774 23112
rect 14185 23103 14243 23109
rect 14185 23100 14197 23103
rect 12768 23072 14197 23100
rect 12768 23060 12774 23072
rect 14185 23069 14197 23072
rect 14231 23069 14243 23103
rect 14185 23063 14243 23069
rect 9815 23035 9873 23041
rect 9815 23001 9827 23035
rect 9861 23032 9873 23035
rect 12802 23032 12808 23044
rect 9861 23004 12808 23032
rect 9861 23001 9873 23004
rect 9815 22995 9873 23001
rect 12802 22992 12808 23004
rect 12860 22992 12866 23044
rect 1535 22967 1593 22973
rect 1535 22933 1547 22967
rect 1581 22964 1593 22967
rect 2590 22964 2596 22976
rect 1581 22936 2596 22964
rect 1581 22933 1593 22936
rect 1535 22927 1593 22933
rect 2590 22924 2596 22936
rect 2648 22924 2654 22976
rect 11287 22967 11345 22973
rect 11287 22933 11299 22967
rect 11333 22964 11345 22967
rect 12894 22964 12900 22976
rect 11333 22936 12900 22964
rect 11333 22933 11345 22936
rect 11287 22927 11345 22933
rect 12894 22924 12900 22936
rect 12952 22924 12958 22976
rect 13170 22924 13176 22976
rect 13228 22964 13234 22976
rect 13311 22967 13369 22973
rect 13311 22964 13323 22967
rect 13228 22936 13323 22964
rect 13228 22924 13234 22936
rect 13311 22933 13323 22936
rect 13357 22933 13369 22967
rect 13311 22927 13369 22933
rect 14734 22924 14740 22976
rect 14792 22964 14798 22976
rect 15427 22967 15485 22973
rect 15427 22964 15439 22967
rect 14792 22936 15439 22964
rect 14792 22924 14798 22936
rect 15427 22933 15439 22936
rect 15473 22933 15485 22967
rect 15427 22927 15485 22933
rect 16022 22924 16028 22976
rect 16080 22964 16086 22976
rect 16439 22967 16497 22973
rect 16439 22964 16451 22967
rect 16080 22936 16451 22964
rect 16080 22924 16086 22936
rect 16439 22933 16451 22936
rect 16485 22933 16497 22967
rect 16439 22927 16497 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1578 22760 1584 22772
rect 1539 22732 1584 22760
rect 1578 22720 1584 22732
rect 1636 22720 1642 22772
rect 7653 22763 7711 22769
rect 7653 22729 7665 22763
rect 7699 22760 7711 22763
rect 8110 22760 8116 22772
rect 7699 22732 8116 22760
rect 7699 22729 7711 22732
rect 7653 22723 7711 22729
rect 8110 22720 8116 22732
rect 8168 22720 8174 22772
rect 10873 22763 10931 22769
rect 10873 22729 10885 22763
rect 10919 22760 10931 22763
rect 11054 22760 11060 22772
rect 10919 22732 11060 22760
rect 10919 22729 10931 22732
rect 10873 22723 10931 22729
rect 11054 22720 11060 22732
rect 11112 22720 11118 22772
rect 13722 22720 13728 22772
rect 13780 22760 13786 22772
rect 15470 22760 15476 22772
rect 13780 22732 15476 22760
rect 13780 22720 13786 22732
rect 15470 22720 15476 22732
rect 15528 22760 15534 22772
rect 15657 22763 15715 22769
rect 15657 22760 15669 22763
rect 15528 22732 15669 22760
rect 15528 22720 15534 22732
rect 15657 22729 15669 22732
rect 15703 22729 15715 22763
rect 15657 22723 15715 22729
rect 18598 22720 18604 22772
rect 18656 22760 18662 22772
rect 21358 22760 21364 22772
rect 18656 22732 21364 22760
rect 18656 22720 18662 22732
rect 21358 22720 21364 22732
rect 21416 22720 21422 22772
rect 24670 22760 24676 22772
rect 24631 22732 24676 22760
rect 24670 22720 24676 22732
rect 24728 22720 24734 22772
rect 8018 22652 8024 22704
rect 8076 22692 8082 22704
rect 9674 22692 9680 22704
rect 8076 22664 9680 22692
rect 8076 22652 8082 22664
rect 9674 22652 9680 22664
rect 9732 22692 9738 22704
rect 10137 22695 10195 22701
rect 10137 22692 10149 22695
rect 9732 22664 10149 22692
rect 9732 22652 9738 22664
rect 10137 22661 10149 22664
rect 10183 22661 10195 22695
rect 10137 22655 10195 22661
rect 10597 22695 10655 22701
rect 10597 22661 10609 22695
rect 10643 22692 10655 22695
rect 20898 22692 20904 22704
rect 10643 22664 13492 22692
rect 10643 22661 10655 22664
rect 10597 22655 10655 22661
rect 7466 22556 7472 22568
rect 7379 22528 7472 22556
rect 7466 22516 7472 22528
rect 7524 22556 7530 22568
rect 8021 22559 8079 22565
rect 8021 22556 8033 22559
rect 7524 22528 8033 22556
rect 7524 22516 7530 22528
rect 8021 22525 8033 22528
rect 8067 22525 8079 22559
rect 8021 22519 8079 22525
rect 8700 22559 8758 22565
rect 8700 22525 8712 22559
rect 8746 22556 8758 22559
rect 9125 22559 9183 22565
rect 9125 22556 9137 22559
rect 8746 22528 9137 22556
rect 8746 22525 8758 22528
rect 8700 22519 8758 22525
rect 9125 22525 9137 22528
rect 9171 22556 9183 22559
rect 9214 22556 9220 22568
rect 9171 22528 9220 22556
rect 9171 22525 9183 22528
rect 9125 22519 9183 22525
rect 7834 22448 7840 22500
rect 7892 22488 7898 22500
rect 8715 22488 8743 22519
rect 9214 22516 9220 22528
rect 9272 22516 9278 22568
rect 9744 22559 9802 22565
rect 9744 22525 9756 22559
rect 9790 22556 9802 22559
rect 10612 22556 10640 22655
rect 11054 22584 11060 22636
rect 11112 22624 11118 22636
rect 13354 22624 13360 22636
rect 11112 22596 13360 22624
rect 11112 22584 11118 22596
rect 13354 22584 13360 22596
rect 13412 22584 13418 22636
rect 13464 22624 13492 22664
rect 13694 22664 20904 22692
rect 13694 22624 13722 22664
rect 20898 22652 20904 22664
rect 20956 22652 20962 22704
rect 13464 22596 13722 22624
rect 14458 22584 14464 22636
rect 14516 22624 14522 22636
rect 15335 22627 15393 22633
rect 15335 22624 15347 22627
rect 14516 22596 15347 22624
rect 14516 22584 14522 22596
rect 15335 22593 15347 22596
rect 15381 22593 15393 22627
rect 15335 22587 15393 22593
rect 15838 22584 15844 22636
rect 15896 22624 15902 22636
rect 16347 22627 16405 22633
rect 16347 22624 16359 22627
rect 15896 22596 16359 22624
rect 15896 22584 15902 22596
rect 16347 22593 16359 22596
rect 16393 22593 16405 22627
rect 16347 22587 16405 22593
rect 9790 22528 10640 22556
rect 10689 22559 10747 22565
rect 9790 22525 9802 22528
rect 9744 22519 9802 22525
rect 10689 22525 10701 22559
rect 10735 22556 10747 22559
rect 10778 22556 10784 22568
rect 10735 22528 10784 22556
rect 10735 22525 10747 22528
rect 10689 22519 10747 22525
rect 10778 22516 10784 22528
rect 10836 22516 10842 22568
rect 12872 22559 12930 22565
rect 12872 22525 12884 22559
rect 12918 22556 12930 22559
rect 12986 22556 12992 22568
rect 12918 22528 12992 22556
rect 12918 22525 12930 22528
rect 12872 22519 12930 22525
rect 12986 22516 12992 22528
rect 13044 22556 13050 22568
rect 13725 22559 13783 22565
rect 13044 22528 13400 22556
rect 13044 22516 13050 22528
rect 7892 22460 8743 22488
rect 8803 22491 8861 22497
rect 7892 22448 7898 22460
rect 8803 22457 8815 22491
rect 8849 22488 8861 22491
rect 9306 22488 9312 22500
rect 8849 22460 9312 22488
rect 8849 22457 8861 22460
rect 8803 22451 8861 22457
rect 9306 22448 9312 22460
rect 9364 22448 9370 22500
rect 13372 22432 13400 22528
rect 13725 22525 13737 22559
rect 13771 22556 13783 22559
rect 13906 22556 13912 22568
rect 13771 22528 13912 22556
rect 13771 22525 13783 22528
rect 13725 22519 13783 22525
rect 13906 22516 13912 22528
rect 13964 22516 13970 22568
rect 14252 22559 14310 22565
rect 14252 22525 14264 22559
rect 14298 22556 14310 22559
rect 15248 22559 15306 22565
rect 14298 22528 14504 22556
rect 14298 22525 14310 22528
rect 14252 22519 14310 22525
rect 9490 22380 9496 22432
rect 9548 22420 9554 22432
rect 9815 22423 9873 22429
rect 9815 22420 9827 22423
rect 9548 22392 9827 22420
rect 9548 22380 9554 22392
rect 9815 22389 9827 22392
rect 9861 22389 9873 22423
rect 11330 22420 11336 22432
rect 11243 22392 11336 22420
rect 9815 22383 9873 22389
rect 11330 22380 11336 22392
rect 11388 22420 11394 22432
rect 12434 22420 12440 22432
rect 11388 22392 12440 22420
rect 11388 22380 11394 22392
rect 12434 22380 12440 22392
rect 12492 22380 12498 22432
rect 12943 22423 13001 22429
rect 12943 22389 12955 22423
rect 12989 22420 13001 22423
rect 13170 22420 13176 22432
rect 12989 22392 13176 22420
rect 12989 22389 13001 22392
rect 12943 22383 13001 22389
rect 13170 22380 13176 22392
rect 13228 22380 13234 22432
rect 13354 22420 13360 22432
rect 13315 22392 13360 22420
rect 13354 22380 13360 22392
rect 13412 22380 13418 22432
rect 13906 22380 13912 22432
rect 13964 22420 13970 22432
rect 14323 22423 14381 22429
rect 14323 22420 14335 22423
rect 13964 22392 14335 22420
rect 13964 22380 13970 22392
rect 14323 22389 14335 22392
rect 14369 22389 14381 22423
rect 14476 22420 14504 22528
rect 15248 22525 15260 22559
rect 15294 22556 15306 22559
rect 16114 22556 16120 22568
rect 15294 22528 16120 22556
rect 15294 22525 15306 22528
rect 15248 22519 15306 22525
rect 16114 22516 16120 22528
rect 16172 22516 16178 22568
rect 16244 22559 16302 22565
rect 16244 22525 16256 22559
rect 16290 22525 16302 22559
rect 16244 22519 16302 22525
rect 14550 22448 14556 22500
rect 14608 22488 14614 22500
rect 16259 22488 16287 22519
rect 16669 22491 16727 22497
rect 16669 22488 16681 22491
rect 14608 22460 16681 22488
rect 14608 22448 14614 22460
rect 16669 22457 16681 22460
rect 16715 22457 16727 22491
rect 16669 22451 16727 22457
rect 14737 22423 14795 22429
rect 14737 22420 14749 22423
rect 14476 22392 14749 22420
rect 14323 22383 14381 22389
rect 14737 22389 14749 22392
rect 14783 22420 14795 22423
rect 14826 22420 14832 22432
rect 14783 22392 14832 22420
rect 14783 22389 14795 22392
rect 14737 22383 14795 22389
rect 14826 22380 14832 22392
rect 14884 22380 14890 22432
rect 16114 22420 16120 22432
rect 16075 22392 16120 22420
rect 16114 22380 16120 22392
rect 16172 22380 16178 22432
rect 16758 22380 16764 22432
rect 16816 22420 16822 22432
rect 17037 22423 17095 22429
rect 17037 22420 17049 22423
rect 16816 22392 17049 22420
rect 16816 22380 16822 22392
rect 17037 22389 17049 22392
rect 17083 22389 17095 22423
rect 17037 22383 17095 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 6871 22219 6929 22225
rect 6871 22185 6883 22219
rect 6917 22216 6929 22219
rect 7466 22216 7472 22228
rect 6917 22188 7472 22216
rect 6917 22185 6929 22188
rect 6871 22179 6929 22185
rect 7466 22176 7472 22188
rect 7524 22176 7530 22228
rect 12986 22176 12992 22228
rect 13044 22216 13050 22228
rect 13998 22216 14004 22228
rect 13044 22188 13216 22216
rect 13959 22188 14004 22216
rect 13044 22176 13050 22188
rect 13078 22148 13084 22160
rect 13039 22120 13084 22148
rect 13078 22108 13084 22120
rect 13136 22108 13142 22160
rect 13188 22157 13216 22188
rect 13998 22176 14004 22188
rect 14056 22176 14062 22228
rect 14826 22176 14832 22228
rect 14884 22216 14890 22228
rect 14884 22188 17724 22216
rect 14884 22176 14890 22188
rect 13173 22151 13231 22157
rect 13173 22117 13185 22151
rect 13219 22117 13231 22151
rect 13173 22111 13231 22117
rect 15286 22108 15292 22160
rect 15344 22148 15350 22160
rect 17543 22151 17601 22157
rect 17543 22148 17555 22151
rect 15344 22120 17555 22148
rect 15344 22108 15350 22120
rect 17543 22117 17555 22120
rect 17589 22117 17601 22151
rect 17543 22111 17601 22117
rect 6800 22083 6858 22089
rect 6800 22049 6812 22083
rect 6846 22080 6858 22083
rect 7098 22080 7104 22092
rect 6846 22052 7104 22080
rect 6846 22049 6858 22052
rect 6800 22043 6858 22049
rect 7098 22040 7104 22052
rect 7156 22040 7162 22092
rect 7996 22083 8054 22089
rect 7996 22049 8008 22083
rect 8042 22080 8054 22083
rect 8570 22080 8576 22092
rect 8042 22052 8576 22080
rect 8042 22049 8054 22052
rect 7996 22043 8054 22049
rect 8570 22040 8576 22052
rect 8628 22040 8634 22092
rect 9712 22083 9770 22089
rect 9712 22080 9724 22083
rect 9692 22049 9724 22080
rect 9758 22049 9770 22083
rect 10778 22080 10784 22092
rect 10739 22052 10784 22080
rect 9692 22043 9770 22049
rect 9692 21956 9720 22043
rect 10778 22040 10784 22052
rect 10836 22040 10842 22092
rect 12044 22083 12102 22089
rect 12044 22049 12056 22083
rect 12090 22080 12102 22083
rect 12526 22080 12532 22092
rect 12090 22052 12532 22080
rect 12090 22049 12102 22052
rect 12044 22043 12102 22049
rect 12526 22040 12532 22052
rect 12584 22040 12590 22092
rect 15378 22080 15384 22092
rect 15339 22052 15384 22080
rect 15378 22040 15384 22052
rect 15436 22040 15442 22092
rect 16393 22083 16451 22089
rect 16393 22049 16405 22083
rect 16439 22080 16451 22083
rect 16482 22080 16488 22092
rect 16439 22052 16488 22080
rect 16439 22049 16451 22052
rect 16393 22043 16451 22049
rect 16482 22040 16488 22052
rect 16540 22040 16546 22092
rect 17218 22040 17224 22092
rect 17276 22080 17282 22092
rect 17440 22083 17498 22089
rect 17440 22080 17452 22083
rect 17276 22052 17452 22080
rect 17276 22040 17282 22052
rect 17440 22049 17452 22052
rect 17486 22049 17498 22083
rect 17696 22080 17724 22188
rect 18484 22083 18542 22089
rect 18484 22080 18496 22083
rect 17696 22052 18496 22080
rect 17440 22043 17498 22049
rect 18484 22049 18496 22052
rect 18530 22080 18542 22083
rect 18598 22080 18604 22092
rect 18530 22052 18604 22080
rect 18530 22049 18542 22052
rect 18484 22043 18542 22049
rect 18598 22040 18604 22052
rect 18656 22040 18662 22092
rect 20952 22083 21010 22089
rect 20952 22049 20964 22083
rect 20998 22080 21010 22083
rect 21266 22080 21272 22092
rect 20998 22052 21272 22080
rect 20998 22049 21010 22052
rect 20952 22043 21010 22049
rect 21266 22040 21272 22052
rect 21324 22040 21330 22092
rect 12544 22012 12572 22040
rect 14826 22012 14832 22024
rect 12544 21984 14832 22012
rect 14826 21972 14832 21984
rect 14884 21972 14890 22024
rect 17586 21972 17592 22024
rect 17644 22012 17650 22024
rect 21039 22015 21097 22021
rect 21039 22012 21051 22015
rect 17644 21984 21051 22012
rect 17644 21972 17650 21984
rect 21039 21981 21051 21984
rect 21085 21981 21097 22015
rect 21039 21975 21097 21981
rect 9674 21904 9680 21956
rect 9732 21904 9738 21956
rect 10870 21944 10876 21956
rect 10831 21916 10876 21944
rect 10870 21904 10876 21916
rect 10928 21904 10934 21956
rect 12250 21904 12256 21956
rect 12308 21944 12314 21956
rect 13633 21947 13691 21953
rect 13633 21944 13645 21947
rect 12308 21916 13645 21944
rect 12308 21904 12314 21916
rect 13633 21913 13645 21916
rect 13679 21913 13691 21947
rect 13633 21907 13691 21913
rect 17126 21904 17132 21956
rect 17184 21944 17190 21956
rect 18555 21947 18613 21953
rect 18555 21944 18567 21947
rect 17184 21916 18567 21944
rect 17184 21904 17190 21916
rect 18555 21913 18567 21916
rect 18601 21913 18613 21947
rect 18555 21907 18613 21913
rect 8067 21879 8125 21885
rect 8067 21845 8079 21879
rect 8113 21876 8125 21879
rect 8202 21876 8208 21888
rect 8113 21848 8208 21876
rect 8113 21845 8125 21848
rect 8067 21839 8125 21845
rect 8202 21836 8208 21848
rect 8260 21836 8266 21888
rect 8662 21876 8668 21888
rect 8623 21848 8668 21876
rect 8662 21836 8668 21848
rect 8720 21836 8726 21888
rect 9030 21876 9036 21888
rect 8991 21848 9036 21876
rect 9030 21836 9036 21848
rect 9088 21836 9094 21888
rect 9122 21836 9128 21888
rect 9180 21876 9186 21888
rect 9815 21879 9873 21885
rect 9815 21876 9827 21879
rect 9180 21848 9827 21876
rect 9180 21836 9186 21848
rect 9815 21845 9827 21848
rect 9861 21845 9873 21879
rect 9815 21839 9873 21845
rect 11103 21879 11161 21885
rect 11103 21845 11115 21879
rect 11149 21876 11161 21879
rect 11974 21876 11980 21888
rect 11149 21848 11980 21876
rect 11149 21845 11161 21848
rect 11103 21839 11161 21845
rect 11974 21836 11980 21848
rect 12032 21836 12038 21888
rect 12115 21879 12173 21885
rect 12115 21845 12127 21879
rect 12161 21876 12173 21879
rect 12342 21876 12348 21888
rect 12161 21848 12348 21876
rect 12161 21845 12173 21848
rect 12115 21839 12173 21845
rect 12342 21836 12348 21848
rect 12400 21836 12406 21888
rect 15470 21836 15476 21888
rect 15528 21876 15534 21888
rect 15565 21879 15623 21885
rect 15565 21876 15577 21879
rect 15528 21848 15577 21876
rect 15528 21836 15534 21848
rect 15565 21845 15577 21848
rect 15611 21845 15623 21879
rect 15565 21839 15623 21845
rect 16298 21836 16304 21888
rect 16356 21876 16362 21888
rect 16531 21879 16589 21885
rect 16531 21876 16543 21879
rect 16356 21848 16543 21876
rect 16356 21836 16362 21848
rect 16531 21845 16543 21848
rect 16577 21845 16589 21879
rect 16531 21839 16589 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 9030 21632 9036 21684
rect 9088 21672 9094 21684
rect 10275 21675 10333 21681
rect 10275 21672 10287 21675
rect 9088 21644 10287 21672
rect 9088 21632 9094 21644
rect 10275 21641 10287 21644
rect 10321 21641 10333 21675
rect 10275 21635 10333 21641
rect 13078 21632 13084 21684
rect 13136 21672 13142 21684
rect 14369 21675 14427 21681
rect 14369 21672 14381 21675
rect 13136 21644 14381 21672
rect 13136 21632 13142 21644
rect 14369 21641 14381 21644
rect 14415 21641 14427 21675
rect 14369 21635 14427 21641
rect 16482 21632 16488 21684
rect 16540 21672 16546 21684
rect 16761 21675 16819 21681
rect 16761 21672 16773 21675
rect 16540 21644 16773 21672
rect 16540 21632 16546 21644
rect 16761 21641 16773 21644
rect 16807 21641 16819 21675
rect 19337 21675 19395 21681
rect 19337 21672 19349 21675
rect 16761 21635 16819 21641
rect 18023 21644 19349 21672
rect 8481 21607 8539 21613
rect 8481 21573 8493 21607
rect 8527 21604 8539 21607
rect 8570 21604 8576 21616
rect 8527 21576 8576 21604
rect 8527 21573 8539 21576
rect 8481 21567 8539 21573
rect 8570 21564 8576 21576
rect 8628 21564 8634 21616
rect 8665 21539 8723 21545
rect 8665 21505 8677 21539
rect 8711 21536 8723 21539
rect 9048 21536 9076 21632
rect 9674 21564 9680 21616
rect 9732 21604 9738 21616
rect 9732 21576 9777 21604
rect 9732 21564 9738 21576
rect 10870 21564 10876 21616
rect 10928 21604 10934 21616
rect 11057 21607 11115 21613
rect 11057 21604 11069 21607
rect 10928 21576 11069 21604
rect 10928 21564 10934 21576
rect 11057 21573 11069 21576
rect 11103 21604 11115 21607
rect 13630 21604 13636 21616
rect 11103 21576 13636 21604
rect 11103 21573 11115 21576
rect 11057 21567 11115 21573
rect 13630 21564 13636 21576
rect 13688 21564 13694 21616
rect 13998 21604 14004 21616
rect 13786 21576 14004 21604
rect 8711 21508 9076 21536
rect 13449 21539 13507 21545
rect 8711 21505 8723 21508
rect 8665 21499 8723 21505
rect 13449 21505 13461 21539
rect 13495 21536 13507 21539
rect 13786 21536 13814 21576
rect 13998 21564 14004 21576
rect 14056 21564 14062 21616
rect 14090 21564 14096 21616
rect 14148 21604 14154 21616
rect 15059 21607 15117 21613
rect 15059 21604 15071 21607
rect 14148 21576 15071 21604
rect 14148 21564 14154 21576
rect 15059 21573 15071 21576
rect 15105 21573 15117 21607
rect 15059 21567 15117 21573
rect 16393 21607 16451 21613
rect 16393 21573 16405 21607
rect 16439 21604 16451 21607
rect 18023 21604 18051 21644
rect 19337 21641 19349 21644
rect 19383 21641 19395 21675
rect 20898 21672 20904 21684
rect 20859 21644 20904 21672
rect 19337 21635 19395 21641
rect 20898 21632 20904 21644
rect 20956 21632 20962 21684
rect 21266 21672 21272 21684
rect 21227 21644 21272 21672
rect 21266 21632 21272 21644
rect 21324 21672 21330 21684
rect 22002 21672 22008 21684
rect 21324 21644 22008 21672
rect 21324 21632 21330 21644
rect 22002 21632 22008 21644
rect 22060 21632 22066 21684
rect 16439 21576 18051 21604
rect 16439 21573 16451 21576
rect 16393 21567 16451 21573
rect 13495 21508 13814 21536
rect 13495 21505 13507 21508
rect 13449 21499 13507 21505
rect 14642 21496 14648 21548
rect 14700 21536 14706 21548
rect 15378 21536 15384 21548
rect 14700 21508 15384 21536
rect 14700 21496 14706 21508
rect 15378 21496 15384 21508
rect 15436 21536 15442 21548
rect 15749 21539 15807 21545
rect 15749 21536 15761 21539
rect 15436 21508 15761 21536
rect 15436 21496 15442 21508
rect 15749 21505 15761 21508
rect 15795 21505 15807 21539
rect 16408 21536 16436 21567
rect 18322 21564 18328 21616
rect 18380 21604 18386 21616
rect 19199 21607 19257 21613
rect 19199 21604 19211 21607
rect 18380 21576 19211 21604
rect 18380 21564 18386 21576
rect 19199 21573 19211 21576
rect 19245 21573 19257 21607
rect 19199 21567 19257 21573
rect 15749 21499 15807 21505
rect 16015 21508 16436 21536
rect 17865 21539 17923 21545
rect 2130 21428 2136 21480
rect 2188 21468 2194 21480
rect 7628 21471 7686 21477
rect 7628 21468 7640 21471
rect 2188 21440 7640 21468
rect 2188 21428 2194 21440
rect 7628 21437 7640 21440
rect 7674 21468 7686 21471
rect 10204 21471 10262 21477
rect 7674 21440 8156 21468
rect 7674 21437 7686 21440
rect 7628 21431 7686 21437
rect 8128 21344 8156 21440
rect 10204 21437 10216 21471
rect 10250 21468 10262 21471
rect 10597 21471 10655 21477
rect 10597 21468 10609 21471
rect 10250 21440 10609 21468
rect 10250 21437 10262 21440
rect 10204 21431 10262 21437
rect 10597 21437 10609 21440
rect 10643 21468 10655 21471
rect 11054 21468 11060 21480
rect 10643 21440 11060 21468
rect 10643 21437 10655 21440
rect 10597 21431 10655 21437
rect 11054 21428 11060 21440
rect 11112 21428 11118 21480
rect 11216 21471 11274 21477
rect 11216 21437 11228 21471
rect 11262 21468 11274 21471
rect 11698 21468 11704 21480
rect 11262 21440 11704 21468
rect 11262 21437 11274 21440
rect 11216 21431 11274 21437
rect 11698 21428 11704 21440
rect 11756 21428 11762 21480
rect 14826 21428 14832 21480
rect 14884 21468 14890 21480
rect 16015 21477 16043 21508
rect 17865 21505 17877 21539
rect 17911 21536 17923 21539
rect 17911 21508 18552 21536
rect 17911 21505 17923 21508
rect 17865 21499 17923 21505
rect 14956 21471 15014 21477
rect 14956 21468 14968 21471
rect 14884 21440 14968 21468
rect 14884 21428 14890 21440
rect 14956 21437 14968 21440
rect 15002 21468 15014 21471
rect 15473 21471 15531 21477
rect 15473 21468 15485 21471
rect 15002 21440 15485 21468
rect 15002 21437 15014 21440
rect 14956 21431 15014 21437
rect 15473 21437 15485 21440
rect 15519 21437 15531 21471
rect 15473 21431 15531 21437
rect 16000 21471 16058 21477
rect 16000 21437 16012 21471
rect 16046 21437 16058 21471
rect 16000 21431 16058 21437
rect 16114 21428 16120 21480
rect 16172 21468 16178 21480
rect 16996 21471 17054 21477
rect 16996 21468 17008 21471
rect 16172 21440 17008 21468
rect 16172 21428 16178 21440
rect 16996 21437 17008 21440
rect 17042 21468 17054 21471
rect 17880 21468 17908 21499
rect 17042 21440 17908 21468
rect 18049 21471 18107 21477
rect 17042 21437 17054 21440
rect 16996 21431 17054 21437
rect 18049 21437 18061 21471
rect 18095 21468 18107 21471
rect 18414 21468 18420 21480
rect 18095 21440 18420 21468
rect 18095 21437 18107 21440
rect 18049 21431 18107 21437
rect 18414 21428 18420 21440
rect 18472 21428 18478 21480
rect 8662 21360 8668 21412
rect 8720 21400 8726 21412
rect 8757 21403 8815 21409
rect 8757 21400 8769 21403
rect 8720 21372 8769 21400
rect 8720 21360 8726 21372
rect 8757 21369 8769 21372
rect 8803 21369 8815 21403
rect 8757 21363 8815 21369
rect 9309 21403 9367 21409
rect 9309 21369 9321 21403
rect 9355 21369 9367 21403
rect 9309 21363 9367 21369
rect 5721 21335 5779 21341
rect 5721 21301 5733 21335
rect 5767 21332 5779 21335
rect 6914 21332 6920 21344
rect 5767 21304 6920 21332
rect 5767 21301 5779 21304
rect 5721 21295 5779 21301
rect 6914 21292 6920 21304
rect 6972 21292 6978 21344
rect 7098 21332 7104 21344
rect 7059 21304 7104 21332
rect 7098 21292 7104 21304
rect 7156 21292 7162 21344
rect 7699 21335 7757 21341
rect 7699 21301 7711 21335
rect 7745 21332 7757 21335
rect 7926 21332 7932 21344
rect 7745 21304 7932 21332
rect 7745 21301 7757 21304
rect 7699 21295 7757 21301
rect 7926 21292 7932 21304
rect 7984 21292 7990 21344
rect 8110 21332 8116 21344
rect 8071 21304 8116 21332
rect 8110 21292 8116 21304
rect 8168 21292 8174 21344
rect 8478 21292 8484 21344
rect 8536 21332 8542 21344
rect 9324 21332 9352 21363
rect 10042 21332 10048 21344
rect 8536 21304 10048 21332
rect 8536 21292 8542 21304
rect 10042 21292 10048 21304
rect 10100 21292 10106 21344
rect 11054 21292 11060 21344
rect 11112 21332 11118 21344
rect 11716 21341 11744 21428
rect 13541 21403 13599 21409
rect 13541 21369 13553 21403
rect 13587 21369 13599 21403
rect 13541 21363 13599 21369
rect 14093 21403 14151 21409
rect 14093 21369 14105 21403
rect 14139 21400 14151 21403
rect 14366 21400 14372 21412
rect 14139 21372 14372 21400
rect 14139 21369 14151 21372
rect 14093 21363 14151 21369
rect 11287 21335 11345 21341
rect 11287 21332 11299 21335
rect 11112 21304 11299 21332
rect 11112 21292 11118 21304
rect 11287 21301 11299 21304
rect 11333 21301 11345 21335
rect 11287 21295 11345 21301
rect 11701 21335 11759 21341
rect 11701 21301 11713 21335
rect 11747 21332 11759 21335
rect 11790 21332 11796 21344
rect 11747 21304 11796 21332
rect 11747 21301 11759 21304
rect 11701 21295 11759 21301
rect 11790 21292 11796 21304
rect 11848 21292 11854 21344
rect 12069 21335 12127 21341
rect 12069 21301 12081 21335
rect 12115 21332 12127 21335
rect 12526 21332 12532 21344
rect 12115 21304 12532 21332
rect 12115 21301 12127 21304
rect 12069 21295 12127 21301
rect 12526 21292 12532 21304
rect 12584 21292 12590 21344
rect 12897 21335 12955 21341
rect 12897 21301 12909 21335
rect 12943 21332 12955 21335
rect 12986 21332 12992 21344
rect 12943 21304 12992 21332
rect 12943 21301 12955 21304
rect 12897 21295 12955 21301
rect 12986 21292 12992 21304
rect 13044 21292 13050 21344
rect 13078 21292 13084 21344
rect 13136 21332 13142 21344
rect 13173 21335 13231 21341
rect 13173 21332 13185 21335
rect 13136 21304 13185 21332
rect 13136 21292 13142 21304
rect 13173 21301 13185 21304
rect 13219 21332 13231 21335
rect 13556 21332 13584 21363
rect 14366 21360 14372 21372
rect 14424 21360 14430 21412
rect 17083 21403 17141 21409
rect 17083 21369 17095 21403
rect 17129 21400 17141 21403
rect 17954 21400 17960 21412
rect 17129 21372 17960 21400
rect 17129 21369 17141 21372
rect 17083 21363 17141 21369
rect 17954 21360 17960 21372
rect 18012 21360 18018 21412
rect 18524 21400 18552 21508
rect 18598 21496 18604 21548
rect 18656 21536 18662 21548
rect 20916 21536 20944 21632
rect 18656 21508 18701 21536
rect 20523 21508 20944 21536
rect 18656 21496 18662 21508
rect 20523 21477 20551 21508
rect 19128 21471 19186 21477
rect 19128 21437 19140 21471
rect 19174 21468 19186 21471
rect 19337 21471 19395 21477
rect 19337 21468 19349 21471
rect 19174 21440 19349 21468
rect 19174 21437 19186 21440
rect 19128 21431 19186 21437
rect 19337 21437 19349 21440
rect 19383 21437 19395 21471
rect 19337 21431 19395 21437
rect 20492 21471 20551 21477
rect 20492 21437 20504 21471
rect 20538 21440 20551 21471
rect 20579 21471 20637 21477
rect 20538 21437 20550 21440
rect 20492 21431 20550 21437
rect 20579 21437 20591 21471
rect 20625 21468 20637 21471
rect 20898 21468 20904 21480
rect 20625 21440 20904 21468
rect 20625 21437 20637 21440
rect 20579 21431 20637 21437
rect 20898 21428 20904 21440
rect 20956 21428 20962 21480
rect 22830 21400 22836 21412
rect 18524 21372 22836 21400
rect 22830 21360 22836 21372
rect 22888 21360 22894 21412
rect 13219 21304 13584 21332
rect 13219 21301 13231 21304
rect 13173 21295 13231 21301
rect 15562 21292 15568 21344
rect 15620 21332 15626 21344
rect 16071 21335 16129 21341
rect 16071 21332 16083 21335
rect 15620 21304 16083 21332
rect 15620 21292 15626 21304
rect 16071 21301 16083 21304
rect 16117 21301 16129 21335
rect 16071 21295 16129 21301
rect 17218 21292 17224 21344
rect 17276 21332 17282 21344
rect 17405 21335 17463 21341
rect 17405 21332 17417 21335
rect 17276 21304 17417 21332
rect 17276 21292 17282 21304
rect 17405 21301 17417 21304
rect 17451 21301 17463 21335
rect 17405 21295 17463 21301
rect 18046 21292 18052 21344
rect 18104 21332 18110 21344
rect 18233 21335 18291 21341
rect 18233 21332 18245 21335
rect 18104 21304 18245 21332
rect 18104 21292 18110 21304
rect 18233 21301 18245 21304
rect 18279 21301 18291 21335
rect 18233 21295 18291 21301
rect 18598 21292 18604 21344
rect 18656 21332 18662 21344
rect 18877 21335 18935 21341
rect 18877 21332 18889 21335
rect 18656 21304 18889 21332
rect 18656 21292 18662 21304
rect 18877 21301 18889 21304
rect 18923 21301 18935 21335
rect 18877 21295 18935 21301
rect 19337 21335 19395 21341
rect 19337 21301 19349 21335
rect 19383 21332 19395 21335
rect 19613 21335 19671 21341
rect 19613 21332 19625 21335
rect 19383 21304 19625 21332
rect 19383 21301 19395 21304
rect 19337 21295 19395 21301
rect 19613 21301 19625 21304
rect 19659 21332 19671 21335
rect 21542 21332 21548 21344
rect 19659 21304 21548 21332
rect 19659 21301 19671 21304
rect 19613 21295 19671 21301
rect 21542 21292 21548 21304
rect 21600 21292 21606 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 13078 21128 13084 21140
rect 11716 21100 13084 21128
rect 11716 21072 11744 21100
rect 13078 21088 13084 21100
rect 13136 21128 13142 21140
rect 13136 21100 13308 21128
rect 13136 21088 13142 21100
rect 6086 21060 6092 21072
rect 5920 21032 6092 21060
rect 1556 20995 1614 21001
rect 1556 20961 1568 20995
rect 1602 20992 1614 20995
rect 2406 20992 2412 21004
rect 1602 20964 2412 20992
rect 1602 20961 1614 20964
rect 1556 20955 1614 20961
rect 2406 20952 2412 20964
rect 2464 20952 2470 21004
rect 4706 20952 4712 21004
rect 4764 20992 4770 21004
rect 5920 21001 5948 21032
rect 6086 21020 6092 21032
rect 6144 21020 6150 21072
rect 7926 21020 7932 21072
rect 7984 21060 7990 21072
rect 8113 21063 8171 21069
rect 8113 21060 8125 21063
rect 7984 21032 8125 21060
rect 7984 21020 7990 21032
rect 8113 21029 8125 21032
rect 8159 21029 8171 21063
rect 8113 21023 8171 21029
rect 8205 21063 8263 21069
rect 8205 21029 8217 21063
rect 8251 21060 8263 21063
rect 8294 21060 8300 21072
rect 8251 21032 8300 21060
rect 8251 21029 8263 21032
rect 8205 21023 8263 21029
rect 8294 21020 8300 21032
rect 8352 21020 8358 21072
rect 9858 21060 9864 21072
rect 9819 21032 9864 21060
rect 9858 21020 9864 21032
rect 9916 21020 9922 21072
rect 11698 21060 11704 21072
rect 11659 21032 11704 21060
rect 11698 21020 11704 21032
rect 11756 21020 11762 21072
rect 12250 21060 12256 21072
rect 12211 21032 12256 21060
rect 12250 21020 12256 21032
rect 12308 21020 12314 21072
rect 13170 21060 13176 21072
rect 13131 21032 13176 21060
rect 13170 21020 13176 21032
rect 13228 21020 13234 21072
rect 13280 21069 13308 21100
rect 15654 21088 15660 21140
rect 15712 21128 15718 21140
rect 22646 21128 22652 21140
rect 15712 21100 22652 21128
rect 15712 21088 15718 21100
rect 22646 21088 22652 21100
rect 22704 21088 22710 21140
rect 13265 21063 13323 21069
rect 13265 21029 13277 21063
rect 13311 21060 13323 21063
rect 14090 21060 14096 21072
rect 13311 21032 14096 21060
rect 13311 21029 13323 21032
rect 13265 21023 13323 21029
rect 14090 21020 14096 21032
rect 14148 21020 14154 21072
rect 16390 21020 16396 21072
rect 16448 21060 16454 21072
rect 16448 21032 20979 21060
rect 16448 21020 16454 21032
rect 4836 20995 4894 21001
rect 4836 20992 4848 20995
rect 4764 20964 4848 20992
rect 4764 20952 4770 20964
rect 4836 20961 4848 20964
rect 4882 20961 4894 20995
rect 4836 20955 4894 20961
rect 5905 20995 5963 21001
rect 5905 20961 5917 20995
rect 5951 20961 5963 20995
rect 6273 20995 6331 21001
rect 6273 20992 6285 20995
rect 5905 20955 5963 20961
rect 6012 20964 6285 20992
rect 5442 20884 5448 20936
rect 5500 20924 5506 20936
rect 5721 20927 5779 20933
rect 5721 20924 5733 20927
rect 5500 20896 5733 20924
rect 5500 20884 5506 20896
rect 5721 20893 5733 20896
rect 5767 20924 5779 20927
rect 6012 20924 6040 20964
rect 6273 20961 6285 20964
rect 6319 20961 6331 20995
rect 15378 20992 15384 21004
rect 15339 20964 15384 20992
rect 6273 20955 6331 20961
rect 15378 20952 15384 20964
rect 15436 20952 15442 21004
rect 15654 20952 15660 21004
rect 15712 20992 15718 21004
rect 15841 20995 15899 21001
rect 15841 20992 15853 20995
rect 15712 20964 15853 20992
rect 15712 20952 15718 20964
rect 15841 20961 15853 20964
rect 15887 20961 15899 20995
rect 15841 20955 15899 20961
rect 17012 20995 17070 21001
rect 17012 20961 17024 20995
rect 17058 20992 17070 20995
rect 17310 20992 17316 21004
rect 17058 20964 17316 20992
rect 17058 20961 17070 20964
rect 17012 20955 17070 20961
rect 17310 20952 17316 20964
rect 17368 20952 17374 21004
rect 18024 20995 18082 21001
rect 18024 20961 18036 20995
rect 18070 20992 18082 20995
rect 18138 20992 18144 21004
rect 18070 20964 18144 20992
rect 18070 20961 18082 20964
rect 18024 20955 18082 20961
rect 18138 20952 18144 20964
rect 18196 20952 18202 21004
rect 18690 20952 18696 21004
rect 18748 20992 18754 21004
rect 20951 21001 20979 21032
rect 19004 20995 19062 21001
rect 19004 20992 19016 20995
rect 18748 20964 19016 20992
rect 18748 20952 18754 20964
rect 19004 20961 19016 20964
rect 19050 20961 19062 20995
rect 19004 20955 19062 20961
rect 20936 20995 20994 21001
rect 20936 20961 20948 20995
rect 20982 20992 20994 20995
rect 21634 20992 21640 21004
rect 20982 20964 21640 20992
rect 20982 20961 20994 20964
rect 20936 20955 20994 20961
rect 21634 20952 21640 20964
rect 21692 20952 21698 21004
rect 5767 20896 6040 20924
rect 6549 20927 6607 20933
rect 5767 20893 5779 20896
rect 5721 20887 5779 20893
rect 6549 20893 6561 20927
rect 6595 20924 6607 20927
rect 6822 20924 6828 20936
rect 6595 20896 6828 20924
rect 6595 20893 6607 20896
rect 6549 20887 6607 20893
rect 6822 20884 6828 20896
rect 6880 20884 6886 20936
rect 8386 20924 8392 20936
rect 8347 20896 8392 20924
rect 8386 20884 8392 20896
rect 8444 20884 8450 20936
rect 9766 20924 9772 20936
rect 9727 20896 9772 20924
rect 9766 20884 9772 20896
rect 9824 20884 9830 20936
rect 10042 20924 10048 20936
rect 10003 20896 10048 20924
rect 10042 20884 10048 20896
rect 10100 20884 10106 20936
rect 11425 20927 11483 20933
rect 11425 20893 11437 20927
rect 11471 20924 11483 20927
rect 11609 20927 11667 20933
rect 11609 20924 11621 20927
rect 11471 20896 11621 20924
rect 11471 20893 11483 20896
rect 11425 20887 11483 20893
rect 11609 20893 11621 20896
rect 11655 20924 11667 20927
rect 13446 20924 13452 20936
rect 11655 20896 13452 20924
rect 11655 20893 11667 20896
rect 11609 20887 11667 20893
rect 13446 20884 13452 20896
rect 13504 20884 13510 20936
rect 15746 20884 15752 20936
rect 15804 20924 15810 20936
rect 15933 20927 15991 20933
rect 15933 20924 15945 20927
rect 15804 20896 15945 20924
rect 15804 20884 15810 20896
rect 15933 20893 15945 20896
rect 15979 20893 15991 20927
rect 18156 20924 18184 20952
rect 19518 20924 19524 20936
rect 15933 20887 15991 20893
rect 16316 20896 16896 20924
rect 18156 20896 19524 20924
rect 13722 20856 13728 20868
rect 13683 20828 13728 20856
rect 13722 20816 13728 20828
rect 13780 20816 13786 20868
rect 1118 20748 1124 20800
rect 1176 20788 1182 20800
rect 1627 20791 1685 20797
rect 1627 20788 1639 20791
rect 1176 20760 1639 20788
rect 1176 20748 1182 20760
rect 1627 20757 1639 20760
rect 1673 20757 1685 20791
rect 1627 20751 1685 20757
rect 4939 20791 4997 20797
rect 4939 20757 4951 20791
rect 4985 20788 4997 20791
rect 5074 20788 5080 20800
rect 4985 20760 5080 20788
rect 4985 20757 4997 20760
rect 4939 20751 4997 20757
rect 5074 20748 5080 20760
rect 5132 20748 5138 20800
rect 11790 20748 11796 20800
rect 11848 20788 11854 20800
rect 16316 20788 16344 20896
rect 16390 20816 16396 20868
rect 16448 20856 16454 20868
rect 16761 20859 16819 20865
rect 16761 20856 16773 20859
rect 16448 20828 16773 20856
rect 16448 20816 16454 20828
rect 16761 20825 16773 20828
rect 16807 20825 16819 20859
rect 16868 20856 16896 20896
rect 19518 20884 19524 20896
rect 19576 20884 19582 20936
rect 20346 20856 20352 20868
rect 16868 20828 20352 20856
rect 16761 20819 16819 20825
rect 20346 20816 20352 20828
rect 20404 20816 20410 20868
rect 20438 20816 20444 20868
rect 20496 20856 20502 20868
rect 21039 20859 21097 20865
rect 21039 20856 21051 20859
rect 20496 20828 21051 20856
rect 20496 20816 20502 20828
rect 21039 20825 21051 20828
rect 21085 20825 21097 20859
rect 21039 20819 21097 20825
rect 16482 20788 16488 20800
rect 11848 20760 16344 20788
rect 16443 20760 16488 20788
rect 11848 20748 11854 20760
rect 16482 20748 16488 20760
rect 16540 20748 16546 20800
rect 16850 20748 16856 20800
rect 16908 20788 16914 20800
rect 17083 20791 17141 20797
rect 17083 20788 17095 20791
rect 16908 20760 17095 20788
rect 16908 20748 16914 20760
rect 17083 20757 17095 20760
rect 17129 20757 17141 20791
rect 17083 20751 17141 20757
rect 18095 20791 18153 20797
rect 18095 20757 18107 20791
rect 18141 20788 18153 20791
rect 18230 20788 18236 20800
rect 18141 20760 18236 20788
rect 18141 20757 18153 20760
rect 18095 20751 18153 20757
rect 18230 20748 18236 20760
rect 18288 20748 18294 20800
rect 19107 20791 19165 20797
rect 19107 20757 19119 20791
rect 19153 20788 19165 20791
rect 20622 20788 20628 20800
rect 19153 20760 20628 20788
rect 19153 20757 19165 20760
rect 19107 20751 19165 20757
rect 20622 20748 20628 20760
rect 20680 20748 20686 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1578 20584 1584 20596
rect 1539 20556 1584 20584
rect 1578 20544 1584 20556
rect 1636 20544 1642 20596
rect 4706 20584 4712 20596
rect 1964 20556 4712 20584
rect 1302 20340 1308 20392
rect 1360 20380 1366 20392
rect 1964 20389 1992 20556
rect 4706 20544 4712 20556
rect 4764 20544 4770 20596
rect 8113 20587 8171 20593
rect 8113 20553 8125 20587
rect 8159 20584 8171 20587
rect 8294 20584 8300 20596
rect 8159 20556 8300 20584
rect 8159 20553 8171 20556
rect 8113 20547 8171 20553
rect 8294 20544 8300 20556
rect 8352 20544 8358 20596
rect 8757 20587 8815 20593
rect 8757 20553 8769 20587
rect 8803 20584 8815 20587
rect 9030 20584 9036 20596
rect 8803 20556 9036 20584
rect 8803 20553 8815 20556
rect 8757 20547 8815 20553
rect 9030 20544 9036 20556
rect 9088 20584 9094 20596
rect 9858 20584 9864 20596
rect 9088 20556 9864 20584
rect 9088 20544 9094 20556
rect 9858 20544 9864 20556
rect 9916 20584 9922 20596
rect 11425 20587 11483 20593
rect 11425 20584 11437 20587
rect 9916 20556 11437 20584
rect 9916 20544 9922 20556
rect 11425 20553 11437 20556
rect 11471 20553 11483 20587
rect 11425 20547 11483 20553
rect 12158 20544 12164 20596
rect 12216 20584 12222 20596
rect 12897 20587 12955 20593
rect 12897 20584 12909 20587
rect 12216 20556 12909 20584
rect 12216 20544 12222 20556
rect 12897 20553 12909 20556
rect 12943 20553 12955 20587
rect 12897 20547 12955 20553
rect 4065 20519 4123 20525
rect 4065 20485 4077 20519
rect 4111 20516 4123 20519
rect 4154 20516 4160 20528
rect 4111 20488 4160 20516
rect 4111 20485 4123 20488
rect 4065 20479 4123 20485
rect 4154 20476 4160 20488
rect 4212 20516 4218 20528
rect 5442 20516 5448 20528
rect 4212 20488 5448 20516
rect 4212 20476 4218 20488
rect 5442 20476 5448 20488
rect 5500 20476 5506 20528
rect 10137 20519 10195 20525
rect 10137 20516 10149 20519
rect 6701 20488 10149 20516
rect 6701 20448 6729 20488
rect 10137 20485 10149 20488
rect 10183 20516 10195 20519
rect 10229 20519 10287 20525
rect 10229 20516 10241 20519
rect 10183 20488 10241 20516
rect 10183 20485 10195 20488
rect 10137 20479 10195 20485
rect 10229 20485 10241 20488
rect 10275 20485 10287 20519
rect 10229 20479 10287 20485
rect 6822 20448 6828 20460
rect 4908 20420 6729 20448
rect 6783 20420 6828 20448
rect 4908 20389 4936 20420
rect 6822 20408 6828 20420
rect 6880 20408 6886 20460
rect 8938 20448 8944 20460
rect 8851 20420 8944 20448
rect 8938 20408 8944 20420
rect 8996 20448 9002 20460
rect 11054 20448 11060 20460
rect 8996 20420 11060 20448
rect 8996 20408 9002 20420
rect 11054 20408 11060 20420
rect 11112 20408 11118 20460
rect 11698 20408 11704 20460
rect 11756 20448 11762 20460
rect 11885 20451 11943 20457
rect 11885 20448 11897 20451
rect 11756 20420 11897 20448
rect 11756 20408 11762 20420
rect 11885 20417 11897 20420
rect 11931 20448 11943 20451
rect 12161 20451 12219 20457
rect 12161 20448 12173 20451
rect 11931 20420 12173 20448
rect 11931 20417 11943 20420
rect 11885 20411 11943 20417
rect 12161 20417 12173 20420
rect 12207 20417 12219 20451
rect 12912 20448 12940 20547
rect 14366 20544 14372 20596
rect 14424 20584 14430 20596
rect 15654 20584 15660 20596
rect 14424 20556 15056 20584
rect 15615 20556 15660 20584
rect 14424 20544 14430 20556
rect 12986 20476 12992 20528
rect 13044 20516 13050 20528
rect 14093 20519 14151 20525
rect 14093 20516 14105 20519
rect 13044 20488 14105 20516
rect 13044 20476 13050 20488
rect 14093 20485 14105 20488
rect 14139 20516 14151 20519
rect 14461 20519 14519 20525
rect 14461 20516 14473 20519
rect 14139 20488 14473 20516
rect 14139 20485 14151 20488
rect 14093 20479 14151 20485
rect 14461 20485 14473 20488
rect 14507 20516 14519 20519
rect 14826 20516 14832 20528
rect 14507 20488 14832 20516
rect 14507 20485 14519 20488
rect 14461 20479 14519 20485
rect 14826 20476 14832 20488
rect 14884 20476 14890 20528
rect 13173 20451 13231 20457
rect 13173 20448 13185 20451
rect 12912 20420 13185 20448
rect 12161 20411 12219 20417
rect 13173 20417 13185 20420
rect 13219 20417 13231 20451
rect 14734 20448 14740 20460
rect 14695 20420 14740 20448
rect 13173 20411 13231 20417
rect 14734 20408 14740 20420
rect 14792 20408 14798 20460
rect 15028 20457 15056 20556
rect 15654 20544 15660 20556
rect 15712 20584 15718 20596
rect 16666 20584 16672 20596
rect 15712 20556 16672 20584
rect 15712 20544 15718 20556
rect 16666 20544 16672 20556
rect 16724 20544 16730 20596
rect 17310 20584 17316 20596
rect 17271 20556 17316 20584
rect 17310 20544 17316 20556
rect 17368 20584 17374 20596
rect 21634 20584 21640 20596
rect 17368 20556 19334 20584
rect 21595 20556 21640 20584
rect 17368 20544 17374 20556
rect 15378 20476 15384 20528
rect 15436 20516 15442 20528
rect 16117 20519 16175 20525
rect 16117 20516 16129 20519
rect 15436 20488 16129 20516
rect 15436 20476 15442 20488
rect 16117 20485 16129 20488
rect 16163 20516 16175 20519
rect 18966 20516 18972 20528
rect 16163 20488 18972 20516
rect 16163 20485 16175 20488
rect 16117 20479 16175 20485
rect 18966 20476 18972 20488
rect 19024 20476 19030 20528
rect 15013 20451 15071 20457
rect 15013 20417 15025 20451
rect 15059 20417 15071 20451
rect 19306 20448 19334 20556
rect 21634 20544 21640 20556
rect 21692 20544 21698 20596
rect 20346 20476 20352 20528
rect 20404 20516 20410 20528
rect 20806 20516 20812 20528
rect 20404 20488 20812 20516
rect 20404 20476 20410 20488
rect 20806 20476 20812 20488
rect 20864 20516 20870 20528
rect 21652 20516 21680 20544
rect 27614 20516 27620 20528
rect 20864 20488 21404 20516
rect 21652 20488 27620 20516
rect 20864 20476 20870 20488
rect 19306 20420 19907 20448
rect 15013 20411 15071 20417
rect 1397 20383 1455 20389
rect 1397 20380 1409 20383
rect 1360 20352 1409 20380
rect 1360 20340 1366 20352
rect 1397 20349 1409 20352
rect 1443 20380 1455 20383
rect 1949 20383 2007 20389
rect 1949 20380 1961 20383
rect 1443 20352 1961 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 1949 20349 1961 20352
rect 1995 20349 2007 20383
rect 3881 20383 3939 20389
rect 3881 20380 3893 20383
rect 1949 20343 2007 20349
rect 3712 20352 3893 20380
rect 2406 20244 2412 20256
rect 2367 20216 2412 20244
rect 2406 20204 2412 20216
rect 2464 20204 2470 20256
rect 2682 20204 2688 20256
rect 2740 20244 2746 20256
rect 3712 20253 3740 20352
rect 3881 20349 3893 20352
rect 3927 20349 3939 20383
rect 3881 20343 3939 20349
rect 4893 20383 4951 20389
rect 4893 20349 4905 20383
rect 4939 20349 4951 20383
rect 5442 20380 5448 20392
rect 5403 20352 5448 20380
rect 4893 20343 4951 20349
rect 4908 20256 4936 20343
rect 5442 20340 5448 20352
rect 5500 20340 5506 20392
rect 10137 20383 10195 20389
rect 10137 20349 10149 20383
rect 10183 20380 10195 20383
rect 10413 20383 10471 20389
rect 10413 20380 10425 20383
rect 10183 20352 10425 20380
rect 10183 20349 10195 20352
rect 10137 20343 10195 20349
rect 10413 20349 10425 20352
rect 10459 20349 10471 20383
rect 10413 20343 10471 20349
rect 10873 20383 10931 20389
rect 10873 20349 10885 20383
rect 10919 20349 10931 20383
rect 10873 20343 10931 20349
rect 5626 20312 5632 20324
rect 5587 20284 5632 20312
rect 5626 20272 5632 20284
rect 5684 20272 5690 20324
rect 6638 20312 6644 20324
rect 6551 20284 6644 20312
rect 6638 20272 6644 20284
rect 6696 20312 6702 20324
rect 7187 20315 7245 20321
rect 7187 20312 7199 20315
rect 6696 20284 7199 20312
rect 6696 20272 6702 20284
rect 7187 20281 7199 20284
rect 7233 20312 7245 20315
rect 7650 20312 7656 20324
rect 7233 20284 7656 20312
rect 7233 20281 7245 20284
rect 7187 20275 7245 20281
rect 7650 20272 7656 20284
rect 7708 20272 7714 20324
rect 9030 20312 9036 20324
rect 8991 20284 9036 20312
rect 9030 20272 9036 20284
rect 9088 20272 9094 20324
rect 9398 20272 9404 20324
rect 9456 20312 9462 20324
rect 9585 20315 9643 20321
rect 9585 20312 9597 20315
rect 9456 20284 9597 20312
rect 9456 20272 9462 20284
rect 9585 20281 9597 20284
rect 9631 20281 9643 20315
rect 10888 20312 10916 20343
rect 17862 20340 17868 20392
rect 17920 20380 17926 20392
rect 18049 20383 18107 20389
rect 18049 20380 18061 20383
rect 17920 20352 18061 20380
rect 17920 20340 17926 20352
rect 18049 20349 18061 20352
rect 18095 20349 18107 20383
rect 18598 20380 18604 20392
rect 18559 20352 18604 20380
rect 18049 20343 18107 20349
rect 18598 20340 18604 20352
rect 18656 20340 18662 20392
rect 19879 20389 19907 20420
rect 20824 20389 20852 20476
rect 21376 20457 21404 20488
rect 27614 20476 27620 20488
rect 27672 20476 27678 20528
rect 21361 20451 21419 20457
rect 21361 20417 21373 20451
rect 21407 20448 21419 20451
rect 24670 20448 24676 20460
rect 21407 20420 24676 20448
rect 21407 20417 21419 20420
rect 21361 20411 21419 20417
rect 24670 20408 24676 20420
rect 24728 20408 24734 20460
rect 19864 20383 19922 20389
rect 19864 20349 19876 20383
rect 19910 20380 19922 20383
rect 20824 20383 20902 20389
rect 19910 20352 20392 20380
rect 20824 20352 20856 20383
rect 19910 20349 19922 20352
rect 19864 20343 19922 20349
rect 11146 20312 11152 20324
rect 9585 20275 9643 20281
rect 9968 20284 10916 20312
rect 11107 20284 11152 20312
rect 9968 20256 9996 20284
rect 11146 20272 11152 20284
rect 11204 20272 11210 20324
rect 12986 20272 12992 20324
rect 13044 20312 13050 20324
rect 13265 20315 13323 20321
rect 13265 20312 13277 20315
rect 13044 20284 13277 20312
rect 13044 20272 13050 20284
rect 13265 20281 13277 20284
rect 13311 20281 13323 20315
rect 13265 20275 13323 20281
rect 13817 20315 13875 20321
rect 13817 20281 13829 20315
rect 13863 20281 13875 20315
rect 13817 20275 13875 20281
rect 3697 20247 3755 20253
rect 3697 20244 3709 20247
rect 2740 20216 3709 20244
rect 2740 20204 2746 20216
rect 3697 20213 3709 20216
rect 3743 20213 3755 20247
rect 3697 20207 3755 20213
rect 4433 20247 4491 20253
rect 4433 20213 4445 20247
rect 4479 20244 4491 20247
rect 4890 20244 4896 20256
rect 4479 20216 4896 20244
rect 4479 20213 4491 20216
rect 4433 20207 4491 20213
rect 4890 20204 4896 20216
rect 4948 20204 4954 20256
rect 5997 20247 6055 20253
rect 5997 20213 6009 20247
rect 6043 20244 6055 20247
rect 6086 20244 6092 20256
rect 6043 20216 6092 20244
rect 6043 20213 6055 20216
rect 5997 20207 6055 20213
rect 6086 20204 6092 20216
rect 6144 20204 6150 20256
rect 7742 20244 7748 20256
rect 7703 20216 7748 20244
rect 7742 20204 7748 20216
rect 7800 20204 7806 20256
rect 9950 20244 9956 20256
rect 9911 20216 9956 20244
rect 9950 20204 9956 20216
rect 10008 20204 10014 20256
rect 13722 20204 13728 20256
rect 13780 20244 13786 20256
rect 13832 20244 13860 20275
rect 14826 20272 14832 20324
rect 14884 20312 14890 20324
rect 16390 20312 16396 20324
rect 14884 20284 14929 20312
rect 16351 20284 16396 20312
rect 14884 20272 14890 20284
rect 16390 20272 16396 20284
rect 16448 20272 16454 20324
rect 16482 20272 16488 20324
rect 16540 20312 16546 20324
rect 17034 20312 17040 20324
rect 16540 20284 16585 20312
rect 16995 20284 17040 20312
rect 16540 20272 16546 20284
rect 17034 20272 17040 20284
rect 17092 20272 17098 20324
rect 18782 20312 18788 20324
rect 18743 20284 18788 20312
rect 18782 20272 18788 20284
rect 18840 20272 18846 20324
rect 13780 20216 13860 20244
rect 17865 20247 17923 20253
rect 13780 20204 13786 20216
rect 17865 20213 17877 20247
rect 17911 20244 17923 20247
rect 18138 20244 18144 20256
rect 17911 20216 18144 20244
rect 17911 20213 17923 20216
rect 17865 20207 17923 20213
rect 18138 20204 18144 20216
rect 18196 20204 18202 20256
rect 18690 20204 18696 20256
rect 18748 20244 18754 20256
rect 19061 20247 19119 20253
rect 19061 20244 19073 20247
rect 18748 20216 19073 20244
rect 18748 20204 18754 20216
rect 19061 20213 19073 20216
rect 19107 20213 19119 20247
rect 19061 20207 19119 20213
rect 19935 20247 19993 20253
rect 19935 20213 19947 20247
rect 19981 20244 19993 20247
rect 20162 20244 20168 20256
rect 19981 20216 20168 20244
rect 19981 20213 19993 20216
rect 19935 20207 19993 20213
rect 20162 20204 20168 20216
rect 20220 20204 20226 20256
rect 20364 20253 20392 20352
rect 20844 20349 20856 20352
rect 20890 20349 20902 20383
rect 20844 20343 20902 20349
rect 21872 20383 21930 20389
rect 21872 20349 21884 20383
rect 21918 20380 21930 20383
rect 22278 20380 22284 20392
rect 21918 20352 22284 20380
rect 21918 20349 21930 20352
rect 21872 20343 21930 20349
rect 22278 20340 22284 20352
rect 22336 20380 22342 20392
rect 24210 20380 24216 20392
rect 22336 20352 24216 20380
rect 22336 20340 22342 20352
rect 24210 20340 24216 20352
rect 24268 20380 24274 20392
rect 25038 20380 25044 20392
rect 24268 20352 25044 20380
rect 24268 20340 24274 20352
rect 25038 20340 25044 20352
rect 25096 20340 25102 20392
rect 20530 20272 20536 20324
rect 20588 20312 20594 20324
rect 21959 20315 22017 20321
rect 21959 20312 21971 20315
rect 20588 20284 21971 20312
rect 20588 20272 20594 20284
rect 21959 20281 21971 20284
rect 22005 20281 22017 20315
rect 21959 20275 22017 20281
rect 20349 20247 20407 20253
rect 20349 20213 20361 20247
rect 20395 20244 20407 20247
rect 20714 20244 20720 20256
rect 20395 20216 20720 20244
rect 20395 20213 20407 20216
rect 20349 20207 20407 20213
rect 20714 20204 20720 20216
rect 20772 20204 20778 20256
rect 20947 20247 21005 20253
rect 20947 20213 20959 20247
rect 20993 20244 21005 20247
rect 21082 20244 21088 20256
rect 20993 20216 21088 20244
rect 20993 20213 21005 20216
rect 20947 20207 21005 20213
rect 21082 20204 21088 20216
rect 21140 20204 21146 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 5169 20043 5227 20049
rect 5169 20009 5181 20043
rect 5215 20040 5227 20043
rect 5442 20040 5448 20052
rect 5215 20012 5448 20040
rect 5215 20009 5227 20012
rect 5169 20003 5227 20009
rect 5442 20000 5448 20012
rect 5500 20000 5506 20052
rect 7193 20043 7251 20049
rect 7193 20009 7205 20043
rect 7239 20040 7251 20043
rect 7282 20040 7288 20052
rect 7239 20012 7288 20040
rect 7239 20009 7251 20012
rect 7193 20003 7251 20009
rect 7282 20000 7288 20012
rect 7340 20040 7346 20052
rect 7742 20040 7748 20052
rect 7340 20012 7748 20040
rect 7340 20000 7346 20012
rect 7742 20000 7748 20012
rect 7800 20000 7806 20052
rect 7926 20000 7932 20052
rect 7984 20040 7990 20052
rect 8389 20043 8447 20049
rect 8389 20040 8401 20043
rect 7984 20012 8401 20040
rect 7984 20000 7990 20012
rect 8389 20009 8401 20012
rect 8435 20009 8447 20043
rect 8938 20040 8944 20052
rect 8899 20012 8944 20040
rect 8389 20003 8447 20009
rect 8938 20000 8944 20012
rect 8996 20000 9002 20052
rect 9493 20043 9551 20049
rect 9493 20009 9505 20043
rect 9539 20040 9551 20043
rect 9766 20040 9772 20052
rect 9539 20012 9772 20040
rect 9539 20009 9551 20012
rect 9493 20003 9551 20009
rect 9766 20000 9772 20012
rect 9824 20049 9830 20052
rect 9824 20043 9873 20049
rect 9824 20009 9827 20043
rect 9861 20009 9873 20043
rect 9824 20003 9873 20009
rect 9824 20000 9830 20003
rect 11698 20000 11704 20052
rect 11756 20040 11762 20052
rect 11793 20043 11851 20049
rect 11793 20040 11805 20043
rect 11756 20012 11805 20040
rect 11756 20000 11762 20012
rect 11793 20009 11805 20012
rect 11839 20009 11851 20043
rect 11793 20003 11851 20009
rect 12345 20043 12403 20049
rect 12345 20009 12357 20043
rect 12391 20040 12403 20043
rect 12986 20040 12992 20052
rect 12391 20012 12992 20040
rect 12391 20009 12403 20012
rect 12345 20003 12403 20009
rect 12986 20000 12992 20012
rect 13044 20000 13050 20052
rect 13081 20043 13139 20049
rect 13081 20009 13093 20043
rect 13127 20040 13139 20043
rect 13170 20040 13176 20052
rect 13127 20012 13176 20040
rect 13127 20009 13139 20012
rect 13081 20003 13139 20009
rect 13170 20000 13176 20012
rect 13228 20000 13234 20052
rect 13541 20043 13599 20049
rect 13541 20009 13553 20043
rect 13587 20040 13599 20043
rect 13630 20040 13636 20052
rect 13587 20012 13636 20040
rect 13587 20009 13599 20012
rect 13541 20003 13599 20009
rect 13630 20000 13636 20012
rect 13688 20000 13694 20052
rect 14090 20040 14096 20052
rect 14051 20012 14096 20040
rect 14090 20000 14096 20012
rect 14148 20000 14154 20052
rect 14734 20040 14740 20052
rect 14695 20012 14740 20040
rect 14734 20000 14740 20012
rect 14792 20000 14798 20052
rect 16301 20043 16359 20049
rect 16301 20009 16313 20043
rect 16347 20040 16359 20043
rect 16850 20040 16856 20052
rect 16347 20012 16856 20040
rect 16347 20009 16359 20012
rect 16301 20003 16359 20009
rect 16850 20000 16856 20012
rect 16908 20000 16914 20052
rect 17862 20000 17868 20052
rect 17920 20040 17926 20052
rect 18049 20043 18107 20049
rect 18049 20040 18061 20043
rect 17920 20012 18061 20040
rect 17920 20000 17926 20012
rect 18049 20009 18061 20012
rect 18095 20009 18107 20043
rect 18049 20003 18107 20009
rect 1535 19975 1593 19981
rect 1535 19941 1547 19975
rect 1581 19972 1593 19975
rect 5810 19972 5816 19984
rect 1581 19944 5816 19972
rect 1581 19941 1593 19944
rect 1535 19935 1593 19941
rect 5810 19932 5816 19944
rect 5868 19932 5874 19984
rect 5991 19975 6049 19981
rect 5991 19941 6003 19975
rect 6037 19972 6049 19975
rect 6638 19972 6644 19984
rect 6037 19944 6644 19972
rect 6037 19941 6049 19944
rect 5991 19935 6049 19941
rect 6638 19932 6644 19944
rect 6696 19932 6702 19984
rect 6914 19932 6920 19984
rect 6972 19972 6978 19984
rect 7466 19972 7472 19984
rect 6972 19944 7472 19972
rect 6972 19932 6978 19944
rect 7466 19932 7472 19944
rect 7524 19932 7530 19984
rect 7558 19932 7564 19984
rect 7616 19972 7622 19984
rect 8478 19972 8484 19984
rect 7616 19944 8484 19972
rect 7616 19932 7622 19944
rect 8478 19932 8484 19944
rect 8536 19972 8542 19984
rect 8662 19972 8668 19984
rect 8536 19944 8668 19972
rect 8536 19932 8542 19944
rect 8662 19932 8668 19944
rect 8720 19932 8726 19984
rect 15930 19932 15936 19984
rect 15988 19972 15994 19984
rect 16577 19975 16635 19981
rect 16577 19972 16589 19975
rect 15988 19944 16589 19972
rect 15988 19932 15994 19944
rect 16577 19941 16589 19944
rect 16623 19941 16635 19975
rect 16577 19935 16635 19941
rect 1210 19864 1216 19916
rect 1268 19904 1274 19916
rect 1432 19907 1490 19913
rect 1432 19904 1444 19907
rect 1268 19876 1444 19904
rect 1268 19864 1274 19876
rect 1432 19873 1444 19876
rect 1478 19873 1490 19907
rect 1432 19867 1490 19873
rect 4062 19864 4068 19916
rect 4120 19904 4126 19916
rect 4617 19907 4675 19913
rect 4617 19904 4629 19907
rect 4120 19876 4629 19904
rect 4120 19864 4126 19876
rect 4617 19873 4629 19876
rect 4663 19873 4675 19907
rect 5626 19904 5632 19916
rect 5587 19876 5632 19904
rect 4617 19867 4675 19873
rect 5626 19864 5632 19876
rect 5684 19864 5690 19916
rect 9582 19904 9588 19916
rect 9543 19876 9588 19904
rect 9582 19864 9588 19876
rect 9640 19864 9646 19916
rect 11146 19864 11152 19916
rect 11204 19904 11210 19916
rect 11425 19907 11483 19913
rect 11425 19904 11437 19907
rect 11204 19876 11437 19904
rect 11204 19864 11210 19876
rect 11425 19873 11437 19876
rect 11471 19873 11483 19907
rect 11425 19867 11483 19873
rect 14734 19864 14740 19916
rect 14792 19904 14798 19916
rect 15197 19907 15255 19913
rect 15197 19904 15209 19907
rect 14792 19876 15209 19904
rect 14792 19864 14798 19876
rect 15197 19873 15209 19876
rect 15243 19873 15255 19907
rect 15197 19867 15255 19873
rect 18785 19907 18843 19913
rect 18785 19873 18797 19907
rect 18831 19873 18843 19907
rect 18785 19867 18843 19873
rect 5258 19796 5264 19848
rect 5316 19836 5322 19848
rect 5537 19839 5595 19845
rect 5537 19836 5549 19839
rect 5316 19808 5549 19836
rect 5316 19796 5322 19808
rect 5537 19805 5549 19808
rect 5583 19836 5595 19839
rect 8113 19839 8171 19845
rect 8113 19836 8125 19839
rect 5583 19808 8125 19836
rect 5583 19805 5595 19808
rect 5537 19799 5595 19805
rect 8113 19805 8125 19808
rect 8159 19836 8171 19839
rect 9398 19836 9404 19848
rect 8159 19808 9404 19836
rect 8159 19805 8171 19808
rect 8113 19799 8171 19805
rect 9398 19796 9404 19808
rect 9456 19796 9462 19848
rect 12066 19796 12072 19848
rect 12124 19836 12130 19848
rect 12526 19836 12532 19848
rect 12124 19808 12532 19836
rect 12124 19796 12130 19808
rect 12526 19796 12532 19808
rect 12584 19796 12590 19848
rect 13170 19836 13176 19848
rect 13131 19808 13176 19836
rect 13170 19796 13176 19808
rect 13228 19796 13234 19848
rect 15427 19839 15485 19845
rect 15427 19805 15439 19839
rect 15473 19836 15485 19839
rect 16485 19839 16543 19845
rect 16485 19836 16497 19839
rect 15473 19808 16497 19836
rect 15473 19805 15485 19808
rect 15427 19799 15485 19805
rect 16485 19805 16497 19808
rect 16531 19836 16543 19839
rect 16942 19836 16948 19848
rect 16531 19808 16948 19836
rect 16531 19805 16543 19808
rect 16485 19799 16543 19805
rect 16942 19796 16948 19808
rect 17000 19796 17006 19848
rect 6549 19771 6607 19777
rect 6549 19737 6561 19771
rect 6595 19768 6607 19771
rect 7558 19768 7564 19780
rect 6595 19740 7564 19768
rect 6595 19737 6607 19740
rect 6549 19731 6607 19737
rect 7558 19728 7564 19740
rect 7616 19728 7622 19780
rect 13354 19728 13360 19780
rect 13412 19768 13418 19780
rect 16574 19768 16580 19780
rect 13412 19740 16580 19768
rect 13412 19728 13418 19740
rect 16574 19728 16580 19740
rect 16632 19728 16638 19780
rect 17034 19768 17040 19780
rect 16995 19740 17040 19768
rect 17034 19728 17040 19740
rect 17092 19728 17098 19780
rect 18800 19768 18828 19867
rect 18874 19864 18880 19916
rect 18932 19904 18938 19916
rect 19061 19907 19119 19913
rect 19061 19904 19073 19907
rect 18932 19876 19073 19904
rect 18932 19864 18938 19876
rect 19061 19873 19073 19876
rect 19107 19873 19119 19907
rect 19061 19867 19119 19873
rect 20254 19864 20260 19916
rect 20312 19904 20318 19916
rect 20809 19907 20867 19913
rect 20809 19904 20821 19907
rect 20312 19876 20821 19904
rect 20312 19864 20318 19876
rect 20809 19873 20821 19876
rect 20855 19873 20867 19907
rect 20809 19867 20867 19873
rect 19334 19836 19340 19848
rect 19295 19808 19340 19836
rect 19334 19796 19340 19808
rect 19392 19796 19398 19848
rect 22554 19796 22560 19848
rect 22612 19836 22618 19848
rect 22649 19839 22707 19845
rect 22649 19836 22661 19839
rect 22612 19808 22661 19836
rect 22612 19796 22618 19808
rect 22649 19805 22661 19808
rect 22695 19805 22707 19839
rect 23658 19836 23664 19848
rect 23619 19808 23664 19836
rect 22649 19799 22707 19805
rect 23658 19796 23664 19808
rect 23716 19796 23722 19848
rect 24118 19796 24124 19848
rect 24176 19836 24182 19848
rect 24673 19839 24731 19845
rect 24673 19836 24685 19839
rect 24176 19808 24685 19836
rect 24176 19796 24182 19808
rect 24673 19805 24685 19808
rect 24719 19805 24731 19839
rect 24673 19799 24731 19805
rect 19058 19768 19064 19780
rect 18800 19740 19064 19768
rect 19058 19728 19064 19740
rect 19116 19728 19122 19780
rect 2869 19703 2927 19709
rect 2869 19669 2881 19703
rect 2915 19700 2927 19703
rect 2958 19700 2964 19712
rect 2915 19672 2964 19700
rect 2915 19669 2927 19672
rect 2869 19663 2927 19669
rect 2958 19660 2964 19672
rect 3016 19660 3022 19712
rect 3099 19703 3157 19709
rect 3099 19669 3111 19703
rect 3145 19700 3157 19703
rect 3786 19700 3792 19712
rect 3145 19672 3792 19700
rect 3145 19669 3157 19672
rect 3099 19663 3157 19669
rect 3786 19660 3792 19672
rect 3844 19660 3850 19712
rect 3878 19660 3884 19712
rect 3936 19700 3942 19712
rect 4801 19703 4859 19709
rect 4801 19700 4813 19703
rect 3936 19672 4813 19700
rect 3936 19660 3942 19672
rect 4801 19669 4813 19672
rect 4847 19669 4859 19703
rect 4801 19663 4859 19669
rect 9950 19660 9956 19712
rect 10008 19700 10014 19712
rect 10502 19700 10508 19712
rect 10008 19672 10508 19700
rect 10008 19660 10014 19672
rect 10502 19660 10508 19672
rect 10560 19660 10566 19712
rect 12618 19700 12624 19712
rect 12579 19672 12624 19700
rect 12618 19660 12624 19672
rect 12676 19660 12682 19712
rect 18509 19703 18567 19709
rect 18509 19669 18521 19703
rect 18555 19700 18567 19703
rect 18598 19700 18604 19712
rect 18555 19672 18604 19700
rect 18555 19669 18567 19672
rect 18509 19663 18567 19669
rect 18598 19660 18604 19672
rect 18656 19700 18662 19712
rect 19613 19703 19671 19709
rect 19613 19700 19625 19703
rect 18656 19672 19625 19700
rect 18656 19660 18662 19672
rect 19613 19669 19625 19672
rect 19659 19700 19671 19703
rect 19978 19700 19984 19712
rect 19659 19672 19984 19700
rect 19659 19669 19671 19672
rect 19613 19663 19671 19669
rect 19978 19660 19984 19672
rect 20036 19660 20042 19712
rect 20346 19660 20352 19712
rect 20404 19700 20410 19712
rect 21039 19703 21097 19709
rect 21039 19700 21051 19703
rect 20404 19672 21051 19700
rect 20404 19660 20410 19672
rect 21039 19669 21051 19672
rect 21085 19669 21097 19703
rect 21039 19663 21097 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1210 19456 1216 19508
rect 1268 19496 1274 19508
rect 2225 19499 2283 19505
rect 2225 19496 2237 19499
rect 1268 19468 2237 19496
rect 1268 19456 1274 19468
rect 2225 19465 2237 19468
rect 2271 19465 2283 19499
rect 2225 19459 2283 19465
rect 5077 19499 5135 19505
rect 5077 19465 5089 19499
rect 5123 19496 5135 19499
rect 5534 19496 5540 19508
rect 5123 19468 5540 19496
rect 5123 19465 5135 19468
rect 5077 19459 5135 19465
rect 5534 19456 5540 19468
rect 5592 19456 5598 19508
rect 7466 19456 7472 19508
rect 7524 19496 7530 19508
rect 8113 19499 8171 19505
rect 8113 19496 8125 19499
rect 7524 19468 8125 19496
rect 7524 19456 7530 19468
rect 8113 19465 8125 19468
rect 8159 19465 8171 19499
rect 8113 19459 8171 19465
rect 8294 19456 8300 19508
rect 8352 19496 8358 19508
rect 8481 19499 8539 19505
rect 8481 19496 8493 19499
rect 8352 19468 8493 19496
rect 8352 19456 8358 19468
rect 8481 19465 8493 19468
rect 8527 19496 8539 19499
rect 8846 19496 8852 19508
rect 8527 19468 8852 19496
rect 8527 19465 8539 19468
rect 8481 19459 8539 19465
rect 8846 19456 8852 19468
rect 8904 19456 8910 19508
rect 11146 19456 11152 19508
rect 11204 19496 11210 19508
rect 11793 19499 11851 19505
rect 11793 19496 11805 19499
rect 11204 19468 11805 19496
rect 11204 19456 11210 19468
rect 11793 19465 11805 19468
rect 11839 19465 11851 19499
rect 11793 19459 11851 19465
rect 12253 19499 12311 19505
rect 12253 19465 12265 19499
rect 12299 19496 12311 19499
rect 12986 19496 12992 19508
rect 12299 19468 12992 19496
rect 12299 19465 12311 19468
rect 12253 19459 12311 19465
rect 5813 19431 5871 19437
rect 5813 19397 5825 19431
rect 5859 19428 5871 19431
rect 7098 19428 7104 19440
rect 5859 19400 7104 19428
rect 5859 19397 5871 19400
rect 5813 19391 5871 19397
rect 7098 19388 7104 19400
rect 7156 19428 7162 19440
rect 7745 19431 7803 19437
rect 7745 19428 7757 19431
rect 7156 19400 7757 19428
rect 7156 19388 7162 19400
rect 7745 19397 7757 19400
rect 7791 19428 7803 19431
rect 10042 19428 10048 19440
rect 7791 19400 10048 19428
rect 7791 19397 7803 19400
rect 7745 19391 7803 19397
rect 10042 19388 10048 19400
rect 10100 19388 10106 19440
rect 11517 19431 11575 19437
rect 11517 19397 11529 19431
rect 11563 19428 11575 19431
rect 11698 19428 11704 19440
rect 11563 19400 11704 19428
rect 11563 19397 11575 19400
rect 11517 19391 11575 19397
rect 11698 19388 11704 19400
rect 11756 19428 11762 19440
rect 12158 19428 12164 19440
rect 11756 19400 12164 19428
rect 11756 19388 11762 19400
rect 12158 19388 12164 19400
rect 12216 19428 12222 19440
rect 12268 19428 12296 19459
rect 12986 19456 12992 19468
rect 13044 19496 13050 19508
rect 13630 19496 13636 19508
rect 13044 19468 13636 19496
rect 13044 19456 13050 19468
rect 13630 19456 13636 19468
rect 13688 19456 13694 19508
rect 15930 19496 15936 19508
rect 15891 19468 15936 19496
rect 15930 19456 15936 19468
rect 15988 19456 15994 19508
rect 16301 19499 16359 19505
rect 16301 19465 16313 19499
rect 16347 19496 16359 19499
rect 16482 19496 16488 19508
rect 16347 19468 16488 19496
rect 16347 19465 16359 19468
rect 16301 19459 16359 19465
rect 16482 19456 16488 19468
rect 16540 19456 16546 19508
rect 16574 19456 16580 19508
rect 16632 19496 16638 19508
rect 18598 19496 18604 19508
rect 16632 19468 18604 19496
rect 16632 19456 16638 19468
rect 18598 19456 18604 19468
rect 18656 19456 18662 19508
rect 19058 19496 19064 19508
rect 19019 19468 19064 19496
rect 19058 19456 19064 19468
rect 19116 19456 19122 19508
rect 24026 19456 24032 19508
rect 24084 19496 24090 19508
rect 24121 19499 24179 19505
rect 24121 19496 24133 19499
rect 24084 19468 24133 19496
rect 24084 19456 24090 19468
rect 24121 19465 24133 19468
rect 24167 19465 24179 19499
rect 24121 19459 24179 19465
rect 12216 19400 12296 19428
rect 12216 19388 12222 19400
rect 17034 19388 17040 19440
rect 17092 19428 17098 19440
rect 17092 19400 18460 19428
rect 17092 19388 17098 19400
rect 18432 19372 18460 19400
rect 18506 19388 18512 19440
rect 18564 19428 18570 19440
rect 22373 19431 22431 19437
rect 22373 19428 22385 19431
rect 18564 19400 22385 19428
rect 18564 19388 18570 19400
rect 22373 19397 22385 19400
rect 22419 19397 22431 19431
rect 22373 19391 22431 19397
rect 5258 19360 5264 19372
rect 5219 19332 5264 19360
rect 5258 19320 5264 19332
rect 5316 19320 5322 19372
rect 6641 19363 6699 19369
rect 6641 19329 6653 19363
rect 6687 19360 6699 19363
rect 7193 19363 7251 19369
rect 7193 19360 7205 19363
rect 6687 19332 7205 19360
rect 6687 19329 6699 19332
rect 6641 19323 6699 19329
rect 7193 19329 7205 19332
rect 7239 19360 7251 19363
rect 8386 19360 8392 19372
rect 7239 19332 8392 19360
rect 7239 19329 7251 19332
rect 7193 19323 7251 19329
rect 8386 19320 8392 19332
rect 8444 19320 8450 19372
rect 8757 19363 8815 19369
rect 8757 19329 8769 19363
rect 8803 19360 8815 19363
rect 9030 19360 9036 19372
rect 8803 19332 9036 19360
rect 8803 19329 8815 19332
rect 8757 19323 8815 19329
rect 9030 19320 9036 19332
rect 9088 19320 9094 19372
rect 9398 19360 9404 19372
rect 9359 19332 9404 19360
rect 9398 19320 9404 19332
rect 9456 19320 9462 19372
rect 11149 19363 11207 19369
rect 11149 19329 11161 19363
rect 11195 19360 11207 19363
rect 13170 19360 13176 19372
rect 11195 19332 13176 19360
rect 11195 19329 11207 19332
rect 11149 19323 11207 19329
rect 13170 19320 13176 19332
rect 13228 19360 13234 19372
rect 14001 19363 14059 19369
rect 14001 19360 14013 19363
rect 13228 19332 14013 19360
rect 13228 19320 13234 19332
rect 14001 19329 14013 19332
rect 14047 19329 14059 19363
rect 14642 19360 14648 19372
rect 14603 19332 14648 19360
rect 14001 19323 14059 19329
rect 14642 19320 14648 19332
rect 14700 19320 14706 19372
rect 16485 19363 16543 19369
rect 16485 19329 16497 19363
rect 16531 19360 16543 19363
rect 16850 19360 16856 19372
rect 16531 19332 16856 19360
rect 16531 19329 16543 19332
rect 16485 19323 16543 19329
rect 16850 19320 16856 19332
rect 16908 19320 16914 19372
rect 18414 19360 18420 19372
rect 18327 19332 18420 19360
rect 18414 19320 18420 19332
rect 18472 19320 18478 19372
rect 18598 19320 18604 19372
rect 18656 19360 18662 19372
rect 18656 19332 21287 19360
rect 18656 19320 18662 19332
rect 1464 19295 1522 19301
rect 1464 19261 1476 19295
rect 1510 19292 1522 19295
rect 1854 19292 1860 19304
rect 1510 19264 1860 19292
rect 1510 19261 1522 19264
rect 1464 19255 1522 19261
rect 1854 19252 1860 19264
rect 1912 19252 1918 19304
rect 3196 19295 3254 19301
rect 3196 19261 3208 19295
rect 3242 19292 3254 19295
rect 3283 19295 3341 19301
rect 3242 19261 3255 19292
rect 3196 19255 3255 19261
rect 3283 19261 3295 19295
rect 3329 19292 3341 19295
rect 3329 19264 5120 19292
rect 3329 19261 3341 19264
rect 3283 19255 3341 19261
rect 3227 19224 3255 19255
rect 3227 19196 3464 19224
rect 3436 19168 3464 19196
rect 4062 19184 4068 19236
rect 4120 19224 4126 19236
rect 4120 19196 4752 19224
rect 4120 19184 4126 19196
rect 4724 19168 4752 19196
rect 1535 19159 1593 19165
rect 1535 19125 1547 19159
rect 1581 19156 1593 19159
rect 2314 19156 2320 19168
rect 1581 19128 2320 19156
rect 1581 19125 1593 19128
rect 1535 19119 1593 19125
rect 2314 19116 2320 19128
rect 2372 19116 2378 19168
rect 2958 19156 2964 19168
rect 2919 19128 2964 19156
rect 2958 19116 2964 19128
rect 3016 19116 3022 19168
rect 3418 19116 3424 19168
rect 3476 19156 3482 19168
rect 3605 19159 3663 19165
rect 3605 19156 3617 19159
rect 3476 19128 3617 19156
rect 3476 19116 3482 19128
rect 3605 19125 3617 19128
rect 3651 19125 3663 19159
rect 3605 19119 3663 19125
rect 4157 19159 4215 19165
rect 4157 19125 4169 19159
rect 4203 19156 4215 19159
rect 4430 19156 4436 19168
rect 4203 19128 4436 19156
rect 4203 19125 4215 19128
rect 4157 19119 4215 19125
rect 4430 19116 4436 19128
rect 4488 19116 4494 19168
rect 4706 19156 4712 19168
rect 4667 19128 4712 19156
rect 4706 19116 4712 19128
rect 4764 19116 4770 19168
rect 5092 19156 5120 19264
rect 5994 19252 6000 19304
rect 6052 19292 6058 19304
rect 6181 19295 6239 19301
rect 6181 19292 6193 19295
rect 6052 19264 6193 19292
rect 6052 19252 6058 19264
rect 6181 19261 6193 19264
rect 6227 19261 6239 19295
rect 6181 19255 6239 19261
rect 10413 19295 10471 19301
rect 10413 19261 10425 19295
rect 10459 19261 10471 19295
rect 10413 19255 10471 19261
rect 5350 19184 5356 19236
rect 5408 19224 5414 19236
rect 6822 19224 6828 19236
rect 5408 19196 5453 19224
rect 6104 19196 6828 19224
rect 5408 19184 5414 19196
rect 6104 19156 6132 19196
rect 6822 19184 6828 19196
rect 6880 19184 6886 19236
rect 7282 19184 7288 19236
rect 7340 19224 7346 19236
rect 7340 19196 7385 19224
rect 7340 19184 7346 19196
rect 8846 19184 8852 19236
rect 8904 19224 8910 19236
rect 8904 19196 8949 19224
rect 8904 19184 8910 19196
rect 5092 19128 6132 19156
rect 8386 19116 8392 19168
rect 8444 19156 8450 19168
rect 9582 19156 9588 19168
rect 8444 19128 9588 19156
rect 8444 19116 8450 19128
rect 9582 19116 9588 19128
rect 9640 19156 9646 19168
rect 9677 19159 9735 19165
rect 9677 19156 9689 19159
rect 9640 19128 9689 19156
rect 9640 19116 9646 19128
rect 9677 19125 9689 19128
rect 9723 19125 9735 19159
rect 9677 19119 9735 19125
rect 10134 19116 10140 19168
rect 10192 19156 10198 19168
rect 10229 19159 10287 19165
rect 10229 19156 10241 19159
rect 10192 19128 10241 19156
rect 10192 19116 10198 19128
rect 10229 19125 10241 19128
rect 10275 19156 10287 19159
rect 10428 19156 10456 19255
rect 10502 19252 10508 19304
rect 10560 19292 10566 19304
rect 10965 19295 11023 19301
rect 10965 19292 10977 19295
rect 10560 19264 10977 19292
rect 10560 19252 10566 19264
rect 10965 19261 10977 19264
rect 11011 19261 11023 19295
rect 10965 19255 11023 19261
rect 10980 19224 11008 19255
rect 11514 19252 11520 19304
rect 11572 19292 11578 19304
rect 12437 19295 12495 19301
rect 12437 19292 12449 19295
rect 11572 19264 12449 19292
rect 11572 19252 11578 19264
rect 12437 19261 12449 19264
rect 12483 19292 12495 19295
rect 12618 19292 12624 19304
rect 12483 19264 12624 19292
rect 12483 19261 12495 19264
rect 12437 19255 12495 19261
rect 12618 19252 12624 19264
rect 12676 19252 12682 19304
rect 17129 19295 17187 19301
rect 17129 19261 17141 19295
rect 17175 19292 17187 19295
rect 17862 19292 17868 19304
rect 17175 19264 17868 19292
rect 17175 19261 17187 19264
rect 17129 19255 17187 19261
rect 17862 19252 17868 19264
rect 17920 19252 17926 19304
rect 19613 19295 19671 19301
rect 19613 19261 19625 19295
rect 19659 19261 19671 19295
rect 19613 19255 19671 19261
rect 11146 19224 11152 19236
rect 10980 19196 11152 19224
rect 11146 19184 11152 19196
rect 11204 19184 11210 19236
rect 12799 19227 12857 19233
rect 12799 19193 12811 19227
rect 12845 19224 12857 19227
rect 12986 19224 12992 19236
rect 12845 19196 12992 19224
rect 12845 19193 12857 19196
rect 12799 19187 12857 19193
rect 12986 19184 12992 19196
rect 13044 19184 13050 19236
rect 14274 19224 14280 19236
rect 14235 19196 14280 19224
rect 14274 19184 14280 19196
rect 14332 19184 14338 19236
rect 14366 19184 14372 19236
rect 14424 19224 14430 19236
rect 14424 19196 14469 19224
rect 14424 19184 14430 19196
rect 16574 19184 16580 19236
rect 16632 19224 16638 19236
rect 18141 19227 18199 19233
rect 18141 19224 18153 19227
rect 16632 19196 16677 19224
rect 17420 19196 18153 19224
rect 16632 19184 16638 19196
rect 10275 19128 10456 19156
rect 13357 19159 13415 19165
rect 10275 19125 10287 19128
rect 10229 19119 10287 19125
rect 13357 19125 13369 19159
rect 13403 19156 13415 19159
rect 14090 19156 14096 19168
rect 13403 19128 14096 19156
rect 13403 19125 13415 19128
rect 13357 19119 13415 19125
rect 14090 19116 14096 19128
rect 14148 19116 14154 19168
rect 14734 19116 14740 19168
rect 14792 19156 14798 19168
rect 15289 19159 15347 19165
rect 15289 19156 15301 19159
rect 14792 19128 15301 19156
rect 14792 19116 14798 19128
rect 15289 19125 15301 19128
rect 15335 19125 15347 19159
rect 15289 19119 15347 19125
rect 17310 19116 17316 19168
rect 17368 19156 17374 19168
rect 17420 19165 17448 19196
rect 18141 19193 18153 19196
rect 18187 19193 18199 19227
rect 18141 19187 18199 19193
rect 18233 19227 18291 19233
rect 18233 19193 18245 19227
rect 18279 19193 18291 19227
rect 18233 19187 18291 19193
rect 17405 19159 17463 19165
rect 17405 19156 17417 19159
rect 17368 19128 17417 19156
rect 17368 19116 17374 19128
rect 17405 19125 17417 19128
rect 17451 19125 17463 19159
rect 17405 19119 17463 19125
rect 17494 19116 17500 19168
rect 17552 19156 17558 19168
rect 17865 19159 17923 19165
rect 17865 19156 17877 19159
rect 17552 19128 17877 19156
rect 17552 19116 17558 19128
rect 17865 19125 17877 19128
rect 17911 19156 17923 19159
rect 18248 19156 18276 19187
rect 18966 19184 18972 19236
rect 19024 19224 19030 19236
rect 19429 19227 19487 19233
rect 19429 19224 19441 19227
rect 19024 19196 19441 19224
rect 19024 19184 19030 19196
rect 19429 19193 19441 19196
rect 19475 19224 19487 19227
rect 19628 19224 19656 19255
rect 19978 19252 19984 19304
rect 20036 19292 20042 19304
rect 21259 19301 21287 19332
rect 20073 19295 20131 19301
rect 20073 19292 20085 19295
rect 20036 19264 20085 19292
rect 20036 19252 20042 19264
rect 20073 19261 20085 19264
rect 20119 19261 20131 19295
rect 20073 19255 20131 19261
rect 21244 19295 21302 19301
rect 21244 19261 21256 19295
rect 21290 19261 21302 19295
rect 21244 19255 21302 19261
rect 19475 19196 19656 19224
rect 21259 19224 21287 19255
rect 21726 19252 21732 19304
rect 21784 19292 21790 19304
rect 22189 19295 22247 19301
rect 22189 19292 22201 19295
rect 21784 19264 22201 19292
rect 21784 19252 21790 19264
rect 22189 19261 22201 19264
rect 22235 19292 22247 19295
rect 22649 19295 22707 19301
rect 22649 19292 22661 19295
rect 22235 19264 22661 19292
rect 22235 19261 22247 19264
rect 22189 19255 22247 19261
rect 22649 19261 22661 19264
rect 22695 19261 22707 19295
rect 22649 19255 22707 19261
rect 23912 19295 23970 19301
rect 23912 19261 23924 19295
rect 23958 19261 23970 19295
rect 23912 19255 23970 19261
rect 23927 19224 23955 19255
rect 24397 19227 24455 19233
rect 24397 19224 24409 19227
rect 21259 19196 21772 19224
rect 23927 19196 24409 19224
rect 19475 19193 19487 19196
rect 19429 19187 19487 19193
rect 17911 19128 18276 19156
rect 17911 19125 17923 19128
rect 17865 19119 17923 19125
rect 19518 19116 19524 19168
rect 19576 19156 19582 19168
rect 19705 19159 19763 19165
rect 19705 19156 19717 19159
rect 19576 19128 19717 19156
rect 19576 19116 19582 19128
rect 19705 19125 19717 19128
rect 19751 19125 19763 19159
rect 19705 19119 19763 19125
rect 20254 19116 20260 19168
rect 20312 19156 20318 19168
rect 20901 19159 20959 19165
rect 20901 19156 20913 19159
rect 20312 19128 20913 19156
rect 20312 19116 20318 19128
rect 20901 19125 20913 19128
rect 20947 19125 20959 19159
rect 20901 19119 20959 19125
rect 21174 19116 21180 19168
rect 21232 19156 21238 19168
rect 21744 19165 21772 19196
rect 24397 19193 24409 19196
rect 24443 19224 24455 19227
rect 24946 19224 24952 19236
rect 24443 19196 24952 19224
rect 24443 19193 24455 19196
rect 24397 19187 24455 19193
rect 24946 19184 24952 19196
rect 25004 19184 25010 19236
rect 21315 19159 21373 19165
rect 21315 19156 21327 19159
rect 21232 19128 21327 19156
rect 21232 19116 21238 19128
rect 21315 19125 21327 19128
rect 21361 19125 21373 19159
rect 21315 19119 21373 19125
rect 21729 19159 21787 19165
rect 21729 19125 21741 19159
rect 21775 19156 21787 19159
rect 22186 19156 22192 19168
rect 21775 19128 22192 19156
rect 21775 19125 21787 19128
rect 21729 19119 21787 19125
rect 22186 19116 22192 19128
rect 22244 19116 22250 19168
rect 24854 19156 24860 19168
rect 24815 19128 24860 19156
rect 24854 19116 24860 19128
rect 24912 19116 24918 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1578 18952 1584 18964
rect 1539 18924 1584 18952
rect 1578 18912 1584 18924
rect 1636 18912 1642 18964
rect 5813 18955 5871 18961
rect 5813 18921 5825 18955
rect 5859 18952 5871 18955
rect 5994 18952 6000 18964
rect 5859 18924 6000 18952
rect 5859 18921 5871 18924
rect 5813 18915 5871 18921
rect 5994 18912 6000 18924
rect 6052 18912 6058 18964
rect 7469 18955 7527 18961
rect 7469 18921 7481 18955
rect 7515 18952 7527 18955
rect 7558 18952 7564 18964
rect 7515 18924 7564 18952
rect 7515 18921 7527 18924
rect 7469 18915 7527 18921
rect 7558 18912 7564 18924
rect 7616 18912 7622 18964
rect 7929 18955 7987 18961
rect 7929 18921 7941 18955
rect 7975 18952 7987 18955
rect 9122 18952 9128 18964
rect 7975 18924 9128 18952
rect 7975 18921 7987 18924
rect 7929 18915 7987 18921
rect 6178 18884 6184 18896
rect 4515 18856 6184 18884
rect 4515 18828 4543 18856
rect 6178 18844 6184 18856
rect 6236 18844 6242 18896
rect 8128 18893 8156 18924
rect 9122 18912 9128 18924
rect 9180 18912 9186 18964
rect 12250 18912 12256 18964
rect 12308 18952 12314 18964
rect 12308 18924 13814 18952
rect 12308 18912 12314 18924
rect 8113 18887 8171 18893
rect 8113 18853 8125 18887
rect 8159 18853 8171 18887
rect 8113 18847 8171 18853
rect 8205 18887 8263 18893
rect 8205 18853 8217 18887
rect 8251 18884 8263 18887
rect 8478 18884 8484 18896
rect 8251 18856 8484 18884
rect 8251 18853 8263 18856
rect 8205 18847 8263 18853
rect 8478 18844 8484 18856
rect 8536 18844 8542 18896
rect 9858 18884 9864 18896
rect 9819 18856 9864 18884
rect 9858 18844 9864 18856
rect 9916 18844 9922 18896
rect 11882 18884 11888 18896
rect 11843 18856 11888 18884
rect 11882 18844 11888 18856
rect 11940 18884 11946 18896
rect 13449 18887 13507 18893
rect 13449 18884 13461 18887
rect 11940 18856 13461 18884
rect 11940 18844 11946 18856
rect 13449 18853 13461 18856
rect 13495 18884 13507 18887
rect 13630 18884 13636 18896
rect 13495 18856 13636 18884
rect 13495 18853 13507 18856
rect 13449 18847 13507 18853
rect 13630 18844 13636 18856
rect 13688 18844 13694 18896
rect 13786 18884 13814 18924
rect 14090 18912 14096 18964
rect 14148 18952 14154 18964
rect 14366 18952 14372 18964
rect 14148 18924 14372 18952
rect 14148 18912 14154 18924
rect 14366 18912 14372 18924
rect 14424 18912 14430 18964
rect 16574 18912 16580 18964
rect 16632 18952 16638 18964
rect 16669 18955 16727 18961
rect 16669 18952 16681 18955
rect 16632 18924 16681 18952
rect 16632 18912 16638 18924
rect 16669 18921 16681 18924
rect 16715 18921 16727 18955
rect 16942 18952 16948 18964
rect 16903 18924 16948 18952
rect 16669 18915 16727 18921
rect 16942 18912 16948 18924
rect 17000 18912 17006 18964
rect 18693 18955 18751 18961
rect 18693 18921 18705 18955
rect 18739 18952 18751 18955
rect 18874 18952 18880 18964
rect 18739 18924 18880 18952
rect 18739 18921 18751 18924
rect 18693 18915 18751 18921
rect 18874 18912 18880 18924
rect 18932 18912 18938 18964
rect 19150 18952 19156 18964
rect 19111 18924 19156 18952
rect 19150 18912 19156 18924
rect 19208 18912 19214 18964
rect 14274 18884 14280 18896
rect 13786 18856 14280 18884
rect 14274 18844 14280 18856
rect 14332 18884 14338 18896
rect 14645 18887 14703 18893
rect 14645 18884 14657 18887
rect 14332 18856 14657 18884
rect 14332 18844 14338 18856
rect 14645 18853 14657 18856
rect 14691 18853 14703 18887
rect 14645 18847 14703 18853
rect 15378 18844 15384 18896
rect 15436 18884 15442 18896
rect 16070 18887 16128 18893
rect 16070 18884 16082 18887
rect 15436 18856 16082 18884
rect 15436 18844 15442 18856
rect 16070 18853 16082 18856
rect 16116 18853 16128 18887
rect 16070 18847 16128 18853
rect 17402 18844 17408 18896
rect 17460 18884 17466 18896
rect 17681 18887 17739 18893
rect 17681 18884 17693 18887
rect 17460 18856 17693 18884
rect 17460 18844 17466 18856
rect 17681 18853 17693 18856
rect 17727 18853 17739 18887
rect 22094 18884 22100 18896
rect 17681 18847 17739 18853
rect 21560 18856 22100 18884
rect 1210 18776 1216 18828
rect 1268 18816 1274 18828
rect 4515 18825 4528 18828
rect 1397 18819 1455 18825
rect 1397 18816 1409 18819
rect 1268 18788 1409 18816
rect 1268 18776 1274 18788
rect 1397 18785 1409 18788
rect 1443 18785 1455 18819
rect 4500 18819 4528 18825
rect 4500 18816 4512 18819
rect 4435 18788 4512 18816
rect 1397 18779 1455 18785
rect 4500 18785 4512 18788
rect 4500 18779 4528 18785
rect 4522 18776 4528 18779
rect 4580 18776 4586 18828
rect 5350 18816 5356 18828
rect 5263 18788 5356 18816
rect 5350 18776 5356 18788
rect 5408 18816 5414 18828
rect 6365 18819 6423 18825
rect 6365 18816 6377 18819
rect 5408 18788 6377 18816
rect 5408 18776 5414 18788
rect 6365 18785 6377 18788
rect 6411 18785 6423 18819
rect 6365 18779 6423 18785
rect 19061 18819 19119 18825
rect 19061 18785 19073 18819
rect 19107 18785 19119 18819
rect 19061 18779 19119 18785
rect 2869 18751 2927 18757
rect 2869 18717 2881 18751
rect 2915 18748 2927 18751
rect 3050 18748 3056 18760
rect 2915 18720 3056 18748
rect 2915 18717 2927 18720
rect 2869 18711 2927 18717
rect 3050 18708 3056 18720
rect 3108 18708 3114 18760
rect 5442 18748 5448 18760
rect 5403 18720 5448 18748
rect 5442 18708 5448 18720
rect 5500 18708 5506 18760
rect 8757 18751 8815 18757
rect 8757 18717 8769 18751
rect 8803 18748 8815 18751
rect 9766 18748 9772 18760
rect 8803 18720 9772 18748
rect 8803 18717 8815 18720
rect 8757 18711 8815 18717
rect 9766 18708 9772 18720
rect 9824 18708 9830 18760
rect 10042 18748 10048 18760
rect 10003 18720 10048 18748
rect 10042 18708 10048 18720
rect 10100 18708 10106 18760
rect 11790 18748 11796 18760
rect 11703 18720 11796 18748
rect 11790 18708 11796 18720
rect 11848 18748 11854 18760
rect 11848 18720 12480 18748
rect 11848 18708 11854 18720
rect 4571 18683 4629 18689
rect 4571 18649 4583 18683
rect 4617 18680 4629 18683
rect 9214 18680 9220 18692
rect 4617 18652 9220 18680
rect 4617 18649 4629 18652
rect 4571 18643 4629 18649
rect 9214 18640 9220 18652
rect 9272 18640 9278 18692
rect 12250 18640 12256 18692
rect 12308 18680 12314 18692
rect 12345 18683 12403 18689
rect 12345 18680 12357 18683
rect 12308 18652 12357 18680
rect 12308 18640 12314 18652
rect 12345 18649 12357 18652
rect 12391 18649 12403 18683
rect 12452 18680 12480 18720
rect 12894 18708 12900 18760
rect 12952 18748 12958 18760
rect 13354 18748 13360 18760
rect 12952 18720 13360 18748
rect 12952 18708 12958 18720
rect 13354 18708 13360 18720
rect 13412 18708 13418 18760
rect 13722 18748 13728 18760
rect 13683 18720 13728 18748
rect 13722 18708 13728 18720
rect 13780 18708 13786 18760
rect 15749 18751 15807 18757
rect 15749 18717 15761 18751
rect 15795 18748 15807 18751
rect 16114 18748 16120 18760
rect 15795 18720 16120 18748
rect 15795 18717 15807 18720
rect 15749 18711 15807 18717
rect 16114 18708 16120 18720
rect 16172 18708 16178 18760
rect 17586 18748 17592 18760
rect 17547 18720 17592 18748
rect 17586 18708 17592 18720
rect 17644 18708 17650 18760
rect 17862 18748 17868 18760
rect 17823 18720 17868 18748
rect 17862 18708 17868 18720
rect 17920 18708 17926 18760
rect 14458 18680 14464 18692
rect 12452 18652 14464 18680
rect 12345 18643 12403 18649
rect 14458 18640 14464 18652
rect 14516 18640 14522 18692
rect 16390 18640 16396 18692
rect 16448 18680 16454 18692
rect 19076 18680 19104 18779
rect 19426 18776 19432 18828
rect 19484 18816 19490 18828
rect 21560 18825 21588 18856
rect 22094 18844 22100 18856
rect 22152 18844 22158 18896
rect 19521 18819 19579 18825
rect 19521 18816 19533 18819
rect 19484 18788 19533 18816
rect 19484 18776 19490 18788
rect 19521 18785 19533 18788
rect 19567 18785 19579 18819
rect 19521 18779 19579 18785
rect 21545 18819 21603 18825
rect 21545 18785 21557 18819
rect 21591 18785 21603 18819
rect 21545 18779 21603 18785
rect 21634 18776 21640 18828
rect 21692 18816 21698 18828
rect 21729 18819 21787 18825
rect 21729 18816 21741 18819
rect 21692 18788 21741 18816
rect 21692 18776 21698 18788
rect 21729 18785 21741 18788
rect 21775 18785 21787 18819
rect 22830 18816 22836 18828
rect 22791 18788 22836 18816
rect 21729 18779 21787 18785
rect 22830 18776 22836 18788
rect 22888 18776 22894 18828
rect 24464 18819 24522 18825
rect 24464 18785 24476 18819
rect 24510 18816 24522 18819
rect 25038 18816 25044 18828
rect 24510 18788 25044 18816
rect 24510 18785 24522 18788
rect 24464 18779 24522 18785
rect 25038 18776 25044 18788
rect 25096 18776 25102 18828
rect 25409 18819 25467 18825
rect 25409 18785 25421 18819
rect 25455 18816 25467 18819
rect 25498 18816 25504 18828
rect 25455 18788 25504 18816
rect 25455 18785 25467 18788
rect 25409 18779 25467 18785
rect 25498 18776 25504 18788
rect 25556 18776 25562 18828
rect 21818 18748 21824 18760
rect 21779 18720 21824 18748
rect 21818 18708 21824 18720
rect 21876 18708 21882 18760
rect 20714 18680 20720 18692
rect 16448 18652 20720 18680
rect 16448 18640 16454 18652
rect 20714 18640 20720 18652
rect 20772 18640 20778 18692
rect 3099 18615 3157 18621
rect 3099 18581 3111 18615
rect 3145 18612 3157 18615
rect 4338 18612 4344 18624
rect 3145 18584 4344 18612
rect 3145 18581 3157 18584
rect 3099 18575 3157 18581
rect 4338 18572 4344 18584
rect 4396 18572 4402 18624
rect 4982 18612 4988 18624
rect 4895 18584 4988 18612
rect 4982 18572 4988 18584
rect 5040 18612 5046 18624
rect 8570 18612 8576 18624
rect 5040 18584 8576 18612
rect 5040 18572 5046 18584
rect 8570 18572 8576 18584
rect 8628 18572 8634 18624
rect 9122 18612 9128 18624
rect 9083 18584 9128 18612
rect 9122 18572 9128 18584
rect 9180 18572 9186 18624
rect 10873 18615 10931 18621
rect 10873 18581 10885 18615
rect 10919 18612 10931 18615
rect 11146 18612 11152 18624
rect 10919 18584 11152 18612
rect 10919 18581 10931 18584
rect 10873 18575 10931 18581
rect 11146 18572 11152 18584
rect 11204 18572 11210 18624
rect 12618 18572 12624 18624
rect 12676 18612 12682 18624
rect 12713 18615 12771 18621
rect 12713 18612 12725 18615
rect 12676 18584 12725 18612
rect 12676 18572 12682 18584
rect 12713 18581 12725 18584
rect 12759 18581 12771 18615
rect 12713 18575 12771 18581
rect 15657 18615 15715 18621
rect 15657 18581 15669 18615
rect 15703 18612 15715 18615
rect 16206 18612 16212 18624
rect 15703 18584 16212 18612
rect 15703 18581 15715 18584
rect 15657 18575 15715 18581
rect 16206 18572 16212 18584
rect 16264 18572 16270 18624
rect 20070 18612 20076 18624
rect 20031 18584 20076 18612
rect 20070 18572 20076 18584
rect 20128 18572 20134 18624
rect 21177 18615 21235 18621
rect 21177 18581 21189 18615
rect 21223 18612 21235 18615
rect 21266 18612 21272 18624
rect 21223 18584 21272 18612
rect 21223 18581 21235 18584
rect 21177 18575 21235 18581
rect 21266 18572 21272 18584
rect 21324 18572 21330 18624
rect 22278 18572 22284 18624
rect 22336 18612 22342 18624
rect 22971 18615 23029 18621
rect 22971 18612 22983 18615
rect 22336 18584 22983 18612
rect 22336 18572 22342 18584
rect 22971 18581 22983 18584
rect 23017 18581 23029 18615
rect 22971 18575 23029 18581
rect 24535 18615 24593 18621
rect 24535 18581 24547 18615
rect 24581 18612 24593 18615
rect 24670 18612 24676 18624
rect 24581 18584 24676 18612
rect 24581 18581 24593 18584
rect 24535 18575 24593 18581
rect 24670 18572 24676 18584
rect 24728 18572 24734 18624
rect 25130 18572 25136 18624
rect 25188 18612 25194 18624
rect 25547 18615 25605 18621
rect 25547 18612 25559 18615
rect 25188 18584 25559 18612
rect 25188 18572 25194 18584
rect 25547 18581 25559 18584
rect 25593 18581 25605 18615
rect 25547 18575 25605 18581
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1578 18408 1584 18420
rect 1539 18380 1584 18408
rect 1578 18368 1584 18380
rect 1636 18368 1642 18420
rect 2038 18408 2044 18420
rect 1999 18380 2044 18408
rect 2038 18368 2044 18380
rect 2096 18368 2102 18420
rect 8018 18408 8024 18420
rect 4126 18380 8024 18408
rect 3050 18340 3056 18352
rect 2963 18312 3056 18340
rect 3050 18300 3056 18312
rect 3108 18340 3114 18352
rect 4126 18340 4154 18380
rect 8018 18368 8024 18380
rect 8076 18368 8082 18420
rect 8478 18368 8484 18420
rect 8536 18408 8542 18420
rect 8573 18411 8631 18417
rect 8573 18408 8585 18411
rect 8536 18380 8585 18408
rect 8536 18368 8542 18380
rect 8573 18377 8585 18380
rect 8619 18377 8631 18411
rect 8573 18371 8631 18377
rect 8846 18368 8852 18420
rect 8904 18408 8910 18420
rect 8941 18411 8999 18417
rect 8941 18408 8953 18411
rect 8904 18380 8953 18408
rect 8904 18368 8910 18380
rect 8941 18377 8953 18380
rect 8987 18377 8999 18411
rect 10597 18411 10655 18417
rect 10597 18408 10609 18411
rect 8941 18371 8999 18377
rect 9324 18380 10609 18408
rect 4522 18340 4528 18352
rect 3108 18312 4154 18340
rect 4483 18312 4528 18340
rect 3108 18300 3114 18312
rect 4522 18300 4528 18312
rect 4580 18300 4586 18352
rect 6086 18300 6092 18352
rect 6144 18340 6150 18352
rect 9324 18340 9352 18380
rect 10597 18377 10609 18380
rect 10643 18377 10655 18411
rect 11882 18408 11888 18420
rect 11843 18380 11888 18408
rect 10597 18371 10655 18377
rect 9766 18340 9772 18352
rect 6144 18312 9352 18340
rect 9727 18312 9772 18340
rect 6144 18300 6150 18312
rect 9766 18300 9772 18312
rect 9824 18300 9830 18352
rect 4172 18244 5304 18272
rect 4172 18216 4200 18244
rect 5276 18216 5304 18244
rect 5442 18232 5448 18284
rect 5500 18272 5506 18284
rect 5537 18275 5595 18281
rect 5537 18272 5549 18275
rect 5500 18244 5549 18272
rect 5500 18232 5506 18244
rect 5537 18241 5549 18244
rect 5583 18272 5595 18275
rect 6181 18275 6239 18281
rect 6181 18272 6193 18275
rect 5583 18244 6193 18272
rect 5583 18241 5595 18244
rect 5537 18235 5595 18241
rect 6181 18241 6193 18244
rect 6227 18241 6239 18275
rect 6181 18235 6239 18241
rect 6730 18232 6736 18284
rect 6788 18272 6794 18284
rect 9858 18272 9864 18284
rect 6788 18244 9864 18272
rect 6788 18232 6794 18244
rect 9858 18232 9864 18244
rect 9916 18272 9922 18284
rect 10137 18275 10195 18281
rect 10137 18272 10149 18275
rect 9916 18244 10149 18272
rect 9916 18232 9922 18244
rect 10137 18241 10149 18244
rect 10183 18241 10195 18275
rect 10137 18235 10195 18241
rect 1397 18207 1455 18213
rect 1397 18173 1409 18207
rect 1443 18204 1455 18207
rect 2038 18204 2044 18216
rect 1443 18176 2044 18204
rect 1443 18173 1455 18176
rect 1397 18167 1455 18173
rect 2038 18164 2044 18176
rect 2096 18164 2102 18216
rect 3234 18204 3240 18216
rect 2608 18176 3240 18204
rect 1486 18028 1492 18080
rect 1544 18068 1550 18080
rect 2608 18077 2636 18176
rect 3234 18164 3240 18176
rect 3292 18164 3298 18216
rect 3789 18207 3847 18213
rect 3789 18173 3801 18207
rect 3835 18204 3847 18207
rect 4154 18204 4160 18216
rect 3835 18176 4160 18204
rect 3835 18173 3847 18176
rect 3789 18167 3847 18173
rect 4154 18164 4160 18176
rect 4212 18164 4218 18216
rect 4982 18204 4988 18216
rect 4943 18176 4988 18204
rect 4982 18164 4988 18176
rect 5040 18164 5046 18216
rect 5258 18204 5264 18216
rect 5171 18176 5264 18204
rect 5258 18164 5264 18176
rect 5316 18164 5322 18216
rect 7098 18204 7104 18216
rect 6288 18176 7104 18204
rect 3973 18139 4031 18145
rect 3973 18105 3985 18139
rect 4019 18136 4031 18139
rect 6288 18136 6316 18176
rect 7098 18164 7104 18176
rect 7156 18204 7162 18216
rect 7373 18207 7431 18213
rect 7373 18204 7385 18207
rect 7156 18176 7385 18204
rect 7156 18164 7162 18176
rect 7373 18173 7385 18176
rect 7419 18173 7431 18207
rect 7373 18167 7431 18173
rect 8297 18207 8355 18213
rect 8297 18173 8309 18207
rect 8343 18204 8355 18207
rect 8938 18204 8944 18216
rect 8343 18176 8944 18204
rect 8343 18173 8355 18176
rect 8297 18167 8355 18173
rect 8938 18164 8944 18176
rect 8996 18164 9002 18216
rect 10612 18204 10640 18371
rect 11882 18368 11888 18380
rect 11940 18368 11946 18420
rect 13630 18408 13636 18420
rect 13591 18380 13636 18408
rect 13630 18368 13636 18380
rect 13688 18368 13694 18420
rect 15930 18368 15936 18420
rect 15988 18408 15994 18420
rect 16945 18411 17003 18417
rect 16945 18408 16957 18411
rect 15988 18380 16957 18408
rect 15988 18368 15994 18380
rect 16945 18377 16957 18380
rect 16991 18408 17003 18411
rect 17402 18408 17408 18420
rect 16991 18380 17408 18408
rect 16991 18377 17003 18380
rect 16945 18371 17003 18377
rect 17402 18368 17408 18380
rect 17460 18408 17466 18420
rect 17497 18411 17555 18417
rect 17497 18408 17509 18411
rect 17460 18380 17509 18408
rect 17460 18368 17466 18380
rect 17497 18377 17509 18380
rect 17543 18377 17555 18411
rect 17497 18371 17555 18377
rect 17586 18368 17592 18420
rect 17644 18408 17650 18420
rect 18187 18411 18245 18417
rect 18187 18408 18199 18411
rect 17644 18380 18199 18408
rect 17644 18368 17650 18380
rect 18187 18377 18199 18380
rect 18233 18377 18245 18411
rect 18598 18408 18604 18420
rect 18559 18380 18604 18408
rect 18187 18371 18245 18377
rect 18598 18368 18604 18380
rect 18656 18368 18662 18420
rect 18874 18368 18880 18420
rect 18932 18408 18938 18420
rect 20901 18411 20959 18417
rect 20901 18408 20913 18411
rect 18932 18380 20913 18408
rect 18932 18368 18938 18380
rect 20901 18377 20913 18380
rect 20947 18408 20959 18411
rect 21634 18408 21640 18420
rect 20947 18380 21640 18408
rect 20947 18377 20959 18380
rect 20901 18371 20959 18377
rect 21634 18368 21640 18380
rect 21692 18368 21698 18420
rect 24762 18408 24768 18420
rect 24723 18380 24768 18408
rect 24762 18368 24768 18380
rect 24820 18368 24826 18420
rect 18414 18300 18420 18352
rect 18472 18340 18478 18352
rect 20809 18343 20867 18349
rect 20809 18340 20821 18343
rect 18472 18312 20821 18340
rect 18472 18300 18478 18312
rect 20809 18309 20821 18312
rect 20855 18309 20867 18343
rect 20809 18303 20867 18309
rect 11514 18272 11520 18284
rect 11475 18244 11520 18272
rect 11514 18232 11520 18244
rect 11572 18232 11578 18284
rect 13722 18232 13728 18284
rect 13780 18272 13786 18284
rect 13780 18244 14136 18272
rect 13780 18232 13786 18244
rect 10781 18207 10839 18213
rect 10781 18204 10793 18207
rect 10612 18176 10793 18204
rect 10781 18173 10793 18176
rect 10827 18173 10839 18207
rect 10781 18167 10839 18173
rect 11146 18164 11152 18216
rect 11204 18204 11210 18216
rect 11241 18207 11299 18213
rect 11241 18204 11253 18207
rect 11204 18176 11253 18204
rect 11204 18164 11210 18176
rect 11241 18173 11253 18176
rect 11287 18173 11299 18207
rect 11241 18167 11299 18173
rect 11330 18164 11336 18216
rect 11388 18204 11394 18216
rect 12437 18207 12495 18213
rect 12437 18204 12449 18207
rect 11388 18176 12449 18204
rect 11388 18164 11394 18176
rect 12437 18173 12449 18176
rect 12483 18204 12495 18207
rect 12618 18204 12624 18216
rect 12483 18176 12624 18204
rect 12483 18173 12495 18176
rect 12437 18167 12495 18173
rect 12618 18164 12624 18176
rect 12676 18164 12682 18216
rect 13357 18207 13415 18213
rect 13357 18173 13369 18207
rect 13403 18204 13415 18207
rect 14001 18207 14059 18213
rect 14001 18204 14013 18207
rect 13403 18176 14013 18204
rect 13403 18173 13415 18176
rect 13357 18167 13415 18173
rect 14001 18173 14013 18176
rect 14047 18173 14059 18207
rect 14001 18167 14059 18173
rect 7650 18136 7656 18148
rect 4019 18108 6316 18136
rect 7608 18108 7656 18136
rect 4019 18105 4031 18108
rect 3973 18099 4031 18105
rect 7650 18096 7656 18108
rect 7708 18145 7714 18148
rect 7708 18139 7756 18145
rect 7708 18105 7710 18139
rect 7744 18105 7756 18139
rect 9214 18136 9220 18148
rect 9175 18108 9220 18136
rect 7708 18099 7756 18105
rect 7708 18096 7741 18099
rect 9214 18096 9220 18108
rect 9272 18096 9278 18148
rect 9309 18139 9367 18145
rect 9309 18105 9321 18139
rect 9355 18105 9367 18139
rect 12758 18139 12816 18145
rect 12758 18136 12770 18139
rect 9309 18099 9367 18105
rect 12268 18108 12770 18136
rect 2593 18071 2651 18077
rect 2593 18068 2605 18071
rect 1544 18040 2605 18068
rect 1544 18028 1550 18040
rect 2593 18037 2605 18040
rect 2639 18037 2651 18071
rect 2593 18031 2651 18037
rect 5905 18071 5963 18077
rect 5905 18037 5917 18071
rect 5951 18068 5963 18071
rect 5994 18068 6000 18080
rect 5951 18040 6000 18068
rect 5951 18037 5963 18040
rect 5905 18031 5963 18037
rect 5994 18028 6000 18040
rect 6052 18068 6058 18080
rect 6178 18068 6184 18080
rect 6052 18040 6184 18068
rect 6052 18028 6058 18040
rect 6178 18028 6184 18040
rect 6236 18068 6242 18080
rect 7193 18071 7251 18077
rect 7193 18068 7205 18071
rect 6236 18040 7205 18068
rect 6236 18028 6242 18040
rect 7193 18037 7205 18040
rect 7239 18068 7251 18071
rect 7713 18068 7741 18096
rect 7239 18040 7741 18068
rect 7239 18037 7251 18040
rect 7193 18031 7251 18037
rect 8846 18028 8852 18080
rect 8904 18068 8910 18080
rect 9324 18068 9352 18099
rect 12268 18080 12296 18108
rect 12758 18105 12770 18108
rect 12804 18105 12816 18139
rect 12758 18099 12816 18105
rect 12250 18068 12256 18080
rect 8904 18040 9352 18068
rect 12211 18040 12256 18068
rect 8904 18028 8910 18040
rect 12250 18028 12256 18040
rect 12308 18028 12314 18080
rect 13630 18028 13636 18080
rect 13688 18068 13694 18080
rect 13814 18068 13820 18080
rect 13688 18040 13820 18068
rect 13688 18028 13694 18040
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 14016 18068 14044 18167
rect 14108 18136 14136 18244
rect 14366 18232 14372 18284
rect 14424 18272 14430 18284
rect 14642 18272 14648 18284
rect 14424 18244 14648 18272
rect 14424 18232 14430 18244
rect 14642 18232 14648 18244
rect 14700 18272 14706 18284
rect 14921 18275 14979 18281
rect 14921 18272 14933 18275
rect 14700 18244 14933 18272
rect 14700 18232 14706 18244
rect 14921 18241 14933 18244
rect 14967 18272 14979 18275
rect 17678 18272 17684 18284
rect 14967 18244 17684 18272
rect 14967 18241 14979 18244
rect 14921 18235 14979 18241
rect 17678 18232 17684 18244
rect 17736 18232 17742 18284
rect 20257 18275 20315 18281
rect 20257 18241 20269 18275
rect 20303 18272 20315 18275
rect 21453 18275 21511 18281
rect 21453 18272 21465 18275
rect 20303 18244 21465 18272
rect 20303 18241 20315 18244
rect 20257 18235 20315 18241
rect 21453 18241 21465 18244
rect 21499 18272 21511 18275
rect 24946 18272 24952 18284
rect 21499 18244 24952 18272
rect 21499 18241 21511 18244
rect 21453 18235 21511 18241
rect 24946 18232 24952 18244
rect 25004 18232 25010 18284
rect 16025 18207 16083 18213
rect 16025 18173 16037 18207
rect 16071 18204 16083 18207
rect 16206 18204 16212 18216
rect 16071 18176 16212 18204
rect 16071 18173 16083 18176
rect 16025 18167 16083 18173
rect 16206 18164 16212 18176
rect 16264 18164 16270 18216
rect 18116 18207 18174 18213
rect 18116 18173 18128 18207
rect 18162 18204 18174 18207
rect 18598 18204 18604 18216
rect 18162 18176 18604 18204
rect 18162 18173 18174 18176
rect 18116 18167 18174 18173
rect 18598 18164 18604 18176
rect 18656 18164 18662 18216
rect 20625 18207 20683 18213
rect 20625 18173 20637 18207
rect 20671 18204 20683 18207
rect 20714 18204 20720 18216
rect 20671 18176 20720 18204
rect 20671 18173 20683 18176
rect 20625 18167 20683 18173
rect 20714 18164 20720 18176
rect 20772 18164 20778 18216
rect 24121 18207 24179 18213
rect 24121 18173 24133 18207
rect 24167 18204 24179 18207
rect 24581 18207 24639 18213
rect 24581 18204 24593 18207
rect 24167 18176 24593 18204
rect 24167 18173 24179 18176
rect 24121 18167 24179 18173
rect 24581 18173 24593 18176
rect 24627 18204 24639 18207
rect 24670 18204 24676 18216
rect 24627 18176 24676 18204
rect 24627 18173 24639 18176
rect 24581 18167 24639 18173
rect 24670 18164 24676 18176
rect 24728 18164 24734 18216
rect 14274 18136 14280 18148
rect 14108 18108 14280 18136
rect 14274 18096 14280 18108
rect 14332 18096 14338 18148
rect 14369 18139 14427 18145
rect 14369 18105 14381 18139
rect 14415 18105 14427 18139
rect 14369 18099 14427 18105
rect 16346 18139 16404 18145
rect 16346 18105 16358 18139
rect 16392 18105 16404 18139
rect 16346 18099 16404 18105
rect 14384 18068 14412 18099
rect 14016 18040 14412 18068
rect 15378 18028 15384 18080
rect 15436 18068 15442 18080
rect 15473 18071 15531 18077
rect 15473 18068 15485 18071
rect 15436 18040 15485 18068
rect 15436 18028 15442 18040
rect 15473 18037 15485 18040
rect 15519 18068 15531 18071
rect 15841 18071 15899 18077
rect 15841 18068 15853 18071
rect 15519 18040 15853 18068
rect 15519 18037 15531 18040
rect 15473 18031 15531 18037
rect 15841 18037 15853 18040
rect 15887 18068 15899 18071
rect 16361 18068 16389 18099
rect 17862 18096 17868 18148
rect 17920 18136 17926 18148
rect 19613 18139 19671 18145
rect 19613 18136 19625 18139
rect 17920 18108 19625 18136
rect 17920 18096 17926 18108
rect 19613 18105 19625 18108
rect 19659 18105 19671 18139
rect 19613 18099 19671 18105
rect 19705 18139 19763 18145
rect 19705 18105 19717 18139
rect 19751 18136 19763 18139
rect 20070 18136 20076 18148
rect 19751 18108 20076 18136
rect 19751 18105 19763 18108
rect 19705 18099 19763 18105
rect 15887 18040 16389 18068
rect 15887 18037 15899 18040
rect 15841 18031 15899 18037
rect 18598 18028 18604 18080
rect 18656 18068 18662 18080
rect 19061 18071 19119 18077
rect 19061 18068 19073 18071
rect 18656 18040 19073 18068
rect 18656 18028 18662 18040
rect 19061 18037 19073 18040
rect 19107 18068 19119 18071
rect 19426 18068 19432 18080
rect 19107 18040 19432 18068
rect 19107 18037 19119 18040
rect 19061 18031 19119 18037
rect 19426 18028 19432 18040
rect 19484 18028 19490 18080
rect 19628 18068 19656 18099
rect 20070 18096 20076 18108
rect 20128 18096 20134 18148
rect 20809 18139 20867 18145
rect 20809 18105 20821 18139
rect 20855 18136 20867 18139
rect 21177 18139 21235 18145
rect 21177 18136 21189 18139
rect 20855 18108 21189 18136
rect 20855 18105 20867 18108
rect 20809 18099 20867 18105
rect 21177 18105 21189 18108
rect 21223 18105 21235 18139
rect 21177 18099 21235 18105
rect 20254 18068 20260 18080
rect 19628 18040 20260 18068
rect 20254 18028 20260 18040
rect 20312 18028 20318 18080
rect 21192 18068 21220 18099
rect 21266 18096 21272 18148
rect 21324 18136 21330 18148
rect 21324 18108 21369 18136
rect 21324 18096 21330 18108
rect 21358 18068 21364 18080
rect 21192 18040 21364 18068
rect 21358 18028 21364 18040
rect 21416 18028 21422 18080
rect 22094 18068 22100 18080
rect 22055 18040 22100 18068
rect 22094 18028 22100 18040
rect 22152 18028 22158 18080
rect 22830 18068 22836 18080
rect 22791 18040 22836 18068
rect 22830 18028 22836 18040
rect 22888 18028 22894 18080
rect 24489 18071 24547 18077
rect 24489 18037 24501 18071
rect 24535 18068 24547 18071
rect 25038 18068 25044 18080
rect 24535 18040 25044 18068
rect 24535 18037 24547 18040
rect 24489 18031 24547 18037
rect 25038 18028 25044 18040
rect 25096 18028 25102 18080
rect 25498 18068 25504 18080
rect 25459 18040 25504 18068
rect 25498 18028 25504 18040
rect 25556 18028 25562 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 3878 17864 3884 17876
rect 3839 17836 3884 17864
rect 3878 17824 3884 17836
rect 3936 17824 3942 17876
rect 5258 17864 5264 17876
rect 5219 17836 5264 17864
rect 5258 17824 5264 17836
rect 5316 17824 5322 17876
rect 6178 17864 6184 17876
rect 6139 17836 6184 17864
rect 6178 17824 6184 17836
rect 6236 17824 6242 17876
rect 6730 17864 6736 17876
rect 6691 17836 6736 17864
rect 6730 17824 6736 17836
rect 6788 17824 6794 17876
rect 7098 17824 7104 17876
rect 7156 17864 7162 17876
rect 7377 17867 7435 17873
rect 7377 17864 7389 17867
rect 7156 17836 7389 17864
rect 7156 17824 7162 17836
rect 7377 17833 7389 17836
rect 7423 17833 7435 17867
rect 7377 17827 7435 17833
rect 8481 17867 8539 17873
rect 8481 17833 8493 17867
rect 8527 17864 8539 17867
rect 8846 17864 8852 17876
rect 8527 17836 8852 17864
rect 8527 17833 8539 17836
rect 8481 17827 8539 17833
rect 8846 17824 8852 17836
rect 8904 17824 8910 17876
rect 9214 17864 9220 17876
rect 9175 17836 9220 17864
rect 9214 17824 9220 17836
rect 9272 17824 9278 17876
rect 9766 17824 9772 17876
rect 9824 17864 9830 17876
rect 9861 17867 9919 17873
rect 9861 17864 9873 17867
rect 9824 17836 9873 17864
rect 9824 17824 9830 17836
rect 9861 17833 9873 17836
rect 9907 17833 9919 17867
rect 11790 17864 11796 17876
rect 11751 17836 11796 17864
rect 9861 17827 9919 17833
rect 11790 17824 11796 17836
rect 11848 17824 11854 17876
rect 13354 17864 13360 17876
rect 13315 17836 13360 17864
rect 13354 17824 13360 17836
rect 13412 17824 13418 17876
rect 13630 17824 13636 17876
rect 13688 17864 13694 17876
rect 13817 17867 13875 17873
rect 13817 17864 13829 17867
rect 13688 17836 13829 17864
rect 13688 17824 13694 17836
rect 13817 17833 13829 17836
rect 13863 17864 13875 17867
rect 14182 17864 14188 17876
rect 13863 17836 14188 17864
rect 13863 17833 13875 17836
rect 13817 17827 13875 17833
rect 14182 17824 14188 17836
rect 14240 17824 14246 17876
rect 14274 17824 14280 17876
rect 14332 17864 14338 17876
rect 14369 17867 14427 17873
rect 14369 17864 14381 17867
rect 14332 17836 14381 17864
rect 14332 17824 14338 17836
rect 14369 17833 14381 17836
rect 14415 17833 14427 17867
rect 14369 17827 14427 17833
rect 15795 17867 15853 17873
rect 15795 17833 15807 17867
rect 15841 17864 15853 17867
rect 17310 17864 17316 17876
rect 15841 17836 17316 17864
rect 15841 17833 15853 17836
rect 15795 17827 15853 17833
rect 17310 17824 17316 17836
rect 17368 17824 17374 17876
rect 17586 17824 17592 17876
rect 17644 17864 17650 17876
rect 17681 17867 17739 17873
rect 17681 17864 17693 17867
rect 17644 17836 17693 17864
rect 17644 17824 17650 17836
rect 17681 17833 17693 17836
rect 17727 17833 17739 17867
rect 17681 17827 17739 17833
rect 18969 17867 19027 17873
rect 18969 17833 18981 17867
rect 19015 17864 19027 17867
rect 19150 17864 19156 17876
rect 19015 17836 19156 17864
rect 19015 17833 19027 17836
rect 18969 17827 19027 17833
rect 3510 17796 3516 17808
rect 3423 17768 3516 17796
rect 3510 17756 3516 17768
rect 3568 17796 3574 17808
rect 4154 17796 4160 17808
rect 3568 17768 4160 17796
rect 3568 17756 3574 17768
rect 4154 17756 4160 17768
rect 4212 17796 4218 17808
rect 7923 17799 7981 17805
rect 4212 17768 4752 17796
rect 4212 17756 4218 17768
rect 2961 17731 3019 17737
rect 2961 17697 2973 17731
rect 3007 17728 3019 17731
rect 3602 17728 3608 17740
rect 3007 17700 3608 17728
rect 3007 17697 3019 17700
rect 2961 17691 3019 17697
rect 3602 17688 3608 17700
rect 3660 17688 3666 17740
rect 4522 17728 4528 17740
rect 4483 17700 4528 17728
rect 4522 17688 4528 17700
rect 4580 17688 4586 17740
rect 4724 17737 4752 17768
rect 7923 17765 7935 17799
rect 7969 17796 7981 17799
rect 8294 17796 8300 17808
rect 7969 17768 8300 17796
rect 7969 17765 7981 17768
rect 7923 17759 7981 17765
rect 8294 17756 8300 17768
rect 8352 17756 8358 17808
rect 11330 17796 11336 17808
rect 11291 17768 11336 17796
rect 11330 17756 11336 17768
rect 11388 17756 11394 17808
rect 11882 17756 11888 17808
rect 11940 17796 11946 17808
rect 12250 17796 12256 17808
rect 11940 17768 12256 17796
rect 11940 17756 11946 17768
rect 12250 17756 12256 17768
rect 12308 17796 12314 17808
rect 12482 17799 12540 17805
rect 12482 17796 12494 17799
rect 12308 17768 12494 17796
rect 12308 17756 12314 17768
rect 12482 17765 12494 17768
rect 12528 17765 12540 17799
rect 12482 17759 12540 17765
rect 16853 17799 16911 17805
rect 16853 17765 16865 17799
rect 16899 17796 16911 17799
rect 17402 17796 17408 17808
rect 16899 17768 17408 17796
rect 16899 17765 16911 17768
rect 16853 17759 16911 17765
rect 17402 17756 17408 17768
rect 17460 17756 17466 17808
rect 4709 17731 4767 17737
rect 4709 17697 4721 17731
rect 4755 17697 4767 17731
rect 4709 17691 4767 17697
rect 4985 17731 5043 17737
rect 4985 17697 4997 17731
rect 5031 17728 5043 17731
rect 7558 17728 7564 17740
rect 5031 17700 7564 17728
rect 5031 17697 5043 17700
rect 4985 17691 5043 17697
rect 7558 17688 7564 17700
rect 7616 17688 7622 17740
rect 8570 17688 8576 17740
rect 8628 17728 8634 17740
rect 10594 17728 10600 17740
rect 8628 17700 10600 17728
rect 8628 17688 8634 17700
rect 10594 17688 10600 17700
rect 10652 17688 10658 17740
rect 11146 17728 11152 17740
rect 11107 17700 11152 17728
rect 11146 17688 11152 17700
rect 11204 17688 11210 17740
rect 13976 17731 14034 17737
rect 13976 17697 13988 17731
rect 14022 17728 14034 17731
rect 14734 17728 14740 17740
rect 14022 17700 14740 17728
rect 14022 17697 14034 17700
rect 13976 17691 14034 17697
rect 14734 17688 14740 17700
rect 14792 17688 14798 17740
rect 15654 17728 15660 17740
rect 15615 17700 15660 17728
rect 15654 17688 15660 17700
rect 15712 17688 15718 17740
rect 19076 17737 19104 17836
rect 19150 17824 19156 17836
rect 19208 17824 19214 17876
rect 19981 17867 20039 17873
rect 19981 17833 19993 17867
rect 20027 17864 20039 17867
rect 20070 17864 20076 17876
rect 20027 17836 20076 17864
rect 20027 17833 20039 17836
rect 19981 17827 20039 17833
rect 20070 17824 20076 17836
rect 20128 17824 20134 17876
rect 20254 17864 20260 17876
rect 20215 17836 20260 17864
rect 20254 17824 20260 17836
rect 20312 17824 20318 17876
rect 20990 17864 20996 17876
rect 20951 17836 20996 17864
rect 20990 17824 20996 17836
rect 21048 17824 21054 17876
rect 21358 17824 21364 17876
rect 21416 17864 21422 17876
rect 21913 17867 21971 17873
rect 21913 17864 21925 17867
rect 21416 17836 21925 17864
rect 21416 17824 21422 17836
rect 21913 17833 21925 17836
rect 21959 17833 21971 17867
rect 21913 17827 21971 17833
rect 19382 17799 19440 17805
rect 19382 17796 19394 17799
rect 19306 17768 19394 17796
rect 19061 17731 19119 17737
rect 19061 17697 19073 17731
rect 19107 17697 19119 17731
rect 19061 17691 19119 17697
rect 19150 17688 19156 17740
rect 19208 17728 19214 17740
rect 19306 17728 19334 17768
rect 19382 17765 19394 17768
rect 19428 17765 19440 17799
rect 19382 17759 19440 17765
rect 21652 17768 23244 17796
rect 21652 17740 21680 17768
rect 19208 17700 19334 17728
rect 19208 17688 19214 17700
rect 20254 17688 20260 17740
rect 20312 17728 20318 17740
rect 20714 17728 20720 17740
rect 20312 17700 20720 17728
rect 20312 17688 20318 17700
rect 20714 17688 20720 17700
rect 20772 17728 20778 17740
rect 20901 17731 20959 17737
rect 20901 17728 20913 17731
rect 20772 17700 20913 17728
rect 20772 17688 20778 17700
rect 20901 17697 20913 17700
rect 20947 17697 20959 17731
rect 20901 17691 20959 17697
rect 21453 17731 21511 17737
rect 21453 17697 21465 17731
rect 21499 17728 21511 17731
rect 21634 17728 21640 17740
rect 21499 17700 21640 17728
rect 21499 17697 21511 17700
rect 21453 17691 21511 17697
rect 21634 17688 21640 17700
rect 21692 17688 21698 17740
rect 23014 17728 23020 17740
rect 22975 17700 23020 17728
rect 23014 17688 23020 17700
rect 23072 17688 23078 17740
rect 23216 17737 23244 17768
rect 23201 17731 23259 17737
rect 23201 17697 23213 17731
rect 23247 17728 23259 17731
rect 23842 17728 23848 17740
rect 23247 17700 23848 17728
rect 23247 17697 23259 17700
rect 23201 17691 23259 17697
rect 23842 17688 23848 17700
rect 23900 17688 23906 17740
rect 24581 17731 24639 17737
rect 24581 17697 24593 17731
rect 24627 17728 24639 17731
rect 24670 17728 24676 17740
rect 24627 17700 24676 17728
rect 24627 17697 24639 17700
rect 24581 17691 24639 17697
rect 24670 17688 24676 17700
rect 24728 17688 24734 17740
rect 1949 17663 2007 17669
rect 1949 17629 1961 17663
rect 1995 17660 2007 17663
rect 2774 17660 2780 17672
rect 1995 17632 2780 17660
rect 1995 17629 2007 17632
rect 1949 17623 2007 17629
rect 2774 17620 2780 17632
rect 2832 17620 2838 17672
rect 5813 17663 5871 17669
rect 5813 17629 5825 17663
rect 5859 17660 5871 17663
rect 5994 17660 6000 17672
rect 5859 17632 6000 17660
rect 5859 17629 5871 17632
rect 5813 17623 5871 17629
rect 5994 17620 6000 17632
rect 6052 17620 6058 17672
rect 12158 17660 12164 17672
rect 12119 17632 12164 17660
rect 12158 17620 12164 17632
rect 12216 17620 12222 17672
rect 16758 17660 16764 17672
rect 16719 17632 16764 17660
rect 16758 17620 16764 17632
rect 16816 17620 16822 17672
rect 17034 17620 17040 17672
rect 17092 17660 17098 17672
rect 17405 17663 17463 17669
rect 17405 17660 17417 17663
rect 17092 17632 17417 17660
rect 17092 17620 17098 17632
rect 17405 17629 17417 17632
rect 17451 17660 17463 17663
rect 17862 17660 17868 17672
rect 17451 17632 17868 17660
rect 17451 17629 17463 17632
rect 17405 17623 17463 17629
rect 17862 17620 17868 17632
rect 17920 17620 17926 17672
rect 18874 17620 18880 17672
rect 18932 17660 18938 17672
rect 20806 17660 20812 17672
rect 18932 17632 20812 17660
rect 18932 17620 18938 17632
rect 20806 17620 20812 17632
rect 20864 17620 20870 17672
rect 23474 17620 23480 17672
rect 23532 17660 23538 17672
rect 23532 17632 23577 17660
rect 23532 17620 23538 17632
rect 10962 17552 10968 17604
rect 11020 17592 11026 17604
rect 15286 17592 15292 17604
rect 11020 17564 15292 17592
rect 11020 17552 11026 17564
rect 15286 17552 15292 17564
rect 15344 17552 15350 17604
rect 16574 17592 16580 17604
rect 16487 17564 16580 17592
rect 16574 17552 16580 17564
rect 16632 17592 16638 17604
rect 17494 17592 17500 17604
rect 16632 17564 17500 17592
rect 16632 17552 16638 17564
rect 17494 17552 17500 17564
rect 17552 17552 17558 17604
rect 1210 17484 1216 17536
rect 1268 17524 1274 17536
rect 1581 17527 1639 17533
rect 1581 17524 1593 17527
rect 1268 17496 1593 17524
rect 1268 17484 1274 17496
rect 1581 17493 1593 17496
rect 1627 17493 1639 17527
rect 3142 17524 3148 17536
rect 3103 17496 3148 17524
rect 1581 17487 1639 17493
rect 3142 17484 3148 17496
rect 3200 17484 3206 17536
rect 4154 17484 4160 17536
rect 4212 17524 4218 17536
rect 8386 17524 8392 17536
rect 4212 17496 8392 17524
rect 4212 17484 4218 17496
rect 8386 17484 8392 17496
rect 8444 17484 8450 17536
rect 8846 17524 8852 17536
rect 8807 17496 8852 17524
rect 8846 17484 8852 17496
rect 8904 17484 8910 17536
rect 13078 17524 13084 17536
rect 13039 17496 13084 17524
rect 13078 17484 13084 17496
rect 13136 17484 13142 17536
rect 14047 17527 14105 17533
rect 14047 17493 14059 17527
rect 14093 17524 14105 17527
rect 14274 17524 14280 17536
rect 14093 17496 14280 17524
rect 14093 17493 14105 17496
rect 14047 17487 14105 17493
rect 14274 17484 14280 17496
rect 14332 17484 14338 17536
rect 16114 17484 16120 17536
rect 16172 17524 16178 17536
rect 16209 17527 16267 17533
rect 16209 17524 16221 17527
rect 16172 17496 16221 17524
rect 16172 17484 16178 17496
rect 16209 17493 16221 17496
rect 16255 17524 16267 17527
rect 16942 17524 16948 17536
rect 16255 17496 16948 17524
rect 16255 17493 16267 17496
rect 16209 17487 16267 17493
rect 16942 17484 16948 17496
rect 17000 17484 17006 17536
rect 17678 17484 17684 17536
rect 17736 17524 17742 17536
rect 22649 17527 22707 17533
rect 22649 17524 22661 17527
rect 17736 17496 22661 17524
rect 17736 17484 17742 17496
rect 22649 17493 22661 17496
rect 22695 17524 22707 17527
rect 22738 17524 22744 17536
rect 22695 17496 22744 17524
rect 22695 17493 22707 17496
rect 22649 17487 22707 17493
rect 22738 17484 22744 17496
rect 22796 17484 22802 17536
rect 24765 17527 24823 17533
rect 24765 17493 24777 17527
rect 24811 17524 24823 17527
rect 27614 17524 27620 17536
rect 24811 17496 27620 17524
rect 24811 17493 24823 17496
rect 24765 17487 24823 17493
rect 27614 17484 27620 17496
rect 27672 17484 27678 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1578 17320 1584 17332
rect 1539 17292 1584 17320
rect 1578 17280 1584 17292
rect 1636 17280 1642 17332
rect 2041 17323 2099 17329
rect 2041 17289 2053 17323
rect 2087 17320 2099 17323
rect 2130 17320 2136 17332
rect 2087 17292 2136 17320
rect 2087 17289 2099 17292
rect 2041 17283 2099 17289
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17116 1455 17119
rect 2056 17116 2084 17283
rect 2130 17280 2136 17292
rect 2188 17280 2194 17332
rect 2961 17323 3019 17329
rect 2961 17289 2973 17323
rect 3007 17320 3019 17323
rect 3510 17320 3516 17332
rect 3007 17292 3516 17320
rect 3007 17289 3019 17292
rect 2961 17283 3019 17289
rect 3510 17280 3516 17292
rect 3568 17280 3574 17332
rect 8665 17323 8723 17329
rect 8665 17289 8677 17323
rect 8711 17320 8723 17323
rect 8938 17320 8944 17332
rect 8711 17292 8944 17320
rect 8711 17289 8723 17292
rect 8665 17283 8723 17289
rect 8938 17280 8944 17292
rect 8996 17280 9002 17332
rect 10594 17320 10600 17332
rect 10555 17292 10600 17320
rect 10594 17280 10600 17292
rect 10652 17280 10658 17332
rect 11885 17323 11943 17329
rect 11885 17289 11897 17323
rect 11931 17320 11943 17323
rect 12158 17320 12164 17332
rect 11931 17292 12164 17320
rect 11931 17289 11943 17292
rect 11885 17283 11943 17289
rect 4982 17252 4988 17264
rect 3896 17224 4988 17252
rect 1443 17088 2084 17116
rect 3053 17119 3111 17125
rect 1443 17085 1455 17088
rect 1397 17079 1455 17085
rect 3053 17085 3065 17119
rect 3099 17116 3111 17119
rect 3142 17116 3148 17128
rect 3099 17088 3148 17116
rect 3099 17085 3111 17088
rect 3053 17079 3111 17085
rect 3142 17076 3148 17088
rect 3200 17116 3206 17128
rect 3896 17125 3924 17224
rect 4982 17212 4988 17224
rect 5040 17212 5046 17264
rect 5534 17252 5540 17264
rect 5368 17224 5540 17252
rect 5368 17184 5396 17224
rect 5534 17212 5540 17224
rect 5592 17252 5598 17264
rect 5592 17224 10824 17252
rect 5592 17212 5598 17224
rect 5184 17156 5396 17184
rect 5813 17187 5871 17193
rect 3881 17119 3939 17125
rect 3881 17116 3893 17119
rect 3200 17088 3893 17116
rect 3200 17076 3206 17088
rect 3881 17085 3893 17088
rect 3927 17085 3939 17119
rect 3881 17079 3939 17085
rect 3970 17076 3976 17128
rect 4028 17116 4034 17128
rect 5184 17125 5212 17156
rect 5813 17153 5825 17187
rect 5859 17184 5871 17187
rect 5994 17184 6000 17196
rect 5859 17156 6000 17184
rect 5859 17153 5871 17156
rect 5813 17147 5871 17153
rect 5994 17144 6000 17156
rect 6052 17184 6058 17196
rect 6457 17187 6515 17193
rect 6457 17184 6469 17187
rect 6052 17156 6469 17184
rect 6052 17144 6058 17156
rect 6457 17153 6469 17156
rect 6503 17153 6515 17187
rect 6457 17147 6515 17153
rect 9493 17187 9551 17193
rect 9493 17153 9505 17187
rect 9539 17184 9551 17187
rect 9766 17184 9772 17196
rect 9539 17156 9772 17184
rect 9539 17153 9551 17156
rect 9493 17147 9551 17153
rect 9766 17144 9772 17156
rect 9824 17144 9830 17196
rect 10796 17128 10824 17224
rect 11517 17187 11575 17193
rect 11517 17153 11529 17187
rect 11563 17184 11575 17187
rect 11900 17184 11928 17283
rect 12158 17280 12164 17292
rect 12216 17280 12222 17332
rect 13078 17280 13084 17332
rect 13136 17320 13142 17332
rect 13357 17323 13415 17329
rect 13357 17320 13369 17323
rect 13136 17292 13369 17320
rect 13136 17280 13142 17292
rect 13357 17289 13369 17292
rect 13403 17320 13415 17323
rect 13722 17320 13728 17332
rect 13403 17292 13728 17320
rect 13403 17289 13415 17292
rect 13357 17283 13415 17289
rect 13722 17280 13728 17292
rect 13780 17280 13786 17332
rect 17402 17320 17408 17332
rect 17363 17292 17408 17320
rect 17402 17280 17408 17292
rect 17460 17280 17466 17332
rect 17494 17280 17500 17332
rect 17552 17320 17558 17332
rect 18506 17320 18512 17332
rect 17552 17292 18512 17320
rect 17552 17280 17558 17292
rect 18506 17280 18512 17292
rect 18564 17280 18570 17332
rect 18601 17323 18659 17329
rect 18601 17289 18613 17323
rect 18647 17320 18659 17323
rect 18874 17320 18880 17332
rect 18647 17292 18880 17320
rect 18647 17289 18659 17292
rect 18601 17283 18659 17289
rect 12434 17212 12440 17264
rect 12492 17252 12498 17264
rect 14185 17255 14243 17261
rect 12492 17224 13814 17252
rect 12492 17212 12498 17224
rect 13630 17184 13636 17196
rect 11563 17156 11928 17184
rect 13591 17156 13636 17184
rect 11563 17153 11575 17156
rect 11517 17147 11575 17153
rect 13630 17144 13636 17156
rect 13688 17144 13694 17196
rect 13786 17184 13814 17224
rect 14185 17221 14197 17255
rect 14231 17252 14243 17255
rect 14366 17252 14372 17264
rect 14231 17224 14372 17252
rect 14231 17221 14243 17224
rect 14185 17215 14243 17221
rect 14366 17212 14372 17224
rect 14424 17212 14430 17264
rect 15519 17255 15577 17261
rect 15519 17221 15531 17255
rect 15565 17252 15577 17255
rect 16758 17252 16764 17264
rect 15565 17224 16764 17252
rect 15565 17221 15577 17224
rect 15519 17215 15577 17221
rect 16758 17212 16764 17224
rect 16816 17212 16822 17264
rect 17034 17252 17040 17264
rect 16995 17224 17040 17252
rect 17034 17212 17040 17224
rect 17092 17212 17098 17264
rect 16485 17187 16543 17193
rect 13786 17156 15459 17184
rect 4065 17119 4123 17125
rect 4065 17116 4077 17119
rect 4028 17088 4077 17116
rect 4028 17076 4034 17088
rect 4065 17085 4077 17088
rect 4111 17116 4123 17119
rect 4985 17119 5043 17125
rect 4111 17088 4292 17116
rect 4111 17085 4123 17088
rect 4065 17079 4123 17085
rect 4264 17048 4292 17088
rect 4985 17085 4997 17119
rect 5031 17116 5043 17119
rect 5169 17119 5227 17125
rect 5169 17116 5181 17119
rect 5031 17088 5181 17116
rect 5031 17085 5043 17088
rect 4985 17079 5043 17085
rect 5169 17085 5181 17088
rect 5215 17085 5227 17119
rect 5169 17079 5227 17085
rect 5258 17076 5264 17128
rect 5316 17116 5322 17128
rect 5537 17119 5595 17125
rect 5537 17116 5549 17119
rect 5316 17088 5549 17116
rect 5316 17076 5322 17088
rect 5537 17085 5549 17088
rect 5583 17085 5595 17119
rect 5537 17079 5595 17085
rect 7101 17119 7159 17125
rect 7101 17085 7113 17119
rect 7147 17116 7159 17119
rect 7282 17116 7288 17128
rect 7147 17088 7288 17116
rect 7147 17085 7159 17088
rect 7101 17079 7159 17085
rect 7282 17076 7288 17088
rect 7340 17116 7346 17128
rect 7466 17116 7472 17128
rect 7340 17088 7472 17116
rect 7340 17076 7346 17088
rect 7466 17076 7472 17088
rect 7524 17076 7530 17128
rect 7650 17116 7656 17128
rect 7611 17088 7656 17116
rect 7650 17076 7656 17088
rect 7708 17076 7714 17128
rect 10778 17116 10784 17128
rect 10739 17088 10784 17116
rect 10778 17076 10784 17088
rect 10836 17076 10842 17128
rect 11146 17076 11152 17128
rect 11204 17116 11210 17128
rect 15431 17125 15459 17156
rect 16485 17153 16497 17187
rect 16531 17184 16543 17187
rect 17773 17187 17831 17193
rect 17773 17184 17785 17187
rect 16531 17156 17785 17184
rect 16531 17153 16543 17156
rect 16485 17147 16543 17153
rect 17773 17153 17785 17156
rect 17819 17184 17831 17187
rect 18187 17187 18245 17193
rect 18187 17184 18199 17187
rect 17819 17156 18199 17184
rect 17819 17153 17831 17156
rect 17773 17147 17831 17153
rect 18187 17153 18199 17156
rect 18233 17153 18245 17187
rect 18187 17147 18245 17153
rect 11241 17119 11299 17125
rect 11241 17116 11253 17119
rect 11204 17088 11253 17116
rect 11204 17076 11210 17088
rect 11241 17085 11253 17088
rect 11287 17085 11299 17119
rect 11241 17079 11299 17085
rect 12488 17119 12546 17125
rect 12488 17085 12500 17119
rect 12534 17116 12546 17119
rect 15416 17119 15474 17125
rect 12534 17088 13032 17116
rect 12534 17085 12546 17088
rect 12488 17079 12546 17085
rect 6454 17048 6460 17060
rect 4264 17020 6460 17048
rect 6454 17008 6460 17020
rect 6512 17008 6518 17060
rect 7926 17048 7932 17060
rect 7887 17020 7932 17048
rect 7926 17008 7932 17020
rect 7984 17008 7990 17060
rect 8846 17048 8852 17060
rect 8759 17020 8852 17048
rect 8846 17008 8852 17020
rect 8904 17008 8910 17060
rect 8938 17008 8944 17060
rect 8996 17048 9002 17060
rect 12575 17051 12633 17057
rect 12575 17048 12587 17051
rect 8996 17020 9041 17048
rect 9743 17020 12587 17048
rect 8996 17008 9002 17020
rect 3234 16980 3240 16992
rect 3195 16952 3240 16980
rect 3234 16940 3240 16952
rect 3292 16940 3298 16992
rect 3602 16980 3608 16992
rect 3563 16952 3608 16980
rect 3602 16940 3608 16952
rect 3660 16940 3666 16992
rect 3970 16940 3976 16992
rect 4028 16980 4034 16992
rect 4249 16983 4307 16989
rect 4249 16980 4261 16983
rect 4028 16952 4261 16980
rect 4028 16940 4034 16952
rect 4249 16949 4261 16952
rect 4295 16949 4307 16983
rect 4249 16943 4307 16949
rect 4522 16940 4528 16992
rect 4580 16980 4586 16992
rect 4617 16983 4675 16989
rect 4617 16980 4629 16983
rect 4580 16952 4629 16980
rect 4580 16940 4586 16952
rect 4617 16949 4629 16952
rect 4663 16980 4675 16983
rect 5166 16980 5172 16992
rect 4663 16952 5172 16980
rect 4663 16949 4675 16952
rect 4617 16943 4675 16949
rect 5166 16940 5172 16952
rect 5224 16940 5230 16992
rect 6086 16980 6092 16992
rect 6047 16952 6092 16980
rect 6086 16940 6092 16952
rect 6144 16940 6150 16992
rect 8294 16980 8300 16992
rect 8255 16952 8300 16980
rect 8294 16940 8300 16952
rect 8352 16940 8358 16992
rect 8864 16980 8892 17008
rect 9743 16980 9771 17020
rect 12575 17017 12587 17020
rect 12621 17017 12633 17051
rect 12575 17011 12633 17017
rect 9950 16980 9956 16992
rect 8864 16952 9771 16980
rect 9911 16952 9956 16980
rect 9950 16940 9956 16952
rect 10008 16980 10014 16992
rect 10229 16983 10287 16989
rect 10229 16980 10241 16983
rect 10008 16952 10241 16980
rect 10008 16940 10014 16952
rect 10229 16949 10241 16952
rect 10275 16949 10287 16983
rect 10229 16943 10287 16949
rect 11882 16940 11888 16992
rect 11940 16980 11946 16992
rect 13004 16989 13032 17088
rect 15416 17085 15428 17119
rect 15462 17116 15474 17119
rect 15841 17119 15899 17125
rect 15841 17116 15853 17119
rect 15462 17088 15853 17116
rect 15462 17085 15474 17088
rect 15416 17079 15474 17085
rect 15841 17085 15853 17088
rect 15887 17085 15899 17119
rect 15841 17079 15899 17085
rect 18100 17119 18158 17125
rect 18100 17085 18112 17119
rect 18146 17116 18158 17119
rect 18616 17116 18644 17283
rect 18874 17280 18880 17292
rect 18932 17280 18938 17332
rect 19981 17323 20039 17329
rect 19981 17289 19993 17323
rect 20027 17320 20039 17323
rect 21266 17320 21272 17332
rect 20027 17292 21272 17320
rect 20027 17289 20039 17292
rect 19981 17283 20039 17289
rect 21266 17280 21272 17292
rect 21324 17280 21330 17332
rect 23014 17320 23020 17332
rect 22975 17292 23020 17320
rect 23014 17280 23020 17292
rect 23072 17280 23078 17332
rect 25406 17320 25412 17332
rect 25367 17292 25412 17320
rect 25406 17280 25412 17292
rect 25464 17280 25470 17332
rect 20349 17255 20407 17261
rect 20349 17221 20361 17255
rect 20395 17252 20407 17255
rect 21634 17252 21640 17264
rect 20395 17224 21640 17252
rect 20395 17221 20407 17224
rect 20349 17215 20407 17221
rect 21634 17212 21640 17224
rect 21692 17212 21698 17264
rect 22695 17255 22753 17261
rect 22695 17221 22707 17255
rect 22741 17252 22753 17255
rect 24670 17252 24676 17264
rect 22741 17224 24676 17252
rect 22741 17221 22753 17224
rect 22695 17215 22753 17221
rect 24670 17212 24676 17224
rect 24728 17212 24734 17264
rect 19061 17187 19119 17193
rect 19061 17153 19073 17187
rect 19107 17184 19119 17187
rect 19426 17184 19432 17196
rect 19107 17156 19432 17184
rect 19107 17153 19119 17156
rect 19061 17147 19119 17153
rect 19426 17144 19432 17156
rect 19484 17144 19490 17196
rect 20254 17144 20260 17196
rect 20312 17184 20318 17196
rect 20625 17187 20683 17193
rect 20625 17184 20637 17187
rect 20312 17156 20637 17184
rect 20312 17144 20318 17156
rect 20625 17153 20637 17156
rect 20671 17153 20683 17187
rect 20625 17147 20683 17153
rect 20714 17144 20720 17196
rect 20772 17184 20778 17196
rect 20901 17187 20959 17193
rect 20901 17184 20913 17187
rect 20772 17156 20913 17184
rect 20772 17144 20778 17156
rect 20901 17153 20913 17156
rect 20947 17184 20959 17187
rect 21082 17184 21088 17196
rect 20947 17156 21088 17184
rect 20947 17153 20959 17156
rect 20901 17147 20959 17153
rect 21082 17144 21088 17156
rect 21140 17144 21146 17196
rect 21266 17144 21272 17196
rect 21324 17184 21330 17196
rect 21542 17184 21548 17196
rect 21324 17156 21548 17184
rect 21324 17144 21330 17156
rect 21542 17144 21548 17156
rect 21600 17144 21606 17196
rect 18146 17088 18644 17116
rect 22624 17119 22682 17125
rect 18146 17085 18158 17088
rect 18100 17079 18158 17085
rect 22624 17085 22636 17119
rect 22670 17116 22682 17119
rect 22738 17116 22744 17128
rect 22670 17088 22744 17116
rect 22670 17085 22682 17088
rect 22624 17079 22682 17085
rect 22738 17076 22744 17088
rect 22796 17076 22802 17128
rect 22922 17076 22928 17128
rect 22980 17116 22986 17128
rect 23477 17119 23535 17125
rect 23477 17116 23489 17119
rect 22980 17088 23489 17116
rect 22980 17076 22986 17088
rect 23477 17085 23489 17088
rect 23523 17116 23535 17119
rect 23661 17119 23719 17125
rect 23661 17116 23673 17119
rect 23523 17088 23673 17116
rect 23523 17085 23535 17088
rect 23477 17079 23535 17085
rect 23661 17085 23673 17088
rect 23707 17085 23719 17119
rect 24121 17119 24179 17125
rect 24121 17116 24133 17119
rect 23661 17079 23719 17085
rect 23860 17088 24133 17116
rect 23860 17060 23888 17088
rect 24121 17085 24133 17088
rect 24167 17085 24179 17119
rect 25222 17116 25228 17128
rect 25183 17088 25228 17116
rect 24121 17079 24179 17085
rect 25222 17076 25228 17088
rect 25280 17116 25286 17128
rect 25777 17119 25835 17125
rect 25777 17116 25789 17119
rect 25280 17088 25789 17116
rect 25280 17076 25286 17088
rect 25777 17085 25789 17088
rect 25823 17085 25835 17119
rect 25777 17079 25835 17085
rect 13722 17048 13728 17060
rect 13683 17020 13728 17048
rect 13722 17008 13728 17020
rect 13780 17008 13786 17060
rect 15654 17048 15660 17060
rect 14476 17020 15660 17048
rect 12161 16983 12219 16989
rect 12161 16980 12173 16983
rect 11940 16952 12173 16980
rect 11940 16940 11946 16952
rect 12161 16949 12173 16952
rect 12207 16949 12219 16983
rect 12161 16943 12219 16949
rect 12989 16983 13047 16989
rect 12989 16949 13001 16983
rect 13035 16980 13047 16983
rect 13078 16980 13084 16992
rect 13035 16952 13084 16980
rect 13035 16949 13047 16952
rect 12989 16943 13047 16949
rect 13078 16940 13084 16952
rect 13136 16980 13142 16992
rect 14476 16980 14504 17020
rect 15654 17008 15660 17020
rect 15712 17048 15718 17060
rect 16209 17051 16267 17057
rect 16209 17048 16221 17051
rect 15712 17020 16221 17048
rect 15712 17008 15718 17020
rect 16209 17017 16221 17020
rect 16255 17017 16267 17051
rect 16574 17048 16580 17060
rect 16535 17020 16580 17048
rect 16209 17011 16267 17017
rect 16574 17008 16580 17020
rect 16632 17008 16638 17060
rect 19382 17051 19440 17057
rect 19382 17048 19394 17051
rect 19306 17020 19394 17048
rect 13136 16952 14504 16980
rect 14645 16983 14703 16989
rect 13136 16940 13142 16952
rect 14645 16949 14657 16983
rect 14691 16980 14703 16983
rect 14734 16980 14740 16992
rect 14691 16952 14740 16980
rect 14691 16949 14703 16952
rect 14645 16943 14703 16949
rect 14734 16940 14740 16952
rect 14792 16940 14798 16992
rect 18874 16980 18880 16992
rect 18835 16952 18880 16980
rect 18874 16940 18880 16952
rect 18932 16980 18938 16992
rect 19150 16980 19156 16992
rect 18932 16952 19156 16980
rect 18932 16940 18938 16952
rect 19150 16940 19156 16952
rect 19208 16980 19214 16992
rect 19306 16980 19334 17020
rect 19382 17017 19394 17020
rect 19428 17017 19440 17051
rect 19382 17011 19440 17017
rect 20993 17051 21051 17057
rect 20993 17017 21005 17051
rect 21039 17017 21051 17051
rect 20993 17011 21051 17017
rect 21545 17051 21603 17057
rect 21545 17017 21557 17051
rect 21591 17048 21603 17051
rect 21634 17048 21640 17060
rect 21591 17020 21640 17048
rect 21591 17017 21603 17020
rect 21545 17011 21603 17017
rect 19208 16952 19334 16980
rect 19208 16940 19214 16952
rect 20806 16940 20812 16992
rect 20864 16980 20870 16992
rect 21008 16980 21036 17011
rect 21634 17008 21640 17020
rect 21692 17008 21698 17060
rect 22465 17051 22523 17057
rect 22465 17017 22477 17051
rect 22511 17048 22523 17051
rect 23842 17048 23848 17060
rect 22511 17020 23848 17048
rect 22511 17017 22523 17020
rect 22465 17011 22523 17017
rect 23842 17008 23848 17020
rect 23900 17008 23906 17060
rect 21821 16983 21879 16989
rect 21821 16980 21833 16983
rect 20864 16952 21833 16980
rect 20864 16940 20870 16952
rect 21821 16949 21833 16952
rect 21867 16949 21879 16983
rect 21821 16943 21879 16949
rect 23566 16940 23572 16992
rect 23624 16980 23630 16992
rect 23753 16983 23811 16989
rect 23753 16980 23765 16983
rect 23624 16952 23765 16980
rect 23624 16940 23630 16952
rect 23753 16949 23765 16952
rect 23799 16949 23811 16983
rect 23753 16943 23811 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1578 16776 1584 16788
rect 1539 16748 1584 16776
rect 1578 16736 1584 16748
rect 1636 16736 1642 16788
rect 2314 16776 2320 16788
rect 2275 16748 2320 16776
rect 2314 16736 2320 16748
rect 2372 16736 2378 16788
rect 3510 16736 3516 16788
rect 3568 16776 3574 16788
rect 4249 16779 4307 16785
rect 4249 16776 4261 16779
rect 3568 16748 4261 16776
rect 3568 16736 3574 16748
rect 4249 16745 4261 16748
rect 4295 16745 4307 16779
rect 5258 16776 5264 16788
rect 5219 16748 5264 16776
rect 4249 16739 4307 16745
rect 5258 16736 5264 16748
rect 5316 16736 5322 16788
rect 7558 16776 7564 16788
rect 7519 16748 7564 16776
rect 7558 16736 7564 16748
rect 7616 16736 7622 16788
rect 10778 16776 10784 16788
rect 10739 16748 10784 16776
rect 10778 16736 10784 16748
rect 10836 16736 10842 16788
rect 11882 16776 11888 16788
rect 11843 16748 11888 16776
rect 11882 16736 11888 16748
rect 11940 16736 11946 16788
rect 12437 16779 12495 16785
rect 12437 16745 12449 16779
rect 12483 16776 12495 16779
rect 12483 16748 13676 16776
rect 12483 16745 12495 16748
rect 12437 16739 12495 16745
rect 13648 16720 13676 16748
rect 13722 16736 13728 16788
rect 13780 16776 13786 16788
rect 15286 16776 15292 16788
rect 13780 16748 15292 16776
rect 13780 16736 13786 16748
rect 15286 16736 15292 16748
rect 15344 16736 15350 16788
rect 17037 16779 17095 16785
rect 17037 16745 17049 16779
rect 17083 16776 17095 16779
rect 17402 16776 17408 16788
rect 17083 16748 17408 16776
rect 17083 16745 17095 16748
rect 17037 16739 17095 16745
rect 17402 16736 17408 16748
rect 17460 16776 17466 16788
rect 17770 16776 17776 16788
rect 17460 16748 17776 16776
rect 17460 16736 17466 16748
rect 17770 16736 17776 16748
rect 17828 16776 17834 16788
rect 20714 16776 20720 16788
rect 17828 16748 18092 16776
rect 20675 16748 20720 16776
rect 17828 16736 17834 16748
rect 2590 16668 2596 16720
rect 2648 16708 2654 16720
rect 5537 16711 5595 16717
rect 5537 16708 5549 16711
rect 2648 16680 5549 16708
rect 2648 16668 2654 16680
rect 5537 16677 5549 16680
rect 5583 16708 5595 16711
rect 5813 16711 5871 16717
rect 5813 16708 5825 16711
rect 5583 16680 5825 16708
rect 5583 16677 5595 16680
rect 5537 16671 5595 16677
rect 5813 16677 5825 16680
rect 5859 16677 5871 16711
rect 5813 16671 5871 16677
rect 5905 16711 5963 16717
rect 5905 16677 5917 16711
rect 5951 16708 5963 16711
rect 6178 16708 6184 16720
rect 5951 16680 6184 16708
rect 5951 16677 5963 16680
rect 5905 16671 5963 16677
rect 6178 16668 6184 16680
rect 6236 16668 6242 16720
rect 7285 16711 7343 16717
rect 7285 16677 7297 16711
rect 7331 16708 7343 16711
rect 7650 16708 7656 16720
rect 7331 16680 7656 16708
rect 7331 16677 7343 16680
rect 7285 16671 7343 16677
rect 7650 16668 7656 16680
rect 7708 16708 7714 16720
rect 9858 16708 9864 16720
rect 7708 16680 8524 16708
rect 9819 16680 9864 16708
rect 7708 16668 7714 16680
rect 8496 16652 8524 16680
rect 9858 16668 9864 16680
rect 9916 16668 9922 16720
rect 11974 16668 11980 16720
rect 12032 16708 12038 16720
rect 12526 16708 12532 16720
rect 12032 16680 12532 16708
rect 12032 16668 12038 16680
rect 12526 16668 12532 16680
rect 12584 16708 12590 16720
rect 12713 16711 12771 16717
rect 12713 16708 12725 16711
rect 12584 16680 12725 16708
rect 12584 16668 12590 16680
rect 12713 16677 12725 16680
rect 12759 16677 12771 16711
rect 13354 16708 13360 16720
rect 13315 16680 13360 16708
rect 12713 16671 12771 16677
rect 13354 16668 13360 16680
rect 13412 16668 13418 16720
rect 13630 16708 13636 16720
rect 13543 16680 13636 16708
rect 13630 16668 13636 16680
rect 13688 16668 13694 16720
rect 15378 16668 15384 16720
rect 15436 16708 15442 16720
rect 16438 16711 16496 16717
rect 16438 16708 16450 16711
rect 15436 16680 16450 16708
rect 15436 16668 15442 16680
rect 16438 16677 16450 16680
rect 16484 16677 16496 16711
rect 16438 16671 16496 16677
rect 16758 16668 16764 16720
rect 16816 16708 16822 16720
rect 18064 16717 18092 16748
rect 20714 16736 20720 16748
rect 20772 16736 20778 16788
rect 22830 16776 22836 16788
rect 21008 16748 22836 16776
rect 17313 16711 17371 16717
rect 17313 16708 17325 16711
rect 16816 16680 17325 16708
rect 16816 16668 16822 16680
rect 17313 16677 17325 16680
rect 17359 16677 17371 16711
rect 17313 16671 17371 16677
rect 18049 16711 18107 16717
rect 18049 16677 18061 16711
rect 18095 16677 18107 16711
rect 18049 16671 18107 16677
rect 19242 16668 19248 16720
rect 19300 16708 19306 16720
rect 19567 16711 19625 16717
rect 19567 16708 19579 16711
rect 19300 16680 19579 16708
rect 19300 16668 19306 16680
rect 19567 16677 19579 16680
rect 19613 16677 19625 16711
rect 21008 16708 21036 16748
rect 22830 16736 22836 16748
rect 22888 16736 22894 16788
rect 24762 16776 24768 16788
rect 24320 16748 24768 16776
rect 19567 16671 19625 16677
rect 19996 16680 21036 16708
rect 21085 16711 21143 16717
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 3028 16643 3086 16649
rect 3028 16609 3040 16643
rect 3074 16640 3086 16643
rect 4709 16643 4767 16649
rect 3074 16612 3740 16640
rect 3074 16609 3086 16612
rect 3028 16603 3086 16609
rect 3712 16584 3740 16612
rect 4709 16609 4721 16643
rect 4755 16640 4767 16643
rect 4798 16640 4804 16652
rect 4755 16612 4804 16640
rect 4755 16609 4767 16612
rect 4709 16603 4767 16609
rect 4798 16600 4804 16612
rect 4856 16600 4862 16652
rect 7834 16600 7840 16652
rect 7892 16640 7898 16652
rect 8021 16643 8079 16649
rect 8021 16640 8033 16643
rect 7892 16612 8033 16640
rect 7892 16600 7898 16612
rect 8021 16609 8033 16612
rect 8067 16609 8079 16643
rect 8478 16640 8484 16652
rect 8439 16612 8484 16640
rect 8021 16603 8079 16609
rect 8478 16600 8484 16612
rect 8536 16600 8542 16652
rect 3694 16532 3700 16584
rect 3752 16572 3758 16584
rect 3878 16572 3884 16584
rect 3752 16544 3884 16572
rect 3752 16532 3758 16544
rect 3878 16532 3884 16544
rect 3936 16532 3942 16584
rect 6457 16575 6515 16581
rect 6457 16541 6469 16575
rect 6503 16572 6515 16575
rect 7374 16572 7380 16584
rect 6503 16544 7380 16572
rect 6503 16541 6515 16544
rect 6457 16535 6515 16541
rect 7374 16532 7380 16544
rect 7432 16532 7438 16584
rect 8754 16572 8760 16584
rect 8715 16544 8760 16572
rect 8754 16532 8760 16544
rect 8812 16532 8818 16584
rect 9493 16575 9551 16581
rect 9493 16541 9505 16575
rect 9539 16572 9551 16575
rect 9769 16575 9827 16581
rect 9769 16572 9781 16575
rect 9539 16544 9781 16572
rect 9539 16541 9551 16544
rect 9493 16535 9551 16541
rect 9769 16541 9781 16544
rect 9815 16572 9827 16575
rect 11514 16572 11520 16584
rect 9815 16544 10732 16572
rect 11475 16544 11520 16572
rect 9815 16541 9827 16544
rect 9769 16535 9827 16541
rect 3099 16507 3157 16513
rect 3099 16473 3111 16507
rect 3145 16504 3157 16507
rect 4614 16504 4620 16516
rect 3145 16476 4620 16504
rect 3145 16473 3157 16476
rect 3099 16467 3157 16473
rect 4614 16464 4620 16476
rect 4672 16464 4678 16516
rect 4893 16507 4951 16513
rect 4893 16473 4905 16507
rect 4939 16504 4951 16507
rect 9950 16504 9956 16516
rect 4939 16476 9956 16504
rect 4939 16473 4951 16476
rect 4893 16467 4951 16473
rect 9950 16464 9956 16476
rect 10008 16464 10014 16516
rect 10134 16464 10140 16516
rect 10192 16504 10198 16516
rect 10321 16507 10379 16513
rect 10321 16504 10333 16507
rect 10192 16476 10333 16504
rect 10192 16464 10198 16476
rect 10321 16473 10333 16476
rect 10367 16473 10379 16507
rect 10704 16504 10732 16544
rect 11514 16532 11520 16544
rect 11572 16532 11578 16584
rect 13372 16572 13400 16668
rect 19996 16652 20024 16680
rect 21085 16677 21097 16711
rect 21131 16708 21143 16711
rect 21358 16708 21364 16720
rect 21131 16680 21364 16708
rect 21131 16677 21143 16680
rect 21085 16671 21143 16677
rect 21358 16668 21364 16680
rect 21416 16668 21422 16720
rect 21634 16708 21640 16720
rect 21595 16680 21640 16708
rect 21634 16668 21640 16680
rect 21692 16668 21698 16720
rect 23658 16668 23664 16720
rect 23716 16708 23722 16720
rect 24320 16717 24348 16748
rect 24762 16736 24768 16748
rect 24820 16736 24826 16788
rect 24305 16711 24363 16717
rect 24305 16708 24317 16711
rect 23716 16680 24317 16708
rect 23716 16668 23722 16680
rect 24305 16677 24317 16680
rect 24351 16677 24363 16711
rect 24305 16671 24363 16677
rect 24397 16711 24455 16717
rect 24397 16677 24409 16711
rect 24443 16708 24455 16711
rect 24670 16708 24676 16720
rect 24443 16680 24676 16708
rect 24443 16677 24455 16680
rect 24397 16671 24455 16677
rect 24670 16668 24676 16680
rect 24728 16668 24734 16720
rect 19480 16643 19538 16649
rect 19480 16609 19492 16643
rect 19526 16640 19538 16643
rect 19978 16640 19984 16652
rect 19526 16612 19984 16640
rect 19526 16609 19538 16612
rect 19480 16603 19538 16609
rect 19978 16600 19984 16612
rect 20036 16600 20042 16652
rect 22830 16640 22836 16652
rect 22791 16612 22836 16640
rect 22830 16600 22836 16612
rect 22888 16600 22894 16652
rect 23106 16640 23112 16652
rect 23067 16612 23112 16640
rect 23106 16600 23112 16612
rect 23164 16600 23170 16652
rect 13541 16575 13599 16581
rect 13541 16572 13553 16575
rect 13372 16544 13553 16572
rect 13541 16541 13553 16544
rect 13587 16541 13599 16575
rect 13541 16535 13599 16541
rect 13817 16575 13875 16581
rect 13817 16541 13829 16575
rect 13863 16541 13875 16575
rect 16114 16572 16120 16584
rect 16075 16544 16120 16572
rect 13817 16535 13875 16541
rect 13170 16504 13176 16516
rect 10704 16476 13176 16504
rect 10321 16467 10379 16473
rect 13170 16464 13176 16476
rect 13228 16464 13234 16516
rect 1578 16396 1584 16448
rect 1636 16436 1642 16448
rect 1949 16439 2007 16445
rect 1949 16436 1961 16439
rect 1636 16408 1961 16436
rect 1636 16396 1642 16408
rect 1949 16405 1961 16408
rect 1995 16405 2007 16439
rect 1949 16399 2007 16405
rect 3697 16439 3755 16445
rect 3697 16405 3709 16439
rect 3743 16436 3755 16439
rect 4062 16436 4068 16448
rect 3743 16408 4068 16436
rect 3743 16405 3755 16408
rect 3697 16399 3755 16405
rect 4062 16396 4068 16408
rect 4120 16396 4126 16448
rect 4982 16396 4988 16448
rect 5040 16436 5046 16448
rect 10778 16436 10784 16448
rect 5040 16408 10784 16436
rect 5040 16396 5046 16408
rect 10778 16396 10784 16408
rect 10836 16396 10842 16448
rect 13538 16396 13544 16448
rect 13596 16436 13602 16448
rect 13832 16436 13860 16535
rect 16114 16532 16120 16544
rect 16172 16532 16178 16584
rect 17678 16532 17684 16584
rect 17736 16572 17742 16584
rect 17957 16575 18015 16581
rect 17957 16572 17969 16575
rect 17736 16544 17969 16572
rect 17736 16532 17742 16544
rect 17957 16541 17969 16544
rect 18003 16541 18015 16575
rect 18414 16572 18420 16584
rect 18375 16544 18420 16572
rect 17957 16535 18015 16541
rect 18414 16532 18420 16544
rect 18472 16532 18478 16584
rect 20993 16575 21051 16581
rect 20993 16541 21005 16575
rect 21039 16572 21051 16575
rect 22278 16572 22284 16584
rect 21039 16544 22284 16572
rect 21039 16541 21051 16544
rect 20993 16535 21051 16541
rect 22278 16532 22284 16544
rect 22336 16532 22342 16584
rect 23382 16572 23388 16584
rect 23343 16544 23388 16572
rect 23382 16532 23388 16544
rect 23440 16532 23446 16584
rect 24946 16572 24952 16584
rect 24859 16544 24952 16572
rect 24946 16532 24952 16544
rect 25004 16572 25010 16584
rect 25222 16572 25228 16584
rect 25004 16544 25228 16572
rect 25004 16532 25010 16544
rect 25222 16532 25228 16544
rect 25280 16532 25286 16584
rect 17402 16464 17408 16516
rect 17460 16504 17466 16516
rect 18966 16504 18972 16516
rect 17460 16476 18972 16504
rect 17460 16464 17466 16476
rect 18966 16464 18972 16476
rect 19024 16464 19030 16516
rect 19426 16464 19432 16516
rect 19484 16504 19490 16516
rect 19889 16507 19947 16513
rect 19889 16504 19901 16507
rect 19484 16476 19901 16504
rect 19484 16464 19490 16476
rect 19889 16473 19901 16476
rect 19935 16473 19947 16507
rect 19889 16467 19947 16473
rect 13596 16408 13860 16436
rect 13596 16396 13602 16408
rect 14642 16396 14648 16448
rect 14700 16436 14706 16448
rect 18322 16436 18328 16448
rect 14700 16408 18328 16436
rect 14700 16396 14706 16408
rect 18322 16396 18328 16408
rect 18380 16396 18386 16448
rect 18874 16396 18880 16448
rect 18932 16436 18938 16448
rect 19061 16439 19119 16445
rect 19061 16436 19073 16439
rect 18932 16408 19073 16436
rect 18932 16396 18938 16408
rect 19061 16405 19073 16408
rect 19107 16405 19119 16439
rect 23658 16436 23664 16448
rect 23619 16408 23664 16436
rect 19061 16399 19119 16405
rect 23658 16396 23664 16408
rect 23716 16436 23722 16448
rect 23842 16436 23848 16448
rect 23716 16408 23848 16436
rect 23716 16396 23722 16408
rect 23842 16396 23848 16408
rect 23900 16396 23906 16448
rect 24026 16436 24032 16448
rect 23987 16408 24032 16436
rect 24026 16396 24032 16408
rect 24084 16396 24090 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 1394 16192 1400 16244
rect 1452 16232 1458 16244
rect 2409 16235 2467 16241
rect 2409 16232 2421 16235
rect 1452 16204 2421 16232
rect 1452 16192 1458 16204
rect 2409 16201 2421 16204
rect 2455 16232 2467 16235
rect 4154 16232 4160 16244
rect 2455 16204 4160 16232
rect 2455 16201 2467 16204
rect 2409 16195 2467 16201
rect 4154 16192 4160 16204
rect 4212 16192 4218 16244
rect 6178 16232 6184 16244
rect 6139 16204 6184 16232
rect 6178 16192 6184 16204
rect 6236 16192 6242 16244
rect 9950 16232 9956 16244
rect 9911 16204 9956 16232
rect 9950 16192 9956 16204
rect 10008 16192 10014 16244
rect 13078 16192 13084 16244
rect 13136 16232 13142 16244
rect 13538 16232 13544 16244
rect 13136 16204 13544 16232
rect 13136 16192 13142 16204
rect 13538 16192 13544 16204
rect 13596 16192 13602 16244
rect 13630 16192 13636 16244
rect 13688 16232 13694 16244
rect 15013 16235 15071 16241
rect 15013 16232 15025 16235
rect 13688 16204 15025 16232
rect 13688 16192 13694 16204
rect 15013 16201 15025 16204
rect 15059 16201 15071 16235
rect 15013 16195 15071 16201
rect 16574 16192 16580 16244
rect 16632 16232 16638 16244
rect 16945 16235 17003 16241
rect 16945 16232 16957 16235
rect 16632 16204 16957 16232
rect 16632 16192 16638 16204
rect 16945 16201 16957 16204
rect 16991 16201 17003 16235
rect 17770 16232 17776 16244
rect 17731 16204 17776 16232
rect 16945 16195 17003 16201
rect 17770 16192 17776 16204
rect 17828 16192 17834 16244
rect 22278 16232 22284 16244
rect 22239 16204 22284 16232
rect 22278 16192 22284 16204
rect 22336 16192 22342 16244
rect 22741 16235 22799 16241
rect 22741 16201 22753 16235
rect 22787 16232 22799 16235
rect 23106 16232 23112 16244
rect 22787 16204 23112 16232
rect 22787 16201 22799 16204
rect 22741 16195 22799 16201
rect 23106 16192 23112 16204
rect 23164 16192 23170 16244
rect 24581 16235 24639 16241
rect 24581 16201 24593 16235
rect 24627 16232 24639 16235
rect 24670 16232 24676 16244
rect 24627 16204 24676 16232
rect 24627 16201 24639 16204
rect 24581 16195 24639 16201
rect 24670 16192 24676 16204
rect 24728 16232 24734 16244
rect 25225 16235 25283 16241
rect 25225 16232 25237 16235
rect 24728 16204 25237 16232
rect 24728 16192 24734 16204
rect 25225 16201 25237 16204
rect 25271 16201 25283 16235
rect 25590 16232 25596 16244
rect 25551 16204 25596 16232
rect 25225 16195 25283 16201
rect 25590 16192 25596 16204
rect 25648 16192 25654 16244
rect 1670 16124 1676 16176
rect 1728 16164 1734 16176
rect 2866 16164 2872 16176
rect 1728 16136 2872 16164
rect 1728 16124 1734 16136
rect 2866 16124 2872 16136
rect 2924 16124 2930 16176
rect 3881 16167 3939 16173
rect 3881 16133 3893 16167
rect 3927 16164 3939 16167
rect 4062 16164 4068 16176
rect 3927 16136 4068 16164
rect 3927 16133 3939 16136
rect 3881 16127 3939 16133
rect 4062 16124 4068 16136
rect 4120 16124 4126 16176
rect 3752 16099 3810 16105
rect 3752 16065 3764 16099
rect 3798 16065 3810 16099
rect 3752 16059 3810 16065
rect 3973 16099 4031 16105
rect 3973 16065 3985 16099
rect 4019 16096 4031 16099
rect 4154 16096 4160 16108
rect 4019 16068 4160 16096
rect 4019 16065 4031 16068
rect 3973 16059 4031 16065
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 2038 16028 2044 16040
rect 1443 16000 2044 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 2038 15988 2044 16000
rect 2096 15988 2102 16040
rect 2644 16031 2702 16037
rect 2644 15997 2656 16031
rect 2690 16028 2702 16031
rect 2690 15997 2703 16028
rect 2644 15991 2703 15997
rect 106 15852 112 15904
rect 164 15892 170 15904
rect 1581 15895 1639 15901
rect 1581 15892 1593 15895
rect 164 15864 1593 15892
rect 164 15852 170 15864
rect 1581 15861 1593 15864
rect 1627 15861 1639 15895
rect 2038 15892 2044 15904
rect 1999 15864 2044 15892
rect 1581 15855 1639 15861
rect 2038 15852 2044 15864
rect 2096 15852 2102 15904
rect 2675 15892 2703 15991
rect 3510 15988 3516 16040
rect 3568 16028 3574 16040
rect 3605 16031 3663 16037
rect 3605 16028 3617 16031
rect 3568 16000 3617 16028
rect 3568 15988 3574 16000
rect 3605 15997 3617 16000
rect 3651 15997 3663 16031
rect 3605 15991 3663 15997
rect 3758 15972 3786 16059
rect 4154 16056 4160 16068
rect 4212 16056 4218 16108
rect 5166 16056 5172 16108
rect 5224 16096 5230 16108
rect 9968 16096 9996 16192
rect 11882 16124 11888 16176
rect 11940 16164 11946 16176
rect 15378 16164 15384 16176
rect 11940 16136 15384 16164
rect 11940 16124 11946 16136
rect 15378 16124 15384 16136
rect 15436 16164 15442 16176
rect 15473 16167 15531 16173
rect 15473 16164 15485 16167
rect 15436 16136 15485 16164
rect 15436 16124 15442 16136
rect 15473 16133 15485 16136
rect 15519 16164 15531 16167
rect 15841 16167 15899 16173
rect 15841 16164 15853 16167
rect 15519 16136 15853 16164
rect 15519 16133 15531 16136
rect 15473 16127 15531 16133
rect 11146 16096 11152 16108
rect 5224 16068 9628 16096
rect 9968 16068 11152 16096
rect 5224 16056 5230 16068
rect 9600 16040 9628 16068
rect 4617 16031 4675 16037
rect 4617 16028 4629 16031
rect 2731 15963 2789 15969
rect 2731 15929 2743 15963
rect 2777 15960 2789 15963
rect 3326 15960 3332 15972
rect 2777 15932 3332 15960
rect 2777 15929 2789 15932
rect 2731 15923 2789 15929
rect 3326 15920 3332 15932
rect 3384 15920 3390 15972
rect 3694 15920 3700 15972
rect 3752 15960 3786 15972
rect 4080 16000 4629 16028
rect 4080 15960 4108 16000
rect 4617 15997 4629 16000
rect 4663 15997 4675 16031
rect 4617 15991 4675 15997
rect 5077 16031 5135 16037
rect 5077 15997 5089 16031
rect 5123 16028 5135 16031
rect 5350 16028 5356 16040
rect 5123 16000 5356 16028
rect 5123 15997 5135 16000
rect 5077 15991 5135 15997
rect 5350 15988 5356 16000
rect 5408 15988 5414 16040
rect 5721 16031 5779 16037
rect 5721 15997 5733 16031
rect 5767 16028 5779 16031
rect 6362 16028 6368 16040
rect 5767 16000 6368 16028
rect 5767 15997 5779 16000
rect 5721 15991 5779 15997
rect 6362 15988 6368 16000
rect 6420 15988 6426 16040
rect 7193 16031 7251 16037
rect 7193 15997 7205 16031
rect 7239 15997 7251 16031
rect 7193 15991 7251 15997
rect 7377 16031 7435 16037
rect 7377 15997 7389 16031
rect 7423 16028 7435 16031
rect 7653 16031 7711 16037
rect 7423 16000 7604 16028
rect 7423 15997 7435 16000
rect 7377 15991 7435 15997
rect 3752 15932 4108 15960
rect 4341 15963 4399 15969
rect 3752 15920 3758 15932
rect 4341 15929 4353 15963
rect 4387 15960 4399 15963
rect 6270 15960 6276 15972
rect 4387 15932 6276 15960
rect 4387 15929 4399 15932
rect 4341 15923 4399 15929
rect 6270 15920 6276 15932
rect 6328 15920 6334 15972
rect 6641 15963 6699 15969
rect 6641 15929 6653 15963
rect 6687 15960 6699 15963
rect 7208 15960 7236 15991
rect 7576 15972 7604 16000
rect 7653 15997 7665 16031
rect 7699 16028 7711 16031
rect 8481 16031 8539 16037
rect 8481 16028 8493 16031
rect 7699 16000 8493 16028
rect 7699 15997 7711 16000
rect 7653 15991 7711 15997
rect 8481 15997 8493 16000
rect 8527 16028 8539 16031
rect 8662 16028 8668 16040
rect 8527 16000 8668 16028
rect 8527 15997 8539 16000
rect 8481 15991 8539 15997
rect 8662 15988 8668 16000
rect 8720 15988 8726 16040
rect 9582 15988 9588 16040
rect 9640 16028 9646 16040
rect 10980 16037 11008 16068
rect 11146 16056 11152 16068
rect 11204 16056 11210 16108
rect 11241 16099 11299 16105
rect 11241 16065 11253 16099
rect 11287 16096 11299 16099
rect 11514 16096 11520 16108
rect 11287 16068 11520 16096
rect 11287 16065 11299 16068
rect 11241 16059 11299 16065
rect 11514 16056 11520 16068
rect 11572 16056 11578 16108
rect 12526 16096 12532 16108
rect 12487 16068 12532 16096
rect 12526 16056 12532 16068
rect 12584 16056 12590 16108
rect 10321 16031 10379 16037
rect 10321 16028 10333 16031
rect 9640 16000 10333 16028
rect 9640 15988 9646 16000
rect 10321 15997 10333 16000
rect 10367 16028 10379 16031
rect 10505 16031 10563 16037
rect 10505 16028 10517 16031
rect 10367 16000 10517 16028
rect 10367 15997 10379 16000
rect 10321 15991 10379 15997
rect 10505 15997 10517 16000
rect 10551 15997 10563 16031
rect 10505 15991 10563 15997
rect 10965 16031 11023 16037
rect 10965 15997 10977 16031
rect 11011 15997 11023 16031
rect 10965 15991 11023 15997
rect 13909 16031 13967 16037
rect 13909 15997 13921 16031
rect 13955 16028 13967 16031
rect 14182 16028 14188 16040
rect 13955 16000 14188 16028
rect 13955 15997 13967 16000
rect 13909 15991 13967 15997
rect 14182 15988 14188 16000
rect 14240 15988 14246 16040
rect 14461 16031 14519 16037
rect 14461 16028 14473 16031
rect 14384 16000 14473 16028
rect 7466 15960 7472 15972
rect 6687 15932 7472 15960
rect 6687 15929 6699 15932
rect 6641 15923 6699 15929
rect 7466 15920 7472 15932
rect 7524 15920 7530 15972
rect 7558 15920 7564 15972
rect 7616 15960 7622 15972
rect 8386 15960 8392 15972
rect 7616 15932 8392 15960
rect 7616 15920 7622 15932
rect 8386 15920 8392 15932
rect 8444 15920 8450 15972
rect 8802 15963 8860 15969
rect 8802 15929 8814 15963
rect 8848 15960 8860 15963
rect 10042 15960 10048 15972
rect 8848 15932 10048 15960
rect 8848 15929 8860 15932
rect 8802 15923 8860 15929
rect 2958 15892 2964 15904
rect 2675 15864 2964 15892
rect 2958 15852 2964 15864
rect 3016 15892 3022 15904
rect 3053 15895 3111 15901
rect 3053 15892 3065 15895
rect 3016 15864 3065 15892
rect 3016 15852 3022 15864
rect 3053 15861 3065 15864
rect 3099 15861 3111 15895
rect 3053 15855 3111 15861
rect 3513 15895 3571 15901
rect 3513 15861 3525 15895
rect 3559 15892 3571 15895
rect 3878 15892 3884 15904
rect 3559 15864 3884 15892
rect 3559 15861 3571 15864
rect 3513 15855 3571 15861
rect 3878 15852 3884 15864
rect 3936 15852 3942 15904
rect 5258 15892 5264 15904
rect 5219 15864 5264 15892
rect 5258 15852 5264 15864
rect 5316 15852 5322 15904
rect 7834 15852 7840 15904
rect 7892 15892 7898 15904
rect 7929 15895 7987 15901
rect 7929 15892 7941 15895
rect 7892 15864 7941 15892
rect 7892 15852 7898 15864
rect 7929 15861 7941 15864
rect 7975 15861 7987 15895
rect 8294 15892 8300 15904
rect 8255 15864 8300 15892
rect 7929 15855 7987 15861
rect 8294 15852 8300 15864
rect 8352 15892 8358 15904
rect 8817 15892 8845 15923
rect 10042 15920 10048 15932
rect 10100 15920 10106 15972
rect 12621 15963 12679 15969
rect 12621 15929 12633 15963
rect 12667 15929 12679 15963
rect 13170 15960 13176 15972
rect 13131 15932 13176 15960
rect 12621 15923 12679 15929
rect 8352 15864 8845 15892
rect 9401 15895 9459 15901
rect 8352 15852 8358 15864
rect 9401 15861 9413 15895
rect 9447 15892 9459 15895
rect 9766 15892 9772 15904
rect 9447 15864 9772 15892
rect 9447 15861 9459 15864
rect 9401 15855 9459 15861
rect 9766 15852 9772 15864
rect 9824 15852 9830 15904
rect 11609 15895 11667 15901
rect 11609 15861 11621 15895
rect 11655 15892 11667 15895
rect 11882 15892 11888 15904
rect 11655 15864 11888 15892
rect 11655 15861 11667 15864
rect 11609 15855 11667 15861
rect 11882 15852 11888 15864
rect 11940 15852 11946 15904
rect 12250 15892 12256 15904
rect 12163 15864 12256 15892
rect 12250 15852 12256 15864
rect 12308 15892 12314 15904
rect 12636 15892 12664 15923
rect 13170 15920 13176 15932
rect 13228 15920 13234 15972
rect 13541 15963 13599 15969
rect 13541 15929 13553 15963
rect 13587 15960 13599 15963
rect 14384 15960 14412 16000
rect 14461 15997 14473 16000
rect 14507 15997 14519 16031
rect 14461 15991 14519 15997
rect 13587 15932 14412 15960
rect 15672 15960 15700 16136
rect 15841 16133 15853 16136
rect 15887 16133 15899 16167
rect 15841 16127 15899 16133
rect 24762 16124 24768 16176
rect 24820 16164 24826 16176
rect 24857 16167 24915 16173
rect 24857 16164 24869 16167
rect 24820 16136 24869 16164
rect 24820 16124 24826 16136
rect 24857 16133 24869 16136
rect 24903 16133 24915 16167
rect 24857 16127 24915 16133
rect 15746 16056 15752 16108
rect 15804 16096 15810 16108
rect 16025 16099 16083 16105
rect 16025 16096 16037 16099
rect 15804 16068 16037 16096
rect 15804 16056 15810 16068
rect 16025 16065 16037 16068
rect 16071 16096 16083 16099
rect 17221 16099 17279 16105
rect 17221 16096 17233 16099
rect 16071 16068 17233 16096
rect 16071 16065 16083 16068
rect 16025 16059 16083 16065
rect 17221 16065 17233 16068
rect 17267 16065 17279 16099
rect 17221 16059 17279 16065
rect 19334 16056 19340 16108
rect 19392 16096 19398 16108
rect 19429 16099 19487 16105
rect 19429 16096 19441 16099
rect 19392 16068 19441 16096
rect 19392 16056 19398 16068
rect 19429 16065 19441 16068
rect 19475 16065 19487 16099
rect 19429 16059 19487 16065
rect 20898 16056 20904 16108
rect 20956 16096 20962 16108
rect 21269 16099 21327 16105
rect 21269 16096 21281 16099
rect 20956 16068 21281 16096
rect 20956 16056 20962 16068
rect 21269 16065 21281 16068
rect 21315 16096 21327 16099
rect 21542 16096 21548 16108
rect 21315 16068 21548 16096
rect 21315 16065 21327 16068
rect 21269 16059 21327 16065
rect 21542 16056 21548 16068
rect 21600 16056 21606 16108
rect 23661 16099 23719 16105
rect 23661 16096 23673 16099
rect 23446 16068 23673 16096
rect 18049 16031 18107 16037
rect 18049 15997 18061 16031
rect 18095 16028 18107 16031
rect 18509 16031 18567 16037
rect 18509 16028 18521 16031
rect 18095 16000 18521 16028
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 18509 15997 18521 16000
rect 18555 16028 18567 16031
rect 19058 16028 19064 16040
rect 18555 16000 19064 16028
rect 18555 15997 18567 16000
rect 18509 15991 18567 15997
rect 19058 15988 19064 16000
rect 19116 15988 19122 16040
rect 23290 15988 23296 16040
rect 23348 16028 23354 16040
rect 23446 16028 23474 16068
rect 23661 16065 23673 16068
rect 23707 16096 23719 16099
rect 24026 16096 24032 16108
rect 23707 16068 24032 16096
rect 23707 16065 23719 16068
rect 23661 16059 23719 16065
rect 24026 16056 24032 16068
rect 24084 16056 24090 16108
rect 23348 16000 23474 16028
rect 23348 15988 23354 16000
rect 23934 15988 23940 16040
rect 23992 16028 23998 16040
rect 25409 16031 25467 16037
rect 25409 16028 25421 16031
rect 23992 16000 25421 16028
rect 23992 15988 23998 16000
rect 25409 15997 25421 16000
rect 25455 16028 25467 16031
rect 25961 16031 26019 16037
rect 25961 16028 25973 16031
rect 25455 16000 25973 16028
rect 25455 15997 25467 16000
rect 25409 15991 25467 15997
rect 25961 15997 25973 16000
rect 26007 15997 26019 16031
rect 25961 15991 26019 15997
rect 16346 15963 16404 15969
rect 16346 15960 16358 15963
rect 15672 15932 16358 15960
rect 13587 15929 13599 15932
rect 13541 15923 13599 15929
rect 16346 15929 16358 15932
rect 16392 15929 16404 15963
rect 19750 15963 19808 15969
rect 19750 15960 19762 15963
rect 16346 15923 16404 15929
rect 18892 15932 19762 15960
rect 12308 15864 12664 15892
rect 12308 15852 12314 15864
rect 12894 15852 12900 15904
rect 12952 15892 12958 15904
rect 13556 15892 13584 15923
rect 18892 15904 18920 15932
rect 19750 15929 19762 15932
rect 19796 15929 19808 15963
rect 19750 15923 19808 15929
rect 21358 15920 21364 15972
rect 21416 15960 21422 15972
rect 21910 15960 21916 15972
rect 21416 15932 21461 15960
rect 21871 15932 21916 15960
rect 21416 15920 21422 15932
rect 21910 15920 21916 15932
rect 21968 15920 21974 15972
rect 24026 15969 24032 15972
rect 24023 15960 24032 15969
rect 23400 15932 24032 15960
rect 14090 15892 14096 15904
rect 12952 15864 13584 15892
rect 14051 15864 14096 15892
rect 12952 15852 12958 15864
rect 14090 15852 14096 15864
rect 14148 15852 14154 15904
rect 16022 15852 16028 15904
rect 16080 15892 16086 15904
rect 17218 15892 17224 15904
rect 16080 15864 17224 15892
rect 16080 15852 16086 15864
rect 17218 15852 17224 15864
rect 17276 15852 17282 15904
rect 17862 15852 17868 15904
rect 17920 15892 17926 15904
rect 18233 15895 18291 15901
rect 18233 15892 18245 15895
rect 17920 15864 18245 15892
rect 17920 15852 17926 15864
rect 18233 15861 18245 15864
rect 18279 15861 18291 15895
rect 18874 15892 18880 15904
rect 18835 15864 18880 15892
rect 18233 15855 18291 15861
rect 18874 15852 18880 15864
rect 18932 15852 18938 15904
rect 19337 15895 19395 15901
rect 19337 15861 19349 15895
rect 19383 15892 19395 15895
rect 19978 15892 19984 15904
rect 19383 15864 19984 15892
rect 19383 15861 19395 15864
rect 19337 15855 19395 15861
rect 19978 15852 19984 15864
rect 20036 15852 20042 15904
rect 20349 15895 20407 15901
rect 20349 15861 20361 15895
rect 20395 15892 20407 15895
rect 20993 15895 21051 15901
rect 20993 15892 21005 15895
rect 20395 15864 21005 15892
rect 20395 15861 20407 15864
rect 20349 15855 20407 15861
rect 20993 15861 21005 15864
rect 21039 15892 21051 15895
rect 21376 15892 21404 15920
rect 21039 15864 21404 15892
rect 21039 15861 21051 15864
rect 20993 15855 21051 15861
rect 22830 15852 22836 15904
rect 22888 15892 22894 15904
rect 23017 15895 23075 15901
rect 23017 15892 23029 15895
rect 22888 15864 23029 15892
rect 22888 15852 22894 15864
rect 23017 15861 23029 15864
rect 23063 15861 23075 15895
rect 23017 15855 23075 15861
rect 23198 15852 23204 15904
rect 23256 15892 23262 15904
rect 23400 15901 23428 15932
rect 24023 15923 24032 15932
rect 24026 15920 24032 15923
rect 24084 15920 24090 15972
rect 23385 15895 23443 15901
rect 23385 15892 23397 15895
rect 23256 15864 23397 15892
rect 23256 15852 23262 15864
rect 23385 15861 23397 15864
rect 23431 15861 23443 15895
rect 23385 15855 23443 15861
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 2958 15648 2964 15700
rect 3016 15688 3022 15700
rect 3016 15660 3188 15688
rect 3016 15648 3022 15660
rect 1946 15552 1952 15564
rect 1907 15524 1952 15552
rect 1946 15512 1952 15524
rect 2004 15512 2010 15564
rect 2958 15552 2964 15564
rect 2919 15524 2964 15552
rect 2958 15512 2964 15524
rect 3016 15512 3022 15564
rect 3160 15552 3188 15660
rect 3234 15648 3240 15700
rect 3292 15688 3298 15700
rect 5261 15691 5319 15697
rect 5261 15688 5273 15691
rect 3292 15660 5273 15688
rect 3292 15648 3298 15660
rect 5261 15657 5273 15660
rect 5307 15688 5319 15691
rect 5442 15688 5448 15700
rect 5307 15660 5448 15688
rect 5307 15657 5319 15660
rect 5261 15651 5319 15657
rect 5442 15648 5448 15660
rect 5500 15688 5506 15700
rect 5500 15660 6132 15688
rect 5500 15648 5506 15660
rect 3697 15623 3755 15629
rect 3697 15589 3709 15623
rect 3743 15620 3755 15623
rect 4154 15620 4160 15632
rect 3743 15592 4160 15620
rect 3743 15589 3755 15592
rect 3697 15583 3755 15589
rect 4154 15580 4160 15592
rect 4212 15620 4218 15632
rect 4982 15620 4988 15632
rect 4212 15592 4988 15620
rect 4212 15580 4218 15592
rect 4982 15580 4988 15592
rect 5040 15580 5046 15632
rect 5715 15623 5773 15629
rect 5715 15589 5727 15623
rect 5761 15589 5773 15623
rect 6104 15620 6132 15660
rect 6178 15648 6184 15700
rect 6236 15688 6242 15700
rect 6273 15691 6331 15697
rect 6273 15688 6285 15691
rect 6236 15660 6285 15688
rect 6236 15648 6242 15660
rect 6273 15657 6285 15660
rect 6319 15657 6331 15691
rect 6273 15651 6331 15657
rect 6362 15648 6368 15700
rect 6420 15688 6426 15700
rect 7009 15691 7067 15697
rect 7009 15688 7021 15691
rect 6420 15660 7021 15688
rect 6420 15648 6426 15660
rect 7009 15657 7021 15660
rect 7055 15688 7067 15691
rect 7558 15688 7564 15700
rect 7055 15660 7564 15688
rect 7055 15657 7067 15660
rect 7009 15651 7067 15657
rect 7558 15648 7564 15660
rect 7616 15648 7622 15700
rect 8662 15688 8668 15700
rect 8623 15660 8668 15688
rect 8662 15648 8668 15660
rect 8720 15648 8726 15700
rect 9398 15648 9404 15700
rect 9456 15688 9462 15700
rect 9493 15691 9551 15697
rect 9493 15688 9505 15691
rect 9456 15660 9505 15688
rect 9456 15648 9462 15660
rect 9493 15657 9505 15660
rect 9539 15688 9551 15691
rect 9858 15688 9864 15700
rect 9539 15660 9864 15688
rect 9539 15657 9551 15660
rect 9493 15651 9551 15657
rect 9858 15648 9864 15660
rect 9916 15648 9922 15700
rect 11514 15688 11520 15700
rect 11475 15660 11520 15688
rect 11514 15648 11520 15660
rect 11572 15648 11578 15700
rect 12621 15691 12679 15697
rect 12621 15657 12633 15691
rect 12667 15688 12679 15691
rect 13446 15688 13452 15700
rect 12667 15660 13452 15688
rect 12667 15657 12679 15660
rect 12621 15651 12679 15657
rect 13446 15648 13452 15660
rect 13504 15688 13510 15700
rect 13504 15660 13676 15688
rect 13504 15648 13510 15660
rect 6380 15620 6408 15648
rect 6104 15592 6408 15620
rect 7422 15623 7480 15629
rect 5715 15583 5773 15589
rect 7422 15589 7434 15623
rect 7468 15589 7480 15623
rect 7422 15583 7480 15589
rect 3234 15552 3240 15564
rect 3160 15524 3240 15552
rect 3234 15512 3240 15524
rect 3292 15512 3298 15564
rect 3878 15512 3884 15564
rect 3936 15552 3942 15564
rect 4408 15555 4466 15561
rect 4408 15552 4420 15555
rect 3936 15524 4420 15552
rect 3936 15512 3942 15524
rect 4408 15521 4420 15524
rect 4454 15552 4466 15555
rect 4522 15552 4528 15564
rect 4454 15524 4528 15552
rect 4454 15521 4466 15524
rect 4408 15515 4466 15521
rect 4522 15512 4528 15524
rect 4580 15512 4586 15564
rect 5258 15512 5264 15564
rect 5316 15552 5322 15564
rect 5353 15555 5411 15561
rect 5353 15552 5365 15555
rect 5316 15524 5365 15552
rect 5316 15512 5322 15524
rect 5353 15521 5365 15524
rect 5399 15521 5411 15555
rect 5730 15552 5758 15583
rect 6178 15552 6184 15564
rect 5730 15524 6184 15552
rect 5353 15515 5411 15521
rect 6178 15512 6184 15524
rect 6236 15552 6242 15564
rect 7437 15552 7465 15583
rect 10042 15580 10048 15632
rect 10100 15620 10106 15632
rect 10274 15623 10332 15629
rect 10274 15620 10286 15623
rect 10100 15592 10286 15620
rect 10100 15580 10106 15592
rect 10274 15589 10286 15592
rect 10320 15589 10332 15623
rect 10274 15583 10332 15589
rect 11882 15580 11888 15632
rect 11940 15620 11946 15632
rect 12022 15623 12080 15629
rect 12022 15620 12034 15623
rect 11940 15592 12034 15620
rect 11940 15580 11946 15592
rect 12022 15589 12034 15592
rect 12068 15589 12080 15623
rect 13262 15620 13268 15632
rect 13223 15592 13268 15620
rect 12022 15583 12080 15589
rect 13262 15580 13268 15592
rect 13320 15620 13326 15632
rect 13648 15629 13676 15660
rect 13906 15648 13912 15700
rect 13964 15688 13970 15700
rect 14461 15691 14519 15697
rect 14461 15688 14473 15691
rect 13964 15660 14473 15688
rect 13964 15648 13970 15660
rect 14461 15657 14473 15660
rect 14507 15657 14519 15691
rect 14461 15651 14519 15657
rect 16025 15691 16083 15697
rect 16025 15657 16037 15691
rect 16071 15688 16083 15691
rect 16114 15688 16120 15700
rect 16071 15660 16120 15688
rect 16071 15657 16083 15660
rect 16025 15651 16083 15657
rect 16114 15648 16120 15660
rect 16172 15688 16178 15700
rect 16761 15691 16819 15697
rect 16761 15688 16773 15691
rect 16172 15660 16773 15688
rect 16172 15648 16178 15660
rect 16761 15657 16773 15660
rect 16807 15657 16819 15691
rect 16761 15651 16819 15657
rect 19334 15648 19340 15700
rect 19392 15688 19398 15700
rect 19705 15691 19763 15697
rect 19705 15688 19717 15691
rect 19392 15660 19717 15688
rect 19392 15648 19398 15660
rect 19705 15657 19717 15660
rect 19751 15657 19763 15691
rect 19705 15651 19763 15657
rect 21269 15691 21327 15697
rect 21269 15657 21281 15691
rect 21315 15688 21327 15691
rect 21358 15688 21364 15700
rect 21315 15660 21364 15688
rect 21315 15657 21327 15660
rect 21269 15651 21327 15657
rect 21358 15648 21364 15660
rect 21416 15648 21422 15700
rect 21542 15688 21548 15700
rect 21503 15660 21548 15688
rect 21542 15648 21548 15660
rect 21600 15648 21606 15700
rect 24026 15688 24032 15700
rect 23987 15660 24032 15688
rect 24026 15648 24032 15660
rect 24084 15648 24090 15700
rect 13541 15623 13599 15629
rect 13541 15620 13553 15623
rect 13320 15592 13553 15620
rect 13320 15580 13326 15592
rect 13541 15589 13553 15592
rect 13587 15589 13599 15623
rect 13541 15583 13599 15589
rect 13633 15623 13691 15629
rect 13633 15589 13645 15623
rect 13679 15589 13691 15623
rect 13633 15583 13691 15589
rect 17954 15580 17960 15632
rect 18012 15620 18018 15632
rect 18138 15620 18144 15632
rect 18012 15592 18144 15620
rect 18012 15580 18018 15592
rect 18138 15580 18144 15592
rect 18196 15580 18202 15632
rect 18414 15580 18420 15632
rect 18472 15620 18478 15632
rect 18874 15629 18880 15632
rect 18830 15623 18880 15629
rect 18830 15620 18842 15623
rect 18472 15592 18842 15620
rect 18472 15580 18478 15592
rect 18830 15589 18842 15592
rect 18876 15589 18880 15623
rect 18830 15583 18880 15589
rect 18874 15580 18880 15583
rect 18932 15580 18938 15632
rect 22050 15623 22108 15629
rect 22050 15589 22062 15623
rect 22096 15620 22108 15623
rect 23198 15620 23204 15632
rect 22096 15592 23204 15620
rect 22096 15589 22108 15592
rect 22050 15583 22108 15589
rect 6236 15524 7465 15552
rect 6236 15512 6242 15524
rect 8754 15512 8760 15564
rect 8812 15552 8818 15564
rect 9950 15552 9956 15564
rect 8812 15524 9956 15552
rect 8812 15512 8818 15524
rect 9950 15512 9956 15524
rect 10008 15512 10014 15564
rect 10873 15555 10931 15561
rect 10873 15521 10885 15555
rect 10919 15552 10931 15555
rect 11790 15552 11796 15564
rect 10919 15524 11796 15552
rect 10919 15521 10931 15524
rect 10873 15515 10931 15521
rect 11790 15512 11796 15524
rect 11848 15552 11854 15564
rect 12250 15552 12256 15564
rect 11848 15524 12256 15552
rect 11848 15512 11854 15524
rect 12250 15512 12256 15524
rect 12308 15512 12314 15564
rect 14550 15512 14556 15564
rect 14608 15552 14614 15564
rect 15746 15552 15752 15564
rect 14608 15524 15752 15552
rect 14608 15512 14614 15524
rect 15746 15512 15752 15524
rect 15804 15512 15810 15564
rect 16301 15555 16359 15561
rect 16301 15521 16313 15555
rect 16347 15552 16359 15555
rect 16577 15555 16635 15561
rect 16577 15552 16589 15555
rect 16347 15524 16589 15552
rect 16347 15521 16359 15524
rect 16301 15515 16359 15521
rect 16577 15521 16589 15524
rect 16623 15521 16635 15555
rect 16577 15515 16635 15521
rect 16666 15512 16672 15564
rect 16724 15552 16730 15564
rect 17310 15552 17316 15564
rect 16724 15524 17316 15552
rect 16724 15512 16730 15524
rect 17310 15512 17316 15524
rect 17368 15512 17374 15564
rect 19429 15555 19487 15561
rect 19429 15521 19441 15555
rect 19475 15552 19487 15555
rect 20806 15552 20812 15564
rect 19475 15524 20812 15552
rect 19475 15521 19487 15524
rect 19429 15515 19487 15521
rect 20806 15512 20812 15524
rect 20864 15512 20870 15564
rect 21729 15555 21787 15561
rect 21729 15521 21741 15555
rect 21775 15552 21787 15555
rect 21818 15552 21824 15564
rect 21775 15524 21824 15552
rect 21775 15521 21787 15524
rect 21729 15515 21787 15521
rect 21818 15512 21824 15524
rect 21876 15512 21882 15564
rect 2866 15484 2872 15496
rect 2779 15456 2872 15484
rect 2866 15444 2872 15456
rect 2924 15484 2930 15496
rect 3694 15484 3700 15496
rect 2924 15456 3700 15484
rect 2924 15444 2930 15456
rect 3694 15444 3700 15456
rect 3752 15444 3758 15496
rect 7098 15484 7104 15496
rect 7059 15456 7104 15484
rect 7098 15444 7104 15456
rect 7156 15444 7162 15496
rect 11698 15484 11704 15496
rect 11659 15456 11704 15484
rect 11698 15444 11704 15456
rect 11756 15444 11762 15496
rect 13817 15487 13875 15493
rect 13817 15453 13829 15487
rect 13863 15453 13875 15487
rect 13817 15447 13875 15453
rect 18509 15487 18567 15493
rect 18509 15453 18521 15487
rect 18555 15484 18567 15487
rect 19518 15484 19524 15496
rect 18555 15456 19524 15484
rect 18555 15453 18567 15456
rect 18509 15447 18567 15453
rect 4479 15419 4537 15425
rect 4479 15385 4491 15419
rect 4525 15416 4537 15419
rect 7190 15416 7196 15428
rect 4525 15388 7196 15416
rect 4525 15385 4537 15388
rect 4479 15379 4537 15385
rect 7190 15376 7196 15388
rect 7248 15376 7254 15428
rect 8389 15419 8447 15425
rect 8389 15385 8401 15419
rect 8435 15416 8447 15419
rect 8478 15416 8484 15428
rect 8435 15388 8484 15416
rect 8435 15385 8447 15388
rect 8389 15379 8447 15385
rect 8478 15376 8484 15388
rect 8536 15416 8542 15428
rect 12894 15416 12900 15428
rect 8536 15388 12900 15416
rect 8536 15376 8542 15388
rect 12894 15376 12900 15388
rect 12952 15376 12958 15428
rect 13170 15376 13176 15428
rect 13228 15416 13234 15428
rect 13832 15416 13860 15447
rect 19518 15444 19524 15456
rect 19576 15444 19582 15496
rect 21542 15444 21548 15496
rect 21600 15484 21606 15496
rect 22065 15484 22093 15583
rect 23198 15580 23204 15592
rect 23256 15580 23262 15632
rect 23382 15512 23388 15564
rect 23440 15552 23446 15564
rect 23661 15555 23719 15561
rect 23661 15552 23673 15555
rect 23440 15524 23673 15552
rect 23440 15512 23446 15524
rect 23661 15521 23673 15524
rect 23707 15521 23719 15555
rect 23661 15515 23719 15521
rect 24026 15512 24032 15564
rect 24084 15552 24090 15564
rect 24210 15552 24216 15564
rect 24084 15524 24216 15552
rect 24084 15512 24090 15524
rect 24210 15512 24216 15524
rect 24268 15512 24274 15564
rect 25406 15552 25412 15564
rect 25367 15524 25412 15552
rect 25406 15512 25412 15524
rect 25464 15512 25470 15564
rect 21600 15456 22093 15484
rect 21600 15444 21606 15456
rect 13906 15416 13912 15428
rect 13228 15388 13912 15416
rect 13228 15376 13234 15388
rect 13906 15376 13912 15388
rect 13964 15376 13970 15428
rect 16114 15376 16120 15428
rect 16172 15416 16178 15428
rect 17678 15416 17684 15428
rect 16172 15388 17684 15416
rect 16172 15376 16178 15388
rect 17678 15376 17684 15388
rect 17736 15416 17742 15428
rect 17865 15419 17923 15425
rect 17865 15416 17877 15419
rect 17736 15388 17877 15416
rect 17736 15376 17742 15388
rect 17865 15385 17877 15388
rect 17911 15385 17923 15419
rect 17865 15379 17923 15385
rect 1854 15348 1860 15360
rect 1815 15320 1860 15348
rect 1854 15308 1860 15320
rect 1912 15308 1918 15360
rect 2406 15348 2412 15360
rect 2367 15320 2412 15348
rect 2406 15308 2412 15320
rect 2464 15308 2470 15360
rect 2590 15308 2596 15360
rect 2648 15348 2654 15360
rect 3145 15351 3203 15357
rect 3145 15348 3157 15351
rect 2648 15320 3157 15348
rect 2648 15308 2654 15320
rect 3145 15317 3157 15320
rect 3191 15317 3203 15351
rect 4798 15348 4804 15360
rect 4759 15320 4804 15348
rect 3145 15311 3203 15317
rect 4798 15308 4804 15320
rect 4856 15308 4862 15360
rect 6546 15348 6552 15360
rect 6507 15320 6552 15348
rect 6546 15308 6552 15320
rect 6604 15308 6610 15360
rect 7006 15308 7012 15360
rect 7064 15348 7070 15360
rect 8021 15351 8079 15357
rect 8021 15348 8033 15351
rect 7064 15320 8033 15348
rect 7064 15308 7070 15320
rect 8021 15317 8033 15320
rect 8067 15317 8079 15351
rect 8021 15311 8079 15317
rect 16390 15308 16396 15360
rect 16448 15348 16454 15360
rect 16577 15351 16635 15357
rect 16577 15348 16589 15351
rect 16448 15320 16589 15348
rect 16448 15308 16454 15320
rect 16577 15317 16589 15320
rect 16623 15348 16635 15351
rect 17497 15351 17555 15357
rect 17497 15348 17509 15351
rect 16623 15320 17509 15348
rect 16623 15317 16635 15320
rect 16577 15311 16635 15317
rect 17497 15317 17509 15320
rect 17543 15348 17555 15351
rect 18598 15348 18604 15360
rect 17543 15320 18604 15348
rect 17543 15317 17555 15320
rect 17497 15311 17555 15317
rect 18598 15308 18604 15320
rect 18656 15348 18662 15360
rect 19150 15348 19156 15360
rect 18656 15320 19156 15348
rect 18656 15308 18662 15320
rect 19150 15308 19156 15320
rect 19208 15308 19214 15360
rect 22186 15308 22192 15360
rect 22244 15348 22250 15360
rect 22649 15351 22707 15357
rect 22649 15348 22661 15351
rect 22244 15320 22661 15348
rect 22244 15308 22250 15320
rect 22649 15317 22661 15320
rect 22695 15317 22707 15351
rect 22649 15311 22707 15317
rect 24581 15351 24639 15357
rect 24581 15317 24593 15351
rect 24627 15348 24639 15351
rect 24670 15348 24676 15360
rect 24627 15320 24676 15348
rect 24627 15317 24639 15320
rect 24581 15311 24639 15317
rect 24670 15308 24676 15320
rect 24728 15308 24734 15360
rect 24946 15348 24952 15360
rect 24859 15320 24952 15348
rect 24946 15308 24952 15320
rect 25004 15348 25010 15360
rect 25547 15351 25605 15357
rect 25547 15348 25559 15351
rect 25004 15320 25559 15348
rect 25004 15308 25010 15320
rect 25547 15317 25559 15320
rect 25593 15317 25605 15351
rect 25547 15311 25605 15317
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 2114 15147 2172 15153
rect 2114 15113 2126 15147
rect 2160 15144 2172 15147
rect 2498 15144 2504 15156
rect 2160 15116 2504 15144
rect 2160 15113 2172 15116
rect 2114 15107 2172 15113
rect 2498 15104 2504 15116
rect 2556 15144 2562 15156
rect 2866 15144 2872 15156
rect 2556 15116 2872 15144
rect 2556 15104 2562 15116
rect 2866 15104 2872 15116
rect 2924 15104 2930 15156
rect 4522 15144 4528 15156
rect 4483 15116 4528 15144
rect 4522 15104 4528 15116
rect 4580 15104 4586 15156
rect 9398 15144 9404 15156
rect 9359 15116 9404 15144
rect 9398 15104 9404 15116
rect 9456 15104 9462 15156
rect 10042 15144 10048 15156
rect 9955 15116 10048 15144
rect 10042 15104 10048 15116
rect 10100 15144 10106 15156
rect 11882 15144 11888 15156
rect 10100 15116 11888 15144
rect 10100 15104 10106 15116
rect 11882 15104 11888 15116
rect 11940 15104 11946 15156
rect 12986 15144 12992 15156
rect 12947 15116 12992 15144
rect 12986 15104 12992 15116
rect 13044 15104 13050 15156
rect 13446 15144 13452 15156
rect 13407 15116 13452 15144
rect 13446 15104 13452 15116
rect 13504 15104 13510 15156
rect 15746 15104 15752 15156
rect 15804 15144 15810 15156
rect 16669 15147 16727 15153
rect 16669 15144 16681 15147
rect 15804 15116 16681 15144
rect 15804 15104 15810 15116
rect 16669 15113 16681 15116
rect 16715 15113 16727 15147
rect 17310 15144 17316 15156
rect 17271 15116 17316 15144
rect 16669 15107 16727 15113
rect 17310 15104 17316 15116
rect 17368 15104 17374 15156
rect 19518 15104 19524 15156
rect 19576 15144 19582 15156
rect 19613 15147 19671 15153
rect 19613 15144 19625 15147
rect 19576 15116 19625 15144
rect 19576 15104 19582 15116
rect 19613 15113 19625 15116
rect 19659 15113 19671 15147
rect 23106 15144 23112 15156
rect 19613 15107 19671 15113
rect 19720 15116 23112 15144
rect 2222 15076 2228 15088
rect 2183 15048 2228 15076
rect 2222 15036 2228 15048
rect 2280 15076 2286 15088
rect 2961 15079 3019 15085
rect 2961 15076 2973 15079
rect 2280 15048 2973 15076
rect 2280 15036 2286 15048
rect 2961 15045 2973 15048
rect 3007 15045 3019 15079
rect 2961 15039 3019 15045
rect 4430 15036 4436 15088
rect 4488 15076 4494 15088
rect 6549 15079 6607 15085
rect 6549 15076 6561 15079
rect 4488 15048 6561 15076
rect 4488 15036 4494 15048
rect 6549 15045 6561 15048
rect 6595 15076 6607 15079
rect 6914 15076 6920 15088
rect 6595 15048 6920 15076
rect 6595 15045 6607 15048
rect 6549 15039 6607 15045
rect 6914 15036 6920 15048
rect 6972 15036 6978 15088
rect 11698 15036 11704 15088
rect 11756 15076 11762 15088
rect 12253 15079 12311 15085
rect 12253 15076 12265 15079
rect 11756 15048 12265 15076
rect 11756 15036 11762 15048
rect 12253 15045 12265 15048
rect 12299 15076 12311 15079
rect 14090 15076 14096 15088
rect 12299 15048 14096 15076
rect 12299 15045 12311 15048
rect 12253 15039 12311 15045
rect 14090 15036 14096 15048
rect 14148 15036 14154 15088
rect 17034 15076 17040 15088
rect 16086 15048 17040 15076
rect 2314 15008 2320 15020
rect 2275 14980 2320 15008
rect 2314 14968 2320 14980
rect 2372 14968 2378 15020
rect 4249 15011 4307 15017
rect 3804 14980 4200 15008
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14940 2007 14943
rect 2406 14940 2412 14952
rect 1995 14912 2412 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2406 14900 2412 14912
rect 2464 14900 2470 14952
rect 2590 14900 2596 14952
rect 2648 14940 2654 14952
rect 2866 14940 2872 14952
rect 2648 14912 2872 14940
rect 2648 14900 2654 14912
rect 2866 14900 2872 14912
rect 2924 14900 2930 14952
rect 3804 14949 3832 14980
rect 3421 14943 3479 14949
rect 3421 14909 3433 14943
rect 3467 14940 3479 14943
rect 3789 14943 3847 14949
rect 3789 14940 3801 14943
rect 3467 14912 3801 14940
rect 3467 14909 3479 14912
rect 3421 14903 3479 14909
rect 3789 14909 3801 14912
rect 3835 14909 3847 14943
rect 3970 14940 3976 14952
rect 3931 14912 3976 14940
rect 3789 14903 3847 14909
rect 3970 14900 3976 14912
rect 4028 14900 4034 14952
rect 4172 14940 4200 14980
rect 4249 14977 4261 15011
rect 4295 15008 4307 15011
rect 5813 15011 5871 15017
rect 4295 14980 5758 15008
rect 4295 14977 4307 14980
rect 4249 14971 4307 14977
rect 4890 14940 4896 14952
rect 4172 14912 4896 14940
rect 4890 14900 4896 14912
rect 4948 14900 4954 14952
rect 5169 14943 5227 14949
rect 5169 14909 5181 14943
rect 5215 14909 5227 14943
rect 5169 14903 5227 14909
rect 2685 14875 2743 14881
rect 2685 14841 2697 14875
rect 2731 14872 2743 14875
rect 4154 14872 4160 14884
rect 2731 14844 4160 14872
rect 2731 14841 2743 14844
rect 2685 14835 2743 14841
rect 4154 14832 4160 14844
rect 4212 14832 4218 14884
rect 5184 14816 5212 14903
rect 5442 14900 5448 14952
rect 5500 14940 5506 14952
rect 5537 14943 5595 14949
rect 5537 14940 5549 14943
rect 5500 14912 5549 14940
rect 5500 14900 5506 14912
rect 5537 14909 5549 14912
rect 5583 14909 5595 14943
rect 5730 14940 5758 14980
rect 5813 14977 5825 15011
rect 5859 15008 5871 15011
rect 7098 15008 7104 15020
rect 5859 14980 7104 15008
rect 5859 14977 5871 14980
rect 5813 14971 5871 14977
rect 7098 14968 7104 14980
rect 7156 14968 7162 15020
rect 7374 15008 7380 15020
rect 7335 14980 7380 15008
rect 7374 14968 7380 14980
rect 7432 14968 7438 15020
rect 7926 14968 7932 15020
rect 7984 15008 7990 15020
rect 8478 15008 8484 15020
rect 7984 14980 8484 15008
rect 7984 14968 7990 14980
rect 8478 14968 8484 14980
rect 8536 14968 8542 15020
rect 10778 14968 10784 15020
rect 10836 15008 10842 15020
rect 13725 15011 13783 15017
rect 10836 14980 11284 15008
rect 10836 14968 10842 14980
rect 6730 14940 6736 14952
rect 5730 14912 6736 14940
rect 5537 14903 5595 14909
rect 5552 14872 5580 14903
rect 6730 14900 6736 14912
rect 6788 14900 6794 14952
rect 10689 14943 10747 14949
rect 10689 14909 10701 14943
rect 10735 14940 10747 14943
rect 11054 14940 11060 14952
rect 10735 14912 11060 14940
rect 10735 14909 10747 14912
rect 10689 14903 10747 14909
rect 11054 14900 11060 14912
rect 11112 14900 11118 14952
rect 11256 14949 11284 14980
rect 13725 14977 13737 15011
rect 13771 15008 13783 15011
rect 13814 15008 13820 15020
rect 13771 14980 13820 15008
rect 13771 14977 13783 14980
rect 13725 14971 13783 14977
rect 13814 14968 13820 14980
rect 13872 14968 13878 15020
rect 14182 14968 14188 15020
rect 14240 15008 14246 15020
rect 14829 15011 14887 15017
rect 14829 15008 14841 15011
rect 14240 14980 14841 15008
rect 14240 14968 14246 14980
rect 14829 14977 14841 14980
rect 14875 15008 14887 15011
rect 16086 15008 16114 15048
rect 17034 15036 17040 15048
rect 17092 15076 17098 15088
rect 18966 15076 18972 15088
rect 17092 15048 18972 15076
rect 17092 15036 17098 15048
rect 18966 15036 18972 15048
rect 19024 15036 19030 15088
rect 16206 15008 16212 15020
rect 14875 14980 16114 15008
rect 16167 14980 16212 15008
rect 14875 14977 14887 14980
rect 14829 14971 14887 14977
rect 11241 14943 11299 14949
rect 11241 14909 11253 14943
rect 11287 14940 11299 14943
rect 12158 14940 12164 14952
rect 11287 14912 12164 14940
rect 11287 14909 11299 14912
rect 11241 14903 11299 14909
rect 12158 14900 12164 14912
rect 12216 14900 12222 14952
rect 12504 14943 12562 14949
rect 12504 14909 12516 14943
rect 12550 14940 12562 14943
rect 12986 14940 12992 14952
rect 12550 14912 12992 14940
rect 12550 14909 12562 14912
rect 12504 14903 12562 14909
rect 12986 14900 12992 14912
rect 13044 14900 13050 14952
rect 15948 14949 15976 14980
rect 16206 14968 16212 14980
rect 16264 14968 16270 15020
rect 19337 15011 19395 15017
rect 19337 14977 19349 15011
rect 19383 15008 19395 15011
rect 19426 15008 19432 15020
rect 19383 14980 19432 15008
rect 19383 14977 19395 14980
rect 19337 14971 19395 14977
rect 19426 14968 19432 14980
rect 19484 14968 19490 15020
rect 15933 14943 15991 14949
rect 15933 14909 15945 14943
rect 15979 14909 15991 14943
rect 15933 14903 15991 14909
rect 16117 14943 16175 14949
rect 16117 14909 16129 14943
rect 16163 14940 16175 14943
rect 16390 14940 16396 14952
rect 16163 14912 16396 14940
rect 16163 14909 16175 14912
rect 16117 14903 16175 14909
rect 5718 14872 5724 14884
rect 5552 14844 5724 14872
rect 5718 14832 5724 14844
rect 5776 14832 5782 14884
rect 6914 14872 6920 14884
rect 6875 14844 6920 14872
rect 6914 14832 6920 14844
rect 6972 14832 6978 14884
rect 7006 14832 7012 14884
rect 7064 14872 7070 14884
rect 8802 14875 8860 14881
rect 7064 14844 7109 14872
rect 7064 14832 7070 14844
rect 8802 14841 8814 14875
rect 8848 14841 8860 14875
rect 11514 14872 11520 14884
rect 11475 14844 11520 14872
rect 8802 14835 8860 14841
rect 1673 14807 1731 14813
rect 1673 14773 1685 14807
rect 1719 14804 1731 14807
rect 1946 14804 1952 14816
rect 1719 14776 1952 14804
rect 1719 14773 1731 14776
rect 1673 14767 1731 14773
rect 1946 14764 1952 14776
rect 2004 14804 2010 14816
rect 2590 14804 2596 14816
rect 2004 14776 2596 14804
rect 2004 14764 2010 14776
rect 2590 14764 2596 14776
rect 2648 14764 2654 14816
rect 4985 14807 5043 14813
rect 4985 14773 4997 14807
rect 5031 14804 5043 14807
rect 5166 14804 5172 14816
rect 5031 14776 5172 14804
rect 5031 14773 5043 14776
rect 4985 14767 5043 14773
rect 5166 14764 5172 14776
rect 5224 14764 5230 14816
rect 6178 14804 6184 14816
rect 6091 14776 6184 14804
rect 6178 14764 6184 14776
rect 6236 14804 6242 14816
rect 6638 14804 6644 14816
rect 6236 14776 6644 14804
rect 6236 14764 6242 14776
rect 6638 14764 6644 14776
rect 6696 14804 6702 14816
rect 7837 14807 7895 14813
rect 7837 14804 7849 14807
rect 6696 14776 7849 14804
rect 6696 14764 6702 14776
rect 7837 14773 7849 14776
rect 7883 14804 7895 14807
rect 8294 14804 8300 14816
rect 7883 14776 8300 14804
rect 7883 14773 7895 14776
rect 7837 14767 7895 14773
rect 8294 14764 8300 14776
rect 8352 14804 8358 14816
rect 8817 14804 8845 14835
rect 11514 14832 11520 14844
rect 11572 14832 11578 14884
rect 13817 14875 13875 14881
rect 13817 14841 13829 14875
rect 13863 14841 13875 14875
rect 14366 14872 14372 14884
rect 14327 14844 14372 14872
rect 13817 14835 13875 14841
rect 8352 14776 8845 14804
rect 8352 14764 8358 14776
rect 10686 14764 10692 14816
rect 10744 14804 10750 14816
rect 11606 14804 11612 14816
rect 10744 14776 11612 14804
rect 10744 14764 10750 14776
rect 11606 14764 11612 14776
rect 11664 14764 11670 14816
rect 11882 14804 11888 14816
rect 11843 14776 11888 14804
rect 11882 14764 11888 14776
rect 11940 14764 11946 14816
rect 12434 14764 12440 14816
rect 12492 14804 12498 14816
rect 12575 14807 12633 14813
rect 12575 14804 12587 14807
rect 12492 14776 12587 14804
rect 12492 14764 12498 14776
rect 12575 14773 12587 14776
rect 12621 14773 12633 14807
rect 12575 14767 12633 14773
rect 13446 14764 13452 14816
rect 13504 14804 13510 14816
rect 13832 14804 13860 14835
rect 14366 14832 14372 14844
rect 14424 14832 14430 14884
rect 15197 14875 15255 14881
rect 15197 14841 15209 14875
rect 15243 14872 15255 14875
rect 15565 14875 15623 14881
rect 15565 14872 15577 14875
rect 15243 14844 15577 14872
rect 15243 14841 15255 14844
rect 15197 14835 15255 14841
rect 15565 14841 15577 14844
rect 15611 14872 15623 14875
rect 16132 14872 16160 14903
rect 16390 14900 16396 14912
rect 16448 14900 16454 14952
rect 18598 14940 18604 14952
rect 17788 14912 18604 14940
rect 15611 14844 16160 14872
rect 15611 14841 15623 14844
rect 15565 14835 15623 14841
rect 13504 14776 13860 14804
rect 13504 14764 13510 14776
rect 17678 14764 17684 14816
rect 17736 14804 17742 14816
rect 17788 14813 17816 14912
rect 18598 14900 18604 14912
rect 18656 14900 18662 14952
rect 19150 14940 19156 14952
rect 19063 14912 19156 14940
rect 19150 14900 19156 14912
rect 19208 14940 19214 14952
rect 19720 14940 19748 15116
rect 23106 15104 23112 15116
rect 23164 15104 23170 15156
rect 23382 15144 23388 15156
rect 23343 15116 23388 15144
rect 23382 15104 23388 15116
rect 23440 15104 23446 15156
rect 24397 15147 24455 15153
rect 24397 15113 24409 15147
rect 24443 15144 24455 15147
rect 24670 15144 24676 15156
rect 24443 15116 24676 15144
rect 24443 15113 24455 15116
rect 24397 15107 24455 15113
rect 24670 15104 24676 15116
rect 24728 15104 24734 15156
rect 19978 15036 19984 15088
rect 20036 15076 20042 15088
rect 20036 15048 20852 15076
rect 20036 15036 20042 15048
rect 20530 15008 20536 15020
rect 20491 14980 20536 15008
rect 20530 14968 20536 14980
rect 20588 14968 20594 15020
rect 20824 15017 20852 15048
rect 22002 15036 22008 15088
rect 22060 15076 22066 15088
rect 22649 15079 22707 15085
rect 22649 15076 22661 15079
rect 22060 15048 22661 15076
rect 22060 15036 22066 15048
rect 22649 15045 22661 15048
rect 22695 15045 22707 15079
rect 22649 15039 22707 15045
rect 23198 15036 23204 15088
rect 23256 15076 23262 15088
rect 23845 15079 23903 15085
rect 23845 15076 23857 15079
rect 23256 15048 23857 15076
rect 23256 15036 23262 15048
rect 23845 15045 23857 15048
rect 23891 15045 23903 15079
rect 23845 15039 23903 15045
rect 20809 15011 20867 15017
rect 20809 14977 20821 15011
rect 20855 15008 20867 15011
rect 21910 15008 21916 15020
rect 20855 14980 21916 15008
rect 20855 14977 20867 14980
rect 20809 14971 20867 14977
rect 21910 14968 21916 14980
rect 21968 15008 21974 15020
rect 22097 15011 22155 15017
rect 22097 15008 22109 15011
rect 21968 14980 22109 15008
rect 21968 14968 21974 14980
rect 22097 14977 22109 14980
rect 22143 15008 22155 15011
rect 23017 15011 23075 15017
rect 23017 15008 23029 15011
rect 22143 14980 23029 15008
rect 22143 14977 22155 14980
rect 22097 14971 22155 14977
rect 23017 14977 23029 14980
rect 23063 14977 23075 15011
rect 23017 14971 23075 14977
rect 24581 15011 24639 15017
rect 24581 14977 24593 15011
rect 24627 15008 24639 15011
rect 24946 15008 24952 15020
rect 24627 14980 24952 15008
rect 24627 14977 24639 14980
rect 24581 14971 24639 14977
rect 24946 14968 24952 14980
rect 25004 14968 25010 15020
rect 25222 15008 25228 15020
rect 25183 14980 25228 15008
rect 25222 14968 25228 14980
rect 25280 14968 25286 15020
rect 19208 14912 19748 14940
rect 19208 14900 19214 14912
rect 20625 14875 20683 14881
rect 20625 14841 20637 14875
rect 20671 14872 20683 14875
rect 20806 14872 20812 14884
rect 20671 14844 20812 14872
rect 20671 14841 20683 14844
rect 20625 14835 20683 14841
rect 17773 14807 17831 14813
rect 17773 14804 17785 14807
rect 17736 14776 17785 14804
rect 17736 14764 17742 14776
rect 17773 14773 17785 14776
rect 17819 14773 17831 14807
rect 17773 14767 17831 14773
rect 18138 14764 18144 14816
rect 18196 14804 18202 14816
rect 18414 14804 18420 14816
rect 18196 14776 18420 14804
rect 18196 14764 18202 14776
rect 18414 14764 18420 14776
rect 18472 14764 18478 14816
rect 20349 14807 20407 14813
rect 20349 14773 20361 14807
rect 20395 14804 20407 14807
rect 20640 14804 20668 14835
rect 20806 14832 20812 14844
rect 20864 14832 20870 14884
rect 22186 14832 22192 14884
rect 22244 14872 22250 14884
rect 22244 14844 22289 14872
rect 22244 14832 22250 14844
rect 24670 14832 24676 14884
rect 24728 14872 24734 14884
rect 24728 14844 24773 14872
rect 24728 14832 24734 14844
rect 20395 14776 20668 14804
rect 20395 14773 20407 14776
rect 20349 14767 20407 14773
rect 21542 14764 21548 14816
rect 21600 14804 21606 14816
rect 21729 14807 21787 14813
rect 21729 14804 21741 14807
rect 21600 14776 21741 14804
rect 21600 14764 21606 14776
rect 21729 14773 21741 14776
rect 21775 14773 21787 14807
rect 21729 14767 21787 14773
rect 24854 14764 24860 14816
rect 24912 14804 24918 14816
rect 25406 14804 25412 14816
rect 24912 14776 25412 14804
rect 24912 14764 24918 14776
rect 25406 14764 25412 14776
rect 25464 14804 25470 14816
rect 25501 14807 25559 14813
rect 25501 14804 25513 14807
rect 25464 14776 25513 14804
rect 25464 14764 25470 14776
rect 25501 14773 25513 14776
rect 25547 14773 25559 14807
rect 25501 14767 25559 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1765 14603 1823 14609
rect 1765 14569 1777 14603
rect 1811 14600 1823 14603
rect 2314 14600 2320 14612
rect 1811 14572 2320 14600
rect 1811 14569 1823 14572
rect 1765 14563 1823 14569
rect 2314 14560 2320 14572
rect 2372 14560 2378 14612
rect 2958 14600 2964 14612
rect 2919 14572 2964 14600
rect 2958 14560 2964 14572
rect 3016 14560 3022 14612
rect 3605 14603 3663 14609
rect 3605 14569 3617 14603
rect 3651 14600 3663 14603
rect 3878 14600 3884 14612
rect 3651 14572 3884 14600
rect 3651 14569 3663 14572
rect 3605 14563 3663 14569
rect 3878 14560 3884 14572
rect 3936 14560 3942 14612
rect 5258 14560 5264 14612
rect 5316 14600 5322 14612
rect 5445 14603 5503 14609
rect 5445 14600 5457 14603
rect 5316 14572 5457 14600
rect 5316 14560 5322 14572
rect 5445 14569 5457 14572
rect 5491 14569 5503 14603
rect 5445 14563 5503 14569
rect 6917 14603 6975 14609
rect 6917 14569 6929 14603
rect 6963 14600 6975 14603
rect 7006 14600 7012 14612
rect 6963 14572 7012 14600
rect 6963 14569 6975 14572
rect 6917 14563 6975 14569
rect 7006 14560 7012 14572
rect 7064 14560 7070 14612
rect 7098 14560 7104 14612
rect 7156 14600 7162 14612
rect 7193 14603 7251 14609
rect 7193 14600 7205 14603
rect 7156 14572 7205 14600
rect 7156 14560 7162 14572
rect 7193 14569 7205 14572
rect 7239 14569 7251 14603
rect 7193 14563 7251 14569
rect 7374 14560 7380 14612
rect 7432 14600 7438 14612
rect 8478 14600 8484 14612
rect 7432 14572 7966 14600
rect 8439 14572 8484 14600
rect 7432 14560 7438 14572
rect 2038 14532 2044 14544
rect 1999 14504 2044 14532
rect 2038 14492 2044 14504
rect 2096 14492 2102 14544
rect 2774 14492 2780 14544
rect 2832 14532 2838 14544
rect 3970 14532 3976 14544
rect 2832 14504 3976 14532
rect 2832 14492 2838 14504
rect 3970 14492 3976 14504
rect 4028 14532 4034 14544
rect 4157 14535 4215 14541
rect 4157 14532 4169 14535
rect 4028 14504 4169 14532
rect 4028 14492 4034 14504
rect 4157 14501 4169 14504
rect 4203 14501 4215 14535
rect 4157 14495 4215 14501
rect 4249 14535 4307 14541
rect 4249 14501 4261 14535
rect 4295 14532 4307 14535
rect 4522 14532 4528 14544
rect 4295 14504 4528 14532
rect 4295 14501 4307 14504
rect 4249 14495 4307 14501
rect 4522 14492 4528 14504
rect 4580 14532 4586 14544
rect 6546 14532 6552 14544
rect 4580 14504 6552 14532
rect 4580 14492 4586 14504
rect 6546 14492 6552 14504
rect 6604 14492 6610 14544
rect 7650 14532 7656 14544
rect 7611 14504 7656 14532
rect 7650 14492 7656 14504
rect 7708 14492 7714 14544
rect 7938 14532 7966 14572
rect 8478 14560 8484 14572
rect 8536 14560 8542 14612
rect 9490 14600 9496 14612
rect 9451 14572 9496 14600
rect 9490 14560 9496 14572
rect 9548 14560 9554 14612
rect 10134 14600 10140 14612
rect 9692 14572 10140 14600
rect 9692 14532 9720 14572
rect 10134 14560 10140 14572
rect 10192 14600 10198 14612
rect 10778 14600 10784 14612
rect 10192 14572 10456 14600
rect 10739 14572 10784 14600
rect 10192 14560 10198 14572
rect 7938 14504 9720 14532
rect 9766 14492 9772 14544
rect 9824 14532 9830 14544
rect 10428 14541 10456 14572
rect 10778 14560 10784 14572
rect 10836 14560 10842 14612
rect 13446 14560 13452 14612
rect 13504 14600 13510 14612
rect 14185 14603 14243 14609
rect 14185 14600 14197 14603
rect 13504 14572 14197 14600
rect 13504 14560 13510 14572
rect 14185 14569 14197 14572
rect 14231 14569 14243 14603
rect 14185 14563 14243 14569
rect 14274 14560 14280 14612
rect 14332 14600 14338 14612
rect 14645 14603 14703 14609
rect 14645 14600 14657 14603
rect 14332 14572 14657 14600
rect 14332 14560 14338 14572
rect 14645 14569 14657 14572
rect 14691 14600 14703 14603
rect 16942 14600 16948 14612
rect 14691 14572 16114 14600
rect 16903 14572 16948 14600
rect 14691 14569 14703 14572
rect 14645 14563 14703 14569
rect 9861 14535 9919 14541
rect 9861 14532 9873 14535
rect 9824 14504 9873 14532
rect 9824 14492 9830 14504
rect 9861 14501 9873 14504
rect 9907 14501 9919 14535
rect 9861 14495 9919 14501
rect 10413 14535 10471 14541
rect 10413 14501 10425 14535
rect 10459 14501 10471 14535
rect 11790 14532 11796 14544
rect 11751 14504 11796 14532
rect 10413 14495 10471 14501
rect 11790 14492 11796 14504
rect 11848 14492 11854 14544
rect 13357 14535 13415 14541
rect 13357 14501 13369 14535
rect 13403 14532 13415 14535
rect 13630 14532 13636 14544
rect 13403 14504 13636 14532
rect 13403 14501 13415 14504
rect 13357 14495 13415 14501
rect 13630 14492 13636 14504
rect 13688 14492 13694 14544
rect 13906 14532 13912 14544
rect 13867 14504 13912 14532
rect 13906 14492 13912 14504
rect 13964 14492 13970 14544
rect 15378 14492 15384 14544
rect 15436 14532 15442 14544
rect 15473 14535 15531 14541
rect 15473 14532 15485 14535
rect 15436 14504 15485 14532
rect 15436 14492 15442 14504
rect 15473 14501 15485 14504
rect 15519 14501 15531 14535
rect 16086 14532 16114 14572
rect 16942 14560 16948 14572
rect 17000 14560 17006 14612
rect 18782 14560 18788 14612
rect 18840 14600 18846 14612
rect 18969 14603 19027 14609
rect 18969 14600 18981 14603
rect 18840 14572 18981 14600
rect 18840 14560 18846 14572
rect 18969 14569 18981 14572
rect 19015 14569 19027 14603
rect 20530 14600 20536 14612
rect 20491 14572 20536 14600
rect 18969 14563 19027 14569
rect 20530 14560 20536 14572
rect 20588 14560 20594 14612
rect 22097 14603 22155 14609
rect 22097 14569 22109 14603
rect 22143 14600 22155 14603
rect 22186 14600 22192 14612
rect 22143 14572 22192 14600
rect 22143 14569 22155 14572
rect 22097 14563 22155 14569
rect 22186 14560 22192 14572
rect 22244 14560 22250 14612
rect 23474 14560 23480 14612
rect 23532 14600 23538 14612
rect 23661 14603 23719 14609
rect 23661 14600 23673 14603
rect 23532 14572 23673 14600
rect 23532 14560 23538 14572
rect 23661 14569 23673 14572
rect 23707 14569 23719 14603
rect 24762 14600 24768 14612
rect 23661 14563 23719 14569
rect 24228 14572 24768 14600
rect 18230 14532 18236 14544
rect 16086 14504 18236 14532
rect 15473 14495 15531 14501
rect 18230 14492 18236 14504
rect 18288 14492 18294 14544
rect 18693 14535 18751 14541
rect 18693 14501 18705 14535
rect 18739 14532 18751 14535
rect 19150 14532 19156 14544
rect 18739 14504 19156 14532
rect 18739 14501 18751 14504
rect 18693 14495 18751 14501
rect 19150 14492 19156 14504
rect 19208 14492 19214 14544
rect 19426 14532 19432 14544
rect 19387 14504 19432 14532
rect 19426 14492 19432 14504
rect 19484 14492 19490 14544
rect 21082 14532 21088 14544
rect 21043 14504 21088 14532
rect 21082 14492 21088 14504
rect 21140 14492 21146 14544
rect 21634 14532 21640 14544
rect 21595 14504 21640 14532
rect 21634 14492 21640 14504
rect 21692 14492 21698 14544
rect 21818 14492 21824 14544
rect 21876 14532 21882 14544
rect 22373 14535 22431 14541
rect 22373 14532 22385 14535
rect 21876 14504 22385 14532
rect 21876 14492 21882 14504
rect 22373 14501 22385 14504
rect 22419 14501 22431 14535
rect 23290 14532 23296 14544
rect 23251 14504 23296 14532
rect 22373 14495 22431 14501
rect 23290 14492 23296 14504
rect 23348 14492 23354 14544
rect 24228 14541 24256 14572
rect 24762 14560 24768 14572
rect 24820 14560 24826 14612
rect 24213 14535 24271 14541
rect 24213 14501 24225 14535
rect 24259 14501 24271 14535
rect 24213 14495 24271 14501
rect 24305 14535 24363 14541
rect 24305 14501 24317 14535
rect 24351 14532 24363 14535
rect 24670 14532 24676 14544
rect 24351 14504 24676 14532
rect 24351 14501 24363 14504
rect 24305 14495 24363 14501
rect 24670 14492 24676 14504
rect 24728 14492 24734 14544
rect 5534 14424 5540 14476
rect 5592 14464 5598 14476
rect 5629 14467 5687 14473
rect 5629 14464 5641 14467
rect 5592 14436 5641 14464
rect 5592 14424 5598 14436
rect 5629 14433 5641 14436
rect 5675 14433 5687 14467
rect 6086 14464 6092 14476
rect 6047 14436 6092 14464
rect 5629 14427 5687 14433
rect 6086 14424 6092 14436
rect 6144 14424 6150 14476
rect 17129 14467 17187 14473
rect 17129 14433 17141 14467
rect 17175 14433 17187 14467
rect 17310 14464 17316 14476
rect 17271 14436 17316 14464
rect 17129 14427 17187 14433
rect 1949 14399 2007 14405
rect 1949 14365 1961 14399
rect 1995 14396 2007 14399
rect 2130 14396 2136 14408
rect 1995 14368 2136 14396
rect 1995 14365 2007 14368
rect 1949 14359 2007 14365
rect 2130 14356 2136 14368
rect 2188 14356 2194 14408
rect 2593 14399 2651 14405
rect 2593 14365 2605 14399
rect 2639 14396 2651 14399
rect 3050 14396 3056 14408
rect 2639 14368 3056 14396
rect 2639 14365 2651 14368
rect 2593 14359 2651 14365
rect 3050 14356 3056 14368
rect 3108 14396 3114 14408
rect 5169 14399 5227 14405
rect 3108 14368 4154 14396
rect 3108 14356 3114 14368
rect 4126 14328 4154 14368
rect 5169 14365 5181 14399
rect 5215 14396 5227 14399
rect 5718 14396 5724 14408
rect 5215 14368 5724 14396
rect 5215 14365 5227 14368
rect 5169 14359 5227 14365
rect 5718 14356 5724 14368
rect 5776 14356 5782 14408
rect 6362 14396 6368 14408
rect 6323 14368 6368 14396
rect 6362 14356 6368 14368
rect 6420 14356 6426 14408
rect 7561 14399 7619 14405
rect 7561 14365 7573 14399
rect 7607 14396 7619 14399
rect 8570 14396 8576 14408
rect 7607 14368 8576 14396
rect 7607 14365 7619 14368
rect 7561 14359 7619 14365
rect 8570 14356 8576 14368
rect 8628 14356 8634 14408
rect 9769 14399 9827 14405
rect 9769 14396 9781 14399
rect 9692 14368 9781 14396
rect 9692 14340 9720 14368
rect 9769 14365 9781 14368
rect 9815 14396 9827 14399
rect 11698 14396 11704 14408
rect 9815 14368 11376 14396
rect 11659 14368 11704 14396
rect 9815 14365 9827 14368
rect 9769 14359 9827 14365
rect 4709 14331 4767 14337
rect 4709 14328 4721 14331
rect 4126 14300 4721 14328
rect 4709 14297 4721 14300
rect 4755 14328 4767 14331
rect 8113 14331 8171 14337
rect 8113 14328 8125 14331
rect 4755 14300 8125 14328
rect 4755 14297 4767 14300
rect 4709 14291 4767 14297
rect 8113 14297 8125 14300
rect 8159 14328 8171 14331
rect 9214 14328 9220 14340
rect 8159 14300 9220 14328
rect 8159 14297 8171 14300
rect 8113 14291 8171 14297
rect 9214 14288 9220 14300
rect 9272 14288 9278 14340
rect 9674 14288 9680 14340
rect 9732 14288 9738 14340
rect 11348 14328 11376 14368
rect 11698 14356 11704 14368
rect 11756 14356 11762 14408
rect 12345 14399 12403 14405
rect 12345 14365 12357 14399
rect 12391 14396 12403 14399
rect 12526 14396 12532 14408
rect 12391 14368 12532 14396
rect 12391 14365 12403 14368
rect 12345 14359 12403 14365
rect 12360 14328 12388 14359
rect 12526 14356 12532 14368
rect 12584 14356 12590 14408
rect 13262 14396 13268 14408
rect 13223 14368 13268 14396
rect 13262 14356 13268 14368
rect 13320 14356 13326 14408
rect 15381 14399 15439 14405
rect 15381 14365 15393 14399
rect 15427 14365 15439 14399
rect 15654 14396 15660 14408
rect 15615 14368 15660 14396
rect 15381 14359 15439 14365
rect 11348 14300 12388 14328
rect 14826 14288 14832 14340
rect 14884 14328 14890 14340
rect 15396 14328 15424 14359
rect 15654 14356 15660 14368
rect 15712 14356 15718 14408
rect 17144 14396 17172 14427
rect 17310 14424 17316 14436
rect 17368 14424 17374 14476
rect 22833 14467 22891 14473
rect 22833 14433 22845 14467
rect 22879 14464 22891 14467
rect 22922 14464 22928 14476
rect 22879 14436 22928 14464
rect 22879 14433 22891 14436
rect 22833 14427 22891 14433
rect 22922 14424 22928 14436
rect 22980 14424 22986 14476
rect 23106 14464 23112 14476
rect 23067 14436 23112 14464
rect 23106 14424 23112 14436
rect 23164 14424 23170 14476
rect 17586 14396 17592 14408
rect 17144 14368 17592 14396
rect 17586 14356 17592 14368
rect 17644 14356 17650 14408
rect 19337 14399 19395 14405
rect 19337 14365 19349 14399
rect 19383 14365 19395 14399
rect 19978 14396 19984 14408
rect 19939 14368 19984 14396
rect 19337 14359 19395 14365
rect 15562 14328 15568 14340
rect 14884 14300 15568 14328
rect 14884 14288 14890 14300
rect 15562 14288 15568 14300
rect 15620 14288 15626 14340
rect 19352 14328 19380 14359
rect 19978 14356 19984 14368
rect 20036 14356 20042 14408
rect 20162 14356 20168 14408
rect 20220 14396 20226 14408
rect 20993 14399 21051 14405
rect 20993 14396 21005 14399
rect 20220 14368 21005 14396
rect 20220 14356 20226 14368
rect 20993 14365 21005 14368
rect 21039 14396 21051 14399
rect 21910 14396 21916 14408
rect 21039 14368 21916 14396
rect 21039 14365 21051 14368
rect 20993 14359 21051 14365
rect 21910 14356 21916 14368
rect 21968 14356 21974 14408
rect 24857 14399 24915 14405
rect 24857 14365 24869 14399
rect 24903 14396 24915 14399
rect 24946 14396 24952 14408
rect 24903 14368 24952 14396
rect 24903 14365 24915 14368
rect 24857 14359 24915 14365
rect 19518 14328 19524 14340
rect 19352 14300 19524 14328
rect 19518 14288 19524 14300
rect 19576 14328 19582 14340
rect 20438 14328 20444 14340
rect 19576 14300 20444 14328
rect 19576 14288 19582 14300
rect 20438 14288 20444 14300
rect 20496 14288 20502 14340
rect 22002 14288 22008 14340
rect 22060 14328 22066 14340
rect 24872 14328 24900 14359
rect 24946 14356 24952 14368
rect 25004 14356 25010 14408
rect 22060 14300 24900 14328
rect 22060 14288 22066 14300
rect 4338 14220 4344 14272
rect 4396 14260 4402 14272
rect 8386 14260 8392 14272
rect 4396 14232 8392 14260
rect 4396 14220 4402 14232
rect 8386 14220 8392 14232
rect 8444 14220 8450 14272
rect 8846 14260 8852 14272
rect 8807 14232 8852 14260
rect 8846 14220 8852 14232
rect 8904 14220 8910 14272
rect 14458 14220 14464 14272
rect 14516 14260 14522 14272
rect 22830 14260 22836 14272
rect 14516 14232 22836 14260
rect 14516 14220 14522 14232
rect 22830 14220 22836 14232
rect 22888 14220 22894 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 2038 14016 2044 14068
rect 2096 14056 2102 14068
rect 2685 14059 2743 14065
rect 2685 14056 2697 14059
rect 2096 14028 2697 14056
rect 2096 14016 2102 14028
rect 2685 14025 2697 14028
rect 2731 14056 2743 14059
rect 2961 14059 3019 14065
rect 2961 14056 2973 14059
rect 2731 14028 2973 14056
rect 2731 14025 2743 14028
rect 2685 14019 2743 14025
rect 2961 14025 2973 14028
rect 3007 14025 3019 14059
rect 2961 14019 3019 14025
rect 4433 14059 4491 14065
rect 4433 14025 4445 14059
rect 4479 14056 4491 14059
rect 4522 14056 4528 14068
rect 4479 14028 4528 14056
rect 4479 14025 4491 14028
rect 4433 14019 4491 14025
rect 4522 14016 4528 14028
rect 4580 14016 4586 14068
rect 4614 14016 4620 14068
rect 4672 14056 4678 14068
rect 9398 14056 9404 14068
rect 4672 14028 9404 14056
rect 4672 14016 4678 14028
rect 9398 14016 9404 14028
rect 9456 14016 9462 14068
rect 9677 14059 9735 14065
rect 9677 14025 9689 14059
rect 9723 14056 9735 14059
rect 9766 14056 9772 14068
rect 9723 14028 9772 14056
rect 9723 14025 9735 14028
rect 9677 14019 9735 14025
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 9950 14056 9956 14068
rect 9911 14028 9956 14056
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 11514 14016 11520 14068
rect 11572 14056 11578 14068
rect 11793 14059 11851 14065
rect 11793 14056 11805 14059
rect 11572 14028 11805 14056
rect 11572 14016 11578 14028
rect 11793 14025 11805 14028
rect 11839 14025 11851 14059
rect 11793 14019 11851 14025
rect 13357 14059 13415 14065
rect 13357 14025 13369 14059
rect 13403 14056 13415 14059
rect 13814 14056 13820 14068
rect 13403 14028 13820 14056
rect 13403 14025 13415 14028
rect 13357 14019 13415 14025
rect 2314 13948 2320 14000
rect 2372 13988 2378 14000
rect 2774 13988 2780 14000
rect 2372 13960 2780 13988
rect 2372 13948 2378 13960
rect 2774 13948 2780 13960
rect 2832 13948 2838 14000
rect 3694 13948 3700 14000
rect 3752 13988 3758 14000
rect 3878 13988 3884 14000
rect 3752 13960 3884 13988
rect 3752 13948 3758 13960
rect 3878 13948 3884 13960
rect 3936 13988 3942 14000
rect 4709 13991 4767 13997
rect 4709 13988 4721 13991
rect 3936 13960 4721 13988
rect 3936 13948 3942 13960
rect 4709 13957 4721 13960
rect 4755 13957 4767 13991
rect 4709 13951 4767 13957
rect 4890 13948 4896 14000
rect 4948 13988 4954 14000
rect 5445 13991 5503 13997
rect 5445 13988 5457 13991
rect 4948 13960 5457 13988
rect 4948 13948 4954 13960
rect 5445 13957 5457 13960
rect 5491 13957 5503 13991
rect 9214 13988 9220 14000
rect 9175 13960 9220 13988
rect 5445 13951 5503 13957
rect 9214 13948 9220 13960
rect 9272 13948 9278 14000
rect 1578 13880 1584 13932
rect 1636 13920 1642 13932
rect 1765 13923 1823 13929
rect 1765 13920 1777 13923
rect 1636 13892 1777 13920
rect 1636 13880 1642 13892
rect 1765 13889 1777 13892
rect 1811 13920 1823 13923
rect 3326 13920 3332 13932
rect 1811 13892 3332 13920
rect 1811 13889 1823 13892
rect 1765 13883 1823 13889
rect 3326 13880 3332 13892
rect 3384 13880 3390 13932
rect 3970 13880 3976 13932
rect 4028 13920 4034 13932
rect 5077 13923 5135 13929
rect 5077 13920 5089 13923
rect 4028 13892 5089 13920
rect 4028 13880 4034 13892
rect 5077 13889 5089 13892
rect 5123 13889 5135 13923
rect 5077 13883 5135 13889
rect 5166 13880 5172 13932
rect 5224 13920 5230 13932
rect 5224 13892 5856 13920
rect 5224 13880 5230 13892
rect 3513 13855 3571 13861
rect 3513 13821 3525 13855
rect 3559 13852 3571 13855
rect 4614 13852 4620 13864
rect 3559 13824 4620 13852
rect 3559 13821 3571 13824
rect 3513 13815 3571 13821
rect 4614 13812 4620 13824
rect 4672 13812 4678 13864
rect 5184 13852 5212 13880
rect 5828 13861 5856 13892
rect 6362 13880 6368 13932
rect 6420 13920 6426 13932
rect 6825 13923 6883 13929
rect 6825 13920 6837 13923
rect 6420 13892 6837 13920
rect 6420 13880 6426 13892
rect 6825 13889 6837 13892
rect 6871 13920 6883 13923
rect 8021 13923 8079 13929
rect 8021 13920 8033 13923
rect 6871 13892 8033 13920
rect 6871 13889 6883 13892
rect 6825 13883 6883 13889
rect 8021 13889 8033 13892
rect 8067 13889 8079 13923
rect 8021 13883 8079 13889
rect 8665 13923 8723 13929
rect 8665 13889 8677 13923
rect 8711 13920 8723 13923
rect 8846 13920 8852 13932
rect 8711 13892 8852 13920
rect 8711 13889 8723 13892
rect 8665 13883 8723 13889
rect 8846 13880 8852 13892
rect 8904 13920 8910 13932
rect 8904 13892 9444 13920
rect 8904 13880 8910 13892
rect 5253 13855 5311 13861
rect 5253 13852 5265 13855
rect 5184 13824 5265 13852
rect 1673 13787 1731 13793
rect 1673 13753 1685 13787
rect 1719 13784 1731 13787
rect 2086 13787 2144 13793
rect 2086 13784 2098 13787
rect 1719 13756 2098 13784
rect 1719 13753 1731 13756
rect 1673 13747 1731 13753
rect 2086 13753 2098 13756
rect 2132 13784 2144 13787
rect 3329 13787 3387 13793
rect 3329 13784 3341 13787
rect 2132 13756 3341 13784
rect 2132 13753 2144 13756
rect 2086 13747 2144 13753
rect 3329 13753 3341 13756
rect 3375 13784 3387 13787
rect 3834 13787 3892 13793
rect 3834 13784 3846 13787
rect 3375 13756 3846 13784
rect 3375 13753 3387 13756
rect 3329 13747 3387 13753
rect 3834 13753 3846 13756
rect 3880 13753 3892 13787
rect 3834 13747 3892 13753
rect 3849 13716 3877 13747
rect 4338 13744 4344 13796
rect 4396 13784 4402 13796
rect 5184 13784 5212 13824
rect 5253 13821 5265 13824
rect 5299 13821 5311 13855
rect 5253 13815 5311 13821
rect 5813 13855 5871 13861
rect 5813 13821 5825 13855
rect 5859 13852 5871 13855
rect 8294 13852 8300 13864
rect 5859 13824 8300 13852
rect 5859 13821 5871 13824
rect 5813 13815 5871 13821
rect 8294 13812 8300 13824
rect 8352 13812 8358 13864
rect 6546 13784 6552 13796
rect 4396 13756 5212 13784
rect 5368 13756 6552 13784
rect 4396 13744 4402 13756
rect 5368 13716 5396 13756
rect 6546 13744 6552 13756
rect 6604 13784 6610 13796
rect 7146 13787 7204 13793
rect 7146 13784 7158 13787
rect 6604 13756 7158 13784
rect 6604 13744 6610 13756
rect 7146 13753 7158 13756
rect 7192 13753 7204 13787
rect 7146 13747 7204 13753
rect 8757 13787 8815 13793
rect 8757 13753 8769 13787
rect 8803 13753 8815 13787
rect 9416 13784 9444 13892
rect 9490 13880 9496 13932
rect 9548 13920 9554 13932
rect 10229 13923 10287 13929
rect 10229 13920 10241 13923
rect 9548 13892 10241 13920
rect 9548 13880 9554 13892
rect 10229 13889 10241 13892
rect 10275 13889 10287 13923
rect 11808 13920 11836 14019
rect 13814 14016 13820 14028
rect 13872 14056 13878 14068
rect 15378 14056 15384 14068
rect 13872 14028 15384 14056
rect 13872 14016 13878 14028
rect 15378 14016 15384 14028
rect 15436 14016 15442 14068
rect 17221 14059 17279 14065
rect 17221 14025 17233 14059
rect 17267 14056 17279 14059
rect 17310 14056 17316 14068
rect 17267 14028 17316 14056
rect 17267 14025 17279 14028
rect 17221 14019 17279 14025
rect 17310 14016 17316 14028
rect 17368 14016 17374 14068
rect 17586 14056 17592 14068
rect 17547 14028 17592 14056
rect 17586 14016 17592 14028
rect 17644 14016 17650 14068
rect 19426 14016 19432 14068
rect 19484 14056 19490 14068
rect 19521 14059 19579 14065
rect 19521 14056 19533 14059
rect 19484 14028 19533 14056
rect 19484 14016 19490 14028
rect 19521 14025 19533 14028
rect 19567 14056 19579 14059
rect 19889 14059 19947 14065
rect 19889 14056 19901 14059
rect 19567 14028 19901 14056
rect 19567 14025 19579 14028
rect 19521 14019 19579 14025
rect 19889 14025 19901 14028
rect 19935 14056 19947 14059
rect 20809 14059 20867 14065
rect 20809 14056 20821 14059
rect 19935 14028 20821 14056
rect 19935 14025 19947 14028
rect 19889 14019 19947 14025
rect 20809 14025 20821 14028
rect 20855 14056 20867 14059
rect 21082 14056 21088 14068
rect 20855 14028 21088 14056
rect 20855 14025 20867 14028
rect 20809 14019 20867 14025
rect 21082 14016 21088 14028
rect 21140 14016 21146 14068
rect 21910 14056 21916 14068
rect 21871 14028 21916 14056
rect 21910 14016 21916 14028
rect 21968 14016 21974 14068
rect 22922 14056 22928 14068
rect 22883 14028 22928 14056
rect 22922 14016 22928 14028
rect 22980 14056 22986 14068
rect 23382 14056 23388 14068
rect 22980 14028 23388 14056
rect 22980 14016 22986 14028
rect 23382 14016 23388 14028
rect 23440 14016 23446 14068
rect 24581 14059 24639 14065
rect 24581 14025 24593 14059
rect 24627 14056 24639 14059
rect 24670 14056 24676 14068
rect 24627 14028 24676 14056
rect 24627 14025 24639 14028
rect 24581 14019 24639 14025
rect 24670 14016 24676 14028
rect 24728 14016 24734 14068
rect 24762 14016 24768 14068
rect 24820 14056 24826 14068
rect 24857 14059 24915 14065
rect 24857 14056 24869 14059
rect 24820 14028 24869 14056
rect 24820 14016 24826 14028
rect 24857 14025 24869 14028
rect 24903 14025 24915 14059
rect 24857 14019 24915 14025
rect 25406 14016 25412 14068
rect 25464 14056 25470 14068
rect 25547 14059 25605 14065
rect 25547 14056 25559 14059
rect 25464 14028 25559 14056
rect 25464 14016 25470 14028
rect 25547 14025 25559 14028
rect 25593 14025 25605 14059
rect 25547 14019 25605 14025
rect 12526 13948 12532 14000
rect 12584 13988 12590 14000
rect 12584 13960 14412 13988
rect 12584 13948 12590 13960
rect 14384 13932 14412 13960
rect 15286 13948 15292 14000
rect 15344 13988 15350 14000
rect 15344 13960 16252 13988
rect 15344 13948 15350 13960
rect 16224 13932 16252 13960
rect 18322 13948 18328 14000
rect 18380 13988 18386 14000
rect 20070 13988 20076 14000
rect 18380 13960 20076 13988
rect 18380 13948 18386 13960
rect 20070 13948 20076 13960
rect 20128 13948 20134 14000
rect 21634 13988 21640 14000
rect 21008 13960 21640 13988
rect 12437 13923 12495 13929
rect 12437 13920 12449 13923
rect 11808 13892 12449 13920
rect 10229 13883 10287 13889
rect 12437 13889 12449 13892
rect 12483 13889 12495 13923
rect 14274 13920 14280 13932
rect 14235 13892 14280 13920
rect 12437 13883 12495 13889
rect 14274 13880 14280 13892
rect 14332 13880 14338 13932
rect 14366 13880 14372 13932
rect 14424 13920 14430 13932
rect 14921 13923 14979 13929
rect 14921 13920 14933 13923
rect 14424 13892 14933 13920
rect 14424 13880 14430 13892
rect 14921 13889 14933 13892
rect 14967 13920 14979 13923
rect 15654 13920 15660 13932
rect 14967 13892 15660 13920
rect 14967 13889 14979 13892
rect 14921 13883 14979 13889
rect 15654 13880 15660 13892
rect 15712 13880 15718 13932
rect 16206 13920 16212 13932
rect 16119 13892 16212 13920
rect 16206 13880 16212 13892
rect 16264 13880 16270 13932
rect 16482 13920 16488 13932
rect 16443 13892 16488 13920
rect 16482 13880 16488 13892
rect 16540 13880 16546 13932
rect 18601 13923 18659 13929
rect 18601 13889 18613 13923
rect 18647 13920 18659 13923
rect 18782 13920 18788 13932
rect 18647 13892 18788 13920
rect 18647 13889 18659 13892
rect 18601 13883 18659 13889
rect 18782 13880 18788 13892
rect 18840 13880 18846 13932
rect 20714 13880 20720 13932
rect 20772 13920 20778 13932
rect 21008 13929 21036 13960
rect 21634 13948 21640 13960
rect 21692 13948 21698 14000
rect 22373 13991 22431 13997
rect 22373 13957 22385 13991
rect 22419 13988 22431 13991
rect 23106 13988 23112 14000
rect 22419 13960 23112 13988
rect 22419 13957 22431 13960
rect 22373 13951 22431 13957
rect 23106 13948 23112 13960
rect 23164 13948 23170 14000
rect 20993 13923 21051 13929
rect 20993 13920 21005 13923
rect 20772 13892 21005 13920
rect 20772 13880 20778 13892
rect 20993 13889 21005 13892
rect 21039 13889 21051 13923
rect 20993 13883 21051 13889
rect 22646 13880 22652 13932
rect 22704 13920 22710 13932
rect 23014 13920 23020 13932
rect 22704 13892 23020 13920
rect 22704 13880 22710 13892
rect 23014 13880 23020 13892
rect 23072 13880 23078 13932
rect 23474 13880 23480 13932
rect 23532 13920 23538 13932
rect 23661 13923 23719 13929
rect 23661 13920 23673 13923
rect 23532 13892 23673 13920
rect 23532 13880 23538 13892
rect 23661 13889 23673 13892
rect 23707 13889 23719 13923
rect 23661 13883 23719 13889
rect 11517 13855 11575 13861
rect 11517 13821 11529 13855
rect 11563 13852 11575 13855
rect 11790 13852 11796 13864
rect 11563 13824 11796 13852
rect 11563 13821 11575 13824
rect 11517 13815 11575 13821
rect 11790 13812 11796 13824
rect 11848 13812 11854 13864
rect 21637 13855 21695 13861
rect 21637 13821 21649 13855
rect 21683 13852 21695 13855
rect 22002 13852 22008 13864
rect 21683 13824 22008 13852
rect 21683 13821 21695 13824
rect 21637 13815 21695 13821
rect 22002 13812 22008 13824
rect 22060 13812 22066 13864
rect 22370 13812 22376 13864
rect 22428 13852 22434 13864
rect 22465 13855 22523 13861
rect 22465 13852 22477 13855
rect 22428 13824 22477 13852
rect 22428 13812 22434 13824
rect 22465 13821 22477 13824
rect 22511 13821 22523 13855
rect 22465 13815 22523 13821
rect 25222 13812 25228 13864
rect 25280 13852 25286 13864
rect 25444 13855 25502 13861
rect 25444 13852 25456 13855
rect 25280 13824 25456 13852
rect 25280 13812 25286 13824
rect 25444 13821 25456 13824
rect 25490 13852 25502 13855
rect 25869 13855 25927 13861
rect 25869 13852 25881 13855
rect 25490 13824 25881 13852
rect 25490 13821 25502 13824
rect 25444 13815 25502 13821
rect 25869 13821 25881 13824
rect 25915 13821 25927 13855
rect 25869 13815 25927 13821
rect 9950 13784 9956 13796
rect 9416 13756 9956 13784
rect 8757 13747 8815 13753
rect 3849 13688 5396 13716
rect 5442 13676 5448 13728
rect 5500 13716 5506 13728
rect 6181 13719 6239 13725
rect 6181 13716 6193 13719
rect 5500 13688 6193 13716
rect 5500 13676 5506 13688
rect 6181 13685 6193 13688
rect 6227 13716 6239 13719
rect 6270 13716 6276 13728
rect 6227 13688 6276 13716
rect 6227 13685 6239 13688
rect 6181 13679 6239 13685
rect 6270 13676 6276 13688
rect 6328 13676 6334 13728
rect 7745 13719 7803 13725
rect 7745 13685 7757 13719
rect 7791 13716 7803 13719
rect 8389 13719 8447 13725
rect 8389 13716 8401 13719
rect 7791 13688 8401 13716
rect 7791 13685 7803 13688
rect 7745 13679 7803 13685
rect 8389 13685 8401 13688
rect 8435 13716 8447 13719
rect 8772 13716 8800 13747
rect 9950 13744 9956 13756
rect 10008 13744 10014 13796
rect 10042 13744 10048 13796
rect 10100 13784 10106 13796
rect 10321 13787 10379 13793
rect 10321 13784 10333 13787
rect 10100 13756 10333 13784
rect 10100 13744 10106 13756
rect 10321 13753 10333 13756
rect 10367 13784 10379 13787
rect 10686 13784 10692 13796
rect 10367 13756 10692 13784
rect 10367 13753 10379 13756
rect 10321 13747 10379 13753
rect 10686 13744 10692 13756
rect 10744 13744 10750 13796
rect 10873 13787 10931 13793
rect 10873 13753 10885 13787
rect 10919 13753 10931 13787
rect 12758 13787 12816 13793
rect 12758 13784 12770 13787
rect 10873 13747 10931 13753
rect 12176 13756 12770 13784
rect 8435 13688 8800 13716
rect 9968 13716 9996 13744
rect 10888 13716 10916 13747
rect 9968 13688 10916 13716
rect 8435 13685 8447 13688
rect 8389 13679 8447 13685
rect 11882 13676 11888 13728
rect 11940 13716 11946 13728
rect 12176 13725 12204 13756
rect 12758 13753 12770 13756
rect 12804 13753 12816 13787
rect 12758 13747 12816 13753
rect 14369 13787 14427 13793
rect 14369 13753 14381 13787
rect 14415 13753 14427 13787
rect 14369 13747 14427 13753
rect 16025 13787 16083 13793
rect 16025 13753 16037 13787
rect 16071 13784 16083 13787
rect 16301 13787 16359 13793
rect 16301 13784 16313 13787
rect 16071 13756 16313 13784
rect 16071 13753 16083 13756
rect 16025 13747 16083 13753
rect 16301 13753 16313 13756
rect 16347 13784 16359 13787
rect 16574 13784 16580 13796
rect 16347 13756 16580 13784
rect 16347 13753 16359 13756
rect 16301 13747 16359 13753
rect 12161 13719 12219 13725
rect 12161 13716 12173 13719
rect 11940 13688 12173 13716
rect 11940 13676 11946 13688
rect 12161 13685 12173 13688
rect 12207 13685 12219 13719
rect 12161 13679 12219 13685
rect 13170 13676 13176 13728
rect 13228 13716 13234 13728
rect 13630 13716 13636 13728
rect 13228 13688 13636 13716
rect 13228 13676 13234 13688
rect 13630 13676 13636 13688
rect 13688 13716 13694 13728
rect 14001 13719 14059 13725
rect 14001 13716 14013 13719
rect 13688 13688 14013 13716
rect 13688 13676 13694 13688
rect 14001 13685 14013 13688
rect 14047 13716 14059 13719
rect 14384 13716 14412 13747
rect 16574 13744 16580 13756
rect 16632 13744 16638 13796
rect 18922 13787 18980 13793
rect 18922 13784 18934 13787
rect 18432 13756 18934 13784
rect 14047 13688 14412 13716
rect 14047 13685 14059 13688
rect 14001 13679 14059 13685
rect 17402 13676 17408 13728
rect 17460 13716 17466 13728
rect 17586 13716 17592 13728
rect 17460 13688 17592 13716
rect 17460 13676 17466 13688
rect 17586 13676 17592 13688
rect 17644 13676 17650 13728
rect 18138 13676 18144 13728
rect 18196 13716 18202 13728
rect 18432 13725 18460 13756
rect 18922 13753 18934 13756
rect 18968 13753 18980 13787
rect 18922 13747 18980 13753
rect 20441 13787 20499 13793
rect 20441 13753 20453 13787
rect 20487 13784 20499 13787
rect 21082 13784 21088 13796
rect 20487 13756 21088 13784
rect 20487 13753 20499 13756
rect 20441 13747 20499 13753
rect 21082 13744 21088 13756
rect 21140 13744 21146 13796
rect 23982 13787 24040 13793
rect 23982 13753 23994 13787
rect 24028 13753 24040 13787
rect 23982 13747 24040 13753
rect 18417 13719 18475 13725
rect 18417 13716 18429 13719
rect 18196 13688 18429 13716
rect 18196 13676 18202 13688
rect 18417 13685 18429 13688
rect 18463 13685 18475 13719
rect 18417 13679 18475 13685
rect 19058 13676 19064 13728
rect 19116 13716 19122 13728
rect 22649 13719 22707 13725
rect 22649 13716 22661 13719
rect 19116 13688 22661 13716
rect 19116 13676 19122 13688
rect 22649 13685 22661 13688
rect 22695 13685 22707 13719
rect 22649 13679 22707 13685
rect 23290 13676 23296 13728
rect 23348 13716 23354 13728
rect 23385 13719 23443 13725
rect 23385 13716 23397 13719
rect 23348 13688 23397 13716
rect 23348 13676 23354 13688
rect 23385 13685 23397 13688
rect 23431 13716 23443 13719
rect 23997 13716 24025 13747
rect 23431 13688 24025 13716
rect 23431 13685 23443 13688
rect 23385 13679 23443 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1765 13515 1823 13521
rect 1765 13481 1777 13515
rect 1811 13512 1823 13515
rect 2222 13512 2228 13524
rect 1811 13484 2228 13512
rect 1811 13481 1823 13484
rect 1765 13475 1823 13481
rect 2222 13472 2228 13484
rect 2280 13472 2286 13524
rect 2406 13472 2412 13524
rect 2464 13512 2470 13524
rect 2774 13512 2780 13524
rect 2464 13484 2780 13512
rect 2464 13472 2470 13484
rect 2774 13472 2780 13484
rect 2832 13512 2838 13524
rect 3053 13515 3111 13521
rect 3053 13512 3065 13515
rect 2832 13484 3065 13512
rect 2832 13472 2838 13484
rect 3053 13481 3065 13484
rect 3099 13481 3111 13515
rect 3694 13512 3700 13524
rect 3655 13484 3700 13512
rect 3053 13475 3111 13481
rect 3694 13472 3700 13484
rect 3752 13512 3758 13524
rect 4430 13512 4436 13524
rect 3752 13484 4436 13512
rect 3752 13472 3758 13484
rect 4430 13472 4436 13484
rect 4488 13512 4494 13524
rect 5169 13515 5227 13521
rect 5169 13512 5181 13515
rect 4488 13484 5181 13512
rect 4488 13472 4494 13484
rect 5169 13481 5181 13484
rect 5215 13512 5227 13515
rect 5629 13515 5687 13521
rect 5629 13512 5641 13515
rect 5215 13484 5641 13512
rect 5215 13481 5227 13484
rect 5169 13475 5227 13481
rect 5629 13481 5641 13484
rect 5675 13512 5687 13515
rect 6086 13512 6092 13524
rect 5675 13484 6092 13512
rect 5675 13481 5687 13484
rect 5629 13475 5687 13481
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 7285 13515 7343 13521
rect 7285 13481 7297 13515
rect 7331 13512 7343 13515
rect 7650 13512 7656 13524
rect 7331 13484 7656 13512
rect 7331 13481 7343 13484
rect 7285 13475 7343 13481
rect 7650 13472 7656 13484
rect 7708 13472 7714 13524
rect 8294 13512 8300 13524
rect 8255 13484 8300 13512
rect 8294 13472 8300 13484
rect 8352 13472 8358 13524
rect 8570 13472 8576 13524
rect 8628 13512 8634 13524
rect 8941 13515 8999 13521
rect 8941 13512 8953 13515
rect 8628 13484 8953 13512
rect 8628 13472 8634 13484
rect 8941 13481 8953 13484
rect 8987 13481 8999 13515
rect 8941 13475 8999 13481
rect 9493 13515 9551 13521
rect 9493 13481 9505 13515
rect 9539 13512 9551 13515
rect 9674 13512 9680 13524
rect 9539 13484 9680 13512
rect 9539 13481 9551 13484
rect 9493 13475 9551 13481
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 10686 13512 10692 13524
rect 10647 13484 10692 13512
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 11698 13512 11704 13524
rect 11659 13484 11704 13512
rect 11698 13472 11704 13484
rect 11756 13472 11762 13524
rect 11882 13472 11888 13524
rect 11940 13512 11946 13524
rect 12253 13515 12311 13521
rect 12253 13512 12265 13515
rect 11940 13484 12265 13512
rect 11940 13472 11946 13484
rect 12253 13481 12265 13484
rect 12299 13481 12311 13515
rect 12253 13475 12311 13481
rect 12805 13515 12863 13521
rect 12805 13481 12817 13515
rect 12851 13512 12863 13515
rect 13170 13512 13176 13524
rect 12851 13484 13176 13512
rect 12851 13481 12863 13484
rect 12805 13475 12863 13481
rect 13170 13472 13176 13484
rect 13228 13472 13234 13524
rect 13262 13472 13268 13524
rect 13320 13512 13326 13524
rect 13449 13515 13507 13521
rect 13449 13512 13461 13515
rect 13320 13484 13461 13512
rect 13320 13472 13326 13484
rect 13449 13481 13461 13484
rect 13495 13481 13507 13515
rect 13449 13475 13507 13481
rect 14826 13472 14832 13524
rect 14884 13512 14890 13524
rect 15013 13515 15071 13521
rect 15013 13512 15025 13515
rect 14884 13484 15025 13512
rect 14884 13472 14890 13484
rect 15013 13481 15025 13484
rect 15059 13481 15071 13515
rect 16206 13512 16212 13524
rect 16167 13484 16212 13512
rect 15013 13475 15071 13481
rect 16206 13472 16212 13484
rect 16264 13472 16270 13524
rect 16942 13472 16948 13524
rect 17000 13512 17006 13524
rect 18230 13512 18236 13524
rect 17000 13484 18236 13512
rect 17000 13472 17006 13484
rect 18230 13472 18236 13484
rect 18288 13472 18294 13524
rect 19337 13515 19395 13521
rect 19337 13481 19349 13515
rect 19383 13512 19395 13515
rect 19518 13512 19524 13524
rect 19383 13484 19524 13512
rect 19383 13481 19395 13484
rect 19337 13475 19395 13481
rect 19518 13472 19524 13484
rect 19576 13472 19582 13524
rect 21082 13472 21088 13524
rect 21140 13512 21146 13524
rect 21821 13515 21879 13521
rect 21821 13512 21833 13515
rect 21140 13484 21833 13512
rect 21140 13472 21146 13484
rect 21821 13481 21833 13484
rect 21867 13481 21879 13515
rect 24670 13512 24676 13524
rect 24631 13484 24676 13512
rect 21821 13475 21879 13481
rect 24670 13472 24676 13484
rect 24728 13472 24734 13524
rect 25130 13512 25136 13524
rect 25091 13484 25136 13512
rect 25130 13472 25136 13484
rect 25188 13472 25194 13524
rect 1670 13404 1676 13456
rect 1728 13444 1734 13456
rect 1728 13416 2544 13444
rect 1728 13404 1734 13416
rect 1854 13336 1860 13388
rect 1912 13376 1918 13388
rect 2516 13385 2544 13416
rect 2590 13404 2596 13456
rect 2648 13444 2654 13456
rect 2958 13444 2964 13456
rect 2648 13416 2964 13444
rect 2648 13404 2654 13416
rect 2958 13404 2964 13416
rect 3016 13404 3022 13456
rect 6546 13404 6552 13456
rect 6604 13444 6610 13456
rect 6686 13447 6744 13453
rect 6686 13444 6698 13447
rect 6604 13416 6698 13444
rect 6604 13404 6610 13416
rect 6686 13413 6698 13416
rect 6732 13413 6744 13447
rect 6686 13407 6744 13413
rect 7558 13404 7564 13456
rect 7616 13444 7622 13456
rect 9858 13444 9864 13456
rect 7616 13416 8156 13444
rect 9819 13416 9864 13444
rect 7616 13404 7622 13416
rect 1949 13379 2007 13385
rect 1949 13376 1961 13379
rect 1912 13348 1961 13376
rect 1912 13336 1918 13348
rect 1949 13345 1961 13348
rect 1995 13345 2007 13379
rect 1949 13339 2007 13345
rect 2501 13379 2559 13385
rect 2501 13345 2513 13379
rect 2547 13376 2559 13379
rect 2774 13376 2780 13388
rect 2547 13348 2780 13376
rect 2547 13345 2559 13348
rect 2501 13339 2559 13345
rect 2774 13336 2780 13348
rect 2832 13336 2838 13388
rect 4338 13376 4344 13388
rect 4299 13348 4344 13376
rect 4338 13336 4344 13348
rect 4396 13336 4402 13388
rect 4430 13336 4436 13388
rect 4488 13376 4494 13388
rect 4525 13379 4583 13385
rect 4525 13376 4537 13379
rect 4488 13348 4537 13376
rect 4488 13336 4494 13348
rect 4525 13345 4537 13348
rect 4571 13345 4583 13379
rect 4525 13339 4583 13345
rect 4614 13336 4620 13388
rect 4672 13376 4678 13388
rect 8128 13385 8156 13416
rect 9858 13404 9864 13416
rect 9916 13404 9922 13456
rect 9950 13404 9956 13456
rect 10008 13444 10014 13456
rect 10413 13447 10471 13453
rect 10413 13444 10425 13447
rect 10008 13416 10425 13444
rect 10008 13404 10014 13416
rect 10413 13413 10425 13416
rect 10459 13413 10471 13447
rect 10413 13407 10471 13413
rect 13814 13404 13820 13456
rect 13872 13444 13878 13456
rect 13872 13416 13917 13444
rect 13872 13404 13878 13416
rect 16298 13404 16304 13456
rect 16356 13444 16362 13456
rect 16758 13444 16764 13456
rect 16356 13416 16764 13444
rect 16356 13404 16362 13416
rect 16758 13404 16764 13416
rect 16816 13404 16822 13456
rect 16850 13404 16856 13456
rect 16908 13444 16914 13456
rect 16908 13416 16953 13444
rect 16908 13404 16914 13416
rect 17218 13404 17224 13456
rect 17276 13444 17282 13456
rect 17402 13444 17408 13456
rect 17276 13416 17408 13444
rect 17276 13404 17282 13416
rect 17402 13404 17408 13416
rect 17460 13404 17466 13456
rect 17862 13404 17868 13456
rect 17920 13444 17926 13456
rect 18325 13447 18383 13453
rect 18325 13444 18337 13447
rect 17920 13416 18337 13444
rect 17920 13404 17926 13416
rect 18325 13413 18337 13416
rect 18371 13413 18383 13447
rect 18325 13407 18383 13413
rect 18414 13404 18420 13456
rect 18472 13444 18478 13456
rect 18472 13416 18517 13444
rect 18472 13404 18478 13416
rect 18598 13404 18604 13456
rect 18656 13444 18662 13456
rect 21263 13447 21321 13453
rect 18656 13416 21082 13444
rect 18656 13404 18662 13416
rect 4801 13379 4859 13385
rect 4801 13376 4813 13379
rect 4672 13348 4813 13376
rect 4672 13336 4678 13348
rect 4801 13345 4813 13348
rect 4847 13376 4859 13379
rect 7929 13379 7987 13385
rect 7929 13376 7941 13379
rect 4847 13348 7941 13376
rect 4847 13345 4859 13348
rect 4801 13339 4859 13345
rect 7929 13345 7941 13348
rect 7975 13345 7987 13379
rect 7929 13339 7987 13345
rect 8113 13379 8171 13385
rect 8113 13345 8125 13379
rect 8159 13345 8171 13379
rect 15286 13376 15292 13388
rect 15247 13348 15292 13376
rect 8113 13339 8171 13345
rect 15286 13336 15292 13348
rect 15344 13336 15350 13388
rect 19797 13379 19855 13385
rect 19797 13345 19809 13379
rect 19843 13345 19855 13379
rect 21054 13376 21082 13416
rect 21263 13413 21275 13447
rect 21309 13444 21321 13447
rect 21450 13444 21456 13456
rect 21309 13416 21456 13444
rect 21309 13413 21321 13416
rect 21263 13407 21321 13413
rect 21450 13404 21456 13416
rect 21508 13444 21514 13456
rect 23290 13444 23296 13456
rect 21508 13416 23296 13444
rect 21508 13404 21514 13416
rect 23290 13404 23296 13416
rect 23348 13444 23354 13456
rect 23842 13453 23848 13456
rect 23839 13444 23848 13453
rect 23348 13416 23848 13444
rect 23348 13404 23354 13416
rect 23839 13407 23848 13416
rect 23842 13404 23848 13407
rect 23900 13404 23906 13456
rect 23477 13379 23535 13385
rect 21054 13348 21496 13376
rect 19797 13339 19855 13345
rect 2317 13311 2375 13317
rect 2317 13277 2329 13311
rect 2363 13308 2375 13311
rect 3510 13308 3516 13320
rect 2363 13280 3516 13308
rect 2363 13277 2375 13280
rect 2317 13271 2375 13277
rect 3510 13268 3516 13280
rect 3568 13268 3574 13320
rect 6365 13311 6423 13317
rect 6365 13277 6377 13311
rect 6411 13277 6423 13311
rect 6365 13271 6423 13277
rect 3142 13132 3148 13184
rect 3200 13172 3206 13184
rect 3329 13175 3387 13181
rect 3329 13172 3341 13175
rect 3200 13144 3341 13172
rect 3200 13132 3206 13144
rect 3329 13141 3341 13144
rect 3375 13172 3387 13175
rect 3970 13172 3976 13184
rect 3375 13144 3976 13172
rect 3375 13141 3387 13144
rect 3329 13135 3387 13141
rect 3970 13132 3976 13144
rect 4028 13132 4034 13184
rect 6178 13172 6184 13184
rect 6139 13144 6184 13172
rect 6178 13132 6184 13144
rect 6236 13172 6242 13184
rect 6380 13172 6408 13271
rect 6730 13268 6736 13320
rect 6788 13308 6794 13320
rect 8018 13308 8024 13320
rect 6788 13280 8024 13308
rect 6788 13268 6794 13280
rect 8018 13268 8024 13280
rect 8076 13308 8082 13320
rect 8573 13311 8631 13317
rect 8573 13308 8585 13311
rect 8076 13280 8585 13308
rect 8076 13268 8082 13280
rect 8573 13277 8585 13280
rect 8619 13277 8631 13311
rect 8573 13271 8631 13277
rect 9398 13268 9404 13320
rect 9456 13308 9462 13320
rect 9769 13311 9827 13317
rect 9769 13308 9781 13311
rect 9456 13280 9781 13308
rect 9456 13268 9462 13280
rect 9769 13277 9781 13280
rect 9815 13308 9827 13311
rect 10870 13308 10876 13320
rect 9815 13280 10876 13308
rect 9815 13277 9827 13280
rect 9769 13271 9827 13277
rect 10870 13268 10876 13280
rect 10928 13268 10934 13320
rect 11514 13268 11520 13320
rect 11572 13308 11578 13320
rect 11885 13311 11943 13317
rect 11885 13308 11897 13311
rect 11572 13280 11897 13308
rect 11572 13268 11578 13280
rect 11885 13277 11897 13280
rect 11931 13277 11943 13311
rect 11885 13271 11943 13277
rect 12342 13268 12348 13320
rect 12400 13308 12406 13320
rect 13722 13308 13728 13320
rect 12400 13280 13728 13308
rect 12400 13268 12406 13280
rect 13722 13268 13728 13280
rect 13780 13268 13786 13320
rect 13906 13268 13912 13320
rect 13964 13308 13970 13320
rect 14001 13311 14059 13317
rect 14001 13308 14013 13311
rect 13964 13280 14013 13308
rect 13964 13268 13970 13280
rect 14001 13277 14013 13280
rect 14047 13277 14059 13311
rect 14001 13271 14059 13277
rect 16942 13268 16948 13320
rect 17000 13308 17006 13320
rect 17037 13311 17095 13317
rect 17037 13308 17049 13311
rect 17000 13280 17049 13308
rect 17000 13268 17006 13280
rect 17037 13277 17049 13280
rect 17083 13308 17095 13311
rect 17083 13280 18276 13308
rect 17083 13277 17095 13280
rect 17037 13271 17095 13277
rect 14182 13200 14188 13252
rect 14240 13240 14246 13252
rect 15194 13240 15200 13252
rect 14240 13212 15200 13240
rect 14240 13200 14246 13212
rect 15194 13200 15200 13212
rect 15252 13200 15258 13252
rect 15473 13243 15531 13249
rect 15473 13209 15485 13243
rect 15519 13240 15531 13243
rect 17218 13240 17224 13252
rect 15519 13212 17224 13240
rect 15519 13209 15531 13212
rect 15473 13203 15531 13209
rect 17218 13200 17224 13212
rect 17276 13200 17282 13252
rect 18248 13240 18276 13280
rect 18322 13268 18328 13320
rect 18380 13308 18386 13320
rect 19812 13308 19840 13339
rect 20162 13308 20168 13320
rect 18380 13280 20168 13308
rect 18380 13268 18386 13280
rect 20162 13268 20168 13280
rect 20220 13268 20226 13320
rect 20901 13311 20959 13317
rect 20901 13277 20913 13311
rect 20947 13308 20959 13311
rect 20990 13308 20996 13320
rect 20947 13280 20996 13308
rect 20947 13277 20959 13280
rect 20901 13271 20959 13277
rect 20990 13268 20996 13280
rect 21048 13308 21054 13320
rect 21358 13308 21364 13320
rect 21048 13280 21364 13308
rect 21048 13268 21054 13280
rect 21358 13268 21364 13280
rect 21416 13268 21422 13320
rect 21468 13308 21496 13348
rect 23477 13345 23489 13379
rect 23523 13376 23535 13379
rect 23566 13376 23572 13388
rect 23523 13348 23572 13376
rect 23523 13345 23535 13348
rect 23477 13339 23535 13345
rect 23566 13336 23572 13348
rect 23624 13336 23630 13388
rect 23750 13336 23756 13388
rect 23808 13376 23814 13388
rect 25225 13379 25283 13385
rect 25225 13376 25237 13379
rect 23808 13348 25237 13376
rect 23808 13336 23814 13348
rect 25225 13345 25237 13348
rect 25271 13376 25283 13379
rect 25406 13376 25412 13388
rect 25271 13348 25412 13376
rect 25271 13345 25283 13348
rect 25225 13339 25283 13345
rect 25406 13336 25412 13348
rect 25464 13376 25470 13388
rect 27706 13376 27712 13388
rect 25464 13348 27712 13376
rect 25464 13336 25470 13348
rect 27706 13336 27712 13348
rect 27764 13336 27770 13388
rect 21542 13308 21548 13320
rect 21468 13280 21548 13308
rect 21542 13268 21548 13280
rect 21600 13308 21606 13320
rect 22094 13308 22100 13320
rect 21600 13280 22100 13308
rect 21600 13268 21606 13280
rect 22094 13268 22100 13280
rect 22152 13268 22158 13320
rect 18877 13243 18935 13249
rect 18877 13240 18889 13243
rect 18248 13212 18889 13240
rect 18877 13209 18889 13212
rect 18923 13209 18935 13243
rect 18877 13203 18935 13209
rect 19981 13243 20039 13249
rect 19981 13209 19993 13243
rect 20027 13240 20039 13243
rect 23658 13240 23664 13252
rect 20027 13212 23664 13240
rect 20027 13209 20039 13212
rect 19981 13203 20039 13209
rect 6236 13144 6408 13172
rect 6236 13132 6242 13144
rect 7190 13132 7196 13184
rect 7248 13172 7254 13184
rect 12526 13172 12532 13184
rect 7248 13144 12532 13172
rect 7248 13132 7254 13144
rect 12526 13132 12532 13144
rect 12584 13172 12590 13184
rect 13081 13175 13139 13181
rect 13081 13172 13093 13175
rect 12584 13144 13093 13172
rect 12584 13132 12590 13144
rect 13081 13141 13093 13144
rect 13127 13141 13139 13175
rect 15838 13172 15844 13184
rect 15799 13144 15844 13172
rect 13081 13135 13139 13141
rect 15838 13132 15844 13144
rect 15896 13132 15902 13184
rect 18892 13172 18920 13203
rect 23658 13200 23664 13212
rect 23716 13240 23722 13252
rect 24210 13240 24216 13252
rect 23716 13212 24216 13240
rect 23716 13200 23722 13212
rect 24210 13200 24216 13212
rect 24268 13200 24274 13252
rect 20530 13172 20536 13184
rect 18892 13144 20536 13172
rect 20530 13132 20536 13144
rect 20588 13132 20594 13184
rect 20714 13172 20720 13184
rect 20627 13144 20720 13172
rect 20714 13132 20720 13144
rect 20772 13172 20778 13184
rect 21082 13172 21088 13184
rect 20772 13144 21088 13172
rect 20772 13132 20778 13144
rect 21082 13132 21088 13144
rect 21140 13132 21146 13184
rect 22370 13132 22376 13184
rect 22428 13172 22434 13184
rect 22465 13175 22523 13181
rect 22465 13172 22477 13175
rect 22428 13144 22477 13172
rect 22428 13132 22434 13144
rect 22465 13141 22477 13144
rect 22511 13141 22523 13175
rect 22465 13135 22523 13141
rect 24397 13175 24455 13181
rect 24397 13141 24409 13175
rect 24443 13172 24455 13175
rect 24670 13172 24676 13184
rect 24443 13144 24676 13172
rect 24443 13141 24455 13144
rect 24397 13135 24455 13141
rect 24670 13132 24676 13144
rect 24728 13132 24734 13184
rect 25409 13175 25467 13181
rect 25409 13141 25421 13175
rect 25455 13172 25467 13175
rect 25498 13172 25504 13184
rect 25455 13144 25504 13172
rect 25455 13141 25467 13144
rect 25409 13135 25467 13141
rect 25498 13132 25504 13144
rect 25556 13132 25562 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1949 12971 2007 12977
rect 1949 12937 1961 12971
rect 1995 12968 2007 12971
rect 2222 12968 2228 12980
rect 1995 12940 2228 12968
rect 1995 12937 2007 12940
rect 1949 12931 2007 12937
rect 2222 12928 2228 12940
rect 2280 12928 2286 12980
rect 2317 12971 2375 12977
rect 2317 12937 2329 12971
rect 2363 12968 2375 12971
rect 2682 12968 2688 12980
rect 2363 12940 2688 12968
rect 2363 12937 2375 12940
rect 2317 12931 2375 12937
rect 2682 12928 2688 12940
rect 2740 12928 2746 12980
rect 2774 12928 2780 12980
rect 2832 12968 2838 12980
rect 4338 12968 4344 12980
rect 2832 12940 3464 12968
rect 4299 12940 4344 12968
rect 2832 12928 2838 12940
rect 1854 12841 1860 12844
rect 1820 12835 1860 12841
rect 1820 12801 1832 12835
rect 1820 12795 1860 12801
rect 1854 12792 1860 12795
rect 1912 12792 1918 12844
rect 2041 12835 2099 12841
rect 2041 12801 2053 12835
rect 2087 12832 2099 12835
rect 2406 12832 2412 12844
rect 2087 12804 2412 12832
rect 2087 12801 2099 12804
rect 2041 12795 2099 12801
rect 2406 12792 2412 12804
rect 2464 12792 2470 12844
rect 3053 12835 3111 12841
rect 3053 12801 3065 12835
rect 3099 12832 3111 12835
rect 3436 12832 3464 12940
rect 4338 12928 4344 12940
rect 4396 12928 4402 12980
rect 6457 12971 6515 12977
rect 6457 12937 6469 12971
rect 6503 12968 6515 12971
rect 6546 12968 6552 12980
rect 6503 12940 6552 12968
rect 6503 12937 6515 12940
rect 6457 12931 6515 12937
rect 6546 12928 6552 12940
rect 6604 12928 6610 12980
rect 7006 12968 7012 12980
rect 6967 12940 7012 12968
rect 7006 12928 7012 12940
rect 7064 12928 7070 12980
rect 10870 12968 10876 12980
rect 10831 12940 10876 12968
rect 10870 12928 10876 12940
rect 10928 12928 10934 12980
rect 13633 12971 13691 12977
rect 13633 12937 13645 12971
rect 13679 12968 13691 12971
rect 13814 12968 13820 12980
rect 13679 12940 13820 12968
rect 13679 12937 13691 12940
rect 13633 12931 13691 12937
rect 13814 12928 13820 12940
rect 13872 12928 13878 12980
rect 16758 12928 16764 12980
rect 16816 12968 16822 12980
rect 17221 12971 17279 12977
rect 17221 12968 17233 12971
rect 16816 12940 17233 12968
rect 16816 12928 16822 12940
rect 17221 12937 17233 12940
rect 17267 12937 17279 12971
rect 17862 12968 17868 12980
rect 17823 12940 17868 12968
rect 17221 12931 17279 12937
rect 17862 12928 17868 12940
rect 17920 12928 17926 12980
rect 18325 12971 18383 12977
rect 18325 12937 18337 12971
rect 18371 12968 18383 12971
rect 18414 12968 18420 12980
rect 18371 12940 18420 12968
rect 18371 12937 18383 12940
rect 18325 12931 18383 12937
rect 3510 12860 3516 12912
rect 3568 12900 3574 12912
rect 4246 12900 4252 12912
rect 3568 12872 4252 12900
rect 3568 12860 3574 12872
rect 4246 12860 4252 12872
rect 4304 12900 4310 12912
rect 4617 12903 4675 12909
rect 4617 12900 4629 12903
rect 4304 12872 4629 12900
rect 4304 12860 4310 12872
rect 4617 12869 4629 12872
rect 4663 12869 4675 12903
rect 8202 12900 8208 12912
rect 4617 12863 4675 12869
rect 5552 12872 8208 12900
rect 5442 12832 5448 12844
rect 3099 12804 3280 12832
rect 3436 12804 5448 12832
rect 3099 12801 3111 12804
rect 3053 12795 3111 12801
rect 1673 12767 1731 12773
rect 1673 12733 1685 12767
rect 1719 12764 1731 12767
rect 3142 12764 3148 12776
rect 1719 12736 3148 12764
rect 1719 12733 1731 12736
rect 1673 12727 1731 12733
rect 3142 12724 3148 12736
rect 3200 12724 3206 12776
rect 3252 12773 3280 12804
rect 5442 12792 5448 12804
rect 5500 12792 5506 12844
rect 3237 12767 3295 12773
rect 3237 12733 3249 12767
rect 3283 12764 3295 12767
rect 3510 12764 3516 12776
rect 3283 12736 3516 12764
rect 3283 12733 3295 12736
rect 3237 12727 3295 12733
rect 3510 12724 3516 12736
rect 3568 12724 3574 12776
rect 3694 12764 3700 12776
rect 3655 12736 3700 12764
rect 3694 12724 3700 12736
rect 3752 12724 3758 12776
rect 5077 12767 5135 12773
rect 5077 12733 5089 12767
rect 5123 12764 5135 12767
rect 5353 12767 5411 12773
rect 5353 12764 5365 12767
rect 5123 12736 5365 12764
rect 5123 12733 5135 12736
rect 5077 12727 5135 12733
rect 5353 12733 5365 12736
rect 5399 12764 5411 12767
rect 5552 12764 5580 12872
rect 8202 12860 8208 12872
rect 8260 12900 8266 12912
rect 8478 12900 8484 12912
rect 8260 12872 8484 12900
rect 8260 12860 8266 12872
rect 8478 12860 8484 12872
rect 8536 12860 8542 12912
rect 8570 12860 8576 12912
rect 8628 12900 8634 12912
rect 10134 12900 10140 12912
rect 8628 12872 10140 12900
rect 8628 12860 8634 12872
rect 10134 12860 10140 12872
rect 10192 12900 10198 12912
rect 10505 12903 10563 12909
rect 10505 12900 10517 12903
rect 10192 12872 10517 12900
rect 10192 12860 10198 12872
rect 10505 12869 10517 12872
rect 10551 12869 10563 12903
rect 10505 12863 10563 12869
rect 11882 12860 11888 12912
rect 11940 12900 11946 12912
rect 15473 12903 15531 12909
rect 15473 12900 15485 12903
rect 11940 12872 15485 12900
rect 11940 12860 11946 12872
rect 15473 12869 15485 12872
rect 15519 12900 15531 12903
rect 15654 12900 15660 12912
rect 15519 12872 15660 12900
rect 15519 12869 15531 12872
rect 15473 12863 15531 12869
rect 15654 12860 15660 12872
rect 15712 12860 15718 12912
rect 16574 12900 16580 12912
rect 16487 12872 16580 12900
rect 16574 12860 16580 12872
rect 16632 12900 16638 12912
rect 18340 12900 18368 12931
rect 18414 12928 18420 12940
rect 18472 12928 18478 12980
rect 20162 12968 20168 12980
rect 20123 12940 20168 12968
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 21450 12968 21456 12980
rect 20732 12940 21456 12968
rect 20732 12900 20760 12940
rect 21450 12928 21456 12940
rect 21508 12968 21514 12980
rect 21729 12971 21787 12977
rect 21729 12968 21741 12971
rect 21508 12940 21741 12968
rect 21508 12928 21514 12940
rect 21729 12937 21741 12940
rect 21775 12937 21787 12971
rect 21729 12931 21787 12937
rect 23477 12971 23535 12977
rect 23477 12937 23489 12971
rect 23523 12968 23535 12971
rect 23566 12968 23572 12980
rect 23523 12940 23572 12968
rect 23523 12937 23535 12940
rect 23477 12931 23535 12937
rect 23566 12928 23572 12940
rect 23624 12928 23630 12980
rect 23842 12968 23848 12980
rect 23803 12940 23848 12968
rect 23842 12928 23848 12940
rect 23900 12928 23906 12980
rect 25406 12968 25412 12980
rect 25367 12940 25412 12968
rect 25406 12928 25412 12940
rect 25464 12928 25470 12980
rect 22097 12903 22155 12909
rect 22097 12900 22109 12903
rect 16632 12872 18368 12900
rect 19306 12872 20760 12900
rect 20824 12872 22109 12900
rect 16632 12860 16638 12872
rect 5905 12835 5963 12841
rect 5905 12801 5917 12835
rect 5951 12832 5963 12835
rect 6178 12832 6184 12844
rect 5951 12804 6184 12832
rect 5951 12801 5963 12804
rect 5905 12795 5963 12801
rect 6178 12792 6184 12804
rect 6236 12792 6242 12844
rect 6546 12792 6552 12844
rect 6604 12832 6610 12844
rect 7929 12835 7987 12841
rect 7929 12832 7941 12835
rect 6604 12804 7941 12832
rect 6604 12792 6610 12804
rect 7929 12801 7941 12804
rect 7975 12801 7987 12835
rect 7929 12795 7987 12801
rect 5399 12736 5580 12764
rect 5721 12767 5779 12773
rect 5399 12733 5411 12736
rect 5353 12727 5411 12733
rect 5721 12733 5733 12767
rect 5767 12764 5779 12767
rect 6086 12764 6092 12776
rect 5767 12736 6092 12764
rect 5767 12733 5779 12736
rect 5721 12727 5779 12733
rect 6086 12724 6092 12736
rect 6144 12724 6150 12776
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12733 6883 12767
rect 7944 12764 7972 12795
rect 8018 12792 8024 12844
rect 8076 12832 8082 12844
rect 8113 12835 8171 12841
rect 8113 12832 8125 12835
rect 8076 12804 8125 12832
rect 8076 12792 8082 12804
rect 8113 12801 8125 12804
rect 8159 12801 8171 12835
rect 8113 12795 8171 12801
rect 9953 12835 10011 12841
rect 9953 12801 9965 12835
rect 9999 12832 10011 12835
rect 10962 12832 10968 12844
rect 9999 12804 10968 12832
rect 9999 12801 10011 12804
rect 9953 12795 10011 12801
rect 10962 12792 10968 12804
rect 11020 12792 11026 12844
rect 12526 12832 12532 12844
rect 12487 12804 12532 12832
rect 12526 12792 12532 12804
rect 12584 12792 12590 12844
rect 15102 12832 15108 12844
rect 15063 12804 15108 12832
rect 15102 12792 15108 12804
rect 15160 12792 15166 12844
rect 17770 12832 17776 12844
rect 15580 12804 17776 12832
rect 9033 12767 9091 12773
rect 7944 12736 8477 12764
rect 6825 12727 6883 12733
rect 6840 12696 6868 12727
rect 8036 12708 8064 12736
rect 7006 12696 7012 12708
rect 4126 12668 7012 12696
rect 3326 12628 3332 12640
rect 3287 12600 3332 12628
rect 3326 12588 3332 12600
rect 3384 12588 3390 12640
rect 3510 12588 3516 12640
rect 3568 12628 3574 12640
rect 4126 12628 4154 12668
rect 7006 12656 7012 12668
rect 7064 12656 7070 12708
rect 8018 12656 8024 12708
rect 8076 12656 8082 12708
rect 8449 12705 8477 12736
rect 9033 12733 9045 12767
rect 9079 12733 9091 12767
rect 9033 12727 9091 12733
rect 14093 12767 14151 12773
rect 14093 12733 14105 12767
rect 14139 12733 14151 12767
rect 14550 12764 14556 12776
rect 14511 12736 14556 12764
rect 14093 12727 14151 12733
rect 8435 12699 8493 12705
rect 8435 12665 8447 12699
rect 8481 12665 8493 12699
rect 9048 12696 9076 12727
rect 9401 12699 9459 12705
rect 9401 12696 9413 12699
rect 9048 12668 9413 12696
rect 8435 12659 8493 12665
rect 9401 12665 9413 12668
rect 9447 12696 9459 12699
rect 10042 12696 10048 12708
rect 9447 12668 10048 12696
rect 9447 12665 9459 12668
rect 9401 12659 9459 12665
rect 10042 12656 10048 12668
rect 10100 12656 10106 12708
rect 12621 12699 12679 12705
rect 12621 12665 12633 12699
rect 12667 12696 12679 12699
rect 12802 12696 12808 12708
rect 12667 12668 12808 12696
rect 12667 12665 12679 12668
rect 12621 12659 12679 12665
rect 12802 12656 12808 12668
rect 12860 12656 12866 12708
rect 13173 12699 13231 12705
rect 13173 12665 13185 12699
rect 13219 12696 13231 12699
rect 13446 12696 13452 12708
rect 13219 12668 13452 12696
rect 13219 12665 13231 12668
rect 13173 12659 13231 12665
rect 13446 12656 13452 12668
rect 13504 12656 13510 12708
rect 13906 12696 13912 12708
rect 13867 12668 13912 12696
rect 13906 12656 13912 12668
rect 13964 12696 13970 12708
rect 14108 12696 14136 12727
rect 14550 12724 14556 12736
rect 14608 12764 14614 12776
rect 15580 12764 15608 12804
rect 17770 12792 17776 12804
rect 17828 12792 17834 12844
rect 14608 12736 15608 12764
rect 15657 12767 15715 12773
rect 14608 12724 14614 12736
rect 15657 12733 15669 12767
rect 15703 12764 15715 12767
rect 15838 12764 15844 12776
rect 15703 12736 15844 12764
rect 15703 12733 15715 12736
rect 15657 12727 15715 12733
rect 15838 12724 15844 12736
rect 15896 12764 15902 12776
rect 17678 12764 17684 12776
rect 15896 12736 17684 12764
rect 15896 12724 15902 12736
rect 17678 12724 17684 12736
rect 17736 12724 17742 12776
rect 18966 12764 18972 12776
rect 18927 12736 18972 12764
rect 18966 12724 18972 12736
rect 19024 12724 19030 12776
rect 14458 12696 14464 12708
rect 13964 12668 14464 12696
rect 13964 12656 13970 12668
rect 14458 12656 14464 12668
rect 14516 12656 14522 12708
rect 14826 12696 14832 12708
rect 14787 12668 14832 12696
rect 14826 12656 14832 12668
rect 14884 12656 14890 12708
rect 15978 12699 16036 12705
rect 15978 12665 15990 12699
rect 16024 12696 16036 12699
rect 18138 12696 18144 12708
rect 16024 12668 18144 12696
rect 16024 12665 16036 12668
rect 15978 12659 16036 12665
rect 7558 12628 7564 12640
rect 3568 12600 4154 12628
rect 7519 12600 7564 12628
rect 3568 12588 3574 12600
rect 7558 12588 7564 12600
rect 7616 12588 7622 12640
rect 9769 12631 9827 12637
rect 9769 12597 9781 12631
rect 9815 12628 9827 12631
rect 9858 12628 9864 12640
rect 9815 12600 9864 12628
rect 9815 12597 9827 12600
rect 9769 12591 9827 12597
rect 9858 12588 9864 12600
rect 9916 12588 9922 12640
rect 11514 12628 11520 12640
rect 11475 12600 11520 12628
rect 11514 12588 11520 12600
rect 11572 12588 11578 12640
rect 11698 12588 11704 12640
rect 11756 12628 11762 12640
rect 11882 12628 11888 12640
rect 11756 12600 11888 12628
rect 11756 12588 11762 12600
rect 11882 12588 11888 12600
rect 11940 12588 11946 12640
rect 15654 12588 15660 12640
rect 15712 12628 15718 12640
rect 15993 12628 16021 12659
rect 18138 12656 18144 12668
rect 18196 12696 18202 12708
rect 19306 12705 19334 12872
rect 20824 12844 20852 12872
rect 22097 12869 22109 12872
rect 22143 12869 22155 12903
rect 22097 12863 22155 12869
rect 22186 12860 22192 12912
rect 22244 12900 22250 12912
rect 22370 12900 22376 12912
rect 22244 12872 22376 12900
rect 22244 12860 22250 12872
rect 22370 12860 22376 12872
rect 22428 12860 22434 12912
rect 24946 12900 24952 12912
rect 24907 12872 24952 12900
rect 24946 12860 24952 12872
rect 25004 12860 25010 12912
rect 20806 12832 20812 12844
rect 20767 12804 20812 12832
rect 20806 12792 20812 12804
rect 20864 12792 20870 12844
rect 21082 12832 21088 12844
rect 21043 12804 21088 12832
rect 21082 12792 21088 12804
rect 21140 12792 21146 12844
rect 24397 12835 24455 12841
rect 24397 12801 24409 12835
rect 24443 12832 24455 12835
rect 25130 12832 25136 12844
rect 24443 12804 25136 12832
rect 24443 12801 24455 12804
rect 24397 12795 24455 12801
rect 25130 12792 25136 12804
rect 25188 12792 25194 12844
rect 22348 12767 22406 12773
rect 22348 12733 22360 12767
rect 22394 12764 22406 12767
rect 22394 12736 22876 12764
rect 22394 12733 22406 12736
rect 22348 12727 22406 12733
rect 18785 12699 18843 12705
rect 18785 12696 18797 12699
rect 18196 12668 18797 12696
rect 18196 12656 18202 12668
rect 18785 12665 18797 12668
rect 18831 12696 18843 12699
rect 19290 12699 19348 12705
rect 19290 12696 19302 12699
rect 18831 12668 19302 12696
rect 18831 12665 18843 12668
rect 18785 12659 18843 12665
rect 19290 12665 19302 12668
rect 19336 12665 19348 12699
rect 20533 12699 20591 12705
rect 20533 12696 20545 12699
rect 19290 12659 19348 12665
rect 19904 12668 20545 12696
rect 16850 12628 16856 12640
rect 15712 12600 16021 12628
rect 16811 12600 16856 12628
rect 15712 12588 15718 12600
rect 16850 12588 16856 12600
rect 16908 12588 16914 12640
rect 17310 12588 17316 12640
rect 17368 12628 17374 12640
rect 18690 12628 18696 12640
rect 17368 12600 18696 12628
rect 17368 12588 17374 12600
rect 18690 12588 18696 12600
rect 18748 12588 18754 12640
rect 19518 12588 19524 12640
rect 19576 12628 19582 12640
rect 19904 12637 19932 12668
rect 20533 12665 20545 12668
rect 20579 12665 20591 12699
rect 20533 12659 20591 12665
rect 20901 12699 20959 12705
rect 20901 12665 20913 12699
rect 20947 12665 20959 12699
rect 20901 12659 20959 12665
rect 19889 12631 19947 12637
rect 19889 12628 19901 12631
rect 19576 12600 19901 12628
rect 19576 12588 19582 12600
rect 19889 12597 19901 12600
rect 19935 12597 19947 12631
rect 20548 12628 20576 12659
rect 20916 12628 20944 12659
rect 20548 12600 20944 12628
rect 19889 12591 19947 12597
rect 21818 12588 21824 12640
rect 21876 12628 21882 12640
rect 22848 12637 22876 12736
rect 24486 12656 24492 12708
rect 24544 12696 24550 12708
rect 24670 12696 24676 12708
rect 24544 12668 24676 12696
rect 24544 12656 24550 12668
rect 24670 12656 24676 12668
rect 24728 12656 24734 12708
rect 22419 12631 22477 12637
rect 22419 12628 22431 12631
rect 21876 12600 22431 12628
rect 21876 12588 21882 12600
rect 22419 12597 22431 12600
rect 22465 12597 22477 12631
rect 22419 12591 22477 12597
rect 22833 12631 22891 12637
rect 22833 12597 22845 12631
rect 22879 12628 22891 12631
rect 23106 12628 23112 12640
rect 22879 12600 23112 12628
rect 22879 12597 22891 12600
rect 22833 12591 22891 12597
rect 23106 12588 23112 12600
rect 23164 12588 23170 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1946 12384 1952 12436
rect 2004 12424 2010 12436
rect 3237 12427 3295 12433
rect 3237 12424 3249 12427
rect 2004 12396 3249 12424
rect 2004 12384 2010 12396
rect 3237 12393 3249 12396
rect 3283 12424 3295 12427
rect 3326 12424 3332 12436
rect 3283 12396 3332 12424
rect 3283 12393 3295 12396
rect 3237 12387 3295 12393
rect 3326 12384 3332 12396
rect 3384 12384 3390 12436
rect 3602 12384 3608 12436
rect 3660 12424 3666 12436
rect 4709 12427 4767 12433
rect 4709 12424 4721 12427
rect 3660 12396 4721 12424
rect 3660 12384 3666 12396
rect 4709 12393 4721 12396
rect 4755 12393 4767 12427
rect 4709 12387 4767 12393
rect 5074 12384 5080 12436
rect 5132 12424 5138 12436
rect 7006 12424 7012 12436
rect 5132 12396 6729 12424
rect 6967 12396 7012 12424
rect 5132 12384 5138 12396
rect 2133 12359 2191 12365
rect 2133 12325 2145 12359
rect 2179 12356 2191 12359
rect 2222 12356 2228 12368
rect 2179 12328 2228 12356
rect 2179 12325 2191 12328
rect 2133 12319 2191 12325
rect 2222 12316 2228 12328
rect 2280 12316 2286 12368
rect 3786 12316 3792 12368
rect 3844 12356 3850 12368
rect 3970 12356 3976 12368
rect 3844 12328 3976 12356
rect 3844 12316 3850 12328
rect 3970 12316 3976 12328
rect 4028 12356 4034 12368
rect 4065 12359 4123 12365
rect 4065 12356 4077 12359
rect 4028 12328 4077 12356
rect 4028 12316 4034 12328
rect 4065 12325 4077 12328
rect 4111 12356 4123 12359
rect 5534 12356 5540 12368
rect 4111 12328 5540 12356
rect 4111 12325 4123 12328
rect 4065 12319 4123 12325
rect 5534 12316 5540 12328
rect 5592 12356 5598 12368
rect 5721 12359 5779 12365
rect 5721 12356 5733 12359
rect 5592 12328 5733 12356
rect 5592 12316 5598 12328
rect 5721 12325 5733 12328
rect 5767 12325 5779 12359
rect 6701 12356 6729 12396
rect 7006 12384 7012 12396
rect 7064 12384 7070 12436
rect 8018 12424 8024 12436
rect 7979 12396 8024 12424
rect 8018 12384 8024 12396
rect 8076 12384 8082 12436
rect 9306 12384 9312 12436
rect 9364 12424 9370 12436
rect 9401 12427 9459 12433
rect 9401 12424 9413 12427
rect 9364 12396 9413 12424
rect 9364 12384 9370 12396
rect 9401 12393 9413 12396
rect 9447 12393 9459 12427
rect 9401 12387 9459 12393
rect 10781 12427 10839 12433
rect 10781 12393 10793 12427
rect 10827 12424 10839 12427
rect 10962 12424 10968 12436
rect 10827 12396 10968 12424
rect 10827 12393 10839 12396
rect 10781 12387 10839 12393
rect 7469 12359 7527 12365
rect 7469 12356 7481 12359
rect 6701 12328 7481 12356
rect 5721 12319 5779 12325
rect 7469 12325 7481 12328
rect 7515 12356 7527 12359
rect 7742 12356 7748 12368
rect 7515 12328 7748 12356
rect 7515 12325 7527 12328
rect 7469 12319 7527 12325
rect 7742 12316 7748 12328
rect 7800 12316 7806 12368
rect 9416 12356 9444 12387
rect 10962 12384 10968 12396
rect 11020 12384 11026 12436
rect 11514 12424 11520 12436
rect 11475 12396 11520 12424
rect 11514 12384 11520 12396
rect 11572 12384 11578 12436
rect 13722 12384 13728 12436
rect 13780 12424 13786 12436
rect 14461 12427 14519 12433
rect 14461 12424 14473 12427
rect 13780 12396 14473 12424
rect 13780 12384 13786 12396
rect 14461 12393 14473 12396
rect 14507 12393 14519 12427
rect 17678 12424 17684 12436
rect 17639 12396 17684 12424
rect 14461 12387 14519 12393
rect 17678 12384 17684 12396
rect 17736 12384 17742 12436
rect 21039 12427 21097 12433
rect 21039 12424 21051 12427
rect 19306 12396 21051 12424
rect 9769 12359 9827 12365
rect 9769 12356 9781 12359
rect 9416 12328 9781 12356
rect 9769 12325 9781 12328
rect 9815 12325 9827 12359
rect 9769 12319 9827 12325
rect 9858 12316 9864 12368
rect 9916 12356 9922 12368
rect 10226 12356 10232 12368
rect 9916 12328 10232 12356
rect 9916 12316 9922 12328
rect 10226 12316 10232 12328
rect 10284 12316 10290 12368
rect 12989 12359 13047 12365
rect 12989 12325 13001 12359
rect 13035 12356 13047 12359
rect 13630 12356 13636 12368
rect 13035 12328 13636 12356
rect 13035 12325 13047 12328
rect 12989 12319 13047 12325
rect 13630 12316 13636 12328
rect 13688 12316 13694 12368
rect 14185 12359 14243 12365
rect 14185 12325 14197 12359
rect 14231 12356 14243 12359
rect 14550 12356 14556 12368
rect 14231 12328 14556 12356
rect 14231 12325 14243 12328
rect 14185 12319 14243 12325
rect 14550 12316 14556 12328
rect 14608 12316 14614 12368
rect 15654 12316 15660 12368
rect 15712 12356 15718 12368
rect 16162 12359 16220 12365
rect 16162 12356 16174 12359
rect 15712 12328 16174 12356
rect 15712 12316 15718 12328
rect 16162 12325 16174 12328
rect 16208 12325 16220 12359
rect 19306 12356 19334 12396
rect 21039 12393 21051 12396
rect 21085 12393 21097 12427
rect 21358 12424 21364 12436
rect 21319 12396 21364 12424
rect 21039 12387 21097 12393
rect 21358 12384 21364 12396
rect 21416 12384 21422 12436
rect 24397 12427 24455 12433
rect 24397 12393 24409 12427
rect 24443 12424 24455 12427
rect 24486 12424 24492 12436
rect 24443 12396 24492 12424
rect 24443 12393 24455 12396
rect 24397 12387 24455 12393
rect 24486 12384 24492 12396
rect 24544 12384 24550 12436
rect 16162 12319 16220 12325
rect 16316 12328 19334 12356
rect 19429 12359 19487 12365
rect 1762 12248 1768 12300
rect 1820 12288 1826 12300
rect 2317 12291 2375 12297
rect 2317 12288 2329 12291
rect 1820 12260 2329 12288
rect 1820 12248 1826 12260
rect 2317 12257 2329 12260
rect 2363 12257 2375 12291
rect 2317 12251 2375 12257
rect 3694 12248 3700 12300
rect 3752 12288 3758 12300
rect 4982 12288 4988 12300
rect 3752 12260 4988 12288
rect 3752 12248 3758 12260
rect 2498 12180 2504 12232
rect 2556 12220 2562 12232
rect 4448 12229 4476 12260
rect 4982 12248 4988 12260
rect 5040 12248 5046 12300
rect 5350 12288 5356 12300
rect 5311 12260 5356 12288
rect 5350 12248 5356 12260
rect 5408 12248 5414 12300
rect 5994 12288 6000 12300
rect 5955 12260 6000 12288
rect 5994 12248 6000 12260
rect 6052 12248 6058 12300
rect 6086 12248 6092 12300
rect 6144 12288 6150 12300
rect 6457 12291 6515 12297
rect 6457 12288 6469 12291
rect 6144 12260 6469 12288
rect 6144 12248 6150 12260
rect 6457 12257 6469 12260
rect 6503 12257 6515 12291
rect 6457 12251 6515 12257
rect 6822 12248 6828 12300
rect 6880 12288 6886 12300
rect 8754 12288 8760 12300
rect 6880 12260 8760 12288
rect 6880 12248 6886 12260
rect 8754 12248 8760 12260
rect 8812 12288 8818 12300
rect 8849 12291 8907 12297
rect 8849 12288 8861 12291
rect 8812 12260 8861 12288
rect 8812 12248 8818 12260
rect 8849 12257 8861 12260
rect 8895 12257 8907 12291
rect 8849 12251 8907 12257
rect 11517 12291 11575 12297
rect 11517 12257 11529 12291
rect 11563 12257 11575 12291
rect 11517 12251 11575 12257
rect 11793 12291 11851 12297
rect 11793 12257 11805 12291
rect 11839 12288 11851 12291
rect 12158 12288 12164 12300
rect 11839 12260 12164 12288
rect 11839 12257 11851 12260
rect 11793 12251 11851 12257
rect 4212 12223 4270 12229
rect 4212 12220 4224 12223
rect 2556 12192 4224 12220
rect 2556 12180 2562 12192
rect 4212 12189 4224 12192
rect 4258 12189 4270 12223
rect 4212 12183 4270 12189
rect 4433 12223 4491 12229
rect 4433 12189 4445 12223
rect 4479 12189 4491 12223
rect 6638 12220 6644 12232
rect 6599 12192 6644 12220
rect 4433 12183 4491 12189
rect 6638 12180 6644 12192
rect 6696 12180 6702 12232
rect 7374 12180 7380 12232
rect 7432 12220 7438 12232
rect 7653 12223 7711 12229
rect 7653 12220 7665 12223
rect 7432 12192 7665 12220
rect 7432 12180 7438 12192
rect 7653 12189 7665 12192
rect 7699 12189 7711 12223
rect 10134 12220 10140 12232
rect 10095 12192 10140 12220
rect 7653 12183 7711 12189
rect 10134 12180 10140 12192
rect 10192 12180 10198 12232
rect 11532 12220 11560 12251
rect 12158 12248 12164 12260
rect 12216 12248 12222 12300
rect 14366 12248 14372 12300
rect 14424 12288 14430 12300
rect 16316 12288 16344 12328
rect 19429 12325 19441 12359
rect 19475 12356 19487 12359
rect 19518 12356 19524 12368
rect 19475 12328 19524 12356
rect 19475 12325 19487 12328
rect 19429 12319 19487 12325
rect 19518 12316 19524 12328
rect 19576 12316 19582 12368
rect 19978 12356 19984 12368
rect 19939 12328 19984 12356
rect 19978 12316 19984 12328
rect 20036 12316 20042 12368
rect 22462 12356 22468 12368
rect 22423 12328 22468 12356
rect 22462 12316 22468 12328
rect 22520 12316 22526 12368
rect 24673 12359 24731 12365
rect 24673 12325 24685 12359
rect 24719 12356 24731 12359
rect 24762 12356 24768 12368
rect 24719 12328 24768 12356
rect 24719 12325 24731 12328
rect 24673 12319 24731 12325
rect 24762 12316 24768 12328
rect 24820 12316 24826 12368
rect 25038 12316 25044 12368
rect 25096 12356 25102 12368
rect 25225 12359 25283 12365
rect 25225 12356 25237 12359
rect 25096 12328 25237 12356
rect 25096 12316 25102 12328
rect 25225 12325 25237 12328
rect 25271 12325 25283 12359
rect 25225 12319 25283 12325
rect 17586 12288 17592 12300
rect 14424 12260 16344 12288
rect 17547 12260 17592 12288
rect 14424 12248 14430 12260
rect 17586 12248 17592 12260
rect 17644 12248 17650 12300
rect 17678 12248 17684 12300
rect 17736 12288 17742 12300
rect 18141 12291 18199 12297
rect 18141 12288 18153 12291
rect 17736 12260 18153 12288
rect 17736 12248 17742 12260
rect 18141 12257 18153 12260
rect 18187 12288 18199 12291
rect 19058 12288 19064 12300
rect 18187 12260 19064 12288
rect 18187 12257 18199 12260
rect 18141 12251 18199 12257
rect 19058 12248 19064 12260
rect 19116 12248 19122 12300
rect 20968 12291 21026 12297
rect 20968 12257 20980 12291
rect 21014 12288 21026 12291
rect 21450 12288 21456 12300
rect 21014 12260 21456 12288
rect 21014 12257 21026 12260
rect 20968 12251 21026 12257
rect 21450 12248 21456 12260
rect 21508 12248 21514 12300
rect 11882 12220 11888 12232
rect 11532 12192 11888 12220
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 12897 12223 12955 12229
rect 12897 12189 12909 12223
rect 12943 12220 12955 12223
rect 14090 12220 14096 12232
rect 12943 12192 14096 12220
rect 12943 12189 12955 12192
rect 12897 12183 12955 12189
rect 14090 12180 14096 12192
rect 14148 12180 14154 12232
rect 15841 12223 15899 12229
rect 15841 12189 15853 12223
rect 15887 12189 15899 12223
rect 19337 12223 19395 12229
rect 19337 12220 19349 12223
rect 15841 12183 15899 12189
rect 18616 12192 19349 12220
rect 8573 12155 8631 12161
rect 8573 12121 8585 12155
rect 8619 12152 8631 12155
rect 9858 12152 9864 12164
rect 8619 12124 9864 12152
rect 8619 12121 8631 12124
rect 8573 12115 8631 12121
rect 9858 12112 9864 12124
rect 9916 12112 9922 12164
rect 13446 12152 13452 12164
rect 13407 12124 13452 12152
rect 13446 12112 13452 12124
rect 13504 12112 13510 12164
rect 1765 12087 1823 12093
rect 1765 12053 1777 12087
rect 1811 12084 1823 12087
rect 1854 12084 1860 12096
rect 1811 12056 1860 12084
rect 1811 12053 1823 12056
rect 1765 12047 1823 12053
rect 1854 12044 1860 12056
rect 1912 12044 1918 12096
rect 3878 12084 3884 12096
rect 3839 12056 3884 12084
rect 3878 12044 3884 12056
rect 3936 12044 3942 12096
rect 4338 12084 4344 12096
rect 4299 12056 4344 12084
rect 4338 12044 4344 12056
rect 4396 12044 4402 12096
rect 4522 12044 4528 12096
rect 4580 12084 4586 12096
rect 4890 12084 4896 12096
rect 4580 12056 4896 12084
rect 4580 12044 4586 12056
rect 4890 12044 4896 12056
rect 4948 12044 4954 12096
rect 12529 12087 12587 12093
rect 12529 12053 12541 12087
rect 12575 12084 12587 12087
rect 12802 12084 12808 12096
rect 12575 12056 12808 12084
rect 12575 12053 12587 12056
rect 12529 12047 12587 12053
rect 12802 12044 12808 12056
rect 12860 12044 12866 12096
rect 15286 12044 15292 12096
rect 15344 12084 15350 12096
rect 15657 12087 15715 12093
rect 15657 12084 15669 12087
rect 15344 12056 15669 12084
rect 15344 12044 15350 12056
rect 15657 12053 15669 12056
rect 15703 12084 15715 12087
rect 15856 12084 15884 12183
rect 15703 12056 15884 12084
rect 15703 12053 15715 12056
rect 15657 12047 15715 12053
rect 16298 12044 16304 12096
rect 16356 12084 16362 12096
rect 16761 12087 16819 12093
rect 16761 12084 16773 12087
rect 16356 12056 16773 12084
rect 16356 12044 16362 12056
rect 16761 12053 16773 12056
rect 16807 12084 16819 12087
rect 16850 12084 16856 12096
rect 16807 12056 16856 12084
rect 16807 12053 16819 12056
rect 16761 12047 16819 12053
rect 16850 12044 16856 12056
rect 16908 12044 16914 12096
rect 17034 12084 17040 12096
rect 16995 12056 17040 12084
rect 17034 12044 17040 12056
rect 17092 12044 17098 12096
rect 18414 12044 18420 12096
rect 18472 12084 18478 12096
rect 18616 12093 18644 12192
rect 19337 12189 19349 12192
rect 19383 12189 19395 12223
rect 19337 12183 19395 12189
rect 20530 12180 20536 12232
rect 20588 12220 20594 12232
rect 22370 12220 22376 12232
rect 20588 12192 22376 12220
rect 20588 12180 20594 12192
rect 22370 12180 22376 12192
rect 22428 12180 22434 12232
rect 22646 12220 22652 12232
rect 22607 12192 22652 12220
rect 22646 12180 22652 12192
rect 22704 12180 22710 12232
rect 24581 12223 24639 12229
rect 24581 12220 24593 12223
rect 23446 12192 24593 12220
rect 18966 12112 18972 12164
rect 19024 12152 19030 12164
rect 19061 12155 19119 12161
rect 19061 12152 19073 12155
rect 19024 12124 19073 12152
rect 19024 12112 19030 12124
rect 19061 12121 19073 12124
rect 19107 12152 19119 12155
rect 22922 12152 22928 12164
rect 19107 12124 22928 12152
rect 19107 12121 19119 12124
rect 19061 12115 19119 12121
rect 22922 12112 22928 12124
rect 22980 12112 22986 12164
rect 23290 12112 23296 12164
rect 23348 12152 23354 12164
rect 23446 12152 23474 12192
rect 24581 12189 24593 12192
rect 24627 12220 24639 12223
rect 25406 12220 25412 12232
rect 24627 12192 25412 12220
rect 24627 12189 24639 12192
rect 24581 12183 24639 12189
rect 25406 12180 25412 12192
rect 25464 12180 25470 12232
rect 23348 12124 23474 12152
rect 23348 12112 23354 12124
rect 18601 12087 18659 12093
rect 18601 12084 18613 12087
rect 18472 12056 18613 12084
rect 18472 12044 18478 12056
rect 18601 12053 18613 12056
rect 18647 12053 18659 12087
rect 21910 12084 21916 12096
rect 21871 12056 21916 12084
rect 18601 12047 18659 12053
rect 21910 12044 21916 12056
rect 21968 12044 21974 12096
rect 22646 12044 22652 12096
rect 22704 12084 22710 12096
rect 25038 12084 25044 12096
rect 22704 12056 25044 12084
rect 22704 12044 22710 12056
rect 25038 12044 25044 12056
rect 25096 12044 25102 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1762 11840 1768 11892
rect 1820 11880 1826 11892
rect 2041 11883 2099 11889
rect 2041 11880 2053 11883
rect 1820 11852 2053 11880
rect 1820 11840 1826 11852
rect 2041 11849 2053 11852
rect 2087 11849 2099 11883
rect 2041 11843 2099 11849
rect 2222 11840 2228 11892
rect 2280 11880 2286 11892
rect 2501 11883 2559 11889
rect 2501 11880 2513 11883
rect 2280 11852 2513 11880
rect 2280 11840 2286 11852
rect 2501 11849 2513 11852
rect 2547 11849 2559 11883
rect 2866 11880 2872 11892
rect 2827 11852 2872 11880
rect 2501 11843 2559 11849
rect 2516 11812 2544 11843
rect 2866 11840 2872 11852
rect 2924 11840 2930 11892
rect 4065 11883 4123 11889
rect 4065 11880 4077 11883
rect 3252 11852 4077 11880
rect 3252 11821 3280 11852
rect 4065 11849 4077 11852
rect 4111 11880 4123 11883
rect 4338 11880 4344 11892
rect 4111 11852 4344 11880
rect 4111 11849 4123 11852
rect 4065 11843 4123 11849
rect 4338 11840 4344 11852
rect 4396 11840 4402 11892
rect 4433 11883 4491 11889
rect 4433 11849 4445 11883
rect 4479 11880 4491 11883
rect 4798 11880 4804 11892
rect 4479 11852 4804 11880
rect 4479 11849 4491 11852
rect 4433 11843 4491 11849
rect 4798 11840 4804 11852
rect 4856 11840 4862 11892
rect 5534 11840 5540 11892
rect 5592 11880 5598 11892
rect 5629 11883 5687 11889
rect 5629 11880 5641 11883
rect 5592 11852 5641 11880
rect 5592 11840 5598 11852
rect 5629 11849 5641 11852
rect 5675 11849 5687 11883
rect 5629 11843 5687 11849
rect 5994 11840 6000 11892
rect 6052 11880 6058 11892
rect 6549 11883 6607 11889
rect 6549 11880 6561 11883
rect 6052 11852 6561 11880
rect 6052 11840 6058 11852
rect 6549 11849 6561 11852
rect 6595 11880 6607 11883
rect 8662 11880 8668 11892
rect 6595 11852 8668 11880
rect 6595 11849 6607 11852
rect 6549 11843 6607 11849
rect 8662 11840 8668 11852
rect 8720 11840 8726 11892
rect 10226 11880 10232 11892
rect 10187 11852 10232 11880
rect 10226 11840 10232 11852
rect 10284 11840 10290 11892
rect 12158 11880 12164 11892
rect 12119 11852 12164 11880
rect 12158 11840 12164 11852
rect 12216 11840 12222 11892
rect 14090 11880 14096 11892
rect 14003 11852 14096 11880
rect 14090 11840 14096 11852
rect 14148 11880 14154 11892
rect 19518 11880 19524 11892
rect 14148 11852 19334 11880
rect 19479 11852 19524 11880
rect 14148 11840 14154 11852
rect 3237 11815 3295 11821
rect 3237 11812 3249 11815
rect 2516 11784 3249 11812
rect 3237 11781 3249 11784
rect 3283 11781 3295 11815
rect 3237 11775 3295 11781
rect 3326 11772 3332 11824
rect 3384 11812 3390 11824
rect 3694 11812 3700 11824
rect 3384 11784 3700 11812
rect 3384 11772 3390 11784
rect 3694 11772 3700 11784
rect 3752 11812 3758 11824
rect 4893 11815 4951 11821
rect 4893 11812 4905 11815
rect 3752 11784 4905 11812
rect 3752 11772 3758 11784
rect 2372 11747 2430 11753
rect 2372 11713 2384 11747
rect 2418 11744 2430 11747
rect 2498 11744 2504 11756
rect 2418 11716 2504 11744
rect 2418 11713 2430 11716
rect 2372 11707 2430 11713
rect 2498 11704 2504 11716
rect 2556 11704 2562 11756
rect 2593 11747 2651 11753
rect 2593 11713 2605 11747
rect 2639 11744 2651 11747
rect 3344 11744 3372 11772
rect 4172 11753 4200 11784
rect 4893 11781 4905 11784
rect 4939 11812 4951 11815
rect 5810 11812 5816 11824
rect 4939 11784 5816 11812
rect 4939 11781 4951 11784
rect 4893 11775 4951 11781
rect 5810 11772 5816 11784
rect 5868 11772 5874 11824
rect 7834 11772 7840 11824
rect 7892 11812 7898 11824
rect 8757 11815 8815 11821
rect 8757 11812 8769 11815
rect 7892 11784 8769 11812
rect 7892 11772 7898 11784
rect 8757 11781 8769 11784
rect 8803 11812 8815 11815
rect 9858 11812 9864 11824
rect 8803 11784 9864 11812
rect 8803 11781 8815 11784
rect 8757 11775 8815 11781
rect 9858 11772 9864 11784
rect 9916 11772 9922 11824
rect 10686 11772 10692 11824
rect 10744 11812 10750 11824
rect 13722 11812 13728 11824
rect 10744 11784 13728 11812
rect 10744 11772 10750 11784
rect 13722 11772 13728 11784
rect 13780 11772 13786 11824
rect 13998 11772 14004 11824
rect 14056 11812 14062 11824
rect 17034 11812 17040 11824
rect 14056 11784 17040 11812
rect 14056 11772 14062 11784
rect 4157 11747 4215 11753
rect 4157 11744 4169 11747
rect 2639 11716 3372 11744
rect 4135 11716 4169 11744
rect 2639 11713 2651 11716
rect 2593 11707 2651 11713
rect 4157 11713 4169 11716
rect 4203 11713 4215 11747
rect 7742 11744 7748 11756
rect 7703 11716 7748 11744
rect 4157 11707 4215 11713
rect 7742 11704 7748 11716
rect 7800 11704 7806 11756
rect 8110 11704 8116 11756
rect 8168 11744 8174 11756
rect 9306 11744 9312 11756
rect 8168 11716 9312 11744
rect 8168 11704 8174 11716
rect 9306 11704 9312 11716
rect 9364 11704 9370 11756
rect 9950 11744 9956 11756
rect 9911 11716 9956 11744
rect 9950 11704 9956 11716
rect 10008 11704 10014 11756
rect 12434 11704 12440 11756
rect 12492 11744 12498 11756
rect 12713 11747 12771 11753
rect 12713 11744 12725 11747
rect 12492 11716 12725 11744
rect 12492 11704 12498 11716
rect 12713 11713 12725 11716
rect 12759 11713 12771 11747
rect 15286 11744 15292 11756
rect 15247 11716 15292 11744
rect 12713 11707 12771 11713
rect 15286 11704 15292 11716
rect 15344 11704 15350 11756
rect 15654 11704 15660 11756
rect 15712 11744 15718 11756
rect 16224 11753 16252 11784
rect 17034 11772 17040 11784
rect 17092 11772 17098 11824
rect 17313 11815 17371 11821
rect 17313 11781 17325 11815
rect 17359 11812 17371 11815
rect 17678 11812 17684 11824
rect 17359 11784 17684 11812
rect 17359 11781 17371 11784
rect 17313 11775 17371 11781
rect 15841 11747 15899 11753
rect 15841 11744 15853 11747
rect 15712 11716 15853 11744
rect 15712 11704 15718 11716
rect 15841 11713 15853 11716
rect 15887 11713 15899 11747
rect 15841 11707 15899 11713
rect 16209 11747 16267 11753
rect 16209 11713 16221 11747
rect 16255 11713 16267 11747
rect 16482 11744 16488 11756
rect 16443 11716 16488 11744
rect 16209 11707 16267 11713
rect 16482 11704 16488 11716
rect 16540 11704 16546 11756
rect 1765 11679 1823 11685
rect 1765 11645 1777 11679
rect 1811 11676 1823 11679
rect 2222 11676 2228 11688
rect 1811 11648 2228 11676
rect 1811 11645 1823 11648
rect 1765 11639 1823 11645
rect 2222 11636 2228 11648
rect 2280 11636 2286 11688
rect 3878 11636 3884 11688
rect 3936 11685 3942 11688
rect 3936 11679 3994 11685
rect 3936 11645 3948 11679
rect 3982 11645 3994 11679
rect 5350 11676 5356 11688
rect 5311 11648 5356 11676
rect 3936 11639 3994 11645
rect 3936 11636 3942 11639
rect 5350 11636 5356 11648
rect 5408 11636 5414 11688
rect 5442 11636 5448 11688
rect 5500 11676 5506 11688
rect 5537 11679 5595 11685
rect 5537 11676 5549 11679
rect 5500 11648 5549 11676
rect 5500 11636 5506 11648
rect 5537 11645 5549 11648
rect 5583 11676 5595 11679
rect 6181 11679 6239 11685
rect 6181 11676 6193 11679
rect 5583 11648 6193 11676
rect 5583 11645 5595 11648
rect 5537 11639 5595 11645
rect 6181 11645 6193 11648
rect 6227 11645 6239 11679
rect 6181 11639 6239 11645
rect 8389 11679 8447 11685
rect 8389 11645 8401 11679
rect 8435 11676 8447 11679
rect 8570 11676 8576 11688
rect 8435 11648 8576 11676
rect 8435 11645 8447 11648
rect 8389 11639 8447 11645
rect 8570 11636 8576 11648
rect 8628 11676 8634 11688
rect 9122 11676 9128 11688
rect 8628 11648 9128 11676
rect 8628 11636 8634 11648
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 10781 11679 10839 11685
rect 10781 11676 10793 11679
rect 10612 11648 10793 11676
rect 3602 11568 3608 11620
rect 3660 11608 3666 11620
rect 3789 11611 3847 11617
rect 3789 11608 3801 11611
rect 3660 11580 3801 11608
rect 3660 11568 3666 11580
rect 3789 11577 3801 11580
rect 3835 11577 3847 11611
rect 3789 11571 3847 11577
rect 4338 11568 4344 11620
rect 4396 11608 4402 11620
rect 5169 11611 5227 11617
rect 5169 11608 5181 11611
rect 4396 11580 5181 11608
rect 4396 11568 4402 11580
rect 5169 11577 5181 11580
rect 5215 11577 5227 11611
rect 5169 11571 5227 11577
rect 7834 11568 7840 11620
rect 7892 11608 7898 11620
rect 9401 11611 9459 11617
rect 7892 11580 7937 11608
rect 7892 11568 7898 11580
rect 9401 11577 9413 11611
rect 9447 11577 9459 11611
rect 9401 11571 9459 11577
rect 2406 11500 2412 11552
rect 2464 11540 2470 11552
rect 2590 11540 2596 11552
rect 2464 11512 2596 11540
rect 2464 11500 2470 11512
rect 2590 11500 2596 11512
rect 2648 11540 2654 11552
rect 4430 11540 4436 11552
rect 2648 11512 4436 11540
rect 2648 11500 2654 11512
rect 4430 11500 4436 11512
rect 4488 11500 4494 11552
rect 7193 11543 7251 11549
rect 7193 11509 7205 11543
rect 7239 11540 7251 11543
rect 7374 11540 7380 11552
rect 7239 11512 7380 11540
rect 7239 11509 7251 11512
rect 7193 11503 7251 11509
rect 7374 11500 7380 11512
rect 7432 11500 7438 11552
rect 7561 11543 7619 11549
rect 7561 11509 7573 11543
rect 7607 11540 7619 11543
rect 8018 11540 8024 11552
rect 7607 11512 8024 11540
rect 7607 11509 7619 11512
rect 7561 11503 7619 11509
rect 8018 11500 8024 11512
rect 8076 11500 8082 11552
rect 8846 11500 8852 11552
rect 8904 11540 8910 11552
rect 9033 11543 9091 11549
rect 9033 11540 9045 11543
rect 8904 11512 9045 11540
rect 8904 11500 8910 11512
rect 9033 11509 9045 11512
rect 9079 11540 9091 11543
rect 9416 11540 9444 11571
rect 9079 11512 9444 11540
rect 9079 11509 9091 11512
rect 9033 11503 9091 11509
rect 9582 11500 9588 11552
rect 9640 11540 9646 11552
rect 10042 11540 10048 11552
rect 9640 11512 10048 11540
rect 9640 11500 9646 11512
rect 10042 11500 10048 11512
rect 10100 11540 10106 11552
rect 10612 11549 10640 11648
rect 10781 11645 10793 11648
rect 10827 11645 10839 11679
rect 10781 11639 10839 11645
rect 11146 11636 11152 11688
rect 11204 11676 11210 11688
rect 11241 11679 11299 11685
rect 11241 11676 11253 11679
rect 11204 11648 11253 11676
rect 11204 11636 11210 11648
rect 11241 11645 11253 11648
rect 11287 11645 11299 11679
rect 11241 11639 11299 11645
rect 14461 11679 14519 11685
rect 14461 11645 14473 11679
rect 14507 11676 14519 11679
rect 14734 11676 14740 11688
rect 14507 11648 14740 11676
rect 14507 11645 14519 11648
rect 14461 11639 14519 11645
rect 14734 11636 14740 11648
rect 14792 11636 14798 11688
rect 15102 11676 15108 11688
rect 15015 11648 15108 11676
rect 15102 11636 15108 11648
rect 15160 11676 15166 11688
rect 15160 11648 16068 11676
rect 15160 11636 15166 11648
rect 11514 11608 11520 11620
rect 11475 11580 11520 11608
rect 11514 11568 11520 11580
rect 11572 11568 11578 11620
rect 12802 11608 12808 11620
rect 12763 11580 12808 11608
rect 12802 11568 12808 11580
rect 12860 11568 12866 11620
rect 13354 11608 13360 11620
rect 13315 11580 13360 11608
rect 13354 11568 13360 11580
rect 13412 11568 13418 11620
rect 10597 11543 10655 11549
rect 10597 11540 10609 11543
rect 10100 11512 10609 11540
rect 10100 11500 10106 11512
rect 10597 11509 10609 11512
rect 10643 11509 10655 11543
rect 11882 11540 11888 11552
rect 11843 11512 11888 11540
rect 10597 11503 10655 11509
rect 11882 11500 11888 11512
rect 11940 11500 11946 11552
rect 13630 11540 13636 11552
rect 13591 11512 13636 11540
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 16040 11540 16068 11648
rect 16298 11568 16304 11620
rect 16356 11608 16362 11620
rect 16356 11580 16401 11608
rect 16356 11568 16362 11580
rect 17328 11540 17356 11775
rect 17678 11772 17684 11784
rect 17736 11772 17742 11824
rect 19306 11812 19334 11852
rect 19518 11840 19524 11852
rect 19576 11840 19582 11892
rect 22462 11840 22468 11892
rect 22520 11880 22526 11892
rect 22830 11880 22836 11892
rect 22520 11852 22836 11880
rect 22520 11840 22526 11852
rect 22830 11840 22836 11852
rect 22888 11880 22894 11892
rect 22925 11883 22983 11889
rect 22925 11880 22937 11883
rect 22888 11852 22937 11880
rect 22888 11840 22894 11852
rect 22925 11849 22937 11852
rect 22971 11849 22983 11883
rect 22925 11843 22983 11849
rect 24118 11840 24124 11892
rect 24176 11880 24182 11892
rect 24213 11883 24271 11889
rect 24213 11880 24225 11883
rect 24176 11852 24225 11880
rect 24176 11840 24182 11852
rect 24213 11849 24225 11852
rect 24259 11849 24271 11883
rect 25406 11880 25412 11892
rect 25367 11852 25412 11880
rect 24213 11843 24271 11849
rect 20162 11812 20168 11824
rect 19306 11784 20168 11812
rect 20162 11772 20168 11784
rect 20220 11772 20226 11824
rect 20346 11772 20352 11824
rect 20404 11812 20410 11824
rect 20404 11784 20484 11812
rect 20404 11772 20410 11784
rect 17586 11744 17592 11756
rect 17547 11716 17592 11744
rect 17586 11704 17592 11716
rect 17644 11704 17650 11756
rect 20456 11753 20484 11784
rect 22370 11772 22376 11824
rect 22428 11812 22434 11824
rect 23293 11815 23351 11821
rect 23293 11812 23305 11815
rect 22428 11784 23305 11812
rect 22428 11772 22434 11784
rect 23293 11781 23305 11784
rect 23339 11781 23351 11815
rect 23293 11775 23351 11781
rect 20441 11747 20499 11753
rect 20441 11713 20453 11747
rect 20487 11713 20499 11747
rect 20441 11707 20499 11713
rect 20530 11704 20536 11756
rect 20588 11744 20594 11756
rect 20717 11747 20775 11753
rect 20717 11744 20729 11747
rect 20588 11716 20729 11744
rect 20588 11704 20594 11716
rect 20717 11713 20729 11716
rect 20763 11713 20775 11747
rect 22646 11744 22652 11756
rect 22607 11716 22652 11744
rect 20717 11707 20775 11713
rect 22646 11704 22652 11716
rect 22704 11704 22710 11756
rect 24228 11744 24256 11843
rect 25406 11840 25412 11852
rect 25464 11840 25470 11892
rect 25038 11812 25044 11824
rect 24999 11784 25044 11812
rect 25038 11772 25044 11784
rect 25096 11772 25102 11824
rect 24489 11747 24547 11753
rect 24489 11744 24501 11747
rect 24228 11716 24501 11744
rect 24489 11713 24501 11716
rect 24535 11713 24547 11747
rect 24489 11707 24547 11713
rect 18509 11679 18567 11685
rect 18509 11676 18521 11679
rect 18340 11648 18521 11676
rect 16040 11512 17356 11540
rect 18230 11500 18236 11552
rect 18288 11540 18294 11552
rect 18340 11549 18368 11648
rect 18509 11645 18521 11648
rect 18555 11645 18567 11679
rect 18966 11676 18972 11688
rect 18927 11648 18972 11676
rect 18509 11639 18567 11645
rect 18966 11636 18972 11648
rect 19024 11636 19030 11688
rect 20533 11611 20591 11617
rect 20533 11608 20545 11611
rect 20272 11580 20545 11608
rect 20272 11552 20300 11580
rect 20533 11577 20545 11580
rect 20579 11577 20591 11611
rect 22002 11608 22008 11620
rect 21963 11580 22008 11608
rect 20533 11571 20591 11577
rect 22002 11568 22008 11580
rect 22060 11568 22066 11620
rect 22097 11611 22155 11617
rect 22097 11577 22109 11611
rect 22143 11577 22155 11611
rect 22097 11571 22155 11577
rect 18325 11543 18383 11549
rect 18325 11540 18337 11543
rect 18288 11512 18337 11540
rect 18288 11500 18294 11512
rect 18325 11509 18337 11512
rect 18371 11509 18383 11543
rect 18782 11540 18788 11552
rect 18743 11512 18788 11540
rect 18325 11503 18383 11509
rect 18782 11500 18788 11512
rect 18840 11500 18846 11552
rect 20254 11540 20260 11552
rect 20215 11512 20260 11540
rect 20254 11500 20260 11512
rect 20312 11500 20318 11552
rect 21450 11540 21456 11552
rect 21411 11512 21456 11540
rect 21450 11500 21456 11512
rect 21508 11500 21514 11552
rect 21726 11540 21732 11552
rect 21687 11512 21732 11540
rect 21726 11500 21732 11512
rect 21784 11540 21790 11552
rect 22112 11540 22140 11571
rect 24578 11568 24584 11620
rect 24636 11608 24642 11620
rect 24636 11580 24681 11608
rect 24636 11568 24642 11580
rect 21784 11512 22140 11540
rect 23937 11543 23995 11549
rect 21784 11500 21790 11512
rect 23937 11509 23949 11543
rect 23983 11540 23995 11543
rect 24762 11540 24768 11552
rect 23983 11512 24768 11540
rect 23983 11509 23995 11512
rect 23937 11503 23995 11509
rect 24762 11500 24768 11512
rect 24820 11500 24826 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1854 11296 1860 11348
rect 1912 11336 1918 11348
rect 3694 11336 3700 11348
rect 1912 11308 3700 11336
rect 1912 11296 1918 11308
rect 3694 11296 3700 11308
rect 3752 11336 3758 11348
rect 3789 11339 3847 11345
rect 3789 11336 3801 11339
rect 3752 11308 3801 11336
rect 3752 11296 3758 11308
rect 3789 11305 3801 11308
rect 3835 11336 3847 11339
rect 3878 11336 3884 11348
rect 3835 11308 3884 11336
rect 3835 11305 3847 11308
rect 3789 11299 3847 11305
rect 3878 11296 3884 11308
rect 3936 11296 3942 11348
rect 5445 11339 5503 11345
rect 5445 11336 5457 11339
rect 4264 11308 5457 11336
rect 4264 11280 4292 11308
rect 5445 11305 5457 11308
rect 5491 11336 5503 11339
rect 5534 11336 5540 11348
rect 5491 11308 5540 11336
rect 5491 11305 5503 11308
rect 5445 11299 5503 11305
rect 5534 11296 5540 11308
rect 5592 11296 5598 11348
rect 5810 11336 5816 11348
rect 5771 11308 5816 11336
rect 5810 11296 5816 11308
rect 5868 11296 5874 11348
rect 6086 11336 6092 11348
rect 6047 11308 6092 11336
rect 6086 11296 6092 11308
rect 6144 11296 6150 11348
rect 7561 11339 7619 11345
rect 7561 11305 7573 11339
rect 7607 11336 7619 11339
rect 7834 11336 7840 11348
rect 7607 11308 7840 11336
rect 7607 11305 7619 11308
rect 7561 11299 7619 11305
rect 7834 11296 7840 11308
rect 7892 11296 7898 11348
rect 8202 11296 8208 11348
rect 8260 11336 8266 11348
rect 8573 11339 8631 11345
rect 8573 11336 8585 11339
rect 8260 11308 8585 11336
rect 8260 11296 8266 11308
rect 8573 11305 8585 11308
rect 8619 11305 8631 11339
rect 9306 11336 9312 11348
rect 9267 11308 9312 11336
rect 8573 11299 8631 11305
rect 1486 11228 1492 11280
rect 1544 11268 1550 11280
rect 1544 11240 2452 11268
rect 1544 11228 1550 11240
rect 2424 11212 2452 11240
rect 2498 11228 2504 11280
rect 2556 11268 2562 11280
rect 3142 11268 3148 11280
rect 2556 11240 3148 11268
rect 2556 11228 2562 11240
rect 3142 11228 3148 11240
rect 3200 11268 3206 11280
rect 3421 11271 3479 11277
rect 3421 11268 3433 11271
rect 3200 11240 3433 11268
rect 3200 11228 3206 11240
rect 3421 11237 3433 11240
rect 3467 11237 3479 11271
rect 3421 11231 3479 11237
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 1762 11200 1768 11212
rect 1443 11172 1768 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 1762 11160 1768 11172
rect 1820 11160 1826 11212
rect 2406 11200 2412 11212
rect 2319 11172 2412 11200
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 1949 11135 2007 11141
rect 1949 11101 1961 11135
rect 1995 11132 2007 11135
rect 2516 11132 2544 11228
rect 2774 11160 2780 11212
rect 2832 11200 2838 11212
rect 2869 11203 2927 11209
rect 2869 11200 2881 11203
rect 2832 11172 2881 11200
rect 2832 11160 2838 11172
rect 2869 11169 2881 11172
rect 2915 11169 2927 11203
rect 3436 11200 3464 11231
rect 3602 11228 3608 11280
rect 3660 11268 3666 11280
rect 4246 11268 4252 11280
rect 3660 11240 3877 11268
rect 3660 11228 3666 11240
rect 3849 11200 3877 11240
rect 4172 11240 4252 11268
rect 3970 11200 3976 11212
rect 3436 11172 3740 11200
rect 3849 11172 3976 11200
rect 2869 11163 2927 11169
rect 1995 11104 2544 11132
rect 3145 11135 3203 11141
rect 1995 11101 2007 11104
rect 1949 11095 2007 11101
rect 3145 11101 3157 11135
rect 3191 11132 3203 11135
rect 3602 11132 3608 11144
rect 3191 11104 3608 11132
rect 3191 11101 3203 11104
rect 3145 11095 3203 11101
rect 3602 11092 3608 11104
rect 3660 11092 3666 11144
rect 3712 11132 3740 11172
rect 3970 11160 3976 11172
rect 4028 11200 4034 11212
rect 4065 11203 4123 11209
rect 4065 11200 4077 11203
rect 4028 11172 4077 11200
rect 4028 11160 4034 11172
rect 4065 11169 4077 11172
rect 4111 11200 4123 11203
rect 4172 11200 4200 11240
rect 4246 11228 4252 11240
rect 4304 11228 4310 11280
rect 4798 11268 4804 11280
rect 4759 11240 4804 11268
rect 4798 11228 4804 11240
rect 4856 11228 4862 11280
rect 6362 11228 6368 11280
rect 6420 11268 6426 11280
rect 6457 11271 6515 11277
rect 6457 11268 6469 11271
rect 6420 11240 6469 11268
rect 6420 11228 6426 11240
rect 6457 11237 6469 11240
rect 6503 11237 6515 11271
rect 6457 11231 6515 11237
rect 4111 11172 4200 11200
rect 4111 11169 4123 11172
rect 4065 11163 4123 11169
rect 5442 11160 5448 11212
rect 5500 11200 5506 11212
rect 5629 11203 5687 11209
rect 5629 11200 5641 11203
rect 5500 11172 5641 11200
rect 5500 11160 5506 11172
rect 5629 11169 5641 11172
rect 5675 11169 5687 11203
rect 5629 11163 5687 11169
rect 4246 11141 4252 11144
rect 4212 11135 4252 11141
rect 4212 11132 4224 11135
rect 3712 11104 4224 11132
rect 4212 11101 4224 11104
rect 4212 11095 4252 11101
rect 4246 11092 4252 11095
rect 4304 11092 4310 11144
rect 4430 11132 4436 11144
rect 4391 11104 4436 11132
rect 4430 11092 4436 11104
rect 4488 11132 4494 11144
rect 5077 11135 5135 11141
rect 5077 11132 5089 11135
rect 4488 11104 5089 11132
rect 4488 11092 4494 11104
rect 5077 11101 5089 11104
rect 5123 11101 5135 11135
rect 6472 11132 6500 11231
rect 6730 11228 6736 11280
rect 6788 11268 6794 11280
rect 7003 11271 7061 11277
rect 7003 11268 7015 11271
rect 6788 11240 7015 11268
rect 6788 11228 6794 11240
rect 7003 11237 7015 11240
rect 7049 11268 7061 11271
rect 8018 11268 8024 11280
rect 7049 11240 8024 11268
rect 7049 11237 7061 11240
rect 7003 11231 7061 11237
rect 8018 11228 8024 11240
rect 8076 11228 8082 11280
rect 8588 11268 8616 11299
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 14001 11339 14059 11345
rect 14001 11336 14013 11339
rect 12492 11308 14013 11336
rect 12492 11296 12498 11308
rect 14001 11305 14013 11308
rect 14047 11305 14059 11339
rect 14001 11299 14059 11305
rect 14645 11339 14703 11345
rect 14645 11305 14657 11339
rect 14691 11336 14703 11339
rect 15102 11336 15108 11348
rect 14691 11308 15108 11336
rect 14691 11305 14703 11308
rect 14645 11299 14703 11305
rect 15102 11296 15108 11308
rect 15160 11296 15166 11348
rect 15519 11339 15577 11345
rect 15519 11305 15531 11339
rect 15565 11336 15577 11339
rect 16114 11336 16120 11348
rect 15565 11308 16120 11336
rect 15565 11305 15577 11308
rect 15519 11299 15577 11305
rect 16114 11296 16120 11308
rect 16172 11296 16178 11348
rect 16209 11339 16267 11345
rect 16209 11305 16221 11339
rect 16255 11336 16267 11339
rect 16298 11336 16304 11348
rect 16255 11308 16304 11336
rect 16255 11305 16267 11308
rect 16209 11299 16267 11305
rect 16298 11296 16304 11308
rect 16356 11296 16362 11348
rect 18141 11339 18199 11345
rect 18141 11305 18153 11339
rect 18187 11336 18199 11339
rect 18322 11336 18328 11348
rect 18187 11308 18328 11336
rect 18187 11305 18199 11308
rect 18141 11299 18199 11305
rect 18322 11296 18328 11308
rect 18380 11296 18386 11348
rect 18782 11296 18788 11348
rect 18840 11336 18846 11348
rect 18877 11339 18935 11345
rect 18877 11336 18889 11339
rect 18840 11308 18889 11336
rect 18840 11296 18846 11308
rect 18877 11305 18889 11308
rect 18923 11336 18935 11339
rect 19426 11336 19432 11348
rect 18923 11308 19104 11336
rect 19387 11308 19432 11336
rect 18923 11305 18935 11308
rect 18877 11299 18935 11305
rect 9398 11268 9404 11280
rect 8588 11240 9404 11268
rect 9398 11228 9404 11240
rect 9456 11228 9462 11280
rect 9858 11268 9864 11280
rect 9819 11240 9864 11268
rect 9858 11228 9864 11240
rect 9916 11228 9922 11280
rect 11603 11271 11661 11277
rect 11603 11237 11615 11271
rect 11649 11268 11661 11271
rect 11698 11268 11704 11280
rect 11649 11240 11704 11268
rect 11649 11237 11661 11240
rect 11603 11231 11661 11237
rect 11698 11228 11704 11240
rect 11756 11228 11762 11280
rect 12618 11228 12624 11280
rect 12676 11268 12682 11280
rect 13173 11271 13231 11277
rect 13173 11268 13185 11271
rect 12676 11240 13185 11268
rect 12676 11228 12682 11240
rect 13173 11237 13185 11240
rect 13219 11237 13231 11271
rect 13173 11231 13231 11237
rect 13354 11228 13360 11280
rect 13412 11268 13418 11280
rect 13725 11271 13783 11277
rect 13725 11268 13737 11271
rect 13412 11240 13737 11268
rect 13412 11228 13418 11240
rect 13725 11237 13737 11240
rect 13771 11237 13783 11271
rect 16574 11268 16580 11280
rect 16535 11240 16580 11268
rect 13725 11231 13783 11237
rect 16574 11228 16580 11240
rect 16632 11228 16638 11280
rect 17770 11228 17776 11280
rect 17828 11268 17834 11280
rect 18509 11271 18567 11277
rect 18509 11268 18521 11271
rect 17828 11240 18521 11268
rect 17828 11228 17834 11240
rect 18509 11237 18521 11240
rect 18555 11268 18567 11271
rect 18966 11268 18972 11280
rect 18555 11240 18972 11268
rect 18555 11237 18567 11240
rect 18509 11231 18567 11237
rect 18966 11228 18972 11240
rect 19024 11228 19030 11280
rect 6638 11200 6644 11212
rect 6599 11172 6644 11200
rect 6638 11160 6644 11172
rect 6696 11200 6702 11212
rect 8205 11203 8263 11209
rect 8205 11200 8217 11203
rect 6696 11172 8217 11200
rect 6696 11160 6702 11172
rect 8205 11169 8217 11172
rect 8251 11169 8263 11203
rect 8205 11163 8263 11169
rect 8294 11160 8300 11212
rect 8352 11200 8358 11212
rect 8389 11203 8447 11209
rect 8389 11200 8401 11203
rect 8352 11172 8401 11200
rect 8352 11160 8358 11172
rect 8389 11169 8401 11172
rect 8435 11169 8447 11203
rect 15286 11200 15292 11212
rect 15247 11172 15292 11200
rect 8389 11163 8447 11169
rect 15286 11160 15292 11172
rect 15344 11160 15350 11212
rect 17957 11203 18015 11209
rect 17957 11169 17969 11203
rect 18003 11169 18015 11203
rect 17957 11163 18015 11169
rect 6472 11104 7696 11132
rect 5077 11095 5135 11101
rect 1581 11067 1639 11073
rect 1581 11033 1593 11067
rect 1627 11064 1639 11067
rect 2130 11064 2136 11076
rect 1627 11036 2136 11064
rect 1627 11033 1639 11036
rect 1581 11027 1639 11033
rect 2130 11024 2136 11036
rect 2188 11024 2194 11076
rect 2317 11067 2375 11073
rect 2317 11033 2329 11067
rect 2363 11064 2375 11067
rect 2682 11064 2688 11076
rect 2363 11036 2688 11064
rect 2363 11033 2375 11036
rect 2317 11027 2375 11033
rect 2682 11024 2688 11036
rect 2740 11064 2746 11076
rect 3326 11064 3332 11076
rect 2740 11036 3332 11064
rect 2740 11024 2746 11036
rect 3326 11024 3332 11036
rect 3384 11024 3390 11076
rect 7558 11064 7564 11076
rect 4126 11036 7564 11064
rect 3878 10956 3884 11008
rect 3936 10996 3942 11008
rect 4126 10996 4154 11036
rect 7558 11024 7564 11036
rect 7616 11024 7622 11076
rect 7668 11064 7696 11104
rect 8478 11092 8484 11144
rect 8536 11132 8542 11144
rect 9766 11132 9772 11144
rect 8536 11104 9772 11132
rect 8536 11092 8542 11104
rect 9766 11092 9772 11104
rect 9824 11092 9830 11144
rect 9950 11092 9956 11144
rect 10008 11132 10014 11144
rect 10045 11135 10103 11141
rect 10045 11132 10057 11135
rect 10008 11104 10057 11132
rect 10008 11092 10014 11104
rect 10045 11101 10057 11104
rect 10091 11101 10103 11135
rect 10045 11095 10103 11101
rect 11241 11135 11299 11141
rect 11241 11101 11253 11135
rect 11287 11132 11299 11135
rect 11514 11132 11520 11144
rect 11287 11104 11520 11132
rect 11287 11101 11299 11104
rect 11241 11095 11299 11101
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 13081 11135 13139 11141
rect 13081 11101 13093 11135
rect 13127 11132 13139 11135
rect 13998 11132 14004 11144
rect 13127 11104 14004 11132
rect 13127 11101 13139 11104
rect 13081 11095 13139 11101
rect 13998 11092 14004 11104
rect 14056 11092 14062 11144
rect 16485 11135 16543 11141
rect 16485 11101 16497 11135
rect 16531 11101 16543 11135
rect 16942 11132 16948 11144
rect 16903 11104 16948 11132
rect 16485 11095 16543 11101
rect 10781 11067 10839 11073
rect 10781 11064 10793 11067
rect 7668 11036 10793 11064
rect 10781 11033 10793 11036
rect 10827 11064 10839 11067
rect 11146 11064 11152 11076
rect 10827 11036 11152 11064
rect 10827 11033 10839 11036
rect 10781 11027 10839 11033
rect 11146 11024 11152 11036
rect 11204 11024 11210 11076
rect 12161 11067 12219 11073
rect 12161 11033 12173 11067
rect 12207 11064 12219 11067
rect 13630 11064 13636 11076
rect 12207 11036 13636 11064
rect 12207 11033 12219 11036
rect 12161 11027 12219 11033
rect 13630 11024 13636 11036
rect 13688 11024 13694 11076
rect 15378 11064 15384 11076
rect 13786 11036 15384 11064
rect 4338 10996 4344 11008
rect 3936 10968 4154 10996
rect 4299 10968 4344 10996
rect 3936 10956 3942 10968
rect 4338 10956 4344 10968
rect 4396 10956 4402 11008
rect 4982 10956 4988 11008
rect 5040 10996 5046 11008
rect 5166 10996 5172 11008
rect 5040 10968 5172 10996
rect 5040 10956 5046 10968
rect 5166 10956 5172 10968
rect 5224 10956 5230 11008
rect 7834 10996 7840 11008
rect 7795 10968 7840 10996
rect 7834 10956 7840 10968
rect 7892 10956 7898 11008
rect 8846 10996 8852 11008
rect 8807 10968 8852 10996
rect 8846 10956 8852 10968
rect 8904 10956 8910 11008
rect 11790 10956 11796 11008
rect 11848 10996 11854 11008
rect 12621 10999 12679 11005
rect 12621 10996 12633 10999
rect 11848 10968 12633 10996
rect 11848 10956 11854 10968
rect 12621 10965 12633 10968
rect 12667 10996 12679 10999
rect 12802 10996 12808 11008
rect 12667 10968 12808 10996
rect 12667 10965 12679 10968
rect 12621 10959 12679 10965
rect 12802 10956 12808 10968
rect 12860 10956 12866 11008
rect 13078 10956 13084 11008
rect 13136 10996 13142 11008
rect 13786 10996 13814 11036
rect 15378 11024 15384 11036
rect 15436 11024 15442 11076
rect 16500 11064 16528 11095
rect 16942 11092 16948 11104
rect 17000 11092 17006 11144
rect 17862 11092 17868 11144
rect 17920 11132 17926 11144
rect 17972 11132 18000 11163
rect 17920 11104 18000 11132
rect 18984 11132 19012 11228
rect 19076 11209 19104 11308
rect 19426 11296 19432 11308
rect 19484 11296 19490 11348
rect 20346 11336 20352 11348
rect 20307 11308 20352 11336
rect 20346 11296 20352 11308
rect 20404 11296 20410 11348
rect 22186 11296 22192 11348
rect 22244 11336 22250 11348
rect 22281 11339 22339 11345
rect 22281 11336 22293 11339
rect 22244 11308 22293 11336
rect 22244 11296 22250 11308
rect 22281 11305 22293 11308
rect 22327 11305 22339 11339
rect 22830 11336 22836 11348
rect 22791 11308 22836 11336
rect 22281 11299 22339 11305
rect 22296 11268 22324 11299
rect 22830 11296 22836 11308
rect 22888 11296 22894 11348
rect 24578 11296 24584 11348
rect 24636 11336 24642 11348
rect 24857 11339 24915 11345
rect 24857 11336 24869 11339
rect 24636 11308 24869 11336
rect 24636 11296 24642 11308
rect 24857 11305 24869 11308
rect 24903 11305 24915 11339
rect 24857 11299 24915 11305
rect 23474 11268 23480 11280
rect 22296 11240 23480 11268
rect 23474 11228 23480 11240
rect 23532 11268 23538 11280
rect 23982 11271 24040 11277
rect 23982 11268 23994 11271
rect 23532 11240 23994 11268
rect 23532 11228 23538 11240
rect 23982 11237 23994 11240
rect 24028 11237 24040 11271
rect 23982 11231 24040 11237
rect 19061 11203 19119 11209
rect 19061 11169 19073 11203
rect 19107 11169 19119 11203
rect 19061 11163 19119 11169
rect 19242 11160 19248 11212
rect 19300 11200 19306 11212
rect 20070 11200 20076 11212
rect 19300 11172 20076 11200
rect 19300 11160 19306 11172
rect 20070 11160 20076 11172
rect 20128 11160 20134 11212
rect 20806 11200 20812 11212
rect 20767 11172 20812 11200
rect 20806 11160 20812 11172
rect 20864 11200 20870 11212
rect 21266 11200 21272 11212
rect 20864 11172 21272 11200
rect 20864 11160 20870 11172
rect 21266 11160 21272 11172
rect 21324 11160 21330 11212
rect 24581 11203 24639 11209
rect 24581 11169 24593 11203
rect 24627 11200 24639 11203
rect 24762 11200 24768 11212
rect 24627 11172 24768 11200
rect 24627 11169 24639 11172
rect 24581 11163 24639 11169
rect 24762 11160 24768 11172
rect 24820 11160 24826 11212
rect 25444 11203 25502 11209
rect 25444 11169 25456 11203
rect 25490 11169 25502 11203
rect 25444 11163 25502 11169
rect 19610 11132 19616 11144
rect 18984 11104 19616 11132
rect 17920 11092 17926 11104
rect 19610 11092 19616 11104
rect 19668 11092 19674 11144
rect 20254 11132 20260 11144
rect 19996 11104 20260 11132
rect 19996 11073 20024 11104
rect 20254 11092 20260 11104
rect 20312 11132 20318 11144
rect 21082 11132 21088 11144
rect 20312 11104 21088 11132
rect 20312 11092 20318 11104
rect 21082 11092 21088 11104
rect 21140 11092 21146 11144
rect 21913 11135 21971 11141
rect 21913 11101 21925 11135
rect 21959 11132 21971 11135
rect 22278 11132 22284 11144
rect 21959 11104 22284 11132
rect 21959 11101 21971 11104
rect 21913 11095 21971 11101
rect 22278 11092 22284 11104
rect 22336 11092 22342 11144
rect 23658 11132 23664 11144
rect 23619 11104 23664 11132
rect 23658 11092 23664 11104
rect 23716 11092 23722 11144
rect 24026 11092 24032 11144
rect 24084 11132 24090 11144
rect 25222 11132 25228 11144
rect 24084 11104 25228 11132
rect 24084 11092 24090 11104
rect 25222 11092 25228 11104
rect 25280 11132 25286 11144
rect 25459 11132 25487 11163
rect 25280 11104 25487 11132
rect 25280 11092 25286 11104
rect 19981 11067 20039 11073
rect 16500 11036 17540 11064
rect 17512 11005 17540 11036
rect 19981 11033 19993 11067
rect 20027 11033 20039 11067
rect 19981 11027 20039 11033
rect 20162 11024 20168 11076
rect 20220 11064 20226 11076
rect 25547 11067 25605 11073
rect 25547 11064 25559 11067
rect 20220 11036 25559 11064
rect 20220 11024 20226 11036
rect 25547 11033 25559 11036
rect 25593 11033 25605 11067
rect 25547 11027 25605 11033
rect 13136 10968 13814 10996
rect 17497 10999 17555 11005
rect 13136 10956 13142 10968
rect 17497 10965 17509 10999
rect 17543 10996 17555 10999
rect 17586 10996 17592 11008
rect 17543 10968 17592 10996
rect 17543 10965 17555 10968
rect 17497 10959 17555 10965
rect 17586 10956 17592 10968
rect 17644 10956 17650 11008
rect 20070 10956 20076 11008
rect 20128 10996 20134 11008
rect 21039 10999 21097 11005
rect 21039 10996 21051 10999
rect 20128 10968 21051 10996
rect 20128 10956 20134 10968
rect 21039 10965 21051 10968
rect 21085 10965 21097 10999
rect 21358 10996 21364 11008
rect 21319 10968 21364 10996
rect 21039 10959 21097 10965
rect 21358 10956 21364 10968
rect 21416 10956 21422 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1673 10795 1731 10801
rect 1673 10761 1685 10795
rect 1719 10792 1731 10795
rect 1762 10792 1768 10804
rect 1719 10764 1768 10792
rect 1719 10761 1731 10764
rect 1673 10755 1731 10761
rect 1762 10752 1768 10764
rect 1820 10752 1826 10804
rect 2130 10752 2136 10804
rect 2188 10792 2194 10804
rect 2314 10792 2320 10804
rect 2188 10764 2320 10792
rect 2188 10752 2194 10764
rect 2314 10752 2320 10764
rect 2372 10752 2378 10804
rect 3050 10752 3056 10804
rect 3108 10792 3114 10804
rect 4249 10795 4307 10801
rect 4249 10792 4261 10795
rect 3108 10764 4261 10792
rect 3108 10752 3114 10764
rect 4249 10761 4261 10764
rect 4295 10761 4307 10795
rect 4249 10755 4307 10761
rect 4338 10752 4344 10804
rect 4396 10792 4402 10804
rect 4801 10795 4859 10801
rect 4801 10792 4813 10795
rect 4396 10764 4813 10792
rect 4396 10752 4402 10764
rect 4801 10761 4813 10764
rect 4847 10761 4859 10795
rect 4801 10755 4859 10761
rect 5261 10795 5319 10801
rect 5261 10761 5273 10795
rect 5307 10792 5319 10795
rect 5350 10792 5356 10804
rect 5307 10764 5356 10792
rect 5307 10761 5319 10764
rect 5261 10755 5319 10761
rect 5350 10752 5356 10764
rect 5408 10752 5414 10804
rect 6641 10795 6699 10801
rect 6641 10761 6653 10795
rect 6687 10792 6699 10795
rect 6730 10792 6736 10804
rect 6687 10764 6736 10792
rect 6687 10761 6699 10764
rect 6641 10755 6699 10761
rect 6730 10752 6736 10764
rect 6788 10752 6794 10804
rect 13630 10752 13636 10804
rect 13688 10792 13694 10804
rect 14093 10795 14151 10801
rect 14093 10792 14105 10795
rect 13688 10764 14105 10792
rect 13688 10752 13694 10764
rect 14093 10761 14105 10764
rect 14139 10792 14151 10795
rect 14458 10792 14464 10804
rect 14139 10764 14464 10792
rect 14139 10761 14151 10764
rect 14093 10755 14151 10761
rect 14458 10752 14464 10764
rect 14516 10752 14522 10804
rect 15654 10752 15660 10804
rect 15712 10792 15718 10804
rect 15933 10795 15991 10801
rect 15933 10792 15945 10795
rect 15712 10764 15945 10792
rect 15712 10752 15718 10764
rect 15933 10761 15945 10764
rect 15979 10761 15991 10795
rect 17862 10792 17868 10804
rect 17823 10764 17868 10792
rect 15933 10755 15991 10761
rect 17862 10752 17868 10764
rect 17920 10752 17926 10804
rect 21637 10795 21695 10801
rect 21637 10761 21649 10795
rect 21683 10792 21695 10795
rect 21726 10792 21732 10804
rect 21683 10764 21732 10792
rect 21683 10761 21695 10764
rect 21637 10755 21695 10761
rect 21726 10752 21732 10764
rect 21784 10752 21790 10804
rect 23474 10752 23480 10804
rect 23532 10792 23538 10804
rect 24581 10795 24639 10801
rect 23532 10764 23577 10792
rect 23532 10752 23538 10764
rect 24581 10761 24593 10795
rect 24627 10792 24639 10795
rect 24670 10792 24676 10804
rect 24627 10764 24676 10792
rect 24627 10761 24639 10764
rect 24581 10755 24639 10761
rect 24670 10752 24676 10764
rect 24728 10752 24734 10804
rect 25222 10792 25228 10804
rect 25183 10764 25228 10792
rect 25222 10752 25228 10764
rect 25280 10752 25286 10804
rect 25590 10792 25596 10804
rect 25551 10764 25596 10792
rect 25590 10752 25596 10764
rect 25648 10752 25654 10804
rect 3326 10684 3332 10736
rect 3384 10724 3390 10736
rect 3605 10727 3663 10733
rect 3605 10724 3617 10727
rect 3384 10696 3617 10724
rect 3384 10684 3390 10696
rect 3605 10693 3617 10696
rect 3651 10693 3663 10727
rect 3605 10687 3663 10693
rect 2406 10616 2412 10668
rect 2464 10656 2470 10668
rect 3050 10656 3056 10668
rect 2464 10628 3056 10656
rect 2464 10616 2470 10628
rect 3050 10616 3056 10628
rect 3108 10656 3114 10668
rect 3237 10659 3295 10665
rect 3237 10656 3249 10659
rect 3108 10628 3249 10656
rect 3108 10616 3114 10628
rect 3237 10625 3249 10628
rect 3283 10625 3295 10659
rect 3620 10656 3648 10687
rect 3694 10684 3700 10736
rect 3752 10724 3758 10736
rect 3927 10727 3985 10733
rect 3927 10724 3939 10727
rect 3752 10696 3939 10724
rect 3752 10684 3758 10696
rect 3927 10693 3939 10696
rect 3973 10693 3985 10727
rect 4062 10724 4068 10736
rect 4023 10696 4068 10724
rect 3927 10687 3985 10693
rect 4062 10684 4068 10696
rect 4120 10684 4126 10736
rect 13354 10684 13360 10736
rect 13412 10724 13418 10736
rect 13412 10696 14688 10724
rect 13412 10684 13418 10696
rect 4157 10659 4215 10665
rect 3620 10628 3924 10656
rect 3237 10619 3295 10625
rect 14 10548 20 10600
rect 72 10588 78 10600
rect 2041 10591 2099 10597
rect 2041 10588 2053 10591
rect 72 10560 2053 10588
rect 72 10548 78 10560
rect 2041 10557 2053 10560
rect 2087 10588 2099 10591
rect 2314 10588 2320 10600
rect 2087 10560 2320 10588
rect 2087 10557 2099 10560
rect 2041 10551 2099 10557
rect 2314 10548 2320 10560
rect 2372 10548 2378 10600
rect 3786 10588 3792 10600
rect 3747 10560 3792 10588
rect 3786 10548 3792 10560
rect 3844 10548 3850 10600
rect 3896 10588 3924 10628
rect 4157 10625 4169 10659
rect 4203 10625 4215 10659
rect 4157 10619 4215 10625
rect 4172 10588 4200 10619
rect 4982 10616 4988 10668
rect 5040 10656 5046 10668
rect 5442 10656 5448 10668
rect 5040 10628 5448 10656
rect 5040 10616 5046 10628
rect 5442 10616 5448 10628
rect 5500 10656 5506 10668
rect 6181 10659 6239 10665
rect 6181 10656 6193 10659
rect 5500 10628 6193 10656
rect 5500 10616 5506 10628
rect 6181 10625 6193 10628
rect 6227 10625 6239 10659
rect 7098 10656 7104 10668
rect 7011 10628 7104 10656
rect 6181 10619 6239 10625
rect 7098 10616 7104 10628
rect 7156 10656 7162 10668
rect 7834 10656 7840 10668
rect 7156 10628 7840 10656
rect 7156 10616 7162 10628
rect 7834 10616 7840 10628
rect 7892 10616 7898 10668
rect 9122 10616 9128 10668
rect 9180 10656 9186 10668
rect 9217 10659 9275 10665
rect 9217 10656 9229 10659
rect 9180 10628 9229 10656
rect 9180 10616 9186 10628
rect 9217 10625 9229 10628
rect 9263 10625 9275 10659
rect 12802 10656 12808 10668
rect 12763 10628 12808 10656
rect 9217 10619 9275 10625
rect 12802 10616 12808 10628
rect 12860 10616 12866 10668
rect 12894 10616 12900 10668
rect 12952 10656 12958 10668
rect 13633 10659 13691 10665
rect 13633 10656 13645 10659
rect 12952 10628 13645 10656
rect 12952 10616 12958 10628
rect 13633 10625 13645 10628
rect 13679 10625 13691 10659
rect 14366 10656 14372 10668
rect 14327 10628 14372 10656
rect 13633 10619 13691 10625
rect 14366 10616 14372 10628
rect 14424 10616 14430 10668
rect 14660 10665 14688 10696
rect 14918 10684 14924 10736
rect 14976 10724 14982 10736
rect 22603 10727 22661 10733
rect 22603 10724 22615 10727
rect 14976 10696 22615 10724
rect 14976 10684 14982 10696
rect 22603 10693 22615 10696
rect 22649 10693 22661 10727
rect 22603 10687 22661 10693
rect 14645 10659 14703 10665
rect 14645 10625 14657 10659
rect 14691 10625 14703 10659
rect 14645 10619 14703 10625
rect 14826 10616 14832 10668
rect 14884 10656 14890 10668
rect 16114 10656 16120 10668
rect 14884 10628 16120 10656
rect 14884 10616 14890 10628
rect 16114 10616 16120 10628
rect 16172 10616 16178 10668
rect 19889 10659 19947 10665
rect 16776 10628 19840 10656
rect 3896 10560 4200 10588
rect 5258 10548 5264 10600
rect 5316 10588 5322 10600
rect 5537 10591 5595 10597
rect 5537 10588 5549 10591
rect 5316 10560 5549 10588
rect 5316 10548 5322 10560
rect 5537 10557 5549 10560
rect 5583 10557 5595 10591
rect 5537 10551 5595 10557
rect 8021 10591 8079 10597
rect 8021 10557 8033 10591
rect 8067 10588 8079 10591
rect 10134 10588 10140 10600
rect 8067 10560 8708 10588
rect 10047 10560 10140 10588
rect 8067 10557 8079 10560
rect 8021 10551 8079 10557
rect 3804 10520 3832 10548
rect 4062 10520 4068 10532
rect 3804 10492 4068 10520
rect 4062 10480 4068 10492
rect 4120 10480 4126 10532
rect 5350 10520 5356 10532
rect 5311 10492 5356 10520
rect 5350 10480 5356 10492
rect 5408 10480 5414 10532
rect 6730 10480 6736 10532
rect 6788 10520 6794 10532
rect 7190 10520 7196 10532
rect 6788 10492 7196 10520
rect 6788 10480 6794 10492
rect 7190 10480 7196 10492
rect 7248 10520 7254 10532
rect 7422 10523 7480 10529
rect 7422 10520 7434 10523
rect 7248 10492 7434 10520
rect 7248 10480 7254 10492
rect 7422 10489 7434 10492
rect 7468 10489 7480 10523
rect 7422 10483 7480 10489
rect 2498 10452 2504 10464
rect 2459 10424 2504 10452
rect 2498 10412 2504 10424
rect 2556 10412 2562 10464
rect 3694 10412 3700 10464
rect 3752 10452 3758 10464
rect 3970 10452 3976 10464
rect 3752 10424 3976 10452
rect 3752 10412 3758 10424
rect 3970 10412 3976 10424
rect 4028 10412 4034 10464
rect 5626 10452 5632 10464
rect 5587 10424 5632 10452
rect 5626 10412 5632 10424
rect 5684 10412 5690 10464
rect 8294 10412 8300 10464
rect 8352 10452 8358 10464
rect 8389 10455 8447 10461
rect 8389 10452 8401 10455
rect 8352 10424 8401 10452
rect 8352 10412 8358 10424
rect 8389 10421 8401 10424
rect 8435 10421 8447 10455
rect 8680 10452 8708 10560
rect 10134 10548 10140 10560
rect 10192 10588 10198 10600
rect 10597 10591 10655 10597
rect 10597 10588 10609 10591
rect 10192 10560 10609 10588
rect 10192 10548 10198 10560
rect 10597 10557 10609 10560
rect 10643 10557 10655 10591
rect 10597 10551 10655 10557
rect 11517 10591 11575 10597
rect 11517 10557 11529 10591
rect 11563 10588 11575 10591
rect 12161 10591 12219 10597
rect 12161 10588 12173 10591
rect 11563 10560 12173 10588
rect 11563 10557 11575 10560
rect 11517 10551 11575 10557
rect 12161 10557 12173 10560
rect 12207 10557 12219 10591
rect 12161 10551 12219 10557
rect 8754 10480 8760 10532
rect 8812 10520 8818 10532
rect 8941 10523 8999 10529
rect 8941 10520 8953 10523
rect 8812 10492 8953 10520
rect 8812 10480 8818 10492
rect 8941 10489 8953 10492
rect 8987 10489 8999 10523
rect 8941 10483 8999 10489
rect 9033 10523 9091 10529
rect 9033 10489 9045 10523
rect 9079 10489 9091 10523
rect 9033 10483 9091 10489
rect 10505 10523 10563 10529
rect 10505 10489 10517 10523
rect 10551 10520 10563 10523
rect 10918 10523 10976 10529
rect 10918 10520 10930 10523
rect 10551 10492 10930 10520
rect 10551 10489 10563 10492
rect 10505 10483 10563 10489
rect 10918 10489 10930 10492
rect 10964 10520 10976 10523
rect 11698 10520 11704 10532
rect 10964 10492 11704 10520
rect 10964 10489 10976 10492
rect 10918 10483 10976 10489
rect 8846 10452 8852 10464
rect 8680 10424 8852 10452
rect 8389 10415 8447 10421
rect 8846 10412 8852 10424
rect 8904 10452 8910 10464
rect 9048 10452 9076 10483
rect 11698 10480 11704 10492
rect 11756 10520 11762 10532
rect 11793 10523 11851 10529
rect 11793 10520 11805 10523
rect 11756 10492 11805 10520
rect 11756 10480 11762 10492
rect 11793 10489 11805 10492
rect 11839 10489 11851 10523
rect 12176 10520 12204 10551
rect 15286 10548 15292 10600
rect 15344 10588 15350 10600
rect 15473 10591 15531 10597
rect 15473 10588 15485 10591
rect 15344 10560 15485 10588
rect 15344 10548 15350 10560
rect 15473 10557 15485 10560
rect 15519 10588 15531 10591
rect 16776 10588 16804 10628
rect 15519 10560 16804 10588
rect 15519 10557 15531 10560
rect 15473 10551 15531 10557
rect 17954 10548 17960 10600
rect 18012 10588 18018 10600
rect 18176 10591 18234 10597
rect 18176 10588 18188 10591
rect 18012 10560 18188 10588
rect 18012 10548 18018 10560
rect 18176 10557 18188 10560
rect 18222 10588 18234 10591
rect 18601 10591 18659 10597
rect 18601 10588 18613 10591
rect 18222 10560 18613 10588
rect 18222 10557 18234 10560
rect 18176 10551 18234 10557
rect 18601 10557 18613 10560
rect 18647 10557 18659 10591
rect 19242 10588 19248 10600
rect 19203 10560 19248 10588
rect 18601 10551 18659 10557
rect 19242 10548 19248 10560
rect 19300 10548 19306 10600
rect 19610 10588 19616 10600
rect 19571 10560 19616 10588
rect 19610 10548 19616 10560
rect 19668 10548 19674 10600
rect 19812 10588 19840 10628
rect 19889 10625 19901 10659
rect 19935 10656 19947 10659
rect 20717 10659 20775 10665
rect 20717 10656 20729 10659
rect 19935 10628 20729 10656
rect 19935 10625 19947 10628
rect 19889 10619 19947 10625
rect 20717 10625 20729 10628
rect 20763 10656 20775 10659
rect 21358 10656 21364 10668
rect 20763 10628 21364 10656
rect 20763 10625 20775 10628
rect 20717 10619 20775 10625
rect 21358 10616 21364 10628
rect 21416 10616 21422 10668
rect 21450 10588 21456 10600
rect 19812 10560 21456 10588
rect 21450 10548 21456 10560
rect 21508 10548 21514 10600
rect 22532 10591 22590 10597
rect 22532 10557 22544 10591
rect 22578 10588 22590 10591
rect 22830 10588 22836 10600
rect 22578 10560 22836 10588
rect 22578 10557 22590 10560
rect 22532 10551 22590 10557
rect 22830 10548 22836 10560
rect 22888 10588 22894 10600
rect 22925 10591 22983 10597
rect 22925 10588 22937 10591
rect 22888 10560 22937 10588
rect 22888 10548 22894 10560
rect 22925 10557 22937 10560
rect 22971 10557 22983 10591
rect 22925 10551 22983 10557
rect 23661 10591 23719 10597
rect 23661 10557 23673 10591
rect 23707 10588 23719 10591
rect 24578 10588 24584 10600
rect 23707 10560 24584 10588
rect 23707 10557 23719 10560
rect 23661 10551 23719 10557
rect 24578 10548 24584 10560
rect 24636 10588 24642 10600
rect 24857 10591 24915 10597
rect 24857 10588 24869 10591
rect 24636 10560 24869 10588
rect 24636 10548 24642 10560
rect 24857 10557 24869 10560
rect 24903 10557 24915 10591
rect 24857 10551 24915 10557
rect 25409 10591 25467 10597
rect 25409 10557 25421 10591
rect 25455 10588 25467 10591
rect 25590 10588 25596 10600
rect 25455 10560 25596 10588
rect 25455 10557 25467 10560
rect 25409 10551 25467 10557
rect 25590 10548 25596 10560
rect 25648 10588 25654 10600
rect 25961 10591 26019 10597
rect 25961 10588 25973 10591
rect 25648 10560 25973 10588
rect 25648 10548 25654 10560
rect 25961 10557 25973 10560
rect 26007 10557 26019 10591
rect 25961 10551 26019 10557
rect 12618 10520 12624 10532
rect 12176 10492 12624 10520
rect 11793 10483 11851 10489
rect 8904 10424 9076 10452
rect 11808 10452 11836 10483
rect 12618 10480 12624 10492
rect 12676 10520 12682 10532
rect 12897 10523 12955 10529
rect 12897 10520 12909 10523
rect 12676 10492 12909 10520
rect 12676 10480 12682 10492
rect 12897 10489 12909 10492
rect 12943 10489 12955 10523
rect 13446 10520 13452 10532
rect 13407 10492 13452 10520
rect 12897 10483 12955 10489
rect 12434 10452 12440 10464
rect 11808 10424 12440 10452
rect 8904 10412 8910 10424
rect 12434 10412 12440 10424
rect 12492 10412 12498 10464
rect 12912 10452 12940 10483
rect 13446 10480 13452 10492
rect 13504 10480 13510 10532
rect 13725 10523 13783 10529
rect 13725 10520 13737 10523
rect 13556 10492 13737 10520
rect 13556 10452 13584 10492
rect 13725 10489 13737 10492
rect 13771 10489 13783 10523
rect 13725 10483 13783 10489
rect 14458 10480 14464 10532
rect 14516 10520 14522 10532
rect 14516 10492 14561 10520
rect 14516 10480 14522 10492
rect 15654 10480 15660 10532
rect 15712 10520 15718 10532
rect 16438 10523 16496 10529
rect 16438 10520 16450 10523
rect 15712 10492 16450 10520
rect 15712 10480 15718 10492
rect 16438 10489 16450 10492
rect 16484 10520 16496 10523
rect 17218 10520 17224 10532
rect 16484 10492 17224 10520
rect 16484 10489 16496 10492
rect 16438 10483 16496 10489
rect 17218 10480 17224 10492
rect 17276 10520 17282 10532
rect 18969 10523 19027 10529
rect 18969 10520 18981 10523
rect 17276 10492 18981 10520
rect 17276 10480 17282 10492
rect 18969 10489 18981 10492
rect 19015 10520 19027 10523
rect 19426 10520 19432 10532
rect 19015 10492 19432 10520
rect 19015 10489 19027 10492
rect 18969 10483 19027 10489
rect 19426 10480 19432 10492
rect 19484 10520 19490 10532
rect 20165 10523 20223 10529
rect 20165 10520 20177 10523
rect 19484 10492 20177 10520
rect 19484 10480 19490 10492
rect 20165 10489 20177 10492
rect 20211 10520 20223 10523
rect 21038 10523 21096 10529
rect 21038 10520 21050 10523
rect 20211 10492 21050 10520
rect 20211 10489 20223 10492
rect 20165 10483 20223 10489
rect 21038 10489 21050 10492
rect 21084 10520 21096 10523
rect 21913 10523 21971 10529
rect 21913 10520 21925 10523
rect 21084 10492 21925 10520
rect 21084 10489 21096 10492
rect 21038 10483 21096 10489
rect 21913 10489 21925 10492
rect 21959 10520 21971 10523
rect 22186 10520 22192 10532
rect 21959 10492 22192 10520
rect 21959 10489 21971 10492
rect 21913 10483 21971 10489
rect 22186 10480 22192 10492
rect 22244 10480 22250 10532
rect 23474 10480 23480 10532
rect 23532 10520 23538 10532
rect 23750 10520 23756 10532
rect 23532 10492 23756 10520
rect 23532 10480 23538 10492
rect 23750 10480 23756 10492
rect 23808 10520 23814 10532
rect 23982 10523 24040 10529
rect 23982 10520 23994 10523
rect 23808 10492 23994 10520
rect 23808 10480 23814 10492
rect 23982 10489 23994 10492
rect 24028 10489 24040 10523
rect 23982 10483 24040 10489
rect 12912 10424 13584 10452
rect 13633 10455 13691 10461
rect 13633 10421 13645 10455
rect 13679 10452 13691 10455
rect 14734 10452 14740 10464
rect 13679 10424 14740 10452
rect 13679 10421 13691 10424
rect 13633 10415 13691 10421
rect 14734 10412 14740 10424
rect 14792 10412 14798 10464
rect 16574 10412 16580 10464
rect 16632 10452 16638 10464
rect 17037 10455 17095 10461
rect 17037 10452 17049 10455
rect 16632 10424 17049 10452
rect 16632 10412 16638 10424
rect 17037 10421 17049 10424
rect 17083 10452 17095 10455
rect 17313 10455 17371 10461
rect 17313 10452 17325 10455
rect 17083 10424 17325 10452
rect 17083 10421 17095 10424
rect 17037 10415 17095 10421
rect 17313 10421 17325 10424
rect 17359 10421 17371 10455
rect 17313 10415 17371 10421
rect 18279 10455 18337 10461
rect 18279 10421 18291 10455
rect 18325 10452 18337 10455
rect 18506 10452 18512 10464
rect 18325 10424 18512 10452
rect 18325 10421 18337 10424
rect 18279 10415 18337 10421
rect 18506 10412 18512 10424
rect 18564 10412 18570 10464
rect 20625 10455 20683 10461
rect 20625 10421 20637 10455
rect 20671 10452 20683 10455
rect 20806 10452 20812 10464
rect 20671 10424 20812 10452
rect 20671 10421 20683 10424
rect 20625 10415 20683 10421
rect 20806 10412 20812 10424
rect 20864 10452 20870 10464
rect 21726 10452 21732 10464
rect 20864 10424 21732 10452
rect 20864 10412 20870 10424
rect 21726 10412 21732 10424
rect 21784 10412 21790 10464
rect 22278 10452 22284 10464
rect 22239 10424 22284 10452
rect 22278 10412 22284 10424
rect 22336 10412 22342 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 2314 10208 2320 10260
rect 2372 10248 2378 10260
rect 4706 10248 4712 10260
rect 2372 10220 4568 10248
rect 4667 10220 4712 10248
rect 2372 10208 2378 10220
rect 3970 10180 3976 10192
rect 3068 10152 3976 10180
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10112 1455 10115
rect 1946 10112 1952 10124
rect 1443 10084 1952 10112
rect 1443 10081 1455 10084
rect 1397 10075 1455 10081
rect 1946 10072 1952 10084
rect 2004 10072 2010 10124
rect 3068 10121 3096 10152
rect 3970 10140 3976 10152
rect 4028 10140 4034 10192
rect 4540 10180 4568 10220
rect 4706 10208 4712 10220
rect 4764 10208 4770 10260
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 5721 10251 5779 10257
rect 5721 10248 5733 10251
rect 5592 10220 5733 10248
rect 5592 10208 5598 10220
rect 5721 10217 5733 10220
rect 5767 10217 5779 10251
rect 5721 10211 5779 10217
rect 7190 10208 7196 10260
rect 7248 10248 7254 10260
rect 7377 10251 7435 10257
rect 7377 10248 7389 10251
rect 7248 10220 7389 10248
rect 7248 10208 7254 10220
rect 7377 10217 7389 10220
rect 7423 10217 7435 10251
rect 9858 10248 9864 10260
rect 9819 10220 9864 10248
rect 7377 10211 7435 10217
rect 9858 10208 9864 10220
rect 9916 10208 9922 10260
rect 10134 10208 10140 10260
rect 10192 10248 10198 10260
rect 10229 10251 10287 10257
rect 10229 10248 10241 10251
rect 10192 10220 10241 10248
rect 10192 10208 10198 10220
rect 10229 10217 10241 10220
rect 10275 10217 10287 10251
rect 11146 10248 11152 10260
rect 11107 10220 11152 10248
rect 10229 10211 10287 10217
rect 11146 10208 11152 10220
rect 11204 10208 11210 10260
rect 11514 10248 11520 10260
rect 11475 10220 11520 10248
rect 11514 10208 11520 10220
rect 11572 10208 11578 10260
rect 12345 10251 12403 10257
rect 12345 10217 12357 10251
rect 12391 10248 12403 10251
rect 12802 10248 12808 10260
rect 12391 10220 12808 10248
rect 12391 10217 12403 10220
rect 12345 10211 12403 10217
rect 12802 10208 12808 10220
rect 12860 10208 12866 10260
rect 13998 10248 14004 10260
rect 13911 10220 14004 10248
rect 13998 10208 14004 10220
rect 14056 10248 14062 10260
rect 14918 10248 14924 10260
rect 14056 10220 14924 10248
rect 14056 10208 14062 10220
rect 14918 10208 14924 10220
rect 14976 10208 14982 10260
rect 15611 10251 15669 10257
rect 15611 10217 15623 10251
rect 15657 10248 15669 10251
rect 18233 10251 18291 10257
rect 18233 10248 18245 10251
rect 15657 10220 18245 10248
rect 15657 10217 15669 10220
rect 15611 10211 15669 10217
rect 18233 10217 18245 10220
rect 18279 10248 18291 10251
rect 18322 10248 18328 10260
rect 18279 10220 18328 10248
rect 18279 10217 18291 10220
rect 18233 10211 18291 10217
rect 18322 10208 18328 10220
rect 18380 10208 18386 10260
rect 19518 10208 19524 10260
rect 19576 10248 19582 10260
rect 19797 10251 19855 10257
rect 19797 10248 19809 10251
rect 19576 10220 19809 10248
rect 19576 10208 19582 10220
rect 19797 10217 19809 10220
rect 19843 10217 19855 10251
rect 23750 10248 23756 10260
rect 23711 10220 23756 10248
rect 19797 10211 19855 10217
rect 23750 10208 23756 10220
rect 23808 10208 23814 10260
rect 24578 10248 24584 10260
rect 24539 10220 24584 10248
rect 24578 10208 24584 10220
rect 24636 10208 24642 10260
rect 5442 10180 5448 10192
rect 4540 10152 5448 10180
rect 5442 10140 5448 10152
rect 5500 10140 5506 10192
rect 7098 10180 7104 10192
rect 7059 10152 7104 10180
rect 7098 10140 7104 10152
rect 7156 10140 7162 10192
rect 10042 10140 10048 10192
rect 10100 10180 10106 10192
rect 10100 10152 10180 10180
rect 10100 10140 10106 10152
rect 3053 10115 3111 10121
rect 3053 10081 3065 10115
rect 3099 10081 3111 10115
rect 4062 10112 4068 10124
rect 4023 10084 4068 10112
rect 3053 10075 3111 10081
rect 4062 10072 4068 10084
rect 4120 10112 4126 10124
rect 5994 10112 6000 10124
rect 4120 10084 6000 10112
rect 4120 10072 4126 10084
rect 5994 10072 6000 10084
rect 6052 10112 6058 10124
rect 6089 10115 6147 10121
rect 6089 10112 6101 10115
rect 6052 10084 6101 10112
rect 6052 10072 6058 10084
rect 6089 10081 6101 10084
rect 6135 10081 6147 10115
rect 6362 10112 6368 10124
rect 6323 10084 6368 10112
rect 6089 10075 6147 10081
rect 6362 10072 6368 10084
rect 6420 10072 6426 10124
rect 6454 10072 6460 10124
rect 6512 10112 6518 10124
rect 6825 10115 6883 10121
rect 6825 10112 6837 10115
rect 6512 10084 6837 10112
rect 6512 10072 6518 10084
rect 6825 10081 6837 10084
rect 6871 10112 6883 10115
rect 7190 10112 7196 10124
rect 6871 10084 7196 10112
rect 6871 10081 6883 10084
rect 6825 10075 6883 10081
rect 7190 10072 7196 10084
rect 7248 10112 7254 10124
rect 7745 10115 7803 10121
rect 7745 10112 7757 10115
rect 7248 10084 7757 10112
rect 7248 10072 7254 10084
rect 7745 10081 7757 10084
rect 7791 10081 7803 10115
rect 7745 10075 7803 10081
rect 7929 10115 7987 10121
rect 7929 10081 7941 10115
rect 7975 10112 7987 10115
rect 8018 10112 8024 10124
rect 7975 10084 8024 10112
rect 7975 10081 7987 10084
rect 7929 10075 7987 10081
rect 8018 10072 8024 10084
rect 8076 10072 8082 10124
rect 10152 10121 10180 10152
rect 8205 10115 8263 10121
rect 8205 10081 8217 10115
rect 8251 10081 8263 10115
rect 8205 10075 8263 10081
rect 10137 10115 10195 10121
rect 10137 10081 10149 10115
rect 10183 10081 10195 10115
rect 10686 10112 10692 10124
rect 10599 10084 10692 10112
rect 10137 10075 10195 10081
rect 3145 10047 3203 10053
rect 3145 10013 3157 10047
rect 3191 10044 3203 10047
rect 3786 10044 3792 10056
rect 3191 10016 3792 10044
rect 3191 10013 3203 10016
rect 3145 10007 3203 10013
rect 3786 10004 3792 10016
rect 3844 10004 3850 10056
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 4212 10016 4384 10044
rect 4212 10004 4218 10016
rect 4356 9985 4384 10016
rect 4430 10004 4436 10056
rect 4488 10044 4494 10056
rect 4488 10016 4533 10044
rect 4488 10004 4494 10016
rect 7834 10004 7840 10056
rect 7892 10044 7898 10056
rect 8220 10044 8248 10075
rect 10686 10072 10692 10084
rect 10744 10112 10750 10124
rect 11164 10112 11192 10208
rect 12618 10180 12624 10192
rect 12579 10152 12624 10180
rect 12618 10140 12624 10152
rect 12676 10140 12682 10192
rect 13081 10183 13139 10189
rect 13081 10149 13093 10183
rect 13127 10180 13139 10183
rect 13630 10180 13636 10192
rect 13127 10152 13636 10180
rect 13127 10149 13139 10152
rect 13081 10143 13139 10149
rect 13630 10140 13636 10152
rect 13688 10140 13694 10192
rect 14366 10180 14372 10192
rect 14327 10152 14372 10180
rect 14366 10140 14372 10152
rect 14424 10140 14430 10192
rect 16114 10180 16120 10192
rect 16075 10152 16120 10180
rect 16114 10140 16120 10152
rect 16172 10140 16178 10192
rect 16574 10140 16580 10192
rect 16632 10180 16638 10192
rect 16669 10183 16727 10189
rect 16669 10180 16681 10183
rect 16632 10152 16681 10180
rect 16632 10140 16638 10152
rect 16669 10149 16681 10152
rect 16715 10149 16727 10183
rect 18506 10180 18512 10192
rect 18467 10152 18512 10180
rect 16669 10143 16727 10149
rect 18506 10140 18512 10152
rect 18564 10140 18570 10192
rect 18598 10140 18604 10192
rect 18656 10180 18662 10192
rect 21082 10180 21088 10192
rect 18656 10152 18701 10180
rect 21043 10152 21088 10180
rect 18656 10140 18662 10152
rect 21082 10140 21088 10152
rect 21140 10140 21146 10192
rect 23477 10183 23535 10189
rect 23477 10149 23489 10183
rect 23523 10180 23535 10183
rect 23658 10180 23664 10192
rect 23523 10152 23664 10180
rect 23523 10149 23535 10152
rect 23477 10143 23535 10149
rect 23658 10140 23664 10152
rect 23716 10180 23722 10192
rect 24121 10183 24179 10189
rect 24121 10180 24133 10183
rect 23716 10152 24133 10180
rect 23716 10140 23722 10152
rect 24121 10149 24133 10152
rect 24167 10149 24179 10183
rect 24121 10143 24179 10149
rect 11698 10112 11704 10124
rect 10744 10084 11192 10112
rect 11659 10084 11704 10112
rect 10744 10072 10750 10084
rect 11698 10072 11704 10084
rect 11756 10072 11762 10124
rect 15381 10115 15439 10121
rect 15381 10081 15393 10115
rect 15427 10112 15439 10115
rect 15562 10112 15568 10124
rect 15427 10084 15568 10112
rect 15427 10081 15439 10084
rect 15381 10075 15439 10081
rect 15562 10072 15568 10084
rect 15620 10112 15626 10124
rect 16022 10112 16028 10124
rect 15620 10084 16028 10112
rect 15620 10072 15626 10084
rect 16022 10072 16028 10084
rect 16080 10072 16086 10124
rect 22738 10112 22744 10124
rect 22699 10084 22744 10112
rect 22738 10072 22744 10084
rect 22796 10072 22802 10124
rect 23198 10112 23204 10124
rect 23159 10084 23204 10112
rect 23198 10072 23204 10084
rect 23256 10072 23262 10124
rect 23382 10072 23388 10124
rect 23440 10112 23446 10124
rect 24305 10115 24363 10121
rect 24305 10112 24317 10115
rect 23440 10084 24317 10112
rect 23440 10072 23446 10084
rect 24305 10081 24317 10084
rect 24351 10081 24363 10115
rect 24305 10075 24363 10081
rect 24765 10115 24823 10121
rect 24765 10081 24777 10115
rect 24811 10081 24823 10115
rect 24765 10075 24823 10081
rect 8386 10044 8392 10056
rect 7892 10016 8248 10044
rect 8347 10016 8392 10044
rect 7892 10004 7898 10016
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 12989 10047 13047 10053
rect 12989 10013 13001 10047
rect 13035 10044 13047 10047
rect 13262 10044 13268 10056
rect 13035 10016 13268 10044
rect 13035 10013 13047 10016
rect 12989 10007 13047 10013
rect 13262 10004 13268 10016
rect 13320 10044 13326 10056
rect 14274 10044 14280 10056
rect 13320 10016 14280 10044
rect 13320 10004 13326 10016
rect 14274 10004 14280 10016
rect 14332 10004 14338 10056
rect 16577 10047 16635 10053
rect 16577 10013 16589 10047
rect 16623 10044 16635 10047
rect 16942 10044 16948 10056
rect 16623 10016 16948 10044
rect 16623 10013 16635 10016
rect 16577 10007 16635 10013
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 18874 10044 18880 10056
rect 18835 10016 18880 10044
rect 18874 10004 18880 10016
rect 18932 10004 18938 10056
rect 20993 10047 21051 10053
rect 20993 10013 21005 10047
rect 21039 10044 21051 10047
rect 21174 10044 21180 10056
rect 21039 10016 21180 10044
rect 21039 10013 21051 10016
rect 20993 10007 21051 10013
rect 21174 10004 21180 10016
rect 21232 10004 21238 10056
rect 21269 10047 21327 10053
rect 21269 10013 21281 10047
rect 21315 10044 21327 10047
rect 21910 10044 21916 10056
rect 21315 10016 21916 10044
rect 21315 10013 21327 10016
rect 21269 10007 21327 10013
rect 1581 9979 1639 9985
rect 1581 9945 1593 9979
rect 1627 9976 1639 9979
rect 4341 9979 4399 9985
rect 4341 9976 4353 9979
rect 1627 9948 3188 9976
rect 1627 9945 1639 9948
rect 1581 9939 1639 9945
rect 3160 9920 3188 9948
rect 3988 9948 4353 9976
rect 1854 9868 1860 9920
rect 1912 9908 1918 9920
rect 2133 9911 2191 9917
rect 2133 9908 2145 9911
rect 1912 9880 2145 9908
rect 1912 9868 1918 9880
rect 2133 9877 2145 9880
rect 2179 9877 2191 9911
rect 2133 9871 2191 9877
rect 3142 9868 3148 9920
rect 3200 9908 3206 9920
rect 3421 9911 3479 9917
rect 3421 9908 3433 9911
rect 3200 9880 3433 9908
rect 3200 9868 3206 9880
rect 3421 9877 3433 9880
rect 3467 9877 3479 9911
rect 3421 9871 3479 9877
rect 3881 9911 3939 9917
rect 3881 9877 3893 9911
rect 3927 9908 3939 9911
rect 3988 9908 4016 9948
rect 4341 9945 4353 9948
rect 4387 9945 4399 9979
rect 5350 9976 5356 9988
rect 5311 9948 5356 9976
rect 4341 9939 4399 9945
rect 5350 9936 5356 9948
rect 5408 9936 5414 9988
rect 8021 9979 8079 9985
rect 8021 9945 8033 9979
rect 8067 9945 8079 9979
rect 8021 9939 8079 9945
rect 4246 9917 4252 9920
rect 3927 9880 4016 9908
rect 4230 9911 4252 9917
rect 3927 9877 3939 9880
rect 3881 9871 3939 9877
rect 4230 9877 4242 9911
rect 4230 9871 4252 9877
rect 4246 9868 4252 9871
rect 4304 9868 4310 9920
rect 8036 9908 8064 9939
rect 8202 9936 8208 9988
rect 8260 9976 8266 9988
rect 9309 9979 9367 9985
rect 9309 9976 9321 9979
rect 8260 9948 9321 9976
rect 8260 9936 8266 9948
rect 9309 9945 9321 9948
rect 9355 9945 9367 9979
rect 11882 9976 11888 9988
rect 11843 9948 11888 9976
rect 9309 9939 9367 9945
rect 11882 9936 11888 9948
rect 11940 9936 11946 9988
rect 13541 9979 13599 9985
rect 13541 9945 13553 9979
rect 13587 9945 13599 9979
rect 13541 9939 13599 9945
rect 8478 9908 8484 9920
rect 8036 9880 8484 9908
rect 8478 9868 8484 9880
rect 8536 9908 8542 9920
rect 8941 9911 8999 9917
rect 8941 9908 8953 9911
rect 8536 9880 8953 9908
rect 8536 9868 8542 9880
rect 8941 9877 8953 9880
rect 8987 9877 8999 9911
rect 8941 9871 8999 9877
rect 12986 9868 12992 9920
rect 13044 9908 13050 9920
rect 13556 9908 13584 9939
rect 16482 9936 16488 9988
rect 16540 9976 16546 9988
rect 17129 9979 17187 9985
rect 17129 9976 17141 9979
rect 16540 9948 17141 9976
rect 16540 9936 16546 9948
rect 17129 9945 17141 9948
rect 17175 9976 17187 9979
rect 21284 9976 21312 10007
rect 21910 10004 21916 10016
rect 21968 10004 21974 10056
rect 23216 10044 23244 10072
rect 23566 10044 23572 10056
rect 23216 10016 23572 10044
rect 23566 10004 23572 10016
rect 23624 10044 23630 10056
rect 24780 10044 24808 10075
rect 25038 10044 25044 10056
rect 23624 10016 25044 10044
rect 23624 10004 23630 10016
rect 25038 10004 25044 10016
rect 25096 10004 25102 10056
rect 17175 9948 21312 9976
rect 17175 9945 17187 9948
rect 17129 9939 17187 9945
rect 13044 9880 13584 9908
rect 13044 9868 13050 9880
rect 19242 9868 19248 9920
rect 19300 9908 19306 9920
rect 19429 9911 19487 9917
rect 19429 9908 19441 9911
rect 19300 9880 19441 9908
rect 19300 9868 19306 9880
rect 19429 9877 19441 9880
rect 19475 9877 19487 9911
rect 19429 9871 19487 9877
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 2041 9707 2099 9713
rect 2041 9673 2053 9707
rect 2087 9704 2099 9707
rect 2682 9704 2688 9716
rect 2087 9676 2688 9704
rect 2087 9673 2099 9676
rect 2041 9667 2099 9673
rect 1854 9596 1860 9648
rect 1912 9636 1918 9648
rect 2271 9639 2329 9645
rect 2271 9636 2283 9639
rect 1912 9608 2283 9636
rect 1912 9596 1918 9608
rect 2271 9605 2283 9608
rect 2317 9605 2329 9639
rect 2406 9636 2412 9648
rect 2367 9608 2412 9636
rect 2271 9599 2329 9605
rect 2406 9596 2412 9608
rect 2464 9596 2470 9648
rect 106 9528 112 9580
rect 164 9568 170 9580
rect 2516 9577 2544 9676
rect 2682 9664 2688 9676
rect 2740 9664 2746 9716
rect 3421 9707 3479 9713
rect 3421 9673 3433 9707
rect 3467 9704 3479 9707
rect 3835 9707 3893 9713
rect 3835 9704 3847 9707
rect 3467 9676 3847 9704
rect 3467 9673 3479 9676
rect 3421 9667 3479 9673
rect 3835 9673 3847 9676
rect 3881 9673 3893 9707
rect 3835 9667 3893 9673
rect 4154 9664 4160 9716
rect 4212 9704 4218 9716
rect 4709 9707 4767 9713
rect 4709 9704 4721 9707
rect 4212 9676 4721 9704
rect 4212 9664 4218 9676
rect 4709 9673 4721 9676
rect 4755 9673 4767 9707
rect 4709 9667 4767 9673
rect 10042 9664 10048 9716
rect 10100 9704 10106 9716
rect 10137 9707 10195 9713
rect 10137 9704 10149 9707
rect 10100 9676 10149 9704
rect 10100 9664 10106 9676
rect 10137 9673 10149 9676
rect 10183 9673 10195 9707
rect 10137 9667 10195 9673
rect 11422 9664 11428 9716
rect 11480 9704 11486 9716
rect 12161 9707 12219 9713
rect 12161 9704 12173 9707
rect 11480 9676 12173 9704
rect 11480 9664 11486 9676
rect 12161 9673 12173 9676
rect 12207 9673 12219 9707
rect 13630 9704 13636 9716
rect 13591 9676 13636 9704
rect 12161 9667 12219 9673
rect 3973 9639 4031 9645
rect 3973 9605 3985 9639
rect 4019 9636 4031 9639
rect 4019 9608 4200 9636
rect 4019 9605 4031 9608
rect 3973 9599 4031 9605
rect 2501 9571 2559 9577
rect 164 9540 2268 9568
rect 164 9528 170 9540
rect 1673 9503 1731 9509
rect 1673 9469 1685 9503
rect 1719 9500 1731 9503
rect 1946 9500 1952 9512
rect 1719 9472 1952 9500
rect 1719 9469 1731 9472
rect 1673 9463 1731 9469
rect 1946 9460 1952 9472
rect 2004 9460 2010 9512
rect 2130 9500 2136 9512
rect 2091 9472 2136 9500
rect 2130 9460 2136 9472
rect 2188 9460 2194 9512
rect 2240 9432 2268 9540
rect 2501 9537 2513 9571
rect 2547 9537 2559 9571
rect 2501 9531 2559 9537
rect 2590 9528 2596 9580
rect 2648 9568 2654 9580
rect 3421 9571 3479 9577
rect 3421 9568 3433 9571
rect 2648 9540 3433 9568
rect 2648 9528 2654 9540
rect 3421 9537 3433 9540
rect 3467 9537 3479 9571
rect 4062 9568 4068 9580
rect 4023 9540 4068 9568
rect 3421 9531 3479 9537
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 3237 9503 3295 9509
rect 3237 9469 3249 9503
rect 3283 9500 3295 9503
rect 3970 9500 3976 9512
rect 3283 9472 3976 9500
rect 3283 9469 3295 9472
rect 3237 9463 3295 9469
rect 3970 9460 3976 9472
rect 4028 9460 4034 9512
rect 4172 9500 4200 9608
rect 4246 9596 4252 9648
rect 4304 9636 4310 9648
rect 5077 9639 5135 9645
rect 5077 9636 5089 9639
rect 4304 9608 5089 9636
rect 4304 9596 4310 9608
rect 5077 9605 5089 9608
rect 5123 9605 5135 9639
rect 5077 9599 5135 9605
rect 9582 9596 9588 9648
rect 9640 9636 9646 9648
rect 9861 9639 9919 9645
rect 9861 9636 9873 9639
rect 9640 9608 9873 9636
rect 9640 9596 9646 9608
rect 9861 9605 9873 9608
rect 9907 9636 9919 9639
rect 10686 9636 10692 9648
rect 9907 9608 10692 9636
rect 9907 9605 9919 9608
rect 9861 9599 9919 9605
rect 10686 9596 10692 9608
rect 10744 9596 10750 9648
rect 11698 9596 11704 9648
rect 11756 9636 11762 9648
rect 11793 9639 11851 9645
rect 11793 9636 11805 9639
rect 11756 9608 11805 9636
rect 11756 9596 11762 9608
rect 11793 9605 11805 9608
rect 11839 9605 11851 9639
rect 11793 9599 11851 9605
rect 4433 9571 4491 9577
rect 4433 9537 4445 9571
rect 4479 9568 4491 9571
rect 4614 9568 4620 9580
rect 4479 9540 4620 9568
rect 4479 9537 4491 9540
rect 4433 9531 4491 9537
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 6730 9528 6736 9580
rect 6788 9568 6794 9580
rect 7374 9568 7380 9580
rect 6788 9540 6868 9568
rect 7335 9540 7380 9568
rect 6788 9528 6794 9540
rect 4338 9500 4344 9512
rect 4172 9472 4344 9500
rect 4338 9460 4344 9472
rect 4396 9460 4402 9512
rect 5074 9460 5080 9512
rect 5132 9500 5138 9512
rect 6840 9509 6868 9540
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 7558 9528 7564 9580
rect 7616 9568 7622 9580
rect 8294 9568 8300 9580
rect 7616 9540 8300 9568
rect 7616 9528 7622 9540
rect 8294 9528 8300 9540
rect 8352 9568 8358 9580
rect 8849 9571 8907 9577
rect 8849 9568 8861 9571
rect 8352 9540 8861 9568
rect 8352 9528 8358 9540
rect 8849 9537 8861 9540
rect 8895 9537 8907 9571
rect 10704 9568 10732 9596
rect 12176 9568 12204 9667
rect 13630 9664 13636 9676
rect 13688 9664 13694 9716
rect 15654 9664 15660 9716
rect 15712 9704 15718 9716
rect 18230 9704 18236 9716
rect 15712 9676 18236 9704
rect 15712 9664 15718 9676
rect 18230 9664 18236 9676
rect 18288 9664 18294 9716
rect 19518 9664 19524 9716
rect 19576 9704 19582 9716
rect 20993 9707 21051 9713
rect 20993 9704 21005 9707
rect 19576 9676 21005 9704
rect 19576 9664 19582 9676
rect 20993 9673 21005 9676
rect 21039 9673 21051 9707
rect 20993 9667 21051 9673
rect 13354 9596 13360 9648
rect 13412 9636 13418 9648
rect 13412 9608 13814 9636
rect 13412 9596 13418 9608
rect 12713 9571 12771 9577
rect 12713 9568 12725 9571
rect 10704 9540 11284 9568
rect 12176 9540 12725 9568
rect 8849 9531 8907 9537
rect 11256 9512 11284 9540
rect 12713 9537 12725 9540
rect 12759 9537 12771 9571
rect 12986 9568 12992 9580
rect 12947 9540 12992 9568
rect 12713 9531 12771 9537
rect 12986 9528 12992 9540
rect 13044 9528 13050 9580
rect 13786 9568 13814 9608
rect 18874 9596 18880 9648
rect 18932 9636 18938 9648
rect 21008 9636 21036 9667
rect 21910 9664 21916 9716
rect 21968 9704 21974 9716
rect 22738 9704 22744 9716
rect 21968 9676 22744 9704
rect 21968 9664 21974 9676
rect 22738 9664 22744 9676
rect 22796 9664 22802 9716
rect 25038 9704 25044 9716
rect 24999 9676 25044 9704
rect 25038 9664 25044 9676
rect 25096 9664 25102 9716
rect 25406 9704 25412 9716
rect 25367 9676 25412 9704
rect 25406 9664 25412 9676
rect 25464 9664 25470 9716
rect 23198 9636 23204 9648
rect 18932 9608 20392 9636
rect 21008 9608 23204 9636
rect 18932 9596 18938 9608
rect 20364 9580 20392 9608
rect 23198 9596 23204 9608
rect 23256 9596 23262 9648
rect 14277 9571 14335 9577
rect 14277 9568 14289 9571
rect 13786 9540 14289 9568
rect 14277 9537 14289 9540
rect 14323 9568 14335 9571
rect 14550 9568 14556 9580
rect 14323 9540 14556 9568
rect 14323 9537 14335 9540
rect 14277 9531 14335 9537
rect 14550 9528 14556 9540
rect 14608 9528 14614 9580
rect 14734 9568 14740 9580
rect 14695 9540 14740 9568
rect 14734 9528 14740 9540
rect 14792 9528 14798 9580
rect 15470 9528 15476 9580
rect 15528 9568 15534 9580
rect 15933 9571 15991 9577
rect 15933 9568 15945 9571
rect 15528 9540 15945 9568
rect 15528 9528 15534 9540
rect 15933 9537 15945 9540
rect 15979 9568 15991 9571
rect 18322 9568 18328 9580
rect 15979 9540 16896 9568
rect 18283 9540 18328 9568
rect 15979 9537 15991 9540
rect 15933 9531 15991 9537
rect 16868 9512 16896 9540
rect 18322 9528 18328 9540
rect 18380 9528 18386 9580
rect 20070 9568 20076 9580
rect 20031 9540 20076 9568
rect 20070 9528 20076 9540
rect 20128 9528 20134 9580
rect 20346 9568 20352 9580
rect 20259 9540 20352 9568
rect 20346 9528 20352 9540
rect 20404 9528 20410 9580
rect 22278 9568 22284 9580
rect 22239 9540 22284 9568
rect 22278 9528 22284 9540
rect 22336 9528 22342 9580
rect 22922 9528 22928 9580
rect 22980 9568 22986 9580
rect 24213 9571 24271 9577
rect 24213 9568 24225 9571
rect 22980 9540 24225 9568
rect 22980 9528 22986 9540
rect 24213 9537 24225 9540
rect 24259 9537 24271 9571
rect 24213 9531 24271 9537
rect 5261 9503 5319 9509
rect 5261 9500 5273 9503
rect 5132 9472 5273 9500
rect 5132 9460 5138 9472
rect 5261 9469 5273 9472
rect 5307 9500 5319 9503
rect 5813 9503 5871 9509
rect 5813 9500 5825 9503
rect 5307 9472 5825 9500
rect 5307 9469 5319 9472
rect 5261 9463 5319 9469
rect 5813 9469 5825 9472
rect 5859 9469 5871 9503
rect 5813 9463 5871 9469
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9469 6883 9503
rect 6825 9463 6883 9469
rect 7190 9460 7196 9512
rect 7248 9500 7254 9512
rect 7285 9503 7343 9509
rect 7285 9500 7297 9503
rect 7248 9472 7297 9500
rect 7248 9460 7254 9472
rect 7285 9469 7297 9472
rect 7331 9469 7343 9503
rect 7285 9463 7343 9469
rect 8202 9460 8208 9512
rect 8260 9500 8266 9512
rect 8389 9503 8447 9509
rect 8389 9500 8401 9503
rect 8260 9472 8401 9500
rect 8260 9460 8266 9472
rect 8389 9469 8401 9472
rect 8435 9469 8447 9503
rect 8389 9463 8447 9469
rect 8478 9460 8484 9512
rect 8536 9500 8542 9512
rect 8665 9503 8723 9509
rect 8536 9472 8581 9500
rect 8536 9460 8542 9472
rect 8665 9469 8677 9503
rect 8711 9469 8723 9503
rect 8665 9463 8723 9469
rect 10781 9503 10839 9509
rect 10781 9469 10793 9503
rect 10827 9469 10839 9503
rect 11238 9500 11244 9512
rect 11151 9472 11244 9500
rect 10781 9463 10839 9469
rect 2240 9404 3648 9432
rect 2038 9324 2044 9376
rect 2096 9364 2102 9376
rect 2777 9367 2835 9373
rect 2777 9364 2789 9367
rect 2096 9336 2789 9364
rect 2096 9324 2102 9336
rect 2777 9333 2789 9336
rect 2823 9333 2835 9367
rect 2777 9327 2835 9333
rect 3418 9324 3424 9376
rect 3476 9364 3482 9376
rect 3513 9367 3571 9373
rect 3513 9364 3525 9367
rect 3476 9336 3525 9364
rect 3476 9324 3482 9336
rect 3513 9333 3525 9336
rect 3559 9333 3571 9367
rect 3620 9364 3648 9404
rect 3694 9392 3700 9444
rect 3752 9432 3758 9444
rect 3752 9404 3797 9432
rect 4126 9404 5396 9432
rect 3752 9392 3758 9404
rect 4126 9364 4154 9404
rect 3620 9336 4154 9364
rect 5368 9364 5396 9404
rect 8294 9392 8300 9444
rect 8352 9432 8358 9444
rect 8680 9432 8708 9463
rect 9401 9435 9459 9441
rect 9401 9432 9413 9435
rect 8352 9404 9413 9432
rect 8352 9392 8358 9404
rect 9401 9401 9413 9404
rect 9447 9401 9459 9435
rect 9401 9395 9459 9401
rect 10796 9376 10824 9463
rect 11238 9460 11244 9472
rect 11296 9460 11302 9512
rect 15286 9460 15292 9512
rect 15344 9500 15350 9512
rect 16301 9503 16359 9509
rect 16301 9500 16313 9503
rect 15344 9472 16313 9500
rect 15344 9460 15350 9472
rect 16301 9469 16313 9472
rect 16347 9500 16359 9503
rect 16393 9503 16451 9509
rect 16393 9500 16405 9503
rect 16347 9472 16405 9500
rect 16347 9469 16359 9472
rect 16301 9463 16359 9469
rect 16393 9469 16405 9472
rect 16439 9469 16451 9503
rect 16850 9500 16856 9512
rect 16811 9472 16856 9500
rect 16393 9463 16451 9469
rect 16850 9460 16856 9472
rect 16908 9460 16914 9512
rect 21542 9500 21548 9512
rect 21376 9472 21548 9500
rect 11514 9432 11520 9444
rect 11475 9404 11520 9432
rect 11514 9392 11520 9404
rect 11572 9392 11578 9444
rect 12805 9435 12863 9441
rect 12805 9401 12817 9435
rect 12851 9401 12863 9435
rect 12805 9395 12863 9401
rect 14369 9435 14427 9441
rect 14369 9401 14381 9435
rect 14415 9401 14427 9435
rect 15562 9432 15568 9444
rect 15475 9404 15568 9432
rect 14369 9395 14427 9401
rect 5445 9367 5503 9373
rect 5445 9364 5457 9367
rect 5368 9336 5457 9364
rect 3513 9327 3571 9333
rect 5445 9333 5457 9336
rect 5491 9333 5503 9367
rect 5445 9327 5503 9333
rect 6362 9324 6368 9376
rect 6420 9364 6426 9376
rect 6457 9367 6515 9373
rect 6457 9364 6469 9367
rect 6420 9336 6469 9364
rect 6420 9324 6426 9336
rect 6457 9333 6469 9336
rect 6503 9364 6515 9367
rect 7742 9364 7748 9376
rect 6503 9336 7748 9364
rect 6503 9333 6515 9336
rect 6457 9327 6515 9333
rect 7742 9324 7748 9336
rect 7800 9324 7806 9376
rect 8018 9364 8024 9376
rect 7979 9336 8024 9364
rect 8018 9324 8024 9336
rect 8076 9324 8082 9376
rect 10689 9367 10747 9373
rect 10689 9333 10701 9367
rect 10735 9364 10747 9367
rect 10778 9364 10784 9376
rect 10735 9336 10784 9364
rect 10735 9333 10747 9336
rect 10689 9327 10747 9333
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 12618 9324 12624 9376
rect 12676 9364 12682 9376
rect 12820 9364 12848 9395
rect 13998 9364 14004 9376
rect 12676 9336 12848 9364
rect 13959 9336 14004 9364
rect 12676 9324 12682 9336
rect 13998 9324 14004 9336
rect 14056 9364 14062 9376
rect 14384 9364 14412 9395
rect 15562 9392 15568 9404
rect 15620 9432 15626 9444
rect 16482 9432 16488 9444
rect 15620 9404 16488 9432
rect 15620 9392 15626 9404
rect 16482 9392 16488 9404
rect 16540 9392 16546 9444
rect 17129 9435 17187 9441
rect 17129 9401 17141 9435
rect 17175 9432 17187 9435
rect 17770 9432 17776 9444
rect 17175 9404 17776 9432
rect 17175 9401 17187 9404
rect 17129 9395 17187 9401
rect 17770 9392 17776 9404
rect 17828 9392 17834 9444
rect 17865 9435 17923 9441
rect 17865 9401 17877 9435
rect 17911 9432 17923 9435
rect 17954 9432 17960 9444
rect 17911 9404 17960 9432
rect 17911 9401 17923 9404
rect 17865 9395 17923 9401
rect 17954 9392 17960 9404
rect 18012 9432 18018 9444
rect 18417 9435 18475 9441
rect 18417 9432 18429 9435
rect 18012 9404 18429 9432
rect 18012 9392 18018 9404
rect 18417 9401 18429 9404
rect 18463 9401 18475 9435
rect 18966 9432 18972 9444
rect 18927 9404 18972 9432
rect 18417 9395 18475 9401
rect 14056 9336 14412 9364
rect 18432 9364 18460 9395
rect 18966 9392 18972 9404
rect 19024 9392 19030 9444
rect 19889 9435 19947 9441
rect 19889 9401 19901 9435
rect 19935 9432 19947 9435
rect 20165 9435 20223 9441
rect 20165 9432 20177 9435
rect 19935 9404 20177 9432
rect 19935 9401 19947 9404
rect 19889 9395 19947 9401
rect 19996 9376 20024 9404
rect 20165 9401 20177 9404
rect 20211 9401 20223 9435
rect 20165 9395 20223 9401
rect 21376 9376 21404 9472
rect 21542 9460 21548 9472
rect 21600 9460 21606 9512
rect 22097 9503 22155 9509
rect 22097 9469 22109 9503
rect 22143 9500 22155 9503
rect 22738 9500 22744 9512
rect 22143 9472 22744 9500
rect 22143 9469 22155 9472
rect 22097 9463 22155 9469
rect 22738 9460 22744 9472
rect 22796 9460 22802 9512
rect 22830 9460 22836 9512
rect 22888 9500 22894 9512
rect 23385 9503 23443 9509
rect 23385 9500 23397 9503
rect 22888 9472 23397 9500
rect 22888 9460 22894 9472
rect 23385 9469 23397 9472
rect 23431 9500 23443 9503
rect 23661 9503 23719 9509
rect 23661 9500 23673 9503
rect 23431 9472 23673 9500
rect 23431 9469 23443 9472
rect 23385 9463 23443 9469
rect 23661 9469 23673 9472
rect 23707 9469 23719 9503
rect 24118 9500 24124 9512
rect 24079 9472 24124 9500
rect 23661 9463 23719 9469
rect 24118 9460 24124 9472
rect 24176 9460 24182 9512
rect 25130 9460 25136 9512
rect 25188 9500 25194 9512
rect 25225 9503 25283 9509
rect 25225 9500 25237 9503
rect 25188 9472 25237 9500
rect 25188 9460 25194 9472
rect 25225 9469 25237 9472
rect 25271 9500 25283 9503
rect 25777 9503 25835 9509
rect 25777 9500 25789 9503
rect 25271 9472 25789 9500
rect 25271 9469 25283 9472
rect 25225 9463 25283 9469
rect 25777 9469 25789 9472
rect 25823 9469 25835 9503
rect 25777 9463 25835 9469
rect 23474 9392 23480 9444
rect 23532 9432 23538 9444
rect 24673 9435 24731 9441
rect 24673 9432 24685 9435
rect 23532 9404 24685 9432
rect 23532 9392 23538 9404
rect 23676 9376 23704 9404
rect 24673 9401 24685 9404
rect 24719 9401 24731 9435
rect 24673 9395 24731 9401
rect 18598 9364 18604 9376
rect 18432 9336 18604 9364
rect 14056 9324 14062 9336
rect 18598 9324 18604 9336
rect 18656 9364 18662 9376
rect 19245 9367 19303 9373
rect 19245 9364 19257 9367
rect 18656 9336 19257 9364
rect 18656 9324 18662 9336
rect 19245 9333 19257 9336
rect 19291 9333 19303 9367
rect 19245 9327 19303 9333
rect 19978 9324 19984 9376
rect 20036 9324 20042 9376
rect 21358 9364 21364 9376
rect 21319 9336 21364 9364
rect 21358 9324 21364 9336
rect 21416 9324 21422 9376
rect 23658 9324 23664 9376
rect 23716 9324 23722 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 2225 9163 2283 9169
rect 2225 9129 2237 9163
rect 2271 9160 2283 9163
rect 2406 9160 2412 9172
rect 2271 9132 2412 9160
rect 2271 9129 2283 9132
rect 2225 9123 2283 9129
rect 2406 9120 2412 9132
rect 2464 9160 2470 9172
rect 3418 9160 3424 9172
rect 2464 9132 3424 9160
rect 2464 9120 2470 9132
rect 3418 9120 3424 9132
rect 3476 9160 3482 9172
rect 3694 9160 3700 9172
rect 3476 9132 3700 9160
rect 3476 9120 3482 9132
rect 3694 9120 3700 9132
rect 3752 9120 3758 9172
rect 5905 9163 5963 9169
rect 5905 9129 5917 9163
rect 5951 9160 5963 9163
rect 5994 9160 6000 9172
rect 5951 9132 6000 9160
rect 5951 9129 5963 9132
rect 5905 9123 5963 9129
rect 5994 9120 6000 9132
rect 6052 9120 6058 9172
rect 6365 9163 6423 9169
rect 6365 9129 6377 9163
rect 6411 9160 6423 9163
rect 6454 9160 6460 9172
rect 6411 9132 6460 9160
rect 6411 9129 6423 9132
rect 6365 9123 6423 9129
rect 6454 9120 6460 9132
rect 6512 9120 6518 9172
rect 6730 9120 6736 9172
rect 6788 9160 6794 9172
rect 7006 9160 7012 9172
rect 6788 9132 7012 9160
rect 6788 9120 6794 9132
rect 7006 9120 7012 9132
rect 7064 9160 7070 9172
rect 7469 9163 7527 9169
rect 7469 9160 7481 9163
rect 7064 9132 7481 9160
rect 7064 9120 7070 9132
rect 7469 9129 7481 9132
rect 7515 9129 7527 9163
rect 7469 9123 7527 9129
rect 9766 9120 9772 9172
rect 9824 9160 9830 9172
rect 10321 9163 10379 9169
rect 10321 9160 10333 9163
rect 9824 9132 10333 9160
rect 9824 9120 9830 9132
rect 10321 9129 10333 9132
rect 10367 9129 10379 9163
rect 10321 9123 10379 9129
rect 12161 9163 12219 9169
rect 12161 9129 12173 9163
rect 12207 9160 12219 9163
rect 13262 9160 13268 9172
rect 12207 9132 13268 9160
rect 12207 9129 12219 9132
rect 12161 9123 12219 9129
rect 13262 9120 13268 9132
rect 13320 9120 13326 9172
rect 13633 9163 13691 9169
rect 13633 9129 13645 9163
rect 13679 9160 13691 9163
rect 13998 9160 14004 9172
rect 13679 9132 14004 9160
rect 13679 9129 13691 9132
rect 13633 9123 13691 9129
rect 13998 9120 14004 9132
rect 14056 9120 14062 9172
rect 14550 9160 14556 9172
rect 14511 9132 14556 9160
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 16574 9160 16580 9172
rect 16535 9132 16580 9160
rect 16574 9120 16580 9132
rect 16632 9120 16638 9172
rect 17954 9160 17960 9172
rect 17915 9132 17960 9160
rect 17954 9120 17960 9132
rect 18012 9120 18018 9172
rect 18506 9120 18512 9172
rect 18564 9160 18570 9172
rect 18601 9163 18659 9169
rect 18601 9160 18613 9163
rect 18564 9132 18613 9160
rect 18564 9120 18570 9132
rect 18601 9129 18613 9132
rect 18647 9129 18659 9163
rect 21082 9160 21088 9172
rect 21043 9132 21088 9160
rect 18601 9123 18659 9129
rect 21082 9120 21088 9132
rect 21140 9120 21146 9172
rect 22738 9160 22744 9172
rect 22699 9132 22744 9160
rect 22738 9120 22744 9132
rect 22796 9120 22802 9172
rect 23106 9160 23112 9172
rect 23067 9132 23112 9160
rect 23106 9120 23112 9132
rect 23164 9120 23170 9172
rect 24118 9160 24124 9172
rect 24079 9132 24124 9160
rect 24118 9120 24124 9132
rect 24176 9120 24182 9172
rect 3145 9095 3203 9101
rect 3145 9061 3157 9095
rect 3191 9092 3203 9095
rect 3878 9092 3884 9104
rect 3191 9064 3884 9092
rect 3191 9061 3203 9064
rect 3145 9055 3203 9061
rect 3878 9052 3884 9064
rect 3936 9052 3942 9104
rect 4338 9052 4344 9104
rect 4396 9092 4402 9104
rect 10689 9095 10747 9101
rect 10689 9092 10701 9095
rect 4396 9064 10701 9092
rect 4396 9052 4402 9064
rect 10689 9061 10701 9064
rect 10735 9061 10747 9095
rect 10689 9055 10747 9061
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 2038 9024 2044 9036
rect 1443 8996 2044 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2038 8984 2044 8996
rect 2096 8984 2102 9036
rect 2409 9027 2467 9033
rect 2409 8993 2421 9027
rect 2455 8993 2467 9027
rect 2409 8987 2467 8993
rect 2424 8956 2452 8987
rect 2498 8984 2504 9036
rect 2556 9024 2562 9036
rect 2685 9027 2743 9033
rect 2685 9024 2697 9027
rect 2556 8996 2697 9024
rect 2556 8984 2562 8996
rect 2685 8993 2697 8996
rect 2731 8993 2743 9027
rect 2685 8987 2743 8993
rect 6454 8984 6460 9036
rect 6512 9024 6518 9036
rect 6512 8996 6557 9024
rect 6512 8984 6518 8996
rect 6730 8984 6736 9036
rect 6788 9024 6794 9036
rect 8021 9027 8079 9033
rect 6788 8996 6833 9024
rect 6788 8984 6794 8996
rect 8021 8993 8033 9027
rect 8067 9024 8079 9027
rect 8110 9024 8116 9036
rect 8067 8996 8116 9024
rect 8067 8993 8079 8996
rect 8021 8987 8079 8993
rect 8110 8984 8116 8996
rect 8168 8984 8174 9036
rect 8294 9024 8300 9036
rect 8255 8996 8300 9024
rect 8294 8984 8300 8996
rect 8352 8984 8358 9036
rect 9858 9024 9864 9036
rect 9819 8996 9864 9024
rect 9858 8984 9864 8996
rect 9916 8984 9922 9036
rect 10704 9024 10732 9055
rect 10962 9052 10968 9104
rect 11020 9092 11026 9104
rect 11235 9095 11293 9101
rect 11235 9092 11247 9095
rect 11020 9064 11247 9092
rect 11020 9052 11026 9064
rect 11235 9061 11247 9064
rect 11281 9092 11293 9095
rect 12434 9092 12440 9104
rect 11281 9064 12440 9092
rect 11281 9061 11293 9064
rect 11235 9055 11293 9061
rect 12434 9052 12440 9064
rect 12492 9092 12498 9104
rect 13034 9095 13092 9101
rect 13034 9092 13046 9095
rect 12492 9064 13046 9092
rect 12492 9052 12498 9064
rect 13034 9061 13046 9064
rect 13080 9061 13092 9095
rect 13034 9055 13092 9061
rect 13446 9052 13452 9104
rect 13504 9092 13510 9104
rect 14185 9095 14243 9101
rect 14185 9092 14197 9095
rect 13504 9064 14197 9092
rect 13504 9052 13510 9064
rect 14185 9061 14197 9064
rect 14231 9092 14243 9095
rect 14274 9092 14280 9104
rect 14231 9064 14280 9092
rect 14231 9061 14243 9064
rect 14185 9055 14243 9061
rect 14274 9052 14280 9064
rect 14332 9052 14338 9104
rect 17218 9052 17224 9104
rect 17276 9092 17282 9104
rect 19150 9101 19156 9104
rect 17358 9095 17416 9101
rect 17358 9092 17370 9095
rect 17276 9064 17370 9092
rect 17276 9052 17282 9064
rect 17358 9061 17370 9064
rect 17404 9092 17416 9095
rect 19106 9095 19156 9101
rect 19106 9092 19118 9095
rect 17404 9064 19118 9092
rect 17404 9061 17416 9064
rect 17358 9055 17416 9061
rect 19106 9061 19118 9064
rect 19152 9061 19156 9095
rect 19106 9055 19156 9061
rect 19150 9052 19156 9055
rect 19208 9052 19214 9104
rect 20070 9092 20076 9104
rect 20031 9064 20076 9092
rect 20070 9052 20076 9064
rect 20128 9052 20134 9104
rect 20717 9095 20775 9101
rect 20717 9061 20729 9095
rect 20763 9092 20775 9095
rect 21174 9092 21180 9104
rect 20763 9064 21180 9092
rect 20763 9061 20775 9064
rect 20717 9055 20775 9061
rect 21174 9052 21180 9064
rect 21232 9052 21238 9104
rect 21634 9092 21640 9104
rect 21595 9064 21640 9092
rect 21634 9052 21640 9064
rect 21692 9052 21698 9104
rect 23290 9052 23296 9104
rect 23348 9092 23354 9104
rect 24719 9095 24777 9101
rect 24719 9092 24731 9095
rect 23348 9064 24731 9092
rect 23348 9052 23354 9064
rect 24719 9061 24731 9064
rect 24765 9061 24777 9095
rect 24719 9055 24777 9061
rect 10873 9027 10931 9033
rect 10873 9024 10885 9027
rect 10704 8996 10885 9024
rect 10873 8993 10885 8996
rect 10919 8993 10931 9027
rect 11698 9024 11704 9036
rect 10873 8987 10931 8993
rect 11256 8996 11704 9024
rect 3786 8956 3792 8968
rect 2424 8928 3792 8956
rect 3786 8916 3792 8928
rect 3844 8916 3850 8968
rect 3878 8916 3884 8968
rect 3936 8956 3942 8968
rect 4430 8956 4436 8968
rect 3936 8928 3981 8956
rect 4391 8928 4436 8956
rect 3936 8916 3942 8928
rect 4430 8916 4436 8928
rect 4488 8956 4494 8968
rect 5077 8959 5135 8965
rect 5077 8956 5089 8959
rect 4488 8928 5089 8956
rect 4488 8916 4494 8928
rect 5077 8925 5089 8928
rect 5123 8956 5135 8959
rect 5445 8959 5503 8965
rect 5445 8956 5457 8959
rect 5123 8928 5457 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 5445 8925 5457 8928
rect 5491 8925 5503 8959
rect 6914 8956 6920 8968
rect 6875 8928 6920 8956
rect 5445 8919 5503 8925
rect 6914 8916 6920 8928
rect 6972 8916 6978 8968
rect 8757 8959 8815 8965
rect 8757 8925 8769 8959
rect 8803 8956 8815 8959
rect 9674 8956 9680 8968
rect 8803 8928 9680 8956
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 9674 8916 9680 8928
rect 9732 8956 9738 8968
rect 11256 8956 11284 8996
rect 11698 8984 11704 8996
rect 11756 8984 11762 9036
rect 15654 9024 15660 9036
rect 15615 8996 15660 9024
rect 15654 8984 15660 8996
rect 15712 8984 15718 9036
rect 15838 8984 15844 9036
rect 15896 9024 15902 9036
rect 15933 9027 15991 9033
rect 15933 9024 15945 9027
rect 15896 8996 15945 9024
rect 15896 8984 15902 8996
rect 15933 8993 15945 8996
rect 15979 8993 15991 9027
rect 15933 8987 15991 8993
rect 17770 8984 17776 9036
rect 17828 9024 17834 9036
rect 18782 9024 18788 9036
rect 17828 8996 18788 9024
rect 17828 8984 17834 8996
rect 18782 8984 18788 8996
rect 18840 8984 18846 9036
rect 19705 9027 19763 9033
rect 19705 8993 19717 9027
rect 19751 9024 19763 9027
rect 19978 9024 19984 9036
rect 19751 8996 19984 9024
rect 19751 8993 19763 8996
rect 19705 8987 19763 8993
rect 19978 8984 19984 8996
rect 20036 8984 20042 9036
rect 22922 8984 22928 9036
rect 22980 9024 22986 9036
rect 23017 9027 23075 9033
rect 23017 9024 23029 9027
rect 22980 8996 23029 9024
rect 22980 8984 22986 8996
rect 23017 8993 23029 8996
rect 23063 8993 23075 9027
rect 23017 8987 23075 8993
rect 23474 8984 23480 9036
rect 23532 9024 23538 9036
rect 24632 9027 24690 9033
rect 23532 8996 23577 9024
rect 23532 8984 23538 8996
rect 24632 8993 24644 9027
rect 24678 9024 24690 9027
rect 24854 9024 24860 9036
rect 24678 8996 24860 9024
rect 24678 8993 24690 8996
rect 24632 8987 24690 8993
rect 24854 8984 24860 8996
rect 24912 8984 24918 9036
rect 9732 8928 11284 8956
rect 9732 8916 9738 8928
rect 11514 8916 11520 8968
rect 11572 8956 11578 8968
rect 12713 8959 12771 8965
rect 12713 8956 12725 8959
rect 11572 8928 12725 8956
rect 11572 8916 11578 8928
rect 12713 8925 12725 8928
rect 12759 8956 12771 8959
rect 13538 8956 13544 8968
rect 12759 8928 13544 8956
rect 12759 8925 12771 8928
rect 12713 8919 12771 8925
rect 13538 8916 13544 8928
rect 13596 8916 13602 8968
rect 16206 8956 16212 8968
rect 16167 8928 16212 8956
rect 16206 8916 16212 8928
rect 16264 8916 16270 8968
rect 17034 8956 17040 8968
rect 16995 8928 17040 8956
rect 17034 8916 17040 8928
rect 17092 8916 17098 8968
rect 20346 8916 20352 8968
rect 20404 8956 20410 8968
rect 21545 8959 21603 8965
rect 21545 8956 21557 8959
rect 20404 8928 21557 8956
rect 20404 8916 20410 8928
rect 21545 8925 21557 8928
rect 21591 8925 21603 8959
rect 21545 8919 21603 8925
rect 21821 8959 21879 8965
rect 21821 8925 21833 8959
rect 21867 8925 21879 8959
rect 21821 8919 21879 8925
rect 2501 8891 2559 8897
rect 2501 8857 2513 8891
rect 2547 8888 2559 8891
rect 3418 8888 3424 8900
rect 2547 8860 3424 8888
rect 2547 8857 2559 8860
rect 2501 8851 2559 8857
rect 3418 8848 3424 8860
rect 3476 8848 3482 8900
rect 4154 8848 4160 8900
rect 4212 8897 4218 8900
rect 4212 8891 4261 8897
rect 4212 8857 4215 8891
rect 4249 8857 4261 8891
rect 4212 8851 4261 8857
rect 4212 8848 4218 8851
rect 6362 8848 6368 8900
rect 6420 8888 6426 8900
rect 6549 8891 6607 8897
rect 6549 8888 6561 8891
rect 6420 8860 6561 8888
rect 6420 8848 6426 8860
rect 6549 8857 6561 8860
rect 6595 8888 6607 8891
rect 8110 8888 8116 8900
rect 6595 8860 7972 8888
rect 8071 8860 8116 8888
rect 6595 8857 6607 8860
rect 6549 8851 6607 8857
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 1670 8820 1676 8832
rect 1627 8792 1676 8820
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 1670 8780 1676 8792
rect 1728 8780 1734 8832
rect 1854 8780 1860 8832
rect 1912 8820 1918 8832
rect 3697 8823 3755 8829
rect 3697 8820 3709 8823
rect 1912 8792 3709 8820
rect 1912 8780 1918 8792
rect 3697 8789 3709 8792
rect 3743 8820 3755 8823
rect 4062 8820 4068 8832
rect 3743 8792 4068 8820
rect 3743 8789 3755 8792
rect 3697 8783 3755 8789
rect 4062 8780 4068 8792
rect 4120 8780 4126 8832
rect 4338 8820 4344 8832
rect 4299 8792 4344 8820
rect 4338 8780 4344 8792
rect 4396 8780 4402 8832
rect 4522 8820 4528 8832
rect 4483 8792 4528 8820
rect 4522 8780 4528 8792
rect 4580 8780 4586 8832
rect 7834 8820 7840 8832
rect 7795 8792 7840 8820
rect 7834 8780 7840 8792
rect 7892 8780 7898 8832
rect 7944 8820 7972 8860
rect 8110 8848 8116 8860
rect 8168 8848 8174 8900
rect 10045 8891 10103 8897
rect 10045 8857 10057 8891
rect 10091 8888 10103 8891
rect 12894 8888 12900 8900
rect 10091 8860 12900 8888
rect 10091 8857 10103 8860
rect 10045 8851 10103 8857
rect 12894 8848 12900 8860
rect 12952 8848 12958 8900
rect 16942 8888 16948 8900
rect 16855 8860 16948 8888
rect 16942 8848 16948 8860
rect 17000 8888 17006 8900
rect 17000 8860 19334 8888
rect 17000 8848 17006 8860
rect 8478 8820 8484 8832
rect 7944 8792 8484 8820
rect 8478 8780 8484 8792
rect 8536 8820 8542 8832
rect 9033 8823 9091 8829
rect 9033 8820 9045 8823
rect 8536 8792 9045 8820
rect 8536 8780 8542 8792
rect 9033 8789 9045 8792
rect 9079 8789 9091 8823
rect 11790 8820 11796 8832
rect 11751 8792 11796 8820
rect 9033 8783 9091 8789
rect 11790 8780 11796 8792
rect 11848 8780 11854 8832
rect 18322 8820 18328 8832
rect 18283 8792 18328 8820
rect 18322 8780 18328 8792
rect 18380 8780 18386 8832
rect 19306 8820 19334 8860
rect 21174 8848 21180 8900
rect 21232 8888 21238 8900
rect 21836 8888 21864 8919
rect 22738 8916 22744 8968
rect 22796 8956 22802 8968
rect 23566 8956 23572 8968
rect 22796 8928 23572 8956
rect 22796 8916 22802 8928
rect 23566 8916 23572 8928
rect 23624 8916 23630 8968
rect 21232 8860 21864 8888
rect 21232 8848 21238 8860
rect 21266 8820 21272 8832
rect 19306 8792 21272 8820
rect 21266 8780 21272 8792
rect 21324 8780 21330 8832
rect 21836 8820 21864 8860
rect 22462 8848 22468 8900
rect 22520 8888 22526 8900
rect 23014 8888 23020 8900
rect 22520 8860 23020 8888
rect 22520 8848 22526 8860
rect 23014 8848 23020 8860
rect 23072 8848 23078 8900
rect 23934 8820 23940 8832
rect 21836 8792 23940 8820
rect 23934 8780 23940 8792
rect 23992 8780 23998 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 2130 8576 2136 8628
rect 2188 8616 2194 8628
rect 2409 8619 2467 8625
rect 2409 8616 2421 8619
rect 2188 8588 2421 8616
rect 2188 8576 2194 8588
rect 2409 8585 2421 8588
rect 2455 8585 2467 8619
rect 3142 8616 3148 8628
rect 3103 8588 3148 8616
rect 2409 8579 2467 8585
rect 2424 8548 2452 8579
rect 3142 8576 3148 8588
rect 3200 8576 3206 8628
rect 4065 8619 4123 8625
rect 4065 8585 4077 8619
rect 4111 8616 4123 8619
rect 4338 8616 4344 8628
rect 4111 8588 4344 8616
rect 4111 8585 4123 8588
rect 4065 8579 4123 8585
rect 4338 8576 4344 8588
rect 4396 8576 4402 8628
rect 5442 8576 5448 8628
rect 5500 8616 5506 8628
rect 5537 8619 5595 8625
rect 5537 8616 5549 8619
rect 5500 8588 5549 8616
rect 5500 8576 5506 8588
rect 5537 8585 5549 8588
rect 5583 8616 5595 8619
rect 6730 8616 6736 8628
rect 5583 8588 6736 8616
rect 5583 8585 5595 8588
rect 5537 8579 5595 8585
rect 6730 8576 6736 8588
rect 6788 8616 6794 8628
rect 7190 8616 7196 8628
rect 6788 8588 7196 8616
rect 6788 8576 6794 8588
rect 7190 8576 7196 8588
rect 7248 8616 7254 8628
rect 8021 8619 8079 8625
rect 8021 8616 8033 8619
rect 7248 8588 8033 8616
rect 7248 8576 7254 8588
rect 8021 8585 8033 8588
rect 8067 8616 8079 8619
rect 8294 8616 8300 8628
rect 8067 8588 8300 8616
rect 8067 8585 8079 8588
rect 8021 8579 8079 8585
rect 8294 8576 8300 8588
rect 8352 8576 8358 8628
rect 10689 8619 10747 8625
rect 10689 8585 10701 8619
rect 10735 8616 10747 8619
rect 10962 8616 10968 8628
rect 10735 8588 10968 8616
rect 10735 8585 10747 8588
rect 10689 8579 10747 8585
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 12253 8619 12311 8625
rect 12253 8585 12265 8619
rect 12299 8616 12311 8619
rect 12434 8616 12440 8628
rect 12299 8588 12440 8616
rect 12299 8585 12311 8588
rect 12253 8579 12311 8585
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 17218 8616 17224 8628
rect 17179 8588 17224 8616
rect 17218 8576 17224 8588
rect 17276 8576 17282 8628
rect 19150 8616 19156 8628
rect 19111 8588 19156 8616
rect 19150 8576 19156 8588
rect 19208 8576 19214 8628
rect 19613 8619 19671 8625
rect 19613 8585 19625 8619
rect 19659 8616 19671 8619
rect 19978 8616 19984 8628
rect 19659 8588 19984 8616
rect 19659 8585 19671 8588
rect 19613 8579 19671 8585
rect 19978 8576 19984 8588
rect 20036 8576 20042 8628
rect 20901 8619 20959 8625
rect 20901 8585 20913 8619
rect 20947 8616 20959 8619
rect 21634 8616 21640 8628
rect 20947 8588 21640 8616
rect 20947 8585 20959 8588
rect 20901 8579 20959 8585
rect 21634 8576 21640 8588
rect 21692 8616 21698 8628
rect 22281 8619 22339 8625
rect 22281 8616 22293 8619
rect 21692 8588 22293 8616
rect 21692 8576 21698 8588
rect 22281 8585 22293 8588
rect 22327 8585 22339 8619
rect 22281 8579 22339 8585
rect 22649 8619 22707 8625
rect 22649 8585 22661 8619
rect 22695 8616 22707 8619
rect 23106 8616 23112 8628
rect 22695 8588 23112 8616
rect 22695 8585 22707 8588
rect 22649 8579 22707 8585
rect 3878 8548 3884 8560
rect 2424 8520 3884 8548
rect 3878 8508 3884 8520
rect 3936 8508 3942 8560
rect 4154 8508 4160 8560
rect 4212 8548 4218 8560
rect 5169 8551 5227 8557
rect 5169 8548 5181 8551
rect 4212 8520 5181 8548
rect 4212 8508 4218 8520
rect 5169 8517 5181 8520
rect 5215 8517 5227 8551
rect 5169 8511 5227 8517
rect 5905 8551 5963 8557
rect 5905 8517 5917 8551
rect 5951 8548 5963 8551
rect 7650 8548 7656 8560
rect 5951 8520 7656 8548
rect 5951 8517 5963 8520
rect 5905 8511 5963 8517
rect 7650 8508 7656 8520
rect 7708 8508 7714 8560
rect 11425 8551 11483 8557
rect 11425 8517 11437 8551
rect 11471 8548 11483 8551
rect 12986 8548 12992 8560
rect 11471 8520 12992 8548
rect 11471 8517 11483 8520
rect 11425 8511 11483 8517
rect 12986 8508 12992 8520
rect 13044 8508 13050 8560
rect 14458 8508 14464 8560
rect 14516 8548 14522 8560
rect 16114 8548 16120 8560
rect 14516 8520 16120 8548
rect 14516 8508 14522 8520
rect 16114 8508 16120 8520
rect 16172 8548 16178 8560
rect 17678 8548 17684 8560
rect 16172 8520 17684 8548
rect 16172 8508 16178 8520
rect 4249 8483 4307 8489
rect 4249 8449 4261 8483
rect 4295 8480 4307 8483
rect 4706 8480 4712 8492
rect 4295 8452 4712 8480
rect 4295 8449 4307 8452
rect 4249 8443 4307 8449
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 9953 8483 10011 8489
rect 9953 8449 9965 8483
rect 9999 8480 10011 8483
rect 12437 8483 12495 8489
rect 12437 8480 12449 8483
rect 9999 8452 12449 8480
rect 9999 8449 10011 8452
rect 9953 8443 10011 8449
rect 12437 8449 12449 8452
rect 12483 8480 12495 8483
rect 13633 8483 13691 8489
rect 13633 8480 13645 8483
rect 12483 8452 13645 8480
rect 12483 8449 12495 8452
rect 12437 8443 12495 8449
rect 13633 8449 13645 8452
rect 13679 8449 13691 8483
rect 14274 8480 14280 8492
rect 14235 8452 14280 8480
rect 13633 8443 13691 8449
rect 14274 8440 14280 8452
rect 14332 8440 14338 8492
rect 14550 8480 14556 8492
rect 14511 8452 14556 8480
rect 14550 8440 14556 8452
rect 14608 8480 14614 8492
rect 14734 8480 14740 8492
rect 14608 8452 14740 8480
rect 14608 8440 14614 8452
rect 14734 8440 14740 8452
rect 14792 8440 14798 8492
rect 1486 8412 1492 8424
rect 1447 8384 1492 8412
rect 1486 8372 1492 8384
rect 1544 8372 1550 8424
rect 2961 8415 3019 8421
rect 2961 8381 2973 8415
rect 3007 8412 3019 8415
rect 5718 8412 5724 8424
rect 3007 8384 3648 8412
rect 5679 8384 5724 8412
rect 3007 8381 3019 8384
rect 2961 8375 3019 8381
rect 1857 8279 1915 8285
rect 1857 8245 1869 8279
rect 1903 8276 1915 8279
rect 1946 8276 1952 8288
rect 1903 8248 1952 8276
rect 1903 8245 1915 8248
rect 1857 8239 1915 8245
rect 1946 8236 1952 8248
rect 2004 8236 2010 8288
rect 2590 8236 2596 8288
rect 2648 8276 2654 8288
rect 2866 8276 2872 8288
rect 2648 8248 2872 8276
rect 2648 8236 2654 8248
rect 2866 8236 2872 8248
rect 2924 8236 2930 8288
rect 3620 8285 3648 8384
rect 5718 8372 5724 8384
rect 5776 8372 5782 8424
rect 7374 8412 7380 8424
rect 7335 8384 7380 8412
rect 7374 8372 7380 8384
rect 7432 8412 7438 8424
rect 8110 8412 8116 8424
rect 7432 8384 8116 8412
rect 7432 8372 7438 8384
rect 8110 8372 8116 8384
rect 8168 8412 8174 8424
rect 8389 8415 8447 8421
rect 8389 8412 8401 8415
rect 8168 8384 8401 8412
rect 8168 8372 8174 8384
rect 8389 8381 8401 8384
rect 8435 8381 8447 8415
rect 8389 8375 8447 8381
rect 8662 8372 8668 8424
rect 8720 8412 8726 8424
rect 9217 8415 9275 8421
rect 9217 8412 9229 8415
rect 8720 8384 9229 8412
rect 8720 8372 8726 8384
rect 9217 8381 9229 8384
rect 9263 8381 9275 8415
rect 9217 8375 9275 8381
rect 4338 8304 4344 8356
rect 4396 8344 4402 8356
rect 4890 8344 4896 8356
rect 4396 8316 4441 8344
rect 4851 8316 4896 8344
rect 4396 8304 4402 8316
rect 4890 8304 4896 8316
rect 4948 8304 4954 8356
rect 6362 8304 6368 8356
rect 6420 8344 6426 8356
rect 6825 8347 6883 8353
rect 6825 8344 6837 8347
rect 6420 8316 6837 8344
rect 6420 8304 6426 8316
rect 6825 8313 6837 8316
rect 6871 8313 6883 8347
rect 6825 8307 6883 8313
rect 9232 8288 9260 8375
rect 9582 8372 9588 8424
rect 9640 8412 9646 8424
rect 16500 8421 16528 8520
rect 17678 8508 17684 8520
rect 17736 8508 17742 8560
rect 18966 8508 18972 8560
rect 19024 8548 19030 8560
rect 20349 8551 20407 8557
rect 20349 8548 20361 8551
rect 19024 8520 20361 8548
rect 19024 8508 19030 8520
rect 20349 8517 20361 8520
rect 20395 8517 20407 8551
rect 20349 8511 20407 8517
rect 16945 8483 17003 8489
rect 16945 8449 16957 8483
rect 16991 8480 17003 8483
rect 17034 8480 17040 8492
rect 16991 8452 17040 8480
rect 16991 8449 17003 8452
rect 16945 8443 17003 8449
rect 17034 8440 17040 8452
rect 17092 8480 17098 8492
rect 17589 8483 17647 8489
rect 17589 8480 17601 8483
rect 17092 8452 17601 8480
rect 17092 8440 17098 8452
rect 17589 8449 17601 8452
rect 17635 8449 17647 8483
rect 18874 8480 18880 8492
rect 18835 8452 18880 8480
rect 17589 8443 17647 8449
rect 18874 8440 18880 8452
rect 18932 8440 18938 8492
rect 19797 8483 19855 8489
rect 19797 8449 19809 8483
rect 19843 8480 19855 8483
rect 20070 8480 20076 8492
rect 19843 8452 20076 8480
rect 19843 8449 19855 8452
rect 19797 8443 19855 8449
rect 20070 8440 20076 8452
rect 20128 8440 20134 8492
rect 21361 8483 21419 8489
rect 21361 8449 21373 8483
rect 21407 8480 21419 8483
rect 22664 8480 22692 8579
rect 23106 8576 23112 8588
rect 23164 8576 23170 8628
rect 25406 8616 25412 8628
rect 25367 8588 25412 8616
rect 25406 8576 25412 8588
rect 25464 8576 25470 8628
rect 23382 8548 23388 8560
rect 23343 8520 23388 8548
rect 23382 8508 23388 8520
rect 23440 8508 23446 8560
rect 21407 8452 22692 8480
rect 21407 8449 21419 8452
rect 21361 8443 21419 8449
rect 23934 8440 23940 8492
rect 23992 8480 23998 8492
rect 24029 8483 24087 8489
rect 24029 8480 24041 8483
rect 23992 8452 24041 8480
rect 23992 8440 23998 8452
rect 24029 8449 24041 8452
rect 24075 8449 24087 8483
rect 24029 8443 24087 8449
rect 9677 8415 9735 8421
rect 9677 8412 9689 8415
rect 9640 8384 9689 8412
rect 9640 8372 9646 8384
rect 9677 8381 9689 8384
rect 9723 8381 9735 8415
rect 9677 8375 9735 8381
rect 13357 8415 13415 8421
rect 13357 8381 13369 8415
rect 13403 8412 13415 8415
rect 14001 8415 14059 8421
rect 14001 8412 14013 8415
rect 13403 8384 14013 8412
rect 13403 8381 13415 8384
rect 13357 8375 13415 8381
rect 14001 8381 14013 8384
rect 14047 8381 14059 8415
rect 14001 8375 14059 8381
rect 16485 8415 16543 8421
rect 16485 8381 16497 8415
rect 16531 8381 16543 8415
rect 16485 8375 16543 8381
rect 9858 8304 9864 8356
rect 9916 8344 9922 8356
rect 10321 8347 10379 8353
rect 10321 8344 10333 8347
rect 9916 8316 10333 8344
rect 9916 8304 9922 8316
rect 10321 8313 10333 8316
rect 10367 8344 10379 8347
rect 10686 8344 10692 8356
rect 10367 8316 10692 8344
rect 10367 8313 10379 8316
rect 10321 8307 10379 8313
rect 10686 8304 10692 8316
rect 10744 8304 10750 8356
rect 10870 8344 10876 8356
rect 10831 8316 10876 8344
rect 10870 8304 10876 8316
rect 10928 8304 10934 8356
rect 10965 8347 11023 8353
rect 10965 8313 10977 8347
rect 11011 8344 11023 8347
rect 11790 8344 11796 8356
rect 11011 8316 11796 8344
rect 11011 8313 11023 8316
rect 10965 8307 11023 8313
rect 11790 8304 11796 8316
rect 11848 8304 11854 8356
rect 12434 8304 12440 8356
rect 12492 8344 12498 8356
rect 12758 8347 12816 8353
rect 12758 8344 12770 8347
rect 12492 8316 12770 8344
rect 12492 8304 12498 8316
rect 12758 8313 12770 8316
rect 12804 8313 12816 8347
rect 12758 8307 12816 8313
rect 3605 8279 3663 8285
rect 3605 8245 3617 8279
rect 3651 8276 3663 8279
rect 3878 8276 3884 8288
rect 3651 8248 3884 8276
rect 3651 8245 3663 8248
rect 3605 8239 3663 8245
rect 3878 8236 3884 8248
rect 3936 8236 3942 8288
rect 6454 8236 6460 8288
rect 6512 8276 6518 8288
rect 6549 8279 6607 8285
rect 6549 8276 6561 8279
rect 6512 8248 6561 8276
rect 6512 8236 6518 8248
rect 6549 8245 6561 8248
rect 6595 8276 6607 8279
rect 8018 8276 8024 8288
rect 6595 8248 8024 8276
rect 6595 8245 6607 8248
rect 6549 8239 6607 8245
rect 8018 8236 8024 8248
rect 8076 8236 8082 8288
rect 9125 8279 9183 8285
rect 9125 8245 9137 8279
rect 9171 8276 9183 8279
rect 9214 8276 9220 8288
rect 9171 8248 9220 8276
rect 9171 8245 9183 8248
rect 9125 8239 9183 8245
rect 9214 8236 9220 8248
rect 9272 8236 9278 8288
rect 14016 8276 14044 8375
rect 16574 8372 16580 8424
rect 16632 8412 16638 8424
rect 16669 8415 16727 8421
rect 16669 8412 16681 8415
rect 16632 8384 16681 8412
rect 16632 8372 16638 8384
rect 16669 8381 16681 8384
rect 16715 8412 16727 8415
rect 16850 8412 16856 8424
rect 16715 8384 16856 8412
rect 16715 8381 16727 8384
rect 16669 8375 16727 8381
rect 16850 8372 16856 8384
rect 16908 8372 16914 8424
rect 22370 8372 22376 8424
rect 22428 8412 22434 8424
rect 23106 8412 23112 8424
rect 22428 8384 23112 8412
rect 22428 8372 22434 8384
rect 23106 8372 23112 8384
rect 23164 8372 23170 8424
rect 25222 8412 25228 8424
rect 25135 8384 25228 8412
rect 25222 8372 25228 8384
rect 25280 8412 25286 8424
rect 25777 8415 25835 8421
rect 25777 8412 25789 8415
rect 25280 8384 25789 8412
rect 25280 8372 25286 8384
rect 25777 8381 25789 8384
rect 25823 8381 25835 8415
rect 25777 8375 25835 8381
rect 14369 8347 14427 8353
rect 14369 8313 14381 8347
rect 14415 8313 14427 8347
rect 14369 8307 14427 8313
rect 14384 8276 14412 8307
rect 17402 8304 17408 8356
rect 17460 8344 17466 8356
rect 18233 8347 18291 8353
rect 18233 8344 18245 8347
rect 17460 8316 18245 8344
rect 17460 8304 17466 8316
rect 18233 8313 18245 8316
rect 18279 8313 18291 8347
rect 18233 8307 18291 8313
rect 18322 8304 18328 8356
rect 18380 8344 18386 8356
rect 19889 8347 19947 8353
rect 18380 8316 18425 8344
rect 18380 8304 18386 8316
rect 19889 8313 19901 8347
rect 19935 8344 19947 8347
rect 19978 8344 19984 8356
rect 19935 8316 19984 8344
rect 19935 8313 19947 8316
rect 19889 8307 19947 8313
rect 19978 8304 19984 8316
rect 20036 8304 20042 8356
rect 21682 8347 21740 8353
rect 21682 8344 21694 8347
rect 21192 8316 21694 8344
rect 14016 8248 14412 8276
rect 15565 8279 15623 8285
rect 15565 8245 15577 8279
rect 15611 8276 15623 8279
rect 15654 8276 15660 8288
rect 15611 8248 15660 8276
rect 15611 8245 15623 8248
rect 15565 8239 15623 8245
rect 15654 8236 15660 8248
rect 15712 8276 15718 8288
rect 15930 8276 15936 8288
rect 15712 8248 15936 8276
rect 15712 8236 15718 8248
rect 15930 8236 15936 8248
rect 15988 8236 15994 8288
rect 19150 8236 19156 8288
rect 19208 8276 19214 8288
rect 20990 8276 20996 8288
rect 19208 8248 20996 8276
rect 19208 8236 19214 8248
rect 20990 8236 20996 8248
rect 21048 8276 21054 8288
rect 21192 8285 21220 8316
rect 21682 8313 21694 8316
rect 21728 8344 21740 8347
rect 22738 8344 22744 8356
rect 21728 8316 22744 8344
rect 21728 8313 21740 8316
rect 21682 8307 21740 8313
rect 22738 8304 22744 8316
rect 22796 8304 22802 8356
rect 23753 8347 23811 8353
rect 23753 8313 23765 8347
rect 23799 8313 23811 8347
rect 23753 8307 23811 8313
rect 21177 8279 21235 8285
rect 21177 8276 21189 8279
rect 21048 8248 21189 8276
rect 21048 8236 21054 8248
rect 21177 8245 21189 8248
rect 21223 8245 21235 8279
rect 21177 8239 21235 8245
rect 21358 8236 21364 8288
rect 21416 8276 21422 8288
rect 22922 8276 22928 8288
rect 21416 8248 22928 8276
rect 21416 8236 21422 8248
rect 22922 8236 22928 8248
rect 22980 8276 22986 8288
rect 23017 8279 23075 8285
rect 23017 8276 23029 8279
rect 22980 8248 23029 8276
rect 22980 8236 22986 8248
rect 23017 8245 23029 8248
rect 23063 8245 23075 8279
rect 23017 8239 23075 8245
rect 23382 8236 23388 8288
rect 23440 8276 23446 8288
rect 23474 8276 23480 8288
rect 23440 8248 23480 8276
rect 23440 8236 23446 8248
rect 23474 8236 23480 8248
rect 23532 8236 23538 8288
rect 23768 8276 23796 8307
rect 23842 8304 23848 8356
rect 23900 8344 23906 8356
rect 23900 8316 23945 8344
rect 23900 8304 23906 8316
rect 24118 8276 24124 8288
rect 23768 8248 24124 8276
rect 24118 8236 24124 8248
rect 24176 8236 24182 8288
rect 24765 8279 24823 8285
rect 24765 8245 24777 8279
rect 24811 8276 24823 8279
rect 24854 8276 24860 8288
rect 24811 8248 24860 8276
rect 24811 8245 24823 8248
rect 24765 8239 24823 8245
rect 24854 8236 24860 8248
rect 24912 8276 24918 8288
rect 25406 8276 25412 8288
rect 24912 8248 25412 8276
rect 24912 8236 24918 8248
rect 25406 8236 25412 8248
rect 25464 8236 25470 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 1854 8072 1860 8084
rect 1627 8044 1860 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 1854 8032 1860 8044
rect 1912 8032 1918 8084
rect 2038 8032 2044 8084
rect 2096 8072 2102 8084
rect 2225 8075 2283 8081
rect 2225 8072 2237 8075
rect 2096 8044 2237 8072
rect 2096 8032 2102 8044
rect 2225 8041 2237 8044
rect 2271 8041 2283 8075
rect 2225 8035 2283 8041
rect 3142 8032 3148 8084
rect 3200 8072 3206 8084
rect 3510 8072 3516 8084
rect 3200 8044 3516 8072
rect 3200 8032 3206 8044
rect 3510 8032 3516 8044
rect 3568 8072 3574 8084
rect 4062 8072 4068 8084
rect 3568 8044 4068 8072
rect 3568 8032 3574 8044
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 5718 8072 5724 8084
rect 4245 8044 5724 8072
rect 3602 7964 3608 8016
rect 3660 8004 3666 8016
rect 4245 8004 4273 8044
rect 5718 8032 5724 8044
rect 5776 8072 5782 8084
rect 6917 8075 6975 8081
rect 6917 8072 6929 8075
rect 5776 8044 6929 8072
rect 5776 8032 5782 8044
rect 6917 8041 6929 8044
rect 6963 8041 6975 8075
rect 6917 8035 6975 8041
rect 7929 8075 7987 8081
rect 7929 8041 7941 8075
rect 7975 8072 7987 8075
rect 8202 8072 8208 8084
rect 7975 8044 8208 8072
rect 7975 8041 7987 8044
rect 7929 8035 7987 8041
rect 3660 7976 4273 8004
rect 4318 8007 4376 8013
rect 3660 7964 3666 7976
rect 4318 7973 4330 8007
rect 4364 8004 4376 8007
rect 4430 8004 4436 8016
rect 4364 7976 4436 8004
rect 4364 7973 4376 7976
rect 4318 7967 4376 7973
rect 4430 7964 4436 7976
rect 4488 7964 4494 8016
rect 5169 8007 5227 8013
rect 5169 7973 5181 8007
rect 5215 8004 5227 8007
rect 5353 8007 5411 8013
rect 5353 8004 5365 8007
rect 5215 7976 5365 8004
rect 5215 7973 5227 7976
rect 5169 7967 5227 7973
rect 5353 7973 5365 7976
rect 5399 8004 5411 8007
rect 6086 8004 6092 8016
rect 5399 7976 6092 8004
rect 5399 7973 5411 7976
rect 5353 7967 5411 7973
rect 6086 7964 6092 7976
rect 6144 8004 6150 8016
rect 7944 8004 7972 8035
rect 8202 8032 8208 8044
rect 8260 8032 8266 8084
rect 9309 8075 9367 8081
rect 9309 8041 9321 8075
rect 9355 8072 9367 8075
rect 9582 8072 9588 8084
rect 9355 8044 9588 8072
rect 9355 8041 9367 8044
rect 9309 8035 9367 8041
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 13538 8072 13544 8084
rect 13499 8044 13544 8072
rect 13538 8032 13544 8044
rect 13596 8032 13602 8084
rect 15562 8072 15568 8084
rect 15523 8044 15568 8072
rect 15562 8032 15568 8044
rect 15620 8032 15626 8084
rect 17313 8075 17371 8081
rect 17313 8041 17325 8075
rect 17359 8072 17371 8075
rect 17402 8072 17408 8084
rect 17359 8044 17408 8072
rect 17359 8041 17371 8044
rect 17313 8035 17371 8041
rect 17402 8032 17408 8044
rect 17460 8032 17466 8084
rect 18322 8072 18328 8084
rect 18283 8044 18328 8072
rect 18322 8032 18328 8044
rect 18380 8072 18386 8084
rect 18380 8044 19380 8072
rect 18380 8032 18386 8044
rect 6144 7976 7972 8004
rect 8757 8007 8815 8013
rect 6144 7964 6150 7976
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 1946 7936 1952 7948
rect 1443 7908 1952 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 1946 7896 1952 7908
rect 2004 7896 2010 7948
rect 2682 7936 2688 7948
rect 2643 7908 2688 7936
rect 2682 7896 2688 7908
rect 2740 7896 2746 7948
rect 2958 7936 2964 7948
rect 2919 7908 2964 7936
rect 2958 7896 2964 7908
rect 3016 7896 3022 7948
rect 3418 7896 3424 7948
rect 3476 7936 3482 7948
rect 6273 7939 6331 7945
rect 6273 7936 6285 7939
rect 3476 7908 6285 7936
rect 3476 7896 3482 7908
rect 6273 7905 6285 7908
rect 6319 7936 6331 7939
rect 6362 7936 6368 7948
rect 6319 7908 6368 7936
rect 6319 7905 6331 7908
rect 6273 7899 6331 7905
rect 6362 7896 6368 7908
rect 6420 7896 6426 7948
rect 6472 7945 6500 7976
rect 8757 7973 8769 8007
rect 8803 8004 8815 8007
rect 9858 8004 9864 8016
rect 8803 7976 9864 8004
rect 8803 7973 8815 7976
rect 8757 7967 8815 7973
rect 9858 7964 9864 7976
rect 9916 7964 9922 8016
rect 10686 7964 10692 8016
rect 10744 8004 10750 8016
rect 10744 7976 11376 8004
rect 10744 7964 10750 7976
rect 6457 7939 6515 7945
rect 6457 7905 6469 7939
rect 6503 7905 6515 7939
rect 6730 7936 6736 7948
rect 6691 7908 6736 7936
rect 6457 7899 6515 7905
rect 6730 7896 6736 7908
rect 6788 7936 6794 7948
rect 7834 7936 7840 7948
rect 6788 7908 7840 7936
rect 6788 7896 6794 7908
rect 7834 7896 7840 7908
rect 7892 7896 7898 7948
rect 8018 7936 8024 7948
rect 7979 7908 8024 7936
rect 8018 7896 8024 7908
rect 8076 7896 8082 7948
rect 8294 7936 8300 7948
rect 8255 7908 8300 7936
rect 8294 7896 8300 7908
rect 8352 7896 8358 7948
rect 9674 7936 9680 7948
rect 9635 7908 9680 7936
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 10594 7896 10600 7948
rect 10652 7936 10658 7948
rect 10781 7939 10839 7945
rect 10781 7936 10793 7939
rect 10652 7908 10793 7936
rect 10652 7896 10658 7908
rect 10781 7905 10793 7908
rect 10827 7905 10839 7939
rect 11238 7936 11244 7948
rect 11199 7908 11244 7936
rect 10781 7899 10839 7905
rect 11238 7896 11244 7908
rect 11296 7896 11302 7948
rect 11348 7936 11376 7976
rect 12434 7964 12440 8016
rect 12492 8004 12498 8016
rect 12666 8007 12724 8013
rect 12666 8004 12678 8007
rect 12492 7976 12678 8004
rect 12492 7964 12498 7976
rect 12666 7973 12678 7976
rect 12712 7973 12724 8007
rect 12666 7967 12724 7973
rect 12986 7964 12992 8016
rect 13044 8004 13050 8016
rect 13446 8004 13452 8016
rect 13044 7976 13452 8004
rect 13044 7964 13050 7976
rect 13446 7964 13452 7976
rect 13504 8004 13510 8016
rect 13909 8007 13967 8013
rect 13909 8004 13921 8007
rect 13504 7976 13921 8004
rect 13504 7964 13510 7976
rect 13909 7973 13921 7976
rect 13955 7973 13967 8007
rect 13909 7967 13967 7973
rect 17218 7964 17224 8016
rect 17276 8004 17282 8016
rect 17726 8007 17784 8013
rect 17726 8004 17738 8007
rect 17276 7976 17738 8004
rect 17276 7964 17282 7976
rect 17726 7973 17738 7976
rect 17772 7973 17784 8007
rect 18782 8004 18788 8016
rect 18743 7976 18788 8004
rect 17726 7967 17784 7973
rect 18782 7964 18788 7976
rect 18840 7964 18846 8016
rect 19352 8013 19380 8044
rect 20346 8032 20352 8084
rect 20404 8072 20410 8084
rect 20625 8075 20683 8081
rect 20625 8072 20637 8075
rect 20404 8044 20637 8072
rect 20404 8032 20410 8044
rect 20625 8041 20637 8044
rect 20671 8072 20683 8075
rect 20671 8044 21680 8072
rect 20671 8041 20683 8044
rect 20625 8035 20683 8041
rect 19337 8007 19395 8013
rect 19337 7973 19349 8007
rect 19383 8004 19395 8007
rect 19426 8004 19432 8016
rect 19383 7976 19432 8004
rect 19383 7973 19395 7976
rect 19337 7967 19395 7973
rect 19426 7964 19432 7976
rect 19484 7964 19490 8016
rect 21082 8004 21088 8016
rect 21043 7976 21088 8004
rect 21082 7964 21088 7976
rect 21140 7964 21146 8016
rect 21652 8013 21680 8044
rect 24026 8032 24032 8084
rect 24084 8072 24090 8084
rect 24627 8075 24685 8081
rect 24627 8072 24639 8075
rect 24084 8044 24639 8072
rect 24084 8032 24090 8044
rect 24627 8041 24639 8044
rect 24673 8041 24685 8075
rect 24627 8035 24685 8041
rect 21637 8007 21695 8013
rect 21637 7973 21649 8007
rect 21683 7973 21695 8007
rect 21637 7967 21695 7973
rect 22738 7964 22744 8016
rect 22796 8004 22802 8016
rect 23062 8007 23120 8013
rect 23062 8004 23074 8007
rect 22796 7976 23074 8004
rect 22796 7964 22802 7976
rect 23062 7973 23074 7976
rect 23108 7973 23120 8007
rect 23062 7967 23120 7973
rect 14090 7936 14096 7948
rect 11348 7908 14096 7936
rect 14090 7896 14096 7908
rect 14148 7896 14154 7948
rect 15565 7939 15623 7945
rect 15565 7905 15577 7939
rect 15611 7905 15623 7939
rect 15565 7899 15623 7905
rect 15841 7939 15899 7945
rect 15841 7905 15853 7939
rect 15887 7936 15899 7939
rect 16390 7936 16396 7948
rect 15887 7908 16396 7936
rect 15887 7905 15899 7908
rect 15841 7899 15899 7905
rect 3145 7871 3203 7877
rect 3145 7837 3157 7871
rect 3191 7868 3203 7871
rect 3510 7868 3516 7880
rect 3191 7840 3516 7868
rect 3191 7837 3203 7840
rect 3145 7831 3203 7837
rect 3510 7828 3516 7840
rect 3568 7868 3574 7880
rect 4065 7871 4123 7877
rect 4065 7868 4077 7871
rect 3568 7840 4077 7868
rect 3568 7828 3574 7840
rect 4065 7837 4077 7840
rect 4111 7837 4123 7871
rect 4065 7831 4123 7837
rect 4154 7828 4160 7880
rect 4212 7868 4218 7880
rect 4430 7868 4436 7880
rect 4212 7840 4436 7868
rect 4212 7828 4218 7840
rect 4430 7828 4436 7840
rect 4488 7828 4494 7880
rect 11517 7871 11575 7877
rect 11517 7837 11529 7871
rect 11563 7868 11575 7871
rect 12158 7868 12164 7880
rect 11563 7840 12164 7868
rect 11563 7837 11575 7840
rect 11517 7831 11575 7837
rect 12158 7828 12164 7840
rect 12216 7868 12222 7880
rect 12345 7871 12403 7877
rect 12345 7868 12357 7871
rect 12216 7840 12357 7868
rect 12216 7828 12222 7840
rect 12345 7837 12357 7840
rect 12391 7837 12403 7871
rect 15580 7868 15608 7899
rect 16390 7896 16396 7908
rect 16448 7896 16454 7948
rect 23661 7939 23719 7945
rect 23661 7905 23673 7939
rect 23707 7936 23719 7939
rect 23842 7936 23848 7948
rect 23707 7908 23848 7936
rect 23707 7905 23719 7908
rect 23661 7899 23719 7905
rect 23842 7896 23848 7908
rect 23900 7936 23906 7948
rect 24305 7939 24363 7945
rect 24305 7936 24317 7939
rect 23900 7908 24317 7936
rect 23900 7896 23906 7908
rect 24305 7905 24317 7908
rect 24351 7905 24363 7939
rect 24305 7899 24363 7905
rect 24556 7939 24614 7945
rect 24556 7905 24568 7939
rect 24602 7936 24614 7939
rect 24670 7936 24676 7948
rect 24602 7908 24676 7936
rect 24602 7905 24614 7908
rect 24556 7899 24614 7905
rect 24670 7896 24676 7908
rect 24728 7896 24734 7948
rect 16114 7868 16120 7880
rect 15580 7840 16120 7868
rect 12345 7831 12403 7837
rect 16114 7828 16120 7840
rect 16172 7828 16178 7880
rect 17402 7868 17408 7880
rect 17363 7840 17408 7868
rect 17402 7828 17408 7840
rect 17460 7828 17466 7880
rect 19245 7871 19303 7877
rect 19245 7837 19257 7871
rect 19291 7868 19303 7871
rect 19334 7868 19340 7880
rect 19291 7840 19340 7868
rect 19291 7837 19303 7840
rect 19245 7831 19303 7837
rect 19334 7828 19340 7840
rect 19392 7828 19398 7880
rect 19521 7871 19579 7877
rect 19521 7837 19533 7871
rect 19567 7837 19579 7871
rect 19521 7831 19579 7837
rect 842 7760 848 7812
rect 900 7800 906 7812
rect 1486 7800 1492 7812
rect 900 7772 1492 7800
rect 900 7760 906 7772
rect 1486 7760 1492 7772
rect 1544 7800 1550 7812
rect 1857 7803 1915 7809
rect 1857 7800 1869 7803
rect 1544 7772 1869 7800
rect 1544 7760 1550 7772
rect 1857 7769 1869 7772
rect 1903 7769 1915 7803
rect 1857 7763 1915 7769
rect 3694 7760 3700 7812
rect 3752 7800 3758 7812
rect 5169 7803 5227 7809
rect 5169 7800 5181 7803
rect 3752 7772 5181 7800
rect 3752 7760 3758 7772
rect 5169 7769 5181 7772
rect 5215 7769 5227 7803
rect 5169 7763 5227 7769
rect 6362 7760 6368 7812
rect 6420 7800 6426 7812
rect 6549 7803 6607 7809
rect 6549 7800 6561 7803
rect 6420 7772 6561 7800
rect 6420 7760 6426 7772
rect 6549 7769 6561 7772
rect 6595 7800 6607 7803
rect 7374 7800 7380 7812
rect 6595 7772 7380 7800
rect 6595 7769 6607 7772
rect 6549 7763 6607 7769
rect 7374 7760 7380 7772
rect 7432 7800 7438 7812
rect 7469 7803 7527 7809
rect 7469 7800 7481 7803
rect 7432 7772 7481 7800
rect 7432 7760 7438 7772
rect 7469 7769 7481 7772
rect 7515 7800 7527 7803
rect 8113 7803 8171 7809
rect 8113 7800 8125 7803
rect 7515 7772 8125 7800
rect 7515 7769 7527 7772
rect 7469 7763 7527 7769
rect 8113 7769 8125 7772
rect 8159 7800 8171 7803
rect 8202 7800 8208 7812
rect 8159 7772 8208 7800
rect 8159 7769 8171 7772
rect 8113 7763 8171 7769
rect 8202 7760 8208 7772
rect 8260 7760 8266 7812
rect 9766 7760 9772 7812
rect 9824 7800 9830 7812
rect 10597 7803 10655 7809
rect 10597 7800 10609 7803
rect 9824 7772 10609 7800
rect 9824 7760 9830 7772
rect 10597 7769 10609 7772
rect 10643 7800 10655 7803
rect 10870 7800 10876 7812
rect 10643 7772 10876 7800
rect 10643 7769 10655 7772
rect 10597 7763 10655 7769
rect 10870 7760 10876 7772
rect 10928 7760 10934 7812
rect 12250 7760 12256 7812
rect 12308 7800 12314 7812
rect 15013 7803 15071 7809
rect 15013 7800 15025 7803
rect 12308 7772 15025 7800
rect 12308 7760 12314 7772
rect 15013 7769 15025 7772
rect 15059 7800 15071 7803
rect 15838 7800 15844 7812
rect 15059 7772 15844 7800
rect 15059 7769 15071 7772
rect 15013 7763 15071 7769
rect 15838 7760 15844 7772
rect 15896 7760 15902 7812
rect 16482 7760 16488 7812
rect 16540 7800 16546 7812
rect 18782 7800 18788 7812
rect 16540 7772 18788 7800
rect 16540 7760 16546 7772
rect 18782 7760 18788 7772
rect 18840 7760 18846 7812
rect 18966 7760 18972 7812
rect 19024 7800 19030 7812
rect 19536 7800 19564 7831
rect 20714 7828 20720 7880
rect 20772 7868 20778 7880
rect 20993 7871 21051 7877
rect 20993 7868 21005 7871
rect 20772 7840 21005 7868
rect 20772 7828 20778 7840
rect 20993 7837 21005 7840
rect 21039 7837 21051 7871
rect 20993 7831 21051 7837
rect 22741 7871 22799 7877
rect 22741 7837 22753 7871
rect 22787 7837 22799 7871
rect 22741 7831 22799 7837
rect 19024 7772 19564 7800
rect 19024 7760 19030 7772
rect 3881 7735 3939 7741
rect 3881 7701 3893 7735
rect 3927 7732 3939 7735
rect 3970 7732 3976 7744
rect 3927 7704 3976 7732
rect 3927 7701 3939 7704
rect 3881 7695 3939 7701
rect 3970 7692 3976 7704
rect 4028 7692 4034 7744
rect 4338 7692 4344 7744
rect 4396 7732 4402 7744
rect 4985 7735 5043 7741
rect 4985 7732 4997 7735
rect 4396 7704 4997 7732
rect 4396 7692 4402 7704
rect 4985 7701 4997 7704
rect 5031 7701 5043 7735
rect 4985 7695 5043 7701
rect 7742 7692 7748 7744
rect 7800 7732 7806 7744
rect 9861 7735 9919 7741
rect 9861 7732 9873 7735
rect 7800 7704 9873 7732
rect 7800 7692 7806 7704
rect 9861 7701 9873 7704
rect 9907 7732 9919 7735
rect 9950 7732 9956 7744
rect 9907 7704 9956 7732
rect 9907 7701 9919 7704
rect 9861 7695 9919 7701
rect 9950 7692 9956 7704
rect 10008 7692 10014 7744
rect 13262 7732 13268 7744
rect 13223 7704 13268 7732
rect 13262 7692 13268 7704
rect 13320 7692 13326 7744
rect 13538 7692 13544 7744
rect 13596 7732 13602 7744
rect 14277 7735 14335 7741
rect 14277 7732 14289 7735
rect 13596 7704 14289 7732
rect 13596 7692 13602 7704
rect 14277 7701 14289 7704
rect 14323 7701 14335 7735
rect 14277 7695 14335 7701
rect 16393 7735 16451 7741
rect 16393 7701 16405 7735
rect 16439 7732 16451 7735
rect 16574 7732 16580 7744
rect 16439 7704 16580 7732
rect 16439 7701 16451 7704
rect 16393 7695 16451 7701
rect 16574 7692 16580 7704
rect 16632 7692 16638 7744
rect 20070 7692 20076 7744
rect 20128 7732 20134 7744
rect 20165 7735 20223 7741
rect 20165 7732 20177 7735
rect 20128 7704 20177 7732
rect 20128 7692 20134 7704
rect 20165 7701 20177 7704
rect 20211 7701 20223 7735
rect 22002 7732 22008 7744
rect 21963 7704 22008 7732
rect 20165 7695 20223 7701
rect 22002 7692 22008 7704
rect 22060 7692 22066 7744
rect 22649 7735 22707 7741
rect 22649 7701 22661 7735
rect 22695 7732 22707 7735
rect 22756 7732 22784 7831
rect 23750 7732 23756 7744
rect 22695 7704 23756 7732
rect 22695 7701 22707 7704
rect 22649 7695 22707 7701
rect 23750 7692 23756 7704
rect 23808 7692 23814 7744
rect 24029 7735 24087 7741
rect 24029 7701 24041 7735
rect 24075 7732 24087 7735
rect 24118 7732 24124 7744
rect 24075 7704 24124 7732
rect 24075 7701 24087 7704
rect 24029 7695 24087 7701
rect 24118 7692 24124 7704
rect 24176 7692 24182 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1578 7528 1584 7540
rect 1539 7500 1584 7528
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 1946 7528 1952 7540
rect 1907 7500 1952 7528
rect 1946 7488 1952 7500
rect 2004 7488 2010 7540
rect 4062 7488 4068 7540
rect 4120 7528 4126 7540
rect 5905 7531 5963 7537
rect 5905 7528 5917 7531
rect 4120 7500 5917 7528
rect 4120 7488 4126 7500
rect 5905 7497 5917 7500
rect 5951 7497 5963 7531
rect 7190 7528 7196 7540
rect 7151 7500 7196 7528
rect 5905 7491 5963 7497
rect 7190 7488 7196 7500
rect 7248 7488 7254 7540
rect 7282 7488 7288 7540
rect 7340 7528 7346 7540
rect 7469 7531 7527 7537
rect 7469 7528 7481 7531
rect 7340 7500 7481 7528
rect 7340 7488 7346 7500
rect 7469 7497 7481 7500
rect 7515 7497 7527 7531
rect 9674 7528 9680 7540
rect 9635 7500 9680 7528
rect 7469 7491 7527 7497
rect 9674 7488 9680 7500
rect 9732 7488 9738 7540
rect 12158 7528 12164 7540
rect 12119 7500 12164 7528
rect 12158 7488 12164 7500
rect 12216 7488 12222 7540
rect 12434 7488 12440 7540
rect 12492 7528 12498 7540
rect 12621 7531 12679 7537
rect 12621 7528 12633 7531
rect 12492 7500 12633 7528
rect 12492 7488 12498 7500
rect 12621 7497 12633 7500
rect 12667 7497 12679 7531
rect 13262 7528 13268 7540
rect 13223 7500 13268 7528
rect 12621 7491 12679 7497
rect 13262 7488 13268 7500
rect 13320 7488 13326 7540
rect 14090 7488 14096 7540
rect 14148 7528 14154 7540
rect 14369 7531 14427 7537
rect 14369 7528 14381 7531
rect 14148 7500 14381 7528
rect 14148 7488 14154 7500
rect 14369 7497 14381 7500
rect 14415 7497 14427 7531
rect 14369 7491 14427 7497
rect 16025 7531 16083 7537
rect 16025 7497 16037 7531
rect 16071 7528 16083 7531
rect 16114 7528 16120 7540
rect 16071 7500 16120 7528
rect 16071 7497 16083 7500
rect 16025 7491 16083 7497
rect 16114 7488 16120 7500
rect 16172 7488 16178 7540
rect 16390 7528 16396 7540
rect 16303 7500 16396 7528
rect 16390 7488 16396 7500
rect 16448 7528 16454 7540
rect 17494 7528 17500 7540
rect 16448 7500 17500 7528
rect 16448 7488 16454 7500
rect 17494 7488 17500 7500
rect 17552 7488 17558 7540
rect 19426 7528 19432 7540
rect 19387 7500 19432 7528
rect 19426 7488 19432 7500
rect 19484 7488 19490 7540
rect 21082 7488 21088 7540
rect 21140 7528 21146 7540
rect 21453 7531 21511 7537
rect 21453 7528 21465 7531
rect 21140 7500 21465 7528
rect 21140 7488 21146 7500
rect 21453 7497 21465 7500
rect 21499 7497 21511 7531
rect 21453 7491 21511 7497
rect 22738 7488 22744 7540
rect 22796 7528 22802 7540
rect 23017 7531 23075 7537
rect 23017 7528 23029 7531
rect 22796 7500 23029 7528
rect 22796 7488 22802 7500
rect 23017 7497 23029 7500
rect 23063 7497 23075 7531
rect 23017 7491 23075 7497
rect 2501 7463 2559 7469
rect 2501 7429 2513 7463
rect 2547 7460 2559 7463
rect 2682 7460 2688 7472
rect 2547 7432 2688 7460
rect 2547 7429 2559 7432
rect 2501 7423 2559 7429
rect 2682 7420 2688 7432
rect 2740 7460 2746 7472
rect 5350 7460 5356 7472
rect 2740 7432 5356 7460
rect 2740 7420 2746 7432
rect 5350 7420 5356 7432
rect 5408 7420 5414 7472
rect 5629 7463 5687 7469
rect 5629 7429 5641 7463
rect 5675 7460 5687 7463
rect 8386 7460 8392 7472
rect 5675 7432 8392 7460
rect 5675 7429 5687 7432
rect 5629 7423 5687 7429
rect 3694 7352 3700 7404
rect 3752 7392 3758 7404
rect 5442 7392 5448 7404
rect 3752 7364 5448 7392
rect 3752 7352 3758 7364
rect 5442 7352 5448 7364
rect 5500 7352 5506 7404
rect 1118 7284 1124 7336
rect 1176 7324 1182 7336
rect 1397 7327 1455 7333
rect 1397 7324 1409 7327
rect 1176 7296 1409 7324
rect 1176 7284 1182 7296
rect 1397 7293 1409 7296
rect 1443 7293 1455 7327
rect 1397 7287 1455 7293
rect 2869 7327 2927 7333
rect 2869 7293 2881 7327
rect 2915 7293 2927 7327
rect 3142 7324 3148 7336
rect 3103 7296 3148 7324
rect 2869 7287 2927 7293
rect 1762 7216 1768 7268
rect 1820 7256 1826 7268
rect 2884 7256 2912 7287
rect 3142 7284 3148 7296
rect 3200 7284 3206 7336
rect 4246 7324 4252 7336
rect 4207 7296 4252 7324
rect 4246 7284 4252 7296
rect 4304 7284 4310 7336
rect 4709 7327 4767 7333
rect 4709 7293 4721 7327
rect 4755 7324 4767 7327
rect 4798 7324 4804 7336
rect 4755 7296 4804 7324
rect 4755 7293 4767 7296
rect 4709 7287 4767 7293
rect 4798 7284 4804 7296
rect 4856 7284 4862 7336
rect 5736 7333 5764 7432
rect 8386 7420 8392 7432
rect 8444 7420 8450 7472
rect 12894 7420 12900 7472
rect 12952 7460 12958 7472
rect 12952 7432 14872 7460
rect 12952 7420 12958 7432
rect 8202 7352 8208 7404
rect 8260 7392 8266 7404
rect 9309 7395 9367 7401
rect 9309 7392 9321 7395
rect 8260 7364 9321 7392
rect 8260 7352 8266 7364
rect 5721 7327 5779 7333
rect 5721 7293 5733 7327
rect 5767 7293 5779 7327
rect 5721 7287 5779 7293
rect 7285 7327 7343 7333
rect 7285 7293 7297 7327
rect 7331 7324 7343 7327
rect 7558 7324 7564 7336
rect 7331 7296 7564 7324
rect 7331 7293 7343 7296
rect 7285 7287 7343 7293
rect 7558 7284 7564 7296
rect 7616 7284 7622 7336
rect 8018 7284 8024 7336
rect 8076 7324 8082 7336
rect 8113 7327 8171 7333
rect 8113 7324 8125 7327
rect 8076 7296 8125 7324
rect 8076 7284 8082 7296
rect 8113 7293 8125 7296
rect 8159 7324 8171 7327
rect 8294 7324 8300 7336
rect 8159 7296 8300 7324
rect 8159 7293 8171 7296
rect 8113 7287 8171 7293
rect 8294 7284 8300 7296
rect 8352 7284 8358 7336
rect 8404 7333 8432 7364
rect 9309 7361 9321 7364
rect 9355 7361 9367 7395
rect 9309 7355 9367 7361
rect 9398 7352 9404 7404
rect 9456 7392 9462 7404
rect 9950 7392 9956 7404
rect 9456 7364 9956 7392
rect 9456 7352 9462 7364
rect 9950 7352 9956 7364
rect 10008 7392 10014 7404
rect 10594 7392 10600 7404
rect 10008 7364 10600 7392
rect 10008 7352 10014 7364
rect 10594 7352 10600 7364
rect 10652 7352 10658 7404
rect 13446 7392 13452 7404
rect 13407 7364 13452 7392
rect 13446 7352 13452 7364
rect 13504 7352 13510 7404
rect 8389 7327 8447 7333
rect 8389 7293 8401 7327
rect 8435 7293 8447 7327
rect 8389 7287 8447 7293
rect 8573 7327 8631 7333
rect 8573 7293 8585 7327
rect 8619 7293 8631 7327
rect 10778 7324 10784 7336
rect 8573 7287 8631 7293
rect 10244 7296 10784 7324
rect 3326 7256 3332 7268
rect 1820 7228 3332 7256
rect 1820 7216 1826 7228
rect 3326 7216 3332 7228
rect 3384 7216 3390 7268
rect 3697 7259 3755 7265
rect 3697 7225 3709 7259
rect 3743 7256 3755 7259
rect 6270 7256 6276 7268
rect 3743 7228 6276 7256
rect 3743 7225 3755 7228
rect 3697 7219 3755 7225
rect 2130 7148 2136 7200
rect 2188 7188 2194 7200
rect 2685 7191 2743 7197
rect 2685 7188 2697 7191
rect 2188 7160 2697 7188
rect 2188 7148 2194 7160
rect 2685 7157 2697 7160
rect 2731 7157 2743 7191
rect 2685 7151 2743 7157
rect 2958 7148 2964 7200
rect 3016 7188 3022 7200
rect 3712 7188 3740 7219
rect 6270 7216 6276 7228
rect 6328 7216 6334 7268
rect 7834 7216 7840 7268
rect 7892 7256 7898 7268
rect 8588 7256 8616 7287
rect 9030 7256 9036 7268
rect 7892 7228 8616 7256
rect 8991 7228 9036 7256
rect 7892 7216 7898 7228
rect 9030 7216 9036 7228
rect 9088 7216 9094 7268
rect 4062 7188 4068 7200
rect 3016 7160 3740 7188
rect 4023 7160 4068 7188
rect 3016 7148 3022 7160
rect 4062 7148 4068 7160
rect 4120 7148 4126 7200
rect 4430 7188 4436 7200
rect 4391 7160 4436 7188
rect 4430 7148 4436 7160
rect 4488 7148 4494 7200
rect 4706 7148 4712 7200
rect 4764 7188 4770 7200
rect 5169 7191 5227 7197
rect 5169 7188 5181 7191
rect 4764 7160 5181 7188
rect 4764 7148 4770 7160
rect 5169 7157 5181 7160
rect 5215 7157 5227 7191
rect 5169 7151 5227 7157
rect 6362 7148 6368 7200
rect 6420 7188 6426 7200
rect 6457 7191 6515 7197
rect 6457 7188 6469 7191
rect 6420 7160 6469 7188
rect 6420 7148 6426 7160
rect 6457 7157 6469 7160
rect 6503 7157 6515 7191
rect 6457 7151 6515 7157
rect 8018 7148 8024 7200
rect 8076 7188 8082 7200
rect 10244 7197 10272 7296
rect 10778 7284 10784 7296
rect 10836 7284 10842 7336
rect 11054 7284 11060 7336
rect 11112 7324 11118 7336
rect 14844 7333 14872 7432
rect 15010 7352 15016 7404
rect 15068 7392 15074 7404
rect 16408 7392 16436 7488
rect 18230 7420 18236 7472
rect 18288 7460 18294 7472
rect 19153 7463 19211 7469
rect 19153 7460 19165 7463
rect 18288 7432 19165 7460
rect 18288 7420 18294 7432
rect 19153 7429 19165 7432
rect 19199 7460 19211 7463
rect 21100 7460 21128 7488
rect 19199 7432 21128 7460
rect 19199 7429 19211 7432
rect 19153 7423 19211 7429
rect 21266 7420 21272 7472
rect 21324 7460 21330 7472
rect 25363 7463 25421 7469
rect 25363 7460 25375 7463
rect 21324 7432 25375 7460
rect 21324 7420 21330 7432
rect 25363 7429 25375 7432
rect 25409 7429 25421 7463
rect 25363 7423 25421 7429
rect 15068 7364 16436 7392
rect 15068 7352 15074 7364
rect 11241 7327 11299 7333
rect 11241 7324 11253 7327
rect 11112 7296 11253 7324
rect 11112 7284 11118 7296
rect 11241 7293 11253 7296
rect 11287 7324 11299 7327
rect 11793 7327 11851 7333
rect 11793 7324 11805 7327
rect 11287 7296 11805 7324
rect 11287 7293 11299 7296
rect 11241 7287 11299 7293
rect 11793 7293 11805 7296
rect 11839 7293 11851 7327
rect 11793 7287 11851 7293
rect 14829 7327 14887 7333
rect 14829 7293 14841 7327
rect 14875 7324 14887 7327
rect 15197 7327 15255 7333
rect 15197 7324 15209 7327
rect 14875 7296 15209 7324
rect 14875 7293 14887 7296
rect 14829 7287 14887 7293
rect 15197 7293 15209 7296
rect 15243 7324 15255 7327
rect 15286 7324 15292 7336
rect 15243 7296 15292 7324
rect 15243 7293 15255 7296
rect 15197 7287 15255 7293
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 15396 7333 15424 7364
rect 17218 7352 17224 7404
rect 17276 7392 17282 7404
rect 17497 7395 17555 7401
rect 17497 7392 17509 7395
rect 17276 7364 17509 7392
rect 17276 7352 17282 7364
rect 17497 7361 17509 7364
rect 17543 7361 17555 7395
rect 17497 7355 17555 7361
rect 18785 7395 18843 7401
rect 18785 7361 18797 7395
rect 18831 7392 18843 7395
rect 18966 7392 18972 7404
rect 18831 7364 18972 7392
rect 18831 7361 18843 7364
rect 18785 7355 18843 7361
rect 18966 7352 18972 7364
rect 19024 7392 19030 7404
rect 20254 7392 20260 7404
rect 19024 7364 20260 7392
rect 19024 7352 19030 7364
rect 20254 7352 20260 7364
rect 20312 7392 20318 7404
rect 20533 7395 20591 7401
rect 20533 7392 20545 7395
rect 20312 7364 20545 7392
rect 20312 7352 20318 7364
rect 20533 7361 20545 7364
rect 20579 7361 20591 7395
rect 23385 7395 23443 7401
rect 23385 7392 23397 7395
rect 20533 7355 20591 7361
rect 22020 7364 23397 7392
rect 15381 7327 15439 7333
rect 15381 7293 15393 7327
rect 15427 7293 15439 7327
rect 16704 7327 16762 7333
rect 16704 7324 16716 7327
rect 15381 7287 15439 7293
rect 15488 7296 16716 7324
rect 11514 7256 11520 7268
rect 11475 7228 11520 7256
rect 11514 7216 11520 7228
rect 11572 7216 11578 7268
rect 13541 7259 13599 7265
rect 13541 7225 13553 7259
rect 13587 7225 13599 7259
rect 14090 7256 14096 7268
rect 14051 7228 14096 7256
rect 13541 7219 13599 7225
rect 10229 7191 10287 7197
rect 10229 7188 10241 7191
rect 8076 7160 10241 7188
rect 8076 7148 8082 7160
rect 10229 7157 10241 7160
rect 10275 7157 10287 7191
rect 10229 7151 10287 7157
rect 13262 7148 13268 7200
rect 13320 7188 13326 7200
rect 13556 7188 13584 7219
rect 14090 7216 14096 7228
rect 14148 7256 14154 7268
rect 14550 7256 14556 7268
rect 14148 7228 14556 7256
rect 14148 7216 14154 7228
rect 14550 7216 14556 7228
rect 14608 7216 14614 7268
rect 13320 7160 13584 7188
rect 13320 7148 13326 7160
rect 13722 7148 13728 7200
rect 13780 7188 13786 7200
rect 15488 7188 15516 7296
rect 16704 7293 16716 7296
rect 16750 7324 16762 7327
rect 17129 7327 17187 7333
rect 17129 7324 17141 7327
rect 16750 7296 17141 7324
rect 16750 7293 16762 7296
rect 16704 7287 16762 7293
rect 17129 7293 17141 7296
rect 17175 7293 17187 7327
rect 17129 7287 17187 7293
rect 21818 7284 21824 7336
rect 21876 7324 21882 7336
rect 22020 7333 22048 7364
rect 23385 7361 23397 7364
rect 23431 7392 23443 7395
rect 23566 7392 23572 7404
rect 23431 7364 23572 7392
rect 23431 7361 23443 7364
rect 23385 7355 23443 7361
rect 23566 7352 23572 7364
rect 23624 7392 23630 7404
rect 23624 7364 23704 7392
rect 23624 7352 23630 7364
rect 22005 7327 22063 7333
rect 22005 7324 22017 7327
rect 21876 7296 22017 7324
rect 21876 7284 21882 7296
rect 22005 7293 22017 7296
rect 22051 7293 22063 7327
rect 22005 7287 22063 7293
rect 22094 7284 22100 7336
rect 22152 7324 22158 7336
rect 23676 7333 23704 7364
rect 22465 7327 22523 7333
rect 22465 7324 22477 7327
rect 22152 7296 22477 7324
rect 22152 7284 22158 7296
rect 22465 7293 22477 7296
rect 22511 7293 22523 7327
rect 22465 7287 22523 7293
rect 23661 7327 23719 7333
rect 23661 7293 23673 7327
rect 23707 7293 23719 7327
rect 23661 7287 23719 7293
rect 23842 7284 23848 7336
rect 23900 7324 23906 7336
rect 24121 7327 24179 7333
rect 24121 7324 24133 7327
rect 23900 7296 24133 7324
rect 23900 7284 23906 7296
rect 24121 7293 24133 7296
rect 24167 7293 24179 7327
rect 24121 7287 24179 7293
rect 25038 7284 25044 7336
rect 25096 7324 25102 7336
rect 25260 7327 25318 7333
rect 25260 7324 25272 7327
rect 25096 7296 25272 7324
rect 25096 7284 25102 7296
rect 25260 7293 25272 7296
rect 25306 7324 25318 7327
rect 25685 7327 25743 7333
rect 25685 7324 25697 7327
rect 25306 7296 25697 7324
rect 25306 7293 25318 7296
rect 25260 7287 25318 7293
rect 25685 7293 25697 7296
rect 25731 7293 25743 7327
rect 25685 7287 25743 7293
rect 15654 7256 15660 7268
rect 15615 7228 15660 7256
rect 15654 7216 15660 7228
rect 15712 7216 15718 7268
rect 16807 7259 16865 7265
rect 16807 7225 16819 7259
rect 16853 7256 16865 7259
rect 18138 7256 18144 7268
rect 16853 7228 18144 7256
rect 16853 7225 16865 7228
rect 16807 7219 16865 7225
rect 18138 7216 18144 7228
rect 18196 7216 18202 7268
rect 18230 7216 18236 7268
rect 18288 7256 18294 7268
rect 18288 7228 18333 7256
rect 18288 7216 18294 7228
rect 20622 7216 20628 7268
rect 20680 7256 20686 7268
rect 21174 7256 21180 7268
rect 20680 7228 20725 7256
rect 21135 7228 21180 7256
rect 20680 7216 20686 7228
rect 21174 7216 21180 7228
rect 21232 7216 21238 7268
rect 22646 7216 22652 7268
rect 22704 7256 22710 7268
rect 22741 7259 22799 7265
rect 22741 7256 22753 7259
rect 22704 7228 22753 7256
rect 22704 7216 22710 7228
rect 22741 7225 22753 7228
rect 22787 7225 22799 7259
rect 22741 7219 22799 7225
rect 23382 7216 23388 7268
rect 23440 7256 23446 7268
rect 23860 7256 23888 7284
rect 23440 7228 23888 7256
rect 23440 7216 23446 7228
rect 13780 7160 15516 7188
rect 13780 7148 13786 7160
rect 19426 7148 19432 7200
rect 19484 7188 19490 7200
rect 19797 7191 19855 7197
rect 19797 7188 19809 7191
rect 19484 7160 19809 7188
rect 19484 7148 19490 7160
rect 19797 7157 19809 7160
rect 19843 7157 19855 7191
rect 19797 7151 19855 7157
rect 20349 7191 20407 7197
rect 20349 7157 20361 7191
rect 20395 7188 20407 7191
rect 20640 7188 20668 7216
rect 21818 7188 21824 7200
rect 20395 7160 20668 7188
rect 21779 7160 21824 7188
rect 20395 7157 20407 7160
rect 20349 7151 20407 7157
rect 21818 7148 21824 7160
rect 21876 7148 21882 7200
rect 23750 7188 23756 7200
rect 23711 7160 23756 7188
rect 23750 7148 23756 7160
rect 23808 7148 23814 7200
rect 24670 7188 24676 7200
rect 24631 7160 24676 7188
rect 24670 7148 24676 7160
rect 24728 7148 24734 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1670 6984 1676 6996
rect 1583 6956 1676 6984
rect 1670 6944 1676 6956
rect 1728 6984 1734 6996
rect 2958 6984 2964 6996
rect 1728 6956 2964 6984
rect 1728 6944 1734 6956
rect 2958 6944 2964 6956
rect 3016 6944 3022 6996
rect 3418 6944 3424 6996
rect 3476 6984 3482 6996
rect 3697 6987 3755 6993
rect 3697 6984 3709 6987
rect 3476 6956 3709 6984
rect 3476 6944 3482 6956
rect 3697 6953 3709 6956
rect 3743 6953 3755 6987
rect 4246 6984 4252 6996
rect 4207 6956 4252 6984
rect 3697 6947 3755 6953
rect 4246 6944 4252 6956
rect 4304 6944 4310 6996
rect 6086 6984 6092 6996
rect 4632 6956 5948 6984
rect 6047 6956 6092 6984
rect 2406 6916 2412 6928
rect 2367 6888 2412 6916
rect 2406 6876 2412 6888
rect 2464 6876 2470 6928
rect 2498 6876 2504 6928
rect 2556 6916 2562 6928
rect 4632 6916 4660 6956
rect 5166 6916 5172 6928
rect 2556 6888 4660 6916
rect 5127 6888 5172 6916
rect 2556 6876 2562 6888
rect 5166 6876 5172 6888
rect 5224 6876 5230 6928
rect 5920 6916 5948 6956
rect 6086 6944 6092 6956
rect 6144 6944 6150 6996
rect 7466 6944 7472 6996
rect 7524 6984 7530 6996
rect 8297 6987 8355 6993
rect 8297 6984 8309 6987
rect 7524 6956 8309 6984
rect 7524 6944 7530 6956
rect 8297 6953 8309 6956
rect 8343 6953 8355 6987
rect 8297 6947 8355 6953
rect 11238 6944 11244 6996
rect 11296 6984 11302 6996
rect 11425 6987 11483 6993
rect 11425 6984 11437 6987
rect 11296 6956 11437 6984
rect 11296 6944 11302 6956
rect 11425 6953 11437 6956
rect 11471 6953 11483 6987
rect 11425 6947 11483 6953
rect 11514 6944 11520 6996
rect 11572 6984 11578 6996
rect 12434 6984 12440 6996
rect 11572 6956 12440 6984
rect 11572 6944 11578 6956
rect 12434 6944 12440 6956
rect 12492 6984 12498 6996
rect 12621 6987 12679 6993
rect 12621 6984 12633 6987
rect 12492 6956 12633 6984
rect 12492 6944 12498 6956
rect 12621 6953 12633 6956
rect 12667 6953 12679 6987
rect 15010 6984 15016 6996
rect 12621 6947 12679 6953
rect 12728 6956 13492 6984
rect 14971 6956 15016 6984
rect 6365 6919 6423 6925
rect 6365 6916 6377 6919
rect 5920 6888 6377 6916
rect 6365 6885 6377 6888
rect 6411 6916 6423 6919
rect 6730 6916 6736 6928
rect 6411 6888 6736 6916
rect 6411 6885 6423 6888
rect 6365 6879 6423 6885
rect 6730 6876 6736 6888
rect 6788 6916 6794 6928
rect 7558 6916 7564 6928
rect 6788 6888 7144 6916
rect 7519 6888 7564 6916
rect 6788 6876 6794 6888
rect 2130 6848 2136 6860
rect 2091 6820 2136 6848
rect 2130 6808 2136 6820
rect 2188 6808 2194 6860
rect 6270 6808 6276 6860
rect 6328 6848 6334 6860
rect 6549 6851 6607 6857
rect 6549 6848 6561 6851
rect 6328 6820 6561 6848
rect 6328 6808 6334 6820
rect 6549 6817 6561 6820
rect 6595 6817 6607 6851
rect 6549 6811 6607 6817
rect 6822 6808 6828 6860
rect 6880 6848 6886 6860
rect 7006 6848 7012 6860
rect 6880 6820 7012 6848
rect 6880 6808 6886 6820
rect 7006 6808 7012 6820
rect 7064 6808 7070 6860
rect 7116 6848 7144 6888
rect 7558 6876 7564 6888
rect 7616 6876 7622 6928
rect 8202 6876 8208 6928
rect 8260 6916 8266 6928
rect 8941 6919 8999 6925
rect 8941 6916 8953 6919
rect 8260 6888 8953 6916
rect 8260 6876 8266 6888
rect 8941 6885 8953 6888
rect 8987 6885 8999 6919
rect 12728 6916 12756 6956
rect 13354 6916 13360 6928
rect 8941 6879 8999 6885
rect 11900 6888 12756 6916
rect 13315 6888 13360 6916
rect 11900 6860 11928 6888
rect 13354 6876 13360 6888
rect 13412 6876 13418 6928
rect 13464 6916 13492 6956
rect 15010 6944 15016 6956
rect 15068 6944 15074 6996
rect 17218 6944 17224 6996
rect 17276 6984 17282 6996
rect 17957 6987 18015 6993
rect 17957 6984 17969 6987
rect 17276 6956 17969 6984
rect 17276 6944 17282 6956
rect 17957 6953 17969 6956
rect 18003 6953 18015 6987
rect 17957 6947 18015 6953
rect 18138 6944 18144 6996
rect 18196 6984 18202 6996
rect 18785 6987 18843 6993
rect 18785 6984 18797 6987
rect 18196 6956 18797 6984
rect 18196 6944 18202 6956
rect 18785 6953 18797 6956
rect 18831 6953 18843 6987
rect 18785 6947 18843 6953
rect 19659 6987 19717 6993
rect 19659 6953 19671 6987
rect 19705 6984 19717 6987
rect 20070 6984 20076 6996
rect 19705 6956 20076 6984
rect 19705 6953 19717 6956
rect 19659 6947 19717 6953
rect 20070 6944 20076 6956
rect 20128 6944 20134 6996
rect 20622 6944 20628 6996
rect 20680 6984 20686 6996
rect 21821 6987 21879 6993
rect 21821 6984 21833 6987
rect 20680 6956 21833 6984
rect 20680 6944 20686 6956
rect 21821 6953 21833 6956
rect 21867 6953 21879 6987
rect 21821 6947 21879 6953
rect 22554 6944 22560 6996
rect 22612 6984 22618 6996
rect 23569 6987 23627 6993
rect 22612 6956 23474 6984
rect 22612 6944 22618 6956
rect 13906 6916 13912 6928
rect 13464 6888 13912 6916
rect 13906 6876 13912 6888
rect 13964 6916 13970 6928
rect 16390 6916 16396 6928
rect 13964 6888 16396 6916
rect 13964 6876 13970 6888
rect 7929 6851 7987 6857
rect 7929 6848 7941 6851
rect 7116 6820 7941 6848
rect 7929 6817 7941 6820
rect 7975 6817 7987 6851
rect 8110 6848 8116 6860
rect 8071 6820 8116 6848
rect 7929 6811 7987 6817
rect 8110 6808 8116 6820
rect 8168 6808 8174 6860
rect 9950 6808 9956 6860
rect 10008 6848 10014 6860
rect 10045 6851 10103 6857
rect 10045 6848 10057 6851
rect 10008 6820 10057 6848
rect 10008 6808 10014 6820
rect 10045 6817 10057 6820
rect 10091 6817 10103 6851
rect 10045 6811 10103 6817
rect 10597 6851 10655 6857
rect 10597 6817 10609 6851
rect 10643 6848 10655 6851
rect 11054 6848 11060 6860
rect 10643 6820 11060 6848
rect 10643 6817 10655 6820
rect 10597 6811 10655 6817
rect 11054 6808 11060 6820
rect 11112 6808 11118 6860
rect 11882 6848 11888 6860
rect 11795 6820 11888 6848
rect 11882 6808 11888 6820
rect 11940 6808 11946 6860
rect 12161 6851 12219 6857
rect 12161 6817 12173 6851
rect 12207 6848 12219 6851
rect 12250 6848 12256 6860
rect 12207 6820 12256 6848
rect 12207 6817 12219 6820
rect 12161 6811 12219 6817
rect 12250 6808 12256 6820
rect 12308 6808 12314 6860
rect 15580 6857 15608 6888
rect 16390 6876 16396 6888
rect 16448 6916 16454 6928
rect 16448 6888 17724 6916
rect 16448 6876 16454 6888
rect 15565 6851 15623 6857
rect 15565 6817 15577 6851
rect 15611 6817 15623 6851
rect 15565 6811 15623 6817
rect 15749 6851 15807 6857
rect 15749 6817 15761 6851
rect 15795 6848 15807 6851
rect 16114 6848 16120 6860
rect 15795 6820 16120 6848
rect 15795 6817 15807 6820
rect 15749 6811 15807 6817
rect 16114 6808 16120 6820
rect 16172 6808 16178 6860
rect 16206 6808 16212 6860
rect 16264 6848 16270 6860
rect 17586 6848 17592 6860
rect 16264 6820 17592 6848
rect 16264 6808 16270 6820
rect 17586 6808 17592 6820
rect 17644 6808 17650 6860
rect 2041 6783 2099 6789
rect 2041 6749 2053 6783
rect 2087 6780 2099 6783
rect 2498 6780 2504 6792
rect 2087 6752 2504 6780
rect 2087 6749 2099 6752
rect 2041 6743 2099 6749
rect 2498 6740 2504 6752
rect 2556 6740 2562 6792
rect 3418 6740 3424 6792
rect 3476 6780 3482 6792
rect 4246 6780 4252 6792
rect 3476 6752 4252 6780
rect 3476 6740 3482 6752
rect 4246 6740 4252 6752
rect 4304 6740 4310 6792
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6780 5135 6783
rect 5534 6780 5540 6792
rect 5123 6752 5540 6780
rect 5123 6749 5135 6752
rect 5077 6743 5135 6749
rect 5534 6740 5540 6752
rect 5592 6740 5598 6792
rect 7098 6780 7104 6792
rect 7059 6752 7104 6780
rect 7098 6740 7104 6752
rect 7156 6740 7162 6792
rect 10778 6780 10784 6792
rect 10739 6752 10784 6780
rect 10778 6740 10784 6752
rect 10836 6740 10842 6792
rect 12345 6783 12403 6789
rect 12345 6749 12357 6783
rect 12391 6780 12403 6783
rect 13265 6783 13323 6789
rect 12391 6752 13077 6780
rect 12391 6749 12403 6752
rect 12345 6743 12403 6749
rect 3786 6672 3792 6724
rect 3844 6712 3850 6724
rect 4890 6712 4896 6724
rect 3844 6684 4896 6712
rect 3844 6672 3850 6684
rect 4890 6672 4896 6684
rect 4948 6712 4954 6724
rect 5629 6715 5687 6721
rect 5629 6712 5641 6715
rect 4948 6684 5641 6712
rect 4948 6672 4954 6684
rect 5629 6681 5641 6684
rect 5675 6712 5687 6715
rect 6454 6712 6460 6724
rect 5675 6684 6460 6712
rect 5675 6681 5687 6684
rect 5629 6675 5687 6681
rect 6454 6672 6460 6684
rect 6512 6672 6518 6724
rect 3050 6644 3056 6656
rect 3011 6616 3056 6644
rect 3050 6604 3056 6616
rect 3108 6604 3114 6656
rect 3418 6644 3424 6656
rect 3379 6616 3424 6644
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 4709 6647 4767 6653
rect 4709 6613 4721 6647
rect 4755 6644 4767 6647
rect 4798 6644 4804 6656
rect 4755 6616 4804 6644
rect 4755 6613 4767 6616
rect 4709 6607 4767 6613
rect 4798 6604 4804 6616
rect 4856 6644 4862 6656
rect 6178 6644 6184 6656
rect 4856 6616 6184 6644
rect 4856 6604 4862 6616
rect 6178 6604 6184 6616
rect 6236 6644 6242 6656
rect 8018 6644 8024 6656
rect 6236 6616 8024 6644
rect 6236 6604 6242 6616
rect 8018 6604 8024 6616
rect 8076 6604 8082 6656
rect 8294 6604 8300 6656
rect 8352 6644 8358 6656
rect 8665 6647 8723 6653
rect 8665 6644 8677 6647
rect 8352 6616 8677 6644
rect 8352 6604 8358 6616
rect 8665 6613 8677 6616
rect 8711 6644 8723 6647
rect 9306 6644 9312 6656
rect 8711 6616 9312 6644
rect 8711 6613 8723 6616
rect 8665 6607 8723 6613
rect 9306 6604 9312 6616
rect 9364 6604 9370 6656
rect 11054 6644 11060 6656
rect 11015 6616 11060 6644
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 13049 6644 13077 6752
rect 13265 6749 13277 6783
rect 13311 6780 13323 6783
rect 13311 6752 13400 6780
rect 13311 6749 13323 6752
rect 13265 6743 13323 6749
rect 13372 6712 13400 6752
rect 13446 6740 13452 6792
rect 13504 6780 13510 6792
rect 13541 6783 13599 6789
rect 13541 6780 13553 6783
rect 13504 6752 13553 6780
rect 13504 6740 13510 6752
rect 13541 6749 13553 6752
rect 13587 6749 13599 6783
rect 15838 6780 15844 6792
rect 15799 6752 15844 6780
rect 13541 6743 13599 6749
rect 15838 6740 15844 6752
rect 15896 6740 15902 6792
rect 17696 6780 17724 6888
rect 18046 6876 18052 6928
rect 18104 6916 18110 6928
rect 19153 6919 19211 6925
rect 19153 6916 19165 6919
rect 18104 6888 19165 6916
rect 18104 6876 18110 6888
rect 19153 6885 19165 6888
rect 19199 6916 19211 6919
rect 20254 6916 20260 6928
rect 19199 6888 19656 6916
rect 20215 6888 20260 6916
rect 19199 6885 19211 6888
rect 19153 6879 19211 6885
rect 19628 6860 19656 6888
rect 20254 6876 20260 6888
rect 20312 6876 20318 6928
rect 20990 6876 20996 6928
rect 21048 6916 21054 6928
rect 21222 6919 21280 6925
rect 21222 6916 21234 6919
rect 21048 6888 21234 6916
rect 21048 6876 21054 6888
rect 21222 6885 21234 6888
rect 21268 6885 21280 6919
rect 21222 6879 21280 6885
rect 22738 6876 22744 6928
rect 22796 6916 22802 6928
rect 22970 6919 23028 6925
rect 22970 6916 22982 6919
rect 22796 6888 22982 6916
rect 22796 6876 22802 6888
rect 22970 6885 22982 6888
rect 23016 6885 23028 6919
rect 23446 6916 23474 6956
rect 23569 6953 23581 6987
rect 23615 6984 23627 6987
rect 23615 6956 24624 6984
rect 23615 6953 23627 6956
rect 23569 6947 23627 6953
rect 24210 6916 24216 6928
rect 23446 6888 24216 6916
rect 22970 6879 23028 6885
rect 24210 6876 24216 6888
rect 24268 6916 24274 6928
rect 24596 6925 24624 6956
rect 24489 6919 24547 6925
rect 24489 6916 24501 6919
rect 24268 6888 24501 6916
rect 24268 6876 24274 6888
rect 24489 6885 24501 6888
rect 24535 6885 24547 6919
rect 24489 6879 24547 6885
rect 24581 6919 24639 6925
rect 24581 6885 24593 6919
rect 24627 6916 24639 6919
rect 24946 6916 24952 6928
rect 24627 6888 24952 6916
rect 24627 6885 24639 6888
rect 24581 6879 24639 6885
rect 24946 6876 24952 6888
rect 25004 6876 25010 6928
rect 18230 6808 18236 6860
rect 18288 6848 18294 6860
rect 18509 6851 18567 6857
rect 18509 6848 18521 6851
rect 18288 6820 18521 6848
rect 18288 6808 18294 6820
rect 18509 6817 18521 6820
rect 18555 6817 18567 6851
rect 18509 6811 18567 6817
rect 19429 6851 19487 6857
rect 19429 6817 19441 6851
rect 19475 6848 19487 6851
rect 19518 6848 19524 6860
rect 19475 6820 19524 6848
rect 19475 6817 19487 6820
rect 19429 6811 19487 6817
rect 19518 6808 19524 6820
rect 19576 6808 19582 6860
rect 19610 6808 19616 6860
rect 19668 6808 19674 6860
rect 22830 6848 22836 6860
rect 19812 6820 22836 6848
rect 19812 6780 19840 6820
rect 22830 6808 22836 6820
rect 22888 6808 22894 6860
rect 17696 6752 19840 6780
rect 20806 6740 20812 6792
rect 20864 6780 20870 6792
rect 20901 6783 20959 6789
rect 20901 6780 20913 6783
rect 20864 6752 20913 6780
rect 20864 6740 20870 6752
rect 20901 6749 20913 6752
rect 20947 6749 20959 6783
rect 22646 6780 22652 6792
rect 22607 6752 22652 6780
rect 20901 6743 20959 6749
rect 22646 6740 22652 6752
rect 22704 6740 22710 6792
rect 24026 6740 24032 6792
rect 24084 6780 24090 6792
rect 24670 6780 24676 6792
rect 24084 6752 24676 6780
rect 24084 6740 24090 6752
rect 24670 6740 24676 6752
rect 24728 6780 24734 6792
rect 24765 6783 24823 6789
rect 24765 6780 24777 6783
rect 24728 6752 24777 6780
rect 24728 6740 24734 6752
rect 24765 6749 24777 6752
rect 24811 6749 24823 6783
rect 24765 6743 24823 6749
rect 13998 6712 14004 6724
rect 13372 6684 14004 6712
rect 13998 6672 14004 6684
rect 14056 6672 14062 6724
rect 17402 6712 17408 6724
rect 14844 6684 17408 6712
rect 14844 6644 14872 6684
rect 17402 6672 17408 6684
rect 17460 6672 17466 6724
rect 20622 6644 20628 6656
rect 13049 6616 14872 6644
rect 20583 6616 20628 6644
rect 20622 6604 20628 6616
rect 20680 6604 20686 6656
rect 23842 6644 23848 6656
rect 23803 6616 23848 6644
rect 23842 6604 23848 6616
rect 23900 6604 23906 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 1762 6440 1768 6452
rect 1627 6412 1768 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 1762 6400 1768 6412
rect 1820 6400 1826 6452
rect 3050 6400 3056 6452
rect 3108 6440 3114 6452
rect 3421 6443 3479 6449
rect 3421 6440 3433 6443
rect 3108 6412 3433 6440
rect 3108 6400 3114 6412
rect 3421 6409 3433 6412
rect 3467 6409 3479 6443
rect 3421 6403 3479 6409
rect 5166 6400 5172 6452
rect 5224 6440 5230 6452
rect 5261 6443 5319 6449
rect 5261 6440 5273 6443
rect 5224 6412 5273 6440
rect 5224 6400 5230 6412
rect 5261 6409 5273 6412
rect 5307 6409 5319 6443
rect 6270 6440 6276 6452
rect 6231 6412 6276 6440
rect 5261 6403 5319 6409
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 6822 6400 6828 6452
rect 6880 6440 6886 6452
rect 11882 6440 11888 6452
rect 6880 6412 10732 6440
rect 11843 6412 11888 6440
rect 6880 6400 6886 6412
rect 5534 6332 5540 6384
rect 5592 6372 5598 6384
rect 5592 6344 9168 6372
rect 5592 6332 5598 6344
rect 1486 6264 1492 6316
rect 1544 6304 1550 6316
rect 2777 6307 2835 6313
rect 2777 6304 2789 6307
rect 1544 6276 2789 6304
rect 1544 6264 1550 6276
rect 2777 6273 2789 6276
rect 2823 6304 2835 6307
rect 3786 6304 3792 6316
rect 2823 6276 3792 6304
rect 2823 6273 2835 6276
rect 2777 6267 2835 6273
rect 3786 6264 3792 6276
rect 3844 6264 3850 6316
rect 3881 6307 3939 6313
rect 3881 6273 3893 6307
rect 3927 6304 3939 6307
rect 4341 6307 4399 6313
rect 4341 6304 4353 6307
rect 3927 6276 4353 6304
rect 3927 6273 3939 6276
rect 3881 6267 3939 6273
rect 4341 6273 4353 6276
rect 4387 6304 4399 6307
rect 4430 6304 4436 6316
rect 4387 6276 4436 6304
rect 4387 6273 4399 6276
rect 4341 6267 4399 6273
rect 4430 6264 4436 6276
rect 4488 6264 4494 6316
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6304 5963 6307
rect 6822 6304 6828 6316
rect 5951 6276 6828 6304
rect 5951 6273 5963 6276
rect 5905 6267 5963 6273
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 7009 6307 7067 6313
rect 7009 6273 7021 6307
rect 7055 6304 7067 6307
rect 7098 6304 7104 6316
rect 7055 6276 7104 6304
rect 7055 6273 7067 6276
rect 7009 6267 7067 6273
rect 7098 6264 7104 6276
rect 7156 6264 7162 6316
rect 8849 6307 8907 6313
rect 8849 6273 8861 6307
rect 8895 6304 8907 6307
rect 8938 6304 8944 6316
rect 8895 6276 8944 6304
rect 8895 6273 8907 6276
rect 8849 6267 8907 6273
rect 8938 6264 8944 6276
rect 8996 6264 9002 6316
rect 9140 6313 9168 6344
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6304 9183 6307
rect 9858 6304 9864 6316
rect 9171 6276 9864 6304
rect 9171 6273 9183 6276
rect 9125 6267 9183 6273
rect 9858 6264 9864 6276
rect 9916 6264 9922 6316
rect 10704 6304 10732 6412
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 12253 6443 12311 6449
rect 12253 6409 12265 6443
rect 12299 6440 12311 6443
rect 12342 6440 12348 6452
rect 12299 6412 12348 6440
rect 12299 6409 12311 6412
rect 12253 6403 12311 6409
rect 12342 6400 12348 6412
rect 12400 6400 12406 6452
rect 13354 6400 13360 6452
rect 13412 6440 13418 6452
rect 13633 6443 13691 6449
rect 13633 6440 13645 6443
rect 13412 6412 13645 6440
rect 13412 6400 13418 6412
rect 13633 6409 13645 6412
rect 13679 6409 13691 6443
rect 13633 6403 13691 6409
rect 16114 6400 16120 6452
rect 16172 6440 16178 6452
rect 16669 6443 16727 6449
rect 16669 6440 16681 6443
rect 16172 6412 16681 6440
rect 16172 6400 16178 6412
rect 16669 6409 16681 6412
rect 16715 6440 16727 6443
rect 18046 6440 18052 6452
rect 16715 6412 18052 6440
rect 16715 6409 16727 6412
rect 16669 6403 16727 6409
rect 18046 6400 18052 6412
rect 18104 6400 18110 6452
rect 18279 6443 18337 6449
rect 18279 6409 18291 6443
rect 18325 6440 18337 6443
rect 19426 6440 19432 6452
rect 18325 6412 19432 6440
rect 18325 6409 18337 6412
rect 18279 6403 18337 6409
rect 19426 6400 19432 6412
rect 19484 6400 19490 6452
rect 20990 6440 20996 6452
rect 20951 6412 20996 6440
rect 20990 6400 20996 6412
rect 21048 6400 21054 6452
rect 22646 6400 22652 6452
rect 22704 6440 22710 6452
rect 23017 6443 23075 6449
rect 23017 6440 23029 6443
rect 22704 6412 23029 6440
rect 22704 6400 22710 6412
rect 23017 6409 23029 6412
rect 23063 6409 23075 6443
rect 23017 6403 23075 6409
rect 24210 6400 24216 6452
rect 24268 6440 24274 6452
rect 24673 6443 24731 6449
rect 24673 6440 24685 6443
rect 24268 6412 24685 6440
rect 24268 6400 24274 6412
rect 24673 6409 24685 6412
rect 24719 6409 24731 6443
rect 24673 6403 24731 6409
rect 24946 6400 24952 6452
rect 25004 6440 25010 6452
rect 25041 6443 25099 6449
rect 25041 6440 25053 6443
rect 25004 6412 25053 6440
rect 25004 6400 25010 6412
rect 25041 6409 25053 6412
rect 25087 6409 25099 6443
rect 25041 6403 25099 6409
rect 25314 6400 25320 6452
rect 25372 6440 25378 6452
rect 25501 6443 25559 6449
rect 25501 6440 25513 6443
rect 25372 6412 25513 6440
rect 25372 6400 25378 6412
rect 25501 6409 25513 6412
rect 25547 6409 25559 6443
rect 25501 6403 25559 6409
rect 11517 6375 11575 6381
rect 11517 6341 11529 6375
rect 11563 6372 11575 6375
rect 13538 6372 13544 6384
rect 11563 6344 13544 6372
rect 11563 6341 11575 6344
rect 11517 6335 11575 6341
rect 11532 6304 11560 6335
rect 13538 6332 13544 6344
rect 13596 6332 13602 6384
rect 15194 6372 15200 6384
rect 15107 6344 15200 6372
rect 15194 6332 15200 6344
rect 15252 6372 15258 6384
rect 15289 6375 15347 6381
rect 15289 6372 15301 6375
rect 15252 6344 15301 6372
rect 15252 6332 15258 6344
rect 15289 6341 15301 6344
rect 15335 6372 15347 6375
rect 17218 6372 17224 6384
rect 15335 6344 17224 6372
rect 15335 6341 15347 6344
rect 15289 6335 15347 6341
rect 17218 6332 17224 6344
rect 17276 6372 17282 6384
rect 17589 6375 17647 6381
rect 17589 6372 17601 6375
rect 17276 6344 17601 6372
rect 17276 6332 17282 6344
rect 17589 6341 17601 6344
rect 17635 6341 17647 6375
rect 22738 6372 22744 6384
rect 22699 6344 22744 6372
rect 17589 6335 17647 6341
rect 22738 6332 22744 6344
rect 22796 6332 22802 6384
rect 23477 6375 23535 6381
rect 23477 6372 23489 6375
rect 22848 6344 23489 6372
rect 12434 6304 12440 6316
rect 10704 6276 11560 6304
rect 12395 6276 12440 6304
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 1670 6236 1676 6248
rect 1443 6208 1676 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 1670 6196 1676 6208
rect 1728 6196 1734 6248
rect 3326 6196 3332 6248
rect 3384 6236 3390 6248
rect 6914 6236 6920 6248
rect 3384 6208 6920 6236
rect 3384 6196 3390 6208
rect 6914 6196 6920 6208
rect 6972 6236 6978 6248
rect 8110 6236 8116 6248
rect 6972 6208 8116 6236
rect 6972 6196 6978 6208
rect 8110 6196 8116 6208
rect 8168 6236 8174 6248
rect 10704 6245 10732 6276
rect 12434 6264 12440 6276
rect 12492 6264 12498 6316
rect 15381 6307 15439 6313
rect 15381 6273 15393 6307
rect 15427 6304 15439 6307
rect 15654 6304 15660 6316
rect 15427 6276 15660 6304
rect 15427 6273 15439 6276
rect 15381 6267 15439 6273
rect 15654 6264 15660 6276
rect 15712 6304 15718 6316
rect 16945 6307 17003 6313
rect 16945 6304 16957 6307
rect 15712 6276 16957 6304
rect 15712 6264 15718 6276
rect 16945 6273 16957 6276
rect 16991 6273 17003 6307
rect 16945 6267 17003 6273
rect 19061 6307 19119 6313
rect 19061 6273 19073 6307
rect 19107 6304 19119 6307
rect 19242 6304 19248 6316
rect 19107 6276 19248 6304
rect 19107 6273 19119 6276
rect 19061 6267 19119 6273
rect 19242 6264 19248 6276
rect 19300 6304 19306 6316
rect 22848 6304 22876 6344
rect 23477 6341 23489 6344
rect 23523 6372 23535 6375
rect 23523 6344 23704 6372
rect 23523 6341 23535 6344
rect 23477 6335 23535 6341
rect 19300 6276 22876 6304
rect 19300 6264 19306 6276
rect 8205 6239 8263 6245
rect 8205 6236 8217 6239
rect 8168 6208 8217 6236
rect 8168 6196 8174 6208
rect 8205 6205 8217 6208
rect 8251 6205 8263 6239
rect 8205 6199 8263 6205
rect 10689 6239 10747 6245
rect 10689 6205 10701 6239
rect 10735 6205 10747 6239
rect 10689 6199 10747 6205
rect 10873 6239 10931 6245
rect 10873 6205 10885 6239
rect 10919 6236 10931 6239
rect 11054 6236 11060 6248
rect 10919 6208 11060 6236
rect 10919 6205 10931 6208
rect 10873 6199 10931 6205
rect 2498 6168 2504 6180
rect 2459 6140 2504 6168
rect 2498 6128 2504 6140
rect 2556 6128 2562 6180
rect 2593 6171 2651 6177
rect 2593 6137 2605 6171
rect 2639 6168 2651 6171
rect 2958 6168 2964 6180
rect 2639 6140 2964 6168
rect 2639 6137 2651 6140
rect 2593 6131 2651 6137
rect 2958 6128 2964 6140
rect 3016 6128 3022 6180
rect 4662 6171 4720 6177
rect 4662 6168 4674 6171
rect 4172 6140 4674 6168
rect 2225 6103 2283 6109
rect 2225 6069 2237 6103
rect 2271 6100 2283 6103
rect 2406 6100 2412 6112
rect 2271 6072 2412 6100
rect 2271 6069 2283 6072
rect 2225 6063 2283 6069
rect 2406 6060 2412 6072
rect 2464 6100 2470 6112
rect 4062 6100 4068 6112
rect 2464 6072 4068 6100
rect 2464 6060 2470 6072
rect 4062 6060 4068 6072
rect 4120 6100 4126 6112
rect 4172 6109 4200 6140
rect 4662 6137 4674 6140
rect 4708 6168 4720 6171
rect 6549 6171 6607 6177
rect 6549 6168 6561 6171
rect 4708 6140 6561 6168
rect 4708 6137 4720 6140
rect 4662 6131 4720 6137
rect 6549 6137 6561 6140
rect 6595 6168 6607 6171
rect 7330 6171 7388 6177
rect 7330 6168 7342 6171
rect 6595 6140 7342 6168
rect 6595 6137 6607 6140
rect 6549 6131 6607 6137
rect 7330 6137 7342 6140
rect 7376 6137 7388 6171
rect 8573 6171 8631 6177
rect 8573 6168 8585 6171
rect 7330 6131 7388 6137
rect 7944 6140 8585 6168
rect 4157 6103 4215 6109
rect 4157 6100 4169 6103
rect 4120 6072 4169 6100
rect 4120 6060 4126 6072
rect 4157 6069 4169 6072
rect 4203 6069 4215 6103
rect 4157 6063 4215 6069
rect 7834 6060 7840 6112
rect 7892 6100 7898 6112
rect 7944 6109 7972 6140
rect 8573 6137 8585 6140
rect 8619 6137 8631 6171
rect 8573 6131 8631 6137
rect 8941 6171 8999 6177
rect 8941 6137 8953 6171
rect 8987 6137 8999 6171
rect 8941 6131 8999 6137
rect 7929 6103 7987 6109
rect 7929 6100 7941 6103
rect 7892 6072 7941 6100
rect 7892 6060 7898 6072
rect 7929 6069 7941 6072
rect 7975 6069 7987 6103
rect 8588 6100 8616 6131
rect 8956 6100 8984 6131
rect 10134 6128 10140 6180
rect 10192 6168 10198 6180
rect 10888 6168 10916 6199
rect 11054 6196 11060 6208
rect 11112 6196 11118 6248
rect 13722 6196 13728 6248
rect 13780 6236 13786 6248
rect 14220 6239 14278 6245
rect 14220 6236 14232 6239
rect 13780 6208 14232 6236
rect 13780 6196 13786 6208
rect 14220 6205 14232 6208
rect 14266 6236 14278 6239
rect 14645 6239 14703 6245
rect 14645 6236 14657 6239
rect 14266 6208 14657 6236
rect 14266 6205 14278 6208
rect 14220 6199 14278 6205
rect 14645 6205 14657 6208
rect 14691 6205 14703 6239
rect 18208 6239 18266 6245
rect 14645 6199 14703 6205
rect 15626 6208 15884 6236
rect 11146 6168 11152 6180
rect 10192 6140 10916 6168
rect 11107 6140 11152 6168
rect 10192 6128 10198 6140
rect 11146 6128 11152 6140
rect 11204 6128 11210 6180
rect 12342 6128 12348 6180
rect 12400 6168 12406 6180
rect 12758 6171 12816 6177
rect 12758 6168 12770 6171
rect 12400 6140 12770 6168
rect 12400 6128 12406 6140
rect 12758 6137 12770 6140
rect 12804 6137 12816 6171
rect 13998 6168 14004 6180
rect 13911 6140 14004 6168
rect 12758 6131 12816 6137
rect 13998 6128 14004 6140
rect 14056 6168 14062 6180
rect 15626 6168 15654 6208
rect 14056 6140 15654 6168
rect 15702 6171 15760 6177
rect 14056 6128 14062 6140
rect 15702 6137 15714 6171
rect 15748 6137 15760 6171
rect 15856 6168 15884 6208
rect 18208 6205 18220 6239
rect 18254 6236 18266 6239
rect 18693 6239 18751 6245
rect 18693 6236 18705 6239
rect 18254 6208 18705 6236
rect 18254 6205 18266 6208
rect 18208 6199 18266 6205
rect 18693 6205 18705 6208
rect 18739 6236 18751 6239
rect 18966 6236 18972 6248
rect 18739 6208 18972 6236
rect 18739 6205 18751 6208
rect 18693 6199 18751 6205
rect 18966 6196 18972 6208
rect 19024 6196 19030 6248
rect 19352 6245 19380 6276
rect 19337 6239 19395 6245
rect 19337 6205 19349 6239
rect 19383 6205 19395 6239
rect 19610 6236 19616 6248
rect 19571 6208 19616 6236
rect 19337 6199 19395 6205
rect 19610 6196 19616 6208
rect 19668 6236 19674 6248
rect 19978 6236 19984 6248
rect 19668 6208 19984 6236
rect 19668 6196 19674 6208
rect 19978 6196 19984 6208
rect 20036 6196 20042 6248
rect 21453 6239 21511 6245
rect 21453 6205 21465 6239
rect 21499 6236 21511 6239
rect 21821 6239 21879 6245
rect 21821 6236 21833 6239
rect 21499 6208 21833 6236
rect 21499 6205 21511 6208
rect 21453 6199 21511 6205
rect 21821 6205 21833 6208
rect 21867 6236 21879 6239
rect 21910 6236 21916 6248
rect 21867 6208 21916 6236
rect 21867 6205 21879 6208
rect 21821 6199 21879 6205
rect 21910 6196 21916 6208
rect 21968 6196 21974 6248
rect 22002 6196 22008 6248
rect 22060 6236 22066 6248
rect 23676 6245 23704 6344
rect 23661 6239 23719 6245
rect 22060 6208 22105 6236
rect 22060 6196 22066 6208
rect 23661 6205 23673 6239
rect 23707 6205 23719 6239
rect 23661 6199 23719 6205
rect 23842 6196 23848 6248
rect 23900 6236 23906 6248
rect 24213 6239 24271 6245
rect 24213 6236 24225 6239
rect 23900 6208 24225 6236
rect 23900 6196 23906 6208
rect 24213 6205 24225 6208
rect 24259 6236 24271 6239
rect 24302 6236 24308 6248
rect 24259 6208 24308 6236
rect 24259 6205 24271 6208
rect 24213 6199 24271 6205
rect 24302 6196 24308 6208
rect 24360 6196 24366 6248
rect 25130 6196 25136 6248
rect 25188 6236 25194 6248
rect 25260 6239 25318 6245
rect 25260 6236 25272 6239
rect 25188 6208 25272 6236
rect 25188 6196 25194 6208
rect 25260 6205 25272 6208
rect 25306 6236 25318 6239
rect 25685 6239 25743 6245
rect 25685 6236 25697 6239
rect 25306 6208 25697 6236
rect 25306 6205 25318 6208
rect 25260 6199 25318 6205
rect 25685 6205 25697 6208
rect 25731 6205 25743 6239
rect 25685 6199 25743 6205
rect 19426 6168 19432 6180
rect 15856 6140 19432 6168
rect 15702 6131 15760 6137
rect 8588 6072 8984 6100
rect 7929 6063 7987 6069
rect 9950 6060 9956 6112
rect 10008 6100 10014 6112
rect 10045 6103 10103 6109
rect 10045 6100 10057 6103
rect 10008 6072 10057 6100
rect 10008 6060 10014 6072
rect 10045 6069 10057 6072
rect 10091 6069 10103 6103
rect 10045 6063 10103 6069
rect 13357 6103 13415 6109
rect 13357 6069 13369 6103
rect 13403 6100 13415 6103
rect 13538 6100 13544 6112
rect 13403 6072 13544 6100
rect 13403 6069 13415 6072
rect 13357 6063 13415 6069
rect 13538 6060 13544 6072
rect 13596 6060 13602 6112
rect 14090 6060 14096 6112
rect 14148 6100 14154 6112
rect 14323 6103 14381 6109
rect 14323 6100 14335 6103
rect 14148 6072 14335 6100
rect 14148 6060 14154 6072
rect 14323 6069 14335 6072
rect 14369 6069 14381 6103
rect 14323 6063 14381 6069
rect 15194 6060 15200 6112
rect 15252 6100 15258 6112
rect 15717 6100 15745 6131
rect 19426 6128 19432 6140
rect 19484 6128 19490 6180
rect 19889 6171 19947 6177
rect 19889 6137 19901 6171
rect 19935 6168 19947 6171
rect 20070 6168 20076 6180
rect 19935 6140 20076 6168
rect 19935 6137 19947 6140
rect 19889 6131 19947 6137
rect 20070 6128 20076 6140
rect 20128 6128 20134 6180
rect 20625 6171 20683 6177
rect 20625 6137 20637 6171
rect 20671 6168 20683 6171
rect 20806 6168 20812 6180
rect 20671 6140 20812 6168
rect 20671 6137 20683 6140
rect 20625 6131 20683 6137
rect 20806 6128 20812 6140
rect 20864 6168 20870 6180
rect 20864 6140 23704 6168
rect 20864 6128 20870 6140
rect 16298 6100 16304 6112
rect 15252 6072 15745 6100
rect 16259 6072 16304 6100
rect 15252 6060 15258 6072
rect 16298 6060 16304 6072
rect 16356 6060 16362 6112
rect 19518 6060 19524 6112
rect 19576 6100 19582 6112
rect 20165 6103 20223 6109
rect 20165 6100 20177 6103
rect 19576 6072 20177 6100
rect 19576 6060 19582 6072
rect 20165 6069 20177 6072
rect 20211 6069 20223 6103
rect 21818 6100 21824 6112
rect 21779 6072 21824 6100
rect 20165 6063 20223 6069
rect 21818 6060 21824 6072
rect 21876 6060 21882 6112
rect 23676 6100 23704 6140
rect 23753 6103 23811 6109
rect 23753 6100 23765 6103
rect 23676 6072 23765 6100
rect 23753 6069 23765 6072
rect 23799 6069 23811 6103
rect 23753 6063 23811 6069
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1210 5856 1216 5908
rect 1268 5896 1274 5908
rect 1535 5899 1593 5905
rect 1535 5896 1547 5899
rect 1268 5868 1547 5896
rect 1268 5856 1274 5868
rect 1535 5865 1547 5868
rect 1581 5865 1593 5899
rect 2130 5896 2136 5908
rect 2091 5868 2136 5896
rect 1535 5859 1593 5865
rect 2130 5856 2136 5868
rect 2188 5856 2194 5908
rect 2866 5896 2872 5908
rect 2827 5868 2872 5896
rect 2866 5856 2872 5868
rect 2924 5856 2930 5908
rect 3510 5896 3516 5908
rect 3471 5868 3516 5896
rect 3510 5856 3516 5868
rect 3568 5856 3574 5908
rect 3881 5899 3939 5905
rect 3881 5865 3893 5899
rect 3927 5896 3939 5899
rect 4338 5896 4344 5908
rect 3927 5868 4344 5896
rect 3927 5865 3939 5868
rect 3881 5859 3939 5865
rect 4338 5856 4344 5868
rect 4396 5856 4402 5908
rect 5166 5856 5172 5908
rect 5224 5896 5230 5908
rect 5353 5899 5411 5905
rect 5353 5896 5365 5899
rect 5224 5868 5365 5896
rect 5224 5856 5230 5868
rect 5353 5865 5365 5868
rect 5399 5865 5411 5899
rect 5353 5859 5411 5865
rect 5534 5856 5540 5908
rect 5592 5896 5598 5908
rect 5721 5899 5779 5905
rect 5721 5896 5733 5899
rect 5592 5868 5733 5896
rect 5592 5856 5598 5868
rect 5721 5865 5733 5868
rect 5767 5865 5779 5899
rect 7098 5896 7104 5908
rect 7059 5868 7104 5896
rect 5721 5859 5779 5865
rect 7098 5856 7104 5868
rect 7156 5856 7162 5908
rect 8938 5856 8944 5908
rect 8996 5896 9002 5908
rect 9033 5899 9091 5905
rect 9033 5896 9045 5899
rect 8996 5868 9045 5896
rect 8996 5856 9002 5868
rect 9033 5865 9045 5868
rect 9079 5865 9091 5899
rect 9033 5859 9091 5865
rect 11701 5899 11759 5905
rect 11701 5865 11713 5899
rect 11747 5896 11759 5899
rect 12250 5896 12256 5908
rect 11747 5868 12256 5896
rect 11747 5865 11759 5868
rect 11701 5859 11759 5865
rect 12250 5856 12256 5868
rect 12308 5856 12314 5908
rect 12713 5899 12771 5905
rect 12713 5865 12725 5899
rect 12759 5896 12771 5899
rect 15565 5899 15623 5905
rect 12759 5868 13768 5896
rect 12759 5865 12771 5868
rect 12713 5859 12771 5865
rect 13740 5840 13768 5868
rect 15565 5865 15577 5899
rect 15611 5896 15623 5899
rect 16390 5896 16396 5908
rect 15611 5868 16396 5896
rect 15611 5865 15623 5868
rect 15565 5859 15623 5865
rect 16390 5856 16396 5868
rect 16448 5856 16454 5908
rect 17494 5896 17500 5908
rect 17455 5868 17500 5896
rect 17494 5856 17500 5868
rect 17552 5856 17558 5908
rect 17586 5856 17592 5908
rect 17644 5896 17650 5908
rect 18417 5899 18475 5905
rect 18417 5896 18429 5899
rect 17644 5868 18429 5896
rect 17644 5856 17650 5868
rect 18417 5865 18429 5868
rect 18463 5865 18475 5899
rect 19242 5896 19248 5908
rect 19203 5868 19248 5896
rect 18417 5859 18475 5865
rect 19242 5856 19248 5868
rect 19300 5856 19306 5908
rect 20070 5856 20076 5908
rect 20128 5896 20134 5908
rect 20165 5899 20223 5905
rect 20165 5896 20177 5899
rect 20128 5868 20177 5896
rect 20128 5856 20134 5868
rect 20165 5865 20177 5868
rect 20211 5865 20223 5899
rect 24121 5899 24179 5905
rect 24121 5896 24133 5899
rect 20165 5859 20223 5865
rect 22296 5868 24133 5896
rect 4062 5788 4068 5840
rect 4120 5828 4126 5840
rect 4478 5831 4536 5837
rect 4478 5828 4490 5831
rect 4120 5800 4490 5828
rect 4120 5788 4126 5800
rect 4478 5797 4490 5800
rect 4524 5797 4536 5831
rect 5994 5828 6000 5840
rect 4478 5791 4536 5797
rect 5552 5800 6000 5828
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5760 1455 5763
rect 1486 5760 1492 5772
rect 1443 5732 1492 5760
rect 1443 5729 1455 5732
rect 1397 5723 1455 5729
rect 1486 5720 1492 5732
rect 1544 5720 1550 5772
rect 3050 5760 3056 5772
rect 2963 5732 3056 5760
rect 3050 5720 3056 5732
rect 3108 5760 3114 5772
rect 4982 5760 4988 5772
rect 3108 5732 4988 5760
rect 3108 5720 3114 5732
rect 4982 5720 4988 5732
rect 5040 5720 5046 5772
rect 5077 5763 5135 5769
rect 5077 5729 5089 5763
rect 5123 5760 5135 5763
rect 5552 5760 5580 5800
rect 5994 5788 6000 5800
rect 6052 5828 6058 5840
rect 6089 5831 6147 5837
rect 6089 5828 6101 5831
rect 6052 5800 6101 5828
rect 6052 5788 6058 5800
rect 6089 5797 6101 5800
rect 6135 5797 6147 5831
rect 6089 5791 6147 5797
rect 7834 5788 7840 5840
rect 7892 5828 7898 5840
rect 8205 5831 8263 5837
rect 8205 5828 8217 5831
rect 7892 5800 8217 5828
rect 7892 5788 7898 5800
rect 8205 5797 8217 5800
rect 8251 5797 8263 5831
rect 8205 5791 8263 5797
rect 10413 5831 10471 5837
rect 10413 5797 10425 5831
rect 10459 5828 10471 5831
rect 10686 5828 10692 5840
rect 10459 5800 10692 5828
rect 10459 5797 10471 5800
rect 10413 5791 10471 5797
rect 10686 5788 10692 5800
rect 10744 5788 10750 5840
rect 12155 5831 12213 5837
rect 12155 5797 12167 5831
rect 12201 5828 12213 5831
rect 12342 5828 12348 5840
rect 12201 5800 12348 5828
rect 12201 5797 12213 5800
rect 12155 5791 12213 5797
rect 12342 5788 12348 5800
rect 12400 5788 12406 5840
rect 13722 5828 13728 5840
rect 13635 5800 13728 5828
rect 13722 5788 13728 5800
rect 13780 5788 13786 5840
rect 15194 5788 15200 5840
rect 15252 5828 15258 5840
rect 15470 5828 15476 5840
rect 15252 5800 15476 5828
rect 15252 5788 15258 5800
rect 15470 5788 15476 5800
rect 15528 5828 15534 5840
rect 15978 5831 16036 5837
rect 15978 5828 15990 5831
rect 15528 5800 15990 5828
rect 15528 5788 15534 5800
rect 15978 5797 15990 5800
rect 16024 5797 16036 5831
rect 21358 5828 21364 5840
rect 15978 5791 16036 5797
rect 19168 5800 21364 5828
rect 5123 5732 5580 5760
rect 5123 5729 5135 5732
rect 5077 5723 5135 5729
rect 14274 5720 14280 5772
rect 14332 5760 14338 5772
rect 15286 5760 15292 5772
rect 14332 5732 15292 5760
rect 14332 5720 14338 5732
rect 15286 5720 15292 5732
rect 15344 5720 15350 5772
rect 15657 5763 15715 5769
rect 15657 5729 15669 5763
rect 15703 5760 15715 5763
rect 15838 5760 15844 5772
rect 15703 5732 15844 5760
rect 15703 5729 15715 5732
rect 15657 5723 15715 5729
rect 15838 5720 15844 5732
rect 15896 5720 15902 5772
rect 17402 5760 17408 5772
rect 17363 5732 17408 5760
rect 17402 5720 17408 5732
rect 17460 5720 17466 5772
rect 17957 5763 18015 5769
rect 17957 5729 17969 5763
rect 18003 5760 18015 5763
rect 18046 5760 18052 5772
rect 18003 5732 18052 5760
rect 18003 5729 18015 5732
rect 17957 5723 18015 5729
rect 18046 5720 18052 5732
rect 18104 5720 18110 5772
rect 18322 5720 18328 5772
rect 18380 5760 18386 5772
rect 19168 5769 19196 5800
rect 21358 5788 21364 5800
rect 21416 5788 21422 5840
rect 22296 5772 22324 5868
rect 24121 5865 24133 5868
rect 24167 5865 24179 5899
rect 24121 5859 24179 5865
rect 22643 5831 22701 5837
rect 22643 5797 22655 5831
rect 22689 5828 22701 5831
rect 22738 5828 22744 5840
rect 22689 5800 22744 5828
rect 22689 5797 22701 5800
rect 22643 5791 22701 5797
rect 22738 5788 22744 5800
rect 22796 5788 22802 5840
rect 23753 5831 23811 5837
rect 23753 5797 23765 5831
rect 23799 5828 23811 5831
rect 24302 5828 24308 5840
rect 23799 5800 24308 5828
rect 23799 5797 23811 5800
rect 23753 5791 23811 5797
rect 24302 5788 24308 5800
rect 24360 5828 24366 5840
rect 24360 5800 24624 5828
rect 24360 5788 24366 5800
rect 19153 5763 19211 5769
rect 19153 5760 19165 5763
rect 18380 5732 19165 5760
rect 18380 5720 18386 5732
rect 19153 5729 19165 5732
rect 19199 5729 19211 5763
rect 19153 5723 19211 5729
rect 19705 5763 19763 5769
rect 19705 5729 19717 5763
rect 19751 5760 19763 5763
rect 19978 5760 19984 5772
rect 19751 5732 19984 5760
rect 19751 5729 19763 5732
rect 19705 5723 19763 5729
rect 19978 5720 19984 5732
rect 20036 5720 20042 5772
rect 21266 5760 21272 5772
rect 21227 5732 21272 5760
rect 21266 5720 21272 5732
rect 21324 5720 21330 5772
rect 22002 5760 22008 5772
rect 21744 5732 22008 5760
rect 4154 5652 4160 5704
rect 4212 5692 4218 5704
rect 5997 5695 6055 5701
rect 4212 5664 4257 5692
rect 4212 5652 4218 5664
rect 5997 5661 6009 5695
rect 6043 5692 6055 5695
rect 6086 5692 6092 5704
rect 6043 5664 6092 5692
rect 6043 5661 6055 5664
rect 5997 5655 6055 5661
rect 6086 5652 6092 5664
rect 6144 5652 6150 5704
rect 6454 5692 6460 5704
rect 6415 5664 6460 5692
rect 6454 5652 6460 5664
rect 6512 5652 6518 5704
rect 7929 5695 7987 5701
rect 7929 5661 7941 5695
rect 7975 5692 7987 5695
rect 8113 5695 8171 5701
rect 8113 5692 8125 5695
rect 7975 5664 8125 5692
rect 7975 5661 7987 5664
rect 7929 5655 7987 5661
rect 8113 5661 8125 5664
rect 8159 5692 8171 5695
rect 9582 5692 9588 5704
rect 8159 5664 9588 5692
rect 8159 5661 8171 5664
rect 8113 5655 8171 5661
rect 9582 5652 9588 5664
rect 9640 5652 9646 5704
rect 10321 5695 10379 5701
rect 10321 5661 10333 5695
rect 10367 5692 10379 5695
rect 10962 5692 10968 5704
rect 10367 5664 10968 5692
rect 10367 5661 10379 5664
rect 10321 5655 10379 5661
rect 10962 5652 10968 5664
rect 11020 5652 11026 5704
rect 11793 5695 11851 5701
rect 11793 5661 11805 5695
rect 11839 5692 11851 5695
rect 11882 5692 11888 5704
rect 11839 5664 11888 5692
rect 11839 5661 11851 5664
rect 11793 5655 11851 5661
rect 11882 5652 11888 5664
rect 11940 5652 11946 5704
rect 13633 5695 13691 5701
rect 13633 5661 13645 5695
rect 13679 5661 13691 5695
rect 18874 5692 18880 5704
rect 13633 5655 13691 5661
rect 13786 5664 18880 5692
rect 2958 5584 2964 5636
rect 3016 5624 3022 5636
rect 5074 5624 5080 5636
rect 3016 5596 5080 5624
rect 3016 5584 3022 5596
rect 5074 5584 5080 5596
rect 5132 5584 5138 5636
rect 7561 5627 7619 5633
rect 7561 5593 7573 5627
rect 7607 5624 7619 5627
rect 8018 5624 8024 5636
rect 7607 5596 8024 5624
rect 7607 5593 7619 5596
rect 7561 5587 7619 5593
rect 8018 5584 8024 5596
rect 8076 5584 8082 5636
rect 8662 5624 8668 5636
rect 8623 5596 8668 5624
rect 8662 5584 8668 5596
rect 8720 5584 8726 5636
rect 10873 5627 10931 5633
rect 10873 5593 10885 5627
rect 10919 5624 10931 5627
rect 11514 5624 11520 5636
rect 10919 5596 11520 5624
rect 10919 5593 10931 5596
rect 10873 5587 10931 5593
rect 11514 5584 11520 5596
rect 11572 5624 11578 5636
rect 13357 5627 13415 5633
rect 13357 5624 13369 5627
rect 11572 5596 13369 5624
rect 11572 5584 11578 5596
rect 13357 5593 13369 5596
rect 13403 5624 13415 5627
rect 13648 5624 13676 5655
rect 13786 5624 13814 5664
rect 18874 5652 18880 5664
rect 18932 5652 18938 5704
rect 19996 5692 20024 5720
rect 21744 5701 21772 5732
rect 22002 5720 22008 5732
rect 22060 5720 22066 5772
rect 22278 5760 22284 5772
rect 22191 5732 22284 5760
rect 22278 5720 22284 5732
rect 22336 5720 22342 5772
rect 24210 5760 24216 5772
rect 23446 5732 24216 5760
rect 21729 5695 21787 5701
rect 21729 5692 21741 5695
rect 19996 5664 21741 5692
rect 21729 5661 21741 5664
rect 21775 5661 21787 5695
rect 21729 5655 21787 5661
rect 21910 5652 21916 5704
rect 21968 5692 21974 5704
rect 23446 5692 23474 5732
rect 24210 5720 24216 5732
rect 24268 5720 24274 5772
rect 24596 5769 24624 5800
rect 24581 5763 24639 5769
rect 24581 5729 24593 5763
rect 24627 5760 24639 5763
rect 25130 5760 25136 5772
rect 24627 5732 25136 5760
rect 24627 5729 24639 5732
rect 24581 5723 24639 5729
rect 25130 5720 25136 5732
rect 25188 5720 25194 5772
rect 21968 5664 23474 5692
rect 21968 5652 21974 5664
rect 13403 5596 13814 5624
rect 21407 5627 21465 5633
rect 13403 5593 13415 5596
rect 13357 5587 13415 5593
rect 21407 5593 21419 5627
rect 21453 5624 21465 5627
rect 23750 5624 23756 5636
rect 21453 5596 23756 5624
rect 21453 5593 21465 5596
rect 21407 5587 21465 5593
rect 23750 5584 23756 5596
rect 23808 5584 23814 5636
rect 3694 5516 3700 5568
rect 3752 5556 3758 5568
rect 9950 5556 9956 5568
rect 3752 5528 9956 5556
rect 3752 5516 3758 5528
rect 9950 5516 9956 5528
rect 10008 5516 10014 5568
rect 10134 5556 10140 5568
rect 10095 5528 10140 5556
rect 10134 5516 10140 5528
rect 10192 5516 10198 5568
rect 14550 5556 14556 5568
rect 14511 5528 14556 5556
rect 14550 5516 14556 5528
rect 14608 5516 14614 5568
rect 16574 5556 16580 5568
rect 16535 5528 16580 5556
rect 16574 5516 16580 5528
rect 16632 5516 16638 5568
rect 23198 5556 23204 5568
rect 23159 5528 23204 5556
rect 23198 5516 23204 5528
rect 23256 5516 23262 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1578 5352 1584 5364
rect 1539 5324 1584 5352
rect 1578 5312 1584 5324
rect 1636 5312 1642 5364
rect 2406 5312 2412 5364
rect 2464 5352 2470 5364
rect 2501 5355 2559 5361
rect 2501 5352 2513 5355
rect 2464 5324 2513 5352
rect 2464 5312 2470 5324
rect 2501 5321 2513 5324
rect 2547 5352 2559 5355
rect 3050 5352 3056 5364
rect 2547 5324 3056 5352
rect 2547 5321 2559 5324
rect 2501 5315 2559 5321
rect 3050 5312 3056 5324
rect 3108 5312 3114 5364
rect 4617 5355 4675 5361
rect 4617 5321 4629 5355
rect 4663 5352 4675 5355
rect 4890 5352 4896 5364
rect 4663 5324 4896 5352
rect 4663 5321 4675 5324
rect 4617 5315 4675 5321
rect 4890 5312 4896 5324
rect 4948 5312 4954 5364
rect 5994 5352 6000 5364
rect 5955 5324 6000 5352
rect 5994 5312 6000 5324
rect 6052 5312 6058 5364
rect 7834 5352 7840 5364
rect 7795 5324 7840 5352
rect 7834 5312 7840 5324
rect 7892 5312 7898 5364
rect 9030 5312 9036 5364
rect 9088 5352 9094 5364
rect 10873 5355 10931 5361
rect 10873 5352 10885 5355
rect 9088 5324 10885 5352
rect 9088 5312 9094 5324
rect 5353 5287 5411 5293
rect 5353 5253 5365 5287
rect 5399 5284 5411 5287
rect 5534 5284 5540 5296
rect 5399 5256 5540 5284
rect 5399 5253 5411 5256
rect 5353 5247 5411 5253
rect 5534 5244 5540 5256
rect 5592 5244 5598 5296
rect 7469 5287 7527 5293
rect 7469 5284 7481 5287
rect 6967 5256 7481 5284
rect 3881 5219 3939 5225
rect 3881 5185 3893 5219
rect 3927 5216 3939 5219
rect 4154 5216 4160 5228
rect 3927 5188 4160 5216
rect 3927 5185 3939 5188
rect 3881 5179 3939 5185
rect 4154 5176 4160 5188
rect 4212 5176 4218 5228
rect 4614 5176 4620 5228
rect 4672 5216 4678 5228
rect 4801 5219 4859 5225
rect 4801 5216 4813 5219
rect 4672 5188 4813 5216
rect 4672 5176 4678 5188
rect 4801 5185 4813 5188
rect 4847 5216 4859 5219
rect 6273 5219 6331 5225
rect 6273 5216 6285 5219
rect 4847 5188 6285 5216
rect 4847 5185 4859 5188
rect 4801 5179 4859 5185
rect 6273 5185 6285 5188
rect 6319 5185 6331 5219
rect 6273 5179 6331 5185
rect 1394 5148 1400 5160
rect 1355 5120 1400 5148
rect 1394 5108 1400 5120
rect 1452 5148 1458 5160
rect 1949 5151 2007 5157
rect 1949 5148 1961 5151
rect 1452 5120 1961 5148
rect 1452 5108 1458 5120
rect 1949 5117 1961 5120
rect 1995 5117 2007 5151
rect 1949 5111 2007 5117
rect 3053 5151 3111 5157
rect 3053 5117 3065 5151
rect 3099 5148 3111 5151
rect 3418 5148 3424 5160
rect 3099 5120 3424 5148
rect 3099 5117 3111 5120
rect 3053 5111 3111 5117
rect 3418 5108 3424 5120
rect 3476 5108 3482 5160
rect 3694 5148 3700 5160
rect 3655 5120 3700 5148
rect 3694 5108 3700 5120
rect 3752 5108 3758 5160
rect 6967 5157 6995 5256
rect 7469 5253 7481 5256
rect 7515 5284 7527 5287
rect 7926 5284 7932 5296
rect 7515 5256 7932 5284
rect 7515 5253 7527 5256
rect 7469 5247 7527 5253
rect 7926 5244 7932 5256
rect 7984 5284 7990 5296
rect 8570 5284 8576 5296
rect 7984 5256 8576 5284
rect 7984 5244 7990 5256
rect 8570 5244 8576 5256
rect 8628 5244 8634 5296
rect 9122 5244 9128 5296
rect 9180 5284 9186 5296
rect 9180 5256 9904 5284
rect 9180 5244 9186 5256
rect 9876 5228 9904 5256
rect 7055 5219 7113 5225
rect 7055 5185 7067 5219
rect 7101 5216 7113 5219
rect 8941 5219 8999 5225
rect 8941 5216 8953 5219
rect 7101 5188 8953 5216
rect 7101 5185 7113 5188
rect 7055 5179 7113 5185
rect 8941 5185 8953 5188
rect 8987 5216 8999 5219
rect 9585 5219 9643 5225
rect 9585 5216 9597 5219
rect 8987 5188 9597 5216
rect 8987 5185 8999 5188
rect 8941 5179 8999 5185
rect 9585 5185 9597 5188
rect 9631 5185 9643 5219
rect 9858 5216 9864 5228
rect 9819 5188 9864 5216
rect 9585 5179 9643 5185
rect 9858 5176 9864 5188
rect 9916 5176 9922 5228
rect 6952 5151 7010 5157
rect 6952 5117 6964 5151
rect 6998 5117 7010 5151
rect 10704 5148 10732 5324
rect 10873 5321 10885 5324
rect 10919 5321 10931 5355
rect 10873 5315 10931 5321
rect 11885 5355 11943 5361
rect 11885 5321 11897 5355
rect 11931 5352 11943 5355
rect 12161 5355 12219 5361
rect 12161 5352 12173 5355
rect 11931 5324 12173 5352
rect 11931 5321 11943 5324
rect 11885 5315 11943 5321
rect 12161 5321 12173 5324
rect 12207 5352 12219 5355
rect 12342 5352 12348 5364
rect 12207 5324 12348 5352
rect 12207 5321 12219 5324
rect 12161 5315 12219 5321
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 13722 5352 13728 5364
rect 13683 5324 13728 5352
rect 13722 5312 13728 5324
rect 13780 5312 13786 5364
rect 15381 5355 15439 5361
rect 15381 5321 15393 5355
rect 15427 5352 15439 5355
rect 15838 5352 15844 5364
rect 15427 5324 15844 5352
rect 15427 5321 15439 5324
rect 15381 5315 15439 5321
rect 15838 5312 15844 5324
rect 15896 5312 15902 5364
rect 17402 5352 17408 5364
rect 16592 5324 17408 5352
rect 11241 5287 11299 5293
rect 11241 5253 11253 5287
rect 11287 5284 11299 5287
rect 15930 5284 15936 5296
rect 11287 5256 15936 5284
rect 11287 5253 11299 5256
rect 11241 5247 11299 5253
rect 15930 5244 15936 5256
rect 15988 5284 15994 5296
rect 16592 5284 16620 5324
rect 17402 5312 17408 5324
rect 17460 5312 17466 5364
rect 17865 5355 17923 5361
rect 17865 5321 17877 5355
rect 17911 5352 17923 5355
rect 18046 5352 18052 5364
rect 17911 5324 18052 5352
rect 17911 5321 17923 5324
rect 17865 5315 17923 5321
rect 18046 5312 18052 5324
rect 18104 5312 18110 5364
rect 18322 5352 18328 5364
rect 18283 5324 18328 5352
rect 18322 5312 18328 5324
rect 18380 5312 18386 5364
rect 18555 5355 18613 5361
rect 18555 5321 18567 5355
rect 18601 5352 18613 5355
rect 20622 5352 20628 5364
rect 18601 5324 20628 5352
rect 18601 5321 18613 5324
rect 18555 5315 18613 5321
rect 20622 5312 20628 5324
rect 20680 5312 20686 5364
rect 22738 5312 22744 5364
rect 22796 5352 22802 5364
rect 23017 5355 23075 5361
rect 23017 5352 23029 5355
rect 22796 5324 23029 5352
rect 22796 5312 22802 5324
rect 23017 5321 23029 5324
rect 23063 5321 23075 5355
rect 23017 5315 23075 5321
rect 23198 5312 23204 5364
rect 23256 5352 23262 5364
rect 23385 5355 23443 5361
rect 23385 5352 23397 5355
rect 23256 5324 23397 5352
rect 23256 5312 23262 5324
rect 23385 5321 23397 5324
rect 23431 5352 23443 5355
rect 23842 5352 23848 5364
rect 23431 5324 23848 5352
rect 23431 5321 23443 5324
rect 23385 5315 23443 5321
rect 23842 5312 23848 5324
rect 23900 5312 23906 5364
rect 24210 5312 24216 5364
rect 24268 5352 24274 5364
rect 24673 5355 24731 5361
rect 24673 5352 24685 5355
rect 24268 5324 24685 5352
rect 24268 5312 24274 5324
rect 24673 5321 24685 5324
rect 24719 5321 24731 5355
rect 24673 5315 24731 5321
rect 15988 5256 16620 5284
rect 15988 5244 15994 5256
rect 16666 5244 16672 5296
rect 16724 5284 16730 5296
rect 16724 5256 17953 5284
rect 16724 5244 16730 5256
rect 10778 5176 10784 5228
rect 10836 5216 10842 5228
rect 12437 5219 12495 5225
rect 12437 5216 12449 5219
rect 10836 5188 12449 5216
rect 10836 5176 10842 5188
rect 12437 5185 12449 5188
rect 12483 5216 12495 5219
rect 12986 5216 12992 5228
rect 12483 5188 12992 5216
rect 12483 5185 12495 5188
rect 12437 5179 12495 5185
rect 12986 5176 12992 5188
rect 13044 5176 13050 5228
rect 14277 5219 14335 5225
rect 14277 5185 14289 5219
rect 14323 5216 14335 5219
rect 14550 5216 14556 5228
rect 14323 5188 14556 5216
rect 14323 5185 14335 5188
rect 14277 5179 14335 5185
rect 14550 5176 14556 5188
rect 14608 5176 14614 5228
rect 14921 5219 14979 5225
rect 14921 5185 14933 5219
rect 14967 5216 14979 5219
rect 15286 5216 15292 5228
rect 14967 5188 15292 5216
rect 14967 5185 14979 5188
rect 14921 5179 14979 5185
rect 15286 5176 15292 5188
rect 15344 5176 15350 5228
rect 15470 5176 15476 5228
rect 15528 5216 15534 5228
rect 15657 5219 15715 5225
rect 15657 5216 15669 5219
rect 15528 5188 15669 5216
rect 15528 5176 15534 5188
rect 15657 5185 15669 5188
rect 15703 5185 15715 5219
rect 15657 5179 15715 5185
rect 16301 5219 16359 5225
rect 16301 5185 16313 5219
rect 16347 5216 16359 5219
rect 16758 5216 16764 5228
rect 16347 5188 16764 5216
rect 16347 5185 16359 5188
rect 16301 5179 16359 5185
rect 16758 5176 16764 5188
rect 16816 5176 16822 5228
rect 11057 5151 11115 5157
rect 11057 5148 11069 5151
rect 10704 5120 11069 5148
rect 6952 5111 7010 5117
rect 11057 5117 11069 5120
rect 11103 5117 11115 5151
rect 11057 5111 11115 5117
rect 13357 5151 13415 5157
rect 13357 5117 13369 5151
rect 13403 5148 13415 5151
rect 14001 5151 14059 5157
rect 14001 5148 14013 5151
rect 13403 5120 14013 5148
rect 13403 5117 13415 5120
rect 13357 5111 13415 5117
rect 14001 5117 14013 5120
rect 14047 5117 14059 5151
rect 17925 5148 17953 5256
rect 19978 5244 19984 5296
rect 20036 5284 20042 5296
rect 20717 5287 20775 5293
rect 20717 5284 20729 5287
rect 20036 5256 20729 5284
rect 20036 5244 20042 5256
rect 20717 5253 20729 5256
rect 20763 5253 20775 5287
rect 20717 5247 20775 5253
rect 21174 5244 21180 5296
rect 21232 5284 21238 5296
rect 21232 5256 24072 5284
rect 21232 5244 21238 5256
rect 19521 5219 19579 5225
rect 19521 5185 19533 5219
rect 19567 5216 19579 5219
rect 20070 5216 20076 5228
rect 19567 5188 20076 5216
rect 19567 5185 19579 5188
rect 19521 5179 19579 5185
rect 20070 5176 20076 5188
rect 20128 5176 20134 5228
rect 21818 5216 21824 5228
rect 21779 5188 21824 5216
rect 21818 5176 21824 5188
rect 21876 5176 21882 5228
rect 24044 5225 24072 5256
rect 24029 5219 24087 5225
rect 24029 5185 24041 5219
rect 24075 5185 24087 5219
rect 24029 5179 24087 5185
rect 24118 5176 24124 5228
rect 24176 5216 24182 5228
rect 25225 5219 25283 5225
rect 25225 5216 25237 5219
rect 24176 5188 25237 5216
rect 24176 5176 24182 5188
rect 25225 5185 25237 5188
rect 25271 5185 25283 5219
rect 25225 5179 25283 5185
rect 18452 5151 18510 5157
rect 18452 5148 18464 5151
rect 17925 5120 18464 5148
rect 14001 5111 14059 5117
rect 18452 5117 18464 5120
rect 18498 5148 18510 5151
rect 18877 5151 18935 5157
rect 18877 5148 18889 5151
rect 18498 5120 18889 5148
rect 18498 5117 18510 5120
rect 18452 5111 18510 5117
rect 18877 5117 18889 5120
rect 18923 5148 18935 5151
rect 19150 5148 19156 5160
rect 18923 5120 19156 5148
rect 18923 5117 18935 5120
rect 18877 5111 18935 5117
rect 4522 5040 4528 5092
rect 4580 5080 4586 5092
rect 4798 5080 4804 5092
rect 4580 5052 4804 5080
rect 4580 5040 4586 5052
rect 4798 5040 4804 5052
rect 4856 5040 4862 5092
rect 4890 5040 4896 5092
rect 4948 5080 4954 5092
rect 8018 5080 8024 5092
rect 4948 5052 4993 5080
rect 7979 5052 8024 5080
rect 4948 5040 4954 5052
rect 8018 5040 8024 5052
rect 8076 5040 8082 5092
rect 8113 5083 8171 5089
rect 8113 5049 8125 5083
rect 8159 5049 8171 5083
rect 8662 5080 8668 5092
rect 8623 5052 8668 5080
rect 8113 5043 8171 5049
rect 4062 4972 4068 5024
rect 4120 5012 4126 5024
rect 4157 5015 4215 5021
rect 4157 5012 4169 5015
rect 4120 4984 4169 5012
rect 4120 4972 4126 4984
rect 4157 4981 4169 4984
rect 4203 4981 4215 5015
rect 8128 5012 8156 5043
rect 8662 5040 8668 5052
rect 8720 5040 8726 5092
rect 9401 5083 9459 5089
rect 9401 5049 9413 5083
rect 9447 5080 9459 5083
rect 9677 5083 9735 5089
rect 9677 5080 9689 5083
rect 9447 5052 9689 5080
rect 9447 5049 9459 5052
rect 9401 5043 9459 5049
rect 9677 5049 9689 5052
rect 9723 5049 9735 5083
rect 9677 5043 9735 5049
rect 8294 5012 8300 5024
rect 8128 4984 8300 5012
rect 4157 4975 4215 4981
rect 8294 4972 8300 4984
rect 8352 5012 8358 5024
rect 9416 5012 9444 5043
rect 12342 5040 12348 5092
rect 12400 5080 12406 5092
rect 12758 5083 12816 5089
rect 12758 5080 12770 5083
rect 12400 5052 12770 5080
rect 12400 5040 12406 5052
rect 12758 5049 12770 5052
rect 12804 5049 12816 5083
rect 12758 5043 12816 5049
rect 8352 4984 9444 5012
rect 10597 5015 10655 5021
rect 8352 4972 8358 4984
rect 10597 4981 10609 5015
rect 10643 5012 10655 5015
rect 10686 5012 10692 5024
rect 10643 4984 10692 5012
rect 10643 4981 10655 4984
rect 10597 4975 10655 4981
rect 10686 4972 10692 4984
rect 10744 4972 10750 5024
rect 14016 5012 14044 5111
rect 19150 5108 19156 5120
rect 19208 5108 19214 5160
rect 19334 5108 19340 5160
rect 19392 5148 19398 5160
rect 19429 5151 19487 5157
rect 19429 5148 19441 5151
rect 19392 5120 19441 5148
rect 19392 5108 19398 5120
rect 19429 5117 19441 5120
rect 19475 5148 19487 5151
rect 20990 5148 20996 5160
rect 19475 5120 20996 5148
rect 19475 5117 19487 5120
rect 19429 5111 19487 5117
rect 14369 5083 14427 5089
rect 14369 5049 14381 5083
rect 14415 5049 14427 5083
rect 14369 5043 14427 5049
rect 14384 5012 14412 5043
rect 15930 5040 15936 5092
rect 15988 5080 15994 5092
rect 16117 5083 16175 5089
rect 16117 5080 16129 5083
rect 15988 5052 16129 5080
rect 15988 5040 15994 5052
rect 16117 5049 16129 5052
rect 16163 5080 16175 5083
rect 16393 5083 16451 5089
rect 16393 5080 16405 5083
rect 16163 5052 16405 5080
rect 16163 5049 16175 5052
rect 16117 5043 16175 5049
rect 16393 5049 16405 5052
rect 16439 5080 16451 5083
rect 16574 5080 16580 5092
rect 16439 5052 16580 5080
rect 16439 5049 16451 5052
rect 16393 5043 16451 5049
rect 16574 5040 16580 5052
rect 16632 5040 16638 5092
rect 16666 5040 16672 5092
rect 16724 5080 16730 5092
rect 19857 5089 19885 5120
rect 20990 5108 20996 5120
rect 21048 5148 21054 5160
rect 21637 5151 21695 5157
rect 21637 5148 21649 5151
rect 21048 5120 21649 5148
rect 21048 5108 21054 5120
rect 21637 5117 21649 5120
rect 21683 5148 21695 5151
rect 21683 5120 22185 5148
rect 21683 5117 21695 5120
rect 21637 5111 21695 5117
rect 22157 5089 22185 5120
rect 16945 5083 17003 5089
rect 16945 5080 16957 5083
rect 16724 5052 16957 5080
rect 16724 5040 16730 5052
rect 16945 5049 16957 5052
rect 16991 5049 17003 5083
rect 19842 5083 19900 5089
rect 19842 5080 19854 5083
rect 19820 5052 19854 5080
rect 16945 5043 17003 5049
rect 19842 5049 19854 5052
rect 19888 5049 19900 5083
rect 19842 5043 19900 5049
rect 22142 5083 22200 5089
rect 22142 5049 22154 5083
rect 22188 5049 22200 5083
rect 23750 5080 23756 5092
rect 23711 5052 23756 5080
rect 22142 5043 22200 5049
rect 23750 5040 23756 5052
rect 23808 5040 23814 5092
rect 23842 5040 23848 5092
rect 23900 5080 23906 5092
rect 23900 5052 23945 5080
rect 23900 5040 23906 5052
rect 20438 5012 20444 5024
rect 14016 4984 14412 5012
rect 20399 4984 20444 5012
rect 20438 4972 20444 4984
rect 20496 4972 20502 5024
rect 21266 5012 21272 5024
rect 21227 4984 21272 5012
rect 21266 4972 21272 4984
rect 21324 4972 21330 5024
rect 22738 5012 22744 5024
rect 22699 4984 22744 5012
rect 22738 4972 22744 4984
rect 22796 4972 22802 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1118 4768 1124 4820
rect 1176 4808 1182 4820
rect 1581 4811 1639 4817
rect 1581 4808 1593 4811
rect 1176 4780 1593 4808
rect 1176 4768 1182 4780
rect 1581 4777 1593 4780
rect 1627 4777 1639 4811
rect 1581 4771 1639 4777
rect 2087 4811 2145 4817
rect 2087 4777 2099 4811
rect 2133 4808 2145 4811
rect 2498 4808 2504 4820
rect 2133 4780 2504 4808
rect 2133 4777 2145 4780
rect 2087 4771 2145 4777
rect 2498 4768 2504 4780
rect 2556 4768 2562 4820
rect 3513 4811 3571 4817
rect 3513 4777 3525 4811
rect 3559 4808 3571 4811
rect 3694 4808 3700 4820
rect 3559 4780 3700 4808
rect 3559 4777 3571 4780
rect 3513 4771 3571 4777
rect 3694 4768 3700 4780
rect 3752 4768 3758 4820
rect 3881 4811 3939 4817
rect 3881 4777 3893 4811
rect 3927 4808 3939 4811
rect 4154 4808 4160 4820
rect 3927 4780 4160 4808
rect 3927 4777 3939 4780
rect 3881 4771 3939 4777
rect 4154 4768 4160 4780
rect 4212 4768 4218 4820
rect 7190 4768 7196 4820
rect 7248 4808 7254 4820
rect 7377 4811 7435 4817
rect 7377 4808 7389 4811
rect 7248 4780 7389 4808
rect 7248 4768 7254 4780
rect 7377 4777 7389 4780
rect 7423 4777 7435 4811
rect 7377 4771 7435 4777
rect 7929 4811 7987 4817
rect 7929 4777 7941 4811
rect 7975 4808 7987 4811
rect 8294 4808 8300 4820
rect 7975 4780 8300 4808
rect 7975 4777 7987 4780
rect 7929 4771 7987 4777
rect 8294 4768 8300 4780
rect 8352 4768 8358 4820
rect 12986 4808 12992 4820
rect 12947 4780 12992 4808
rect 12986 4768 12992 4780
rect 13044 4768 13050 4820
rect 15657 4811 15715 4817
rect 15657 4777 15669 4811
rect 15703 4808 15715 4811
rect 15746 4808 15752 4820
rect 15703 4780 15752 4808
rect 15703 4777 15715 4780
rect 15657 4771 15715 4777
rect 3099 4743 3157 4749
rect 3099 4709 3111 4743
rect 3145 4740 3157 4743
rect 4614 4740 4620 4752
rect 3145 4712 4620 4740
rect 3145 4709 3157 4712
rect 3099 4703 3157 4709
rect 4614 4700 4620 4712
rect 4672 4700 4678 4752
rect 4890 4740 4896 4752
rect 4851 4712 4896 4740
rect 4890 4700 4896 4712
rect 4948 4700 4954 4752
rect 5445 4743 5503 4749
rect 5445 4709 5457 4743
rect 5491 4740 5503 4743
rect 5997 4743 6055 4749
rect 5997 4740 6009 4743
rect 5491 4712 6009 4740
rect 5491 4709 5503 4712
rect 5445 4703 5503 4709
rect 5997 4709 6009 4712
rect 6043 4740 6055 4743
rect 6086 4740 6092 4752
rect 6043 4712 6092 4740
rect 6043 4709 6055 4712
rect 5997 4703 6055 4709
rect 6086 4700 6092 4712
rect 6144 4740 6150 4752
rect 8662 4740 8668 4752
rect 6144 4712 8668 4740
rect 6144 4700 6150 4712
rect 8662 4700 8668 4712
rect 8720 4700 8726 4752
rect 11790 4749 11796 4752
rect 11787 4740 11796 4749
rect 11703 4712 11796 4740
rect 11787 4703 11796 4712
rect 11848 4740 11854 4752
rect 12342 4740 12348 4752
rect 11848 4712 12348 4740
rect 11790 4700 11796 4703
rect 11848 4700 11854 4712
rect 12342 4700 12348 4712
rect 12400 4700 12406 4752
rect 13446 4740 13452 4752
rect 13407 4712 13452 4740
rect 13446 4700 13452 4712
rect 13504 4700 13510 4752
rect 13538 4700 13544 4752
rect 13596 4740 13602 4752
rect 14093 4743 14151 4749
rect 13596 4712 13641 4740
rect 13596 4700 13602 4712
rect 14093 4709 14105 4743
rect 14139 4740 14151 4743
rect 14274 4740 14280 4752
rect 14139 4712 14280 4740
rect 14139 4709 14151 4712
rect 14093 4703 14151 4709
rect 14274 4700 14280 4712
rect 14332 4700 14338 4752
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4672 1915 4675
rect 1946 4672 1952 4684
rect 1903 4644 1952 4672
rect 1903 4641 1915 4644
rect 1857 4635 1915 4641
rect 1946 4632 1952 4644
rect 2004 4632 2010 4684
rect 2958 4672 2964 4684
rect 2919 4644 2964 4672
rect 2958 4632 2964 4644
rect 3016 4632 3022 4684
rect 7466 4632 7472 4684
rect 7524 4672 7530 4684
rect 9214 4672 9220 4684
rect 7524 4644 9220 4672
rect 7524 4632 7530 4644
rect 9214 4632 9220 4644
rect 9272 4672 9278 4684
rect 9858 4672 9864 4684
rect 9272 4644 9864 4672
rect 9272 4632 9278 4644
rect 9858 4632 9864 4644
rect 9916 4632 9922 4684
rect 10134 4632 10140 4684
rect 10192 4672 10198 4684
rect 10321 4675 10379 4681
rect 10321 4672 10333 4675
rect 10192 4644 10333 4672
rect 10192 4632 10198 4644
rect 10321 4641 10333 4644
rect 10367 4641 10379 4675
rect 10321 4635 10379 4641
rect 10597 4675 10655 4681
rect 10597 4641 10609 4675
rect 10643 4672 10655 4675
rect 11882 4672 11888 4684
rect 10643 4644 11888 4672
rect 10643 4641 10655 4644
rect 10597 4635 10655 4641
rect 11882 4632 11888 4644
rect 11940 4672 11946 4684
rect 12621 4675 12679 4681
rect 12621 4672 12633 4675
rect 11940 4644 12633 4672
rect 11940 4632 11946 4644
rect 12621 4641 12633 4644
rect 12667 4641 12679 4675
rect 12621 4635 12679 4641
rect 4798 4604 4804 4616
rect 4759 4576 4804 4604
rect 4798 4564 4804 4576
rect 4856 4564 4862 4616
rect 6914 4564 6920 4616
rect 6972 4604 6978 4616
rect 7009 4607 7067 4613
rect 7009 4604 7021 4607
rect 6972 4576 7021 4604
rect 6972 4564 6978 4576
rect 7009 4573 7021 4576
rect 7055 4573 7067 4607
rect 7009 4567 7067 4573
rect 11146 4564 11152 4616
rect 11204 4604 11210 4616
rect 11425 4607 11483 4613
rect 11425 4604 11437 4607
rect 11204 4576 11437 4604
rect 11204 4564 11210 4576
rect 11425 4573 11437 4576
rect 11471 4573 11483 4607
rect 15672 4604 15700 4771
rect 15746 4768 15752 4780
rect 15804 4768 15810 4820
rect 16758 4808 16764 4820
rect 16719 4780 16764 4808
rect 16758 4768 16764 4780
rect 16816 4768 16822 4820
rect 19334 4768 19340 4820
rect 19392 4808 19398 4820
rect 19429 4811 19487 4817
rect 19429 4808 19441 4811
rect 19392 4780 19441 4808
rect 19392 4768 19398 4780
rect 19429 4777 19441 4780
rect 19475 4777 19487 4811
rect 19429 4771 19487 4777
rect 19981 4811 20039 4817
rect 19981 4777 19993 4811
rect 20027 4808 20039 4811
rect 20898 4808 20904 4820
rect 20027 4780 20904 4808
rect 20027 4777 20039 4780
rect 19981 4771 20039 4777
rect 20898 4768 20904 4780
rect 20956 4808 20962 4820
rect 20956 4780 21128 4808
rect 20956 4768 20962 4780
rect 15930 4740 15936 4752
rect 15891 4712 15936 4740
rect 15930 4700 15936 4712
rect 15988 4700 15994 4752
rect 17218 4700 17224 4752
rect 17276 4740 17282 4752
rect 17402 4740 17408 4752
rect 17276 4712 17408 4740
rect 17276 4700 17282 4712
rect 17402 4700 17408 4712
rect 17460 4740 17466 4752
rect 21100 4749 21128 4780
rect 21818 4768 21824 4820
rect 21876 4808 21882 4820
rect 21913 4811 21971 4817
rect 21913 4808 21925 4811
rect 21876 4780 21925 4808
rect 21876 4768 21882 4780
rect 21913 4777 21925 4780
rect 21959 4777 21971 4811
rect 22278 4808 22284 4820
rect 22239 4780 22284 4808
rect 21913 4771 21971 4777
rect 22278 4768 22284 4780
rect 22336 4768 22342 4820
rect 23750 4768 23756 4820
rect 23808 4808 23814 4820
rect 24397 4811 24455 4817
rect 24397 4808 24409 4811
rect 23808 4780 24409 4808
rect 23808 4768 23814 4780
rect 24397 4777 24409 4780
rect 24443 4777 24455 4811
rect 24762 4808 24768 4820
rect 24723 4780 24768 4808
rect 24397 4771 24455 4777
rect 24762 4768 24768 4780
rect 24820 4768 24826 4820
rect 17634 4743 17692 4749
rect 17634 4740 17646 4743
rect 17460 4712 17646 4740
rect 17460 4700 17466 4712
rect 17634 4709 17646 4712
rect 17680 4709 17692 4743
rect 17634 4703 17692 4709
rect 21085 4743 21143 4749
rect 21085 4709 21097 4743
rect 21131 4709 21143 4743
rect 21085 4703 21143 4709
rect 22738 4700 22744 4752
rect 22796 4740 22802 4752
rect 23017 4743 23075 4749
rect 23017 4740 23029 4743
rect 22796 4712 23029 4740
rect 22796 4700 22802 4712
rect 23017 4709 23029 4712
rect 23063 4709 23075 4743
rect 23017 4703 23075 4709
rect 17313 4675 17371 4681
rect 17313 4641 17325 4675
rect 17359 4672 17371 4675
rect 17494 4672 17500 4684
rect 17359 4644 17500 4672
rect 17359 4641 17371 4644
rect 17313 4635 17371 4641
rect 17494 4632 17500 4644
rect 17552 4632 17558 4684
rect 19061 4675 19119 4681
rect 19061 4641 19073 4675
rect 19107 4672 19119 4675
rect 19242 4672 19248 4684
rect 19107 4644 19248 4672
rect 19107 4641 19119 4644
rect 19061 4635 19119 4641
rect 19242 4632 19248 4644
rect 19300 4632 19306 4684
rect 24578 4672 24584 4684
rect 24539 4644 24584 4672
rect 24578 4632 24584 4644
rect 24636 4632 24642 4684
rect 15841 4607 15899 4613
rect 15841 4604 15853 4607
rect 11425 4567 11483 4573
rect 13786 4576 14596 4604
rect 15672 4576 15853 4604
rect 10962 4536 10968 4548
rect 10875 4508 10968 4536
rect 10962 4496 10968 4508
rect 11020 4536 11026 4548
rect 13786 4536 13814 4576
rect 11020 4508 13814 4536
rect 11020 4496 11026 4508
rect 4246 4468 4252 4480
rect 4207 4440 4252 4468
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 8846 4468 8852 4480
rect 8807 4440 8852 4468
rect 8846 4428 8852 4440
rect 8904 4428 8910 4480
rect 10686 4428 10692 4480
rect 10744 4468 10750 4480
rect 12345 4471 12403 4477
rect 12345 4468 12357 4471
rect 10744 4440 12357 4468
rect 10744 4428 10750 4440
rect 12345 4437 12357 4440
rect 12391 4468 12403 4471
rect 12894 4468 12900 4480
rect 12391 4440 12900 4468
rect 12391 4437 12403 4440
rect 12345 4431 12403 4437
rect 12894 4428 12900 4440
rect 12952 4468 12958 4480
rect 13354 4468 13360 4480
rect 12952 4440 13360 4468
rect 12952 4428 12958 4440
rect 13354 4428 13360 4440
rect 13412 4428 13418 4480
rect 14458 4468 14464 4480
rect 14419 4440 14464 4468
rect 14458 4428 14464 4440
rect 14516 4428 14522 4480
rect 14568 4468 14596 4576
rect 15841 4573 15853 4576
rect 15887 4573 15899 4607
rect 16206 4604 16212 4616
rect 16167 4576 16212 4604
rect 15841 4567 15899 4573
rect 16206 4564 16212 4576
rect 16264 4564 16270 4616
rect 20990 4604 20996 4616
rect 20951 4576 20996 4604
rect 20990 4564 20996 4576
rect 21048 4564 21054 4616
rect 21266 4604 21272 4616
rect 21227 4576 21272 4604
rect 21266 4564 21272 4576
rect 21324 4564 21330 4616
rect 22922 4604 22928 4616
rect 22883 4576 22928 4604
rect 22922 4564 22928 4576
rect 22980 4564 22986 4616
rect 23201 4607 23259 4613
rect 23201 4573 23213 4607
rect 23247 4604 23259 4607
rect 24026 4604 24032 4616
rect 23247 4576 24032 4604
rect 23247 4573 23259 4576
rect 23201 4567 23259 4573
rect 21284 4536 21312 4564
rect 23216 4536 23244 4567
rect 24026 4564 24032 4576
rect 24084 4564 24090 4616
rect 21284 4508 23244 4536
rect 24210 4496 24216 4548
rect 24268 4536 24274 4548
rect 25590 4536 25596 4548
rect 24268 4508 25596 4536
rect 24268 4496 24274 4508
rect 25590 4496 25596 4508
rect 25648 4496 25654 4548
rect 16758 4468 16764 4480
rect 14568 4440 16764 4468
rect 16758 4428 16764 4440
rect 16816 4428 16822 4480
rect 18230 4468 18236 4480
rect 18191 4440 18236 4468
rect 18230 4428 18236 4440
rect 18288 4428 18294 4480
rect 18598 4468 18604 4480
rect 18559 4440 18604 4468
rect 18598 4428 18604 4440
rect 18656 4428 18662 4480
rect 24121 4471 24179 4477
rect 24121 4437 24133 4471
rect 24167 4468 24179 4471
rect 25130 4468 25136 4480
rect 24167 4440 25136 4468
rect 24167 4437 24179 4440
rect 24121 4431 24179 4437
rect 25130 4428 25136 4440
rect 25188 4428 25194 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1486 4224 1492 4276
rect 1544 4264 1550 4276
rect 1581 4267 1639 4273
rect 1581 4264 1593 4267
rect 1544 4236 1593 4264
rect 1544 4224 1550 4236
rect 1581 4233 1593 4236
rect 1627 4233 1639 4267
rect 1946 4264 1952 4276
rect 1907 4236 1952 4264
rect 1581 4227 1639 4233
rect 1946 4224 1952 4236
rect 2004 4224 2010 4276
rect 2271 4267 2329 4273
rect 2271 4233 2283 4267
rect 2317 4264 2329 4267
rect 2317 4236 4154 4264
rect 2317 4233 2329 4236
rect 2271 4227 2329 4233
rect 2958 4196 2964 4208
rect 2919 4168 2964 4196
rect 2958 4156 2964 4168
rect 3016 4156 3022 4208
rect 4126 4196 4154 4236
rect 4890 4224 4896 4276
rect 4948 4264 4954 4276
rect 5077 4267 5135 4273
rect 5077 4264 5089 4267
rect 4948 4236 5089 4264
rect 4948 4224 4954 4236
rect 5077 4233 5089 4236
rect 5123 4264 5135 4267
rect 5353 4267 5411 4273
rect 5353 4264 5365 4267
rect 5123 4236 5365 4264
rect 5123 4233 5135 4236
rect 5077 4227 5135 4233
rect 5353 4233 5365 4236
rect 5399 4233 5411 4267
rect 5353 4227 5411 4233
rect 11146 4224 11152 4276
rect 11204 4264 11210 4276
rect 12161 4267 12219 4273
rect 12161 4264 12173 4267
rect 11204 4236 12173 4264
rect 11204 4224 11210 4236
rect 12161 4233 12173 4236
rect 12207 4233 12219 4267
rect 13538 4264 13544 4276
rect 13499 4236 13544 4264
rect 12161 4227 12219 4233
rect 13538 4224 13544 4236
rect 13596 4224 13602 4276
rect 14550 4264 14556 4276
rect 13648 4236 14556 4264
rect 13648 4208 13676 4236
rect 14550 4224 14556 4236
rect 14608 4224 14614 4276
rect 15381 4267 15439 4273
rect 15381 4233 15393 4267
rect 15427 4264 15439 4267
rect 15930 4264 15936 4276
rect 15427 4236 15936 4264
rect 15427 4233 15439 4236
rect 15381 4227 15439 4233
rect 15930 4224 15936 4236
rect 15988 4224 15994 4276
rect 17037 4267 17095 4273
rect 17037 4233 17049 4267
rect 17083 4264 17095 4267
rect 17494 4264 17500 4276
rect 17083 4236 17500 4264
rect 17083 4233 17095 4236
rect 17037 4227 17095 4233
rect 17494 4224 17500 4236
rect 17552 4224 17558 4276
rect 17865 4267 17923 4273
rect 17865 4233 17877 4267
rect 17911 4264 17923 4267
rect 18230 4264 18236 4276
rect 17911 4236 18236 4264
rect 17911 4233 17923 4236
rect 17865 4227 17923 4233
rect 18230 4224 18236 4236
rect 18288 4224 18294 4276
rect 19242 4224 19248 4276
rect 19300 4264 19306 4276
rect 19705 4267 19763 4273
rect 19705 4264 19717 4267
rect 19300 4236 19717 4264
rect 19300 4224 19306 4236
rect 19705 4233 19717 4236
rect 19751 4233 19763 4267
rect 20898 4264 20904 4276
rect 20859 4236 20904 4264
rect 19705 4227 19763 4233
rect 20898 4224 20904 4236
rect 20956 4224 20962 4276
rect 22738 4224 22744 4276
rect 22796 4264 22802 4276
rect 23293 4267 23351 4273
rect 23293 4264 23305 4267
rect 22796 4236 23305 4264
rect 22796 4224 22802 4236
rect 23293 4233 23305 4236
rect 23339 4233 23351 4267
rect 23293 4227 23351 4233
rect 24026 4224 24032 4276
rect 24084 4264 24090 4276
rect 24811 4267 24869 4273
rect 24811 4264 24823 4267
rect 24084 4236 24823 4264
rect 24084 4224 24090 4236
rect 24811 4233 24823 4236
rect 24857 4233 24869 4267
rect 25222 4264 25228 4276
rect 25183 4236 25228 4264
rect 24811 4227 24869 4233
rect 25222 4224 25228 4236
rect 25280 4224 25286 4276
rect 9766 4196 9772 4208
rect 4126 4168 9772 4196
rect 9766 4156 9772 4168
rect 9824 4156 9830 4208
rect 9858 4156 9864 4208
rect 9916 4196 9922 4208
rect 13357 4199 13415 4205
rect 9916 4168 9961 4196
rect 9916 4156 9922 4168
rect 13357 4165 13369 4199
rect 13403 4196 13415 4199
rect 13630 4196 13636 4208
rect 13403 4168 13636 4196
rect 13403 4165 13415 4168
rect 13357 4159 13415 4165
rect 13630 4156 13636 4168
rect 13688 4156 13694 4208
rect 16666 4156 16672 4208
rect 16724 4196 16730 4208
rect 19334 4196 19340 4208
rect 16724 4168 18736 4196
rect 19295 4168 19340 4196
rect 16724 4156 16730 4168
rect 2590 4088 2596 4140
rect 2648 4128 2654 4140
rect 2685 4131 2743 4137
rect 2685 4128 2697 4131
rect 2648 4100 2697 4128
rect 2648 4088 2654 4100
rect 2685 4097 2697 4100
rect 2731 4128 2743 4131
rect 3510 4128 3516 4140
rect 2731 4100 3516 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 3510 4088 3516 4100
rect 3568 4088 3574 4140
rect 4062 4128 4068 4140
rect 3988 4100 4068 4128
rect 2200 4063 2258 4069
rect 2200 4029 2212 4063
rect 2246 4060 2258 4063
rect 2608 4060 2636 4088
rect 2246 4032 2636 4060
rect 3145 4063 3203 4069
rect 2246 4029 2258 4032
rect 2200 4023 2258 4029
rect 3145 4029 3157 4063
rect 3191 4060 3203 4063
rect 3602 4060 3608 4072
rect 3191 4032 3608 4060
rect 3191 4029 3203 4032
rect 3145 4023 3203 4029
rect 3602 4020 3608 4032
rect 3660 4020 3666 4072
rect 1762 3952 1768 4004
rect 1820 3992 1826 4004
rect 3988 4001 4016 4100
rect 4062 4088 4068 4100
rect 4120 4088 4126 4140
rect 4157 4131 4215 4137
rect 4157 4097 4169 4131
rect 4203 4128 4215 4131
rect 4246 4128 4252 4140
rect 4203 4100 4252 4128
rect 4203 4097 4215 4100
rect 4157 4091 4215 4097
rect 4246 4088 4252 4100
rect 4304 4088 4310 4140
rect 6270 4088 6276 4140
rect 6328 4128 6334 4140
rect 8846 4128 8852 4140
rect 6328 4100 8852 4128
rect 6328 4088 6334 4100
rect 8846 4088 8852 4100
rect 8904 4088 8910 4140
rect 9122 4128 9128 4140
rect 9083 4100 9128 4128
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 10689 4131 10747 4137
rect 10689 4097 10701 4131
rect 10735 4128 10747 4131
rect 10962 4128 10968 4140
rect 10735 4100 10968 4128
rect 10735 4097 10747 4100
rect 10689 4091 10747 4097
rect 10962 4088 10968 4100
rect 11020 4088 11026 4140
rect 11514 4128 11520 4140
rect 11475 4100 11520 4128
rect 11514 4088 11520 4100
rect 11572 4088 11578 4140
rect 12805 4131 12863 4137
rect 12805 4097 12817 4131
rect 12851 4128 12863 4131
rect 14369 4131 14427 4137
rect 12851 4100 13814 4128
rect 12851 4097 12863 4100
rect 12805 4091 12863 4097
rect 7006 4060 7012 4072
rect 6967 4032 7012 4060
rect 7006 4020 7012 4032
rect 7064 4020 7070 4072
rect 3973 3995 4031 4001
rect 3973 3992 3985 3995
rect 1820 3964 3985 3992
rect 1820 3952 1826 3964
rect 3973 3961 3985 3964
rect 4019 3961 4031 3995
rect 3973 3955 4031 3961
rect 4478 3995 4536 4001
rect 4478 3961 4490 3995
rect 4524 3961 4536 3995
rect 4478 3955 4536 3961
rect 6273 3995 6331 4001
rect 6273 3961 6285 3995
rect 6319 3992 6331 3995
rect 6914 3992 6920 4004
rect 6319 3964 6920 3992
rect 6319 3961 6331 3964
rect 6273 3955 6331 3961
rect 3329 3927 3387 3933
rect 3329 3893 3341 3927
rect 3375 3924 3387 3927
rect 3786 3924 3792 3936
rect 3375 3896 3792 3924
rect 3375 3893 3387 3896
rect 3329 3887 3387 3893
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 4154 3884 4160 3936
rect 4212 3924 4218 3936
rect 4493 3924 4521 3955
rect 6914 3952 6920 3964
rect 6972 3952 6978 4004
rect 7330 3995 7388 4001
rect 7330 3961 7342 3995
rect 7376 3961 7388 3995
rect 7330 3955 7388 3961
rect 8941 3995 8999 4001
rect 8941 3961 8953 3995
rect 8987 3961 8999 3995
rect 10870 3992 10876 4004
rect 10831 3964 10876 3992
rect 8941 3955 8999 3961
rect 6549 3927 6607 3933
rect 6549 3924 6561 3927
rect 4212 3896 6561 3924
rect 4212 3884 4218 3896
rect 6549 3893 6561 3896
rect 6595 3924 6607 3927
rect 7190 3924 7196 3936
rect 6595 3896 7196 3924
rect 6595 3893 6607 3896
rect 6549 3887 6607 3893
rect 7190 3884 7196 3896
rect 7248 3924 7254 3936
rect 7345 3924 7373 3955
rect 7248 3896 7373 3924
rect 7929 3927 7987 3933
rect 7248 3884 7254 3896
rect 7929 3893 7941 3927
rect 7975 3924 7987 3927
rect 8202 3924 8208 3936
rect 7975 3896 8208 3924
rect 7975 3893 7987 3896
rect 7929 3887 7987 3893
rect 8202 3884 8208 3896
rect 8260 3924 8266 3936
rect 8573 3927 8631 3933
rect 8573 3924 8585 3927
rect 8260 3896 8585 3924
rect 8260 3884 8266 3896
rect 8573 3893 8585 3896
rect 8619 3924 8631 3927
rect 8956 3924 8984 3955
rect 10870 3952 10876 3964
rect 10928 3952 10934 4004
rect 10962 3952 10968 4004
rect 11020 3992 11026 4004
rect 12894 3992 12900 4004
rect 11020 3964 11065 3992
rect 12855 3964 12900 3992
rect 11020 3952 11026 3964
rect 12894 3952 12900 3964
rect 12952 3952 12958 4004
rect 8619 3896 8984 3924
rect 8619 3893 8631 3896
rect 8573 3887 8631 3893
rect 10134 3884 10140 3936
rect 10192 3924 10198 3936
rect 10229 3927 10287 3933
rect 10229 3924 10241 3927
rect 10192 3896 10241 3924
rect 10192 3884 10198 3896
rect 10229 3893 10241 3896
rect 10275 3893 10287 3927
rect 11790 3924 11796 3936
rect 11751 3896 11796 3924
rect 10229 3887 10287 3893
rect 11790 3884 11796 3896
rect 11848 3884 11854 3936
rect 13786 3924 13814 4100
rect 14369 4097 14381 4131
rect 14415 4128 14427 4131
rect 14642 4128 14648 4140
rect 14415 4100 14648 4128
rect 14415 4097 14427 4100
rect 14369 4091 14427 4097
rect 14642 4088 14648 4100
rect 14700 4088 14706 4140
rect 15013 4131 15071 4137
rect 15013 4097 15025 4131
rect 15059 4128 15071 4131
rect 16206 4128 16212 4140
rect 15059 4100 16212 4128
rect 15059 4097 15071 4100
rect 15013 4091 15071 4097
rect 16206 4088 16212 4100
rect 16264 4088 16270 4140
rect 17313 4131 17371 4137
rect 17313 4097 17325 4131
rect 17359 4128 17371 4131
rect 17402 4128 17408 4140
rect 17359 4100 17408 4128
rect 17359 4097 17371 4100
rect 17313 4091 17371 4097
rect 17402 4088 17408 4100
rect 17460 4088 17466 4140
rect 18417 4131 18475 4137
rect 18417 4097 18429 4131
rect 18463 4128 18475 4131
rect 18598 4128 18604 4140
rect 18463 4100 18604 4128
rect 18463 4097 18475 4100
rect 18417 4091 18475 4097
rect 18598 4088 18604 4100
rect 18656 4088 18662 4140
rect 18708 4128 18736 4168
rect 19334 4156 19340 4168
rect 19392 4156 19398 4208
rect 19426 4156 19432 4208
rect 19484 4196 19490 4208
rect 21591 4199 21649 4205
rect 21591 4196 21603 4199
rect 19484 4168 21603 4196
rect 19484 4156 19490 4168
rect 21591 4165 21603 4168
rect 21637 4165 21649 4199
rect 24210 4196 24216 4208
rect 24171 4168 24216 4196
rect 21591 4159 21649 4165
rect 24210 4156 24216 4168
rect 24268 4156 24274 4208
rect 24581 4199 24639 4205
rect 24581 4165 24593 4199
rect 24627 4196 24639 4199
rect 24670 4196 24676 4208
rect 24627 4168 24676 4196
rect 24627 4165 24639 4168
rect 24581 4159 24639 4165
rect 24670 4156 24676 4168
rect 24728 4156 24734 4208
rect 20070 4128 20076 4140
rect 18708 4100 19104 4128
rect 19983 4100 20076 4128
rect 14185 3995 14243 4001
rect 14185 3961 14197 3995
rect 14231 3992 14243 3995
rect 14461 3995 14519 4001
rect 14461 3992 14473 3995
rect 14231 3964 14473 3992
rect 14231 3961 14243 3964
rect 14185 3955 14243 3961
rect 14461 3961 14473 3964
rect 14507 3992 14519 3995
rect 15930 3992 15936 4004
rect 14507 3964 15792 3992
rect 15891 3964 15936 3992
rect 14507 3961 14519 3964
rect 14461 3955 14519 3961
rect 14366 3924 14372 3936
rect 13786 3896 14372 3924
rect 14366 3884 14372 3896
rect 14424 3884 14430 3936
rect 15764 3933 15792 3964
rect 15930 3952 15936 3964
rect 15988 3952 15994 4004
rect 16025 3995 16083 4001
rect 16025 3961 16037 3995
rect 16071 3992 16083 3995
rect 16298 3992 16304 4004
rect 16071 3964 16304 3992
rect 16071 3961 16083 3964
rect 16025 3955 16083 3961
rect 15749 3927 15807 3933
rect 15749 3893 15761 3927
rect 15795 3924 15807 3927
rect 16040 3924 16068 3955
rect 16298 3952 16304 3964
rect 16356 3952 16362 4004
rect 16574 3992 16580 4004
rect 16535 3964 16580 3992
rect 16574 3952 16580 3964
rect 16632 3952 16638 4004
rect 18230 3952 18236 4004
rect 18288 3992 18294 4004
rect 19076 4001 19104 4100
rect 20070 4088 20076 4100
rect 20128 4128 20134 4140
rect 20438 4128 20444 4140
rect 20128 4100 20444 4128
rect 20128 4088 20134 4100
rect 20438 4088 20444 4100
rect 20496 4088 20502 4140
rect 20625 4131 20683 4137
rect 20625 4097 20637 4131
rect 20671 4128 20683 4131
rect 21266 4128 21272 4140
rect 20671 4100 21272 4128
rect 20671 4097 20683 4100
rect 20625 4091 20683 4097
rect 21266 4088 21272 4100
rect 21324 4088 21330 4140
rect 22373 4131 22431 4137
rect 22373 4097 22385 4131
rect 22419 4128 22431 4131
rect 22830 4128 22836 4140
rect 22419 4100 22836 4128
rect 22419 4097 22431 4100
rect 22373 4091 22431 4097
rect 22830 4088 22836 4100
rect 22888 4088 22894 4140
rect 21520 4063 21578 4069
rect 21520 4029 21532 4063
rect 21566 4060 21578 4063
rect 21818 4060 21824 4072
rect 21566 4032 21824 4060
rect 21566 4029 21578 4032
rect 21520 4023 21578 4029
rect 21818 4020 21824 4032
rect 21876 4060 21882 4072
rect 21913 4063 21971 4069
rect 21913 4060 21925 4063
rect 21876 4032 21925 4060
rect 21876 4020 21882 4032
rect 21913 4029 21925 4032
rect 21959 4029 21971 4063
rect 21913 4023 21971 4029
rect 22002 4020 22008 4072
rect 22060 4060 22066 4072
rect 22500 4063 22558 4069
rect 22500 4060 22512 4063
rect 22060 4032 22512 4060
rect 22060 4020 22066 4032
rect 22500 4029 22512 4032
rect 22546 4060 22558 4063
rect 22925 4063 22983 4069
rect 22925 4060 22937 4063
rect 22546 4032 22937 4060
rect 22546 4029 22558 4032
rect 22500 4023 22558 4029
rect 22925 4029 22937 4032
rect 22971 4060 22983 4063
rect 23728 4063 23786 4069
rect 23728 4060 23740 4063
rect 22971 4032 23740 4060
rect 22971 4029 22983 4032
rect 22925 4023 22983 4029
rect 23728 4029 23740 4032
rect 23774 4060 23786 4063
rect 24228 4060 24256 4156
rect 23774 4032 24256 4060
rect 24708 4063 24766 4069
rect 23774 4029 23786 4032
rect 23728 4023 23786 4029
rect 24708 4029 24720 4063
rect 24754 4060 24766 4063
rect 25240 4060 25268 4224
rect 24754 4032 25268 4060
rect 24754 4029 24766 4032
rect 24708 4023 24766 4029
rect 18509 3995 18567 4001
rect 18509 3992 18521 3995
rect 18288 3964 18521 3992
rect 18288 3952 18294 3964
rect 18509 3961 18521 3964
rect 18555 3961 18567 3995
rect 18509 3955 18567 3961
rect 19061 3995 19119 4001
rect 19061 3961 19073 3995
rect 19107 3992 19119 3995
rect 19981 3995 20039 4001
rect 19981 3992 19993 3995
rect 19107 3964 19993 3992
rect 19107 3961 19119 3964
rect 19061 3955 19119 3961
rect 19981 3961 19993 3964
rect 20027 3961 20039 3995
rect 19981 3955 20039 3961
rect 15795 3896 16068 3924
rect 19996 3924 20024 3955
rect 20070 3952 20076 4004
rect 20128 3992 20134 4004
rect 20128 3964 20173 3992
rect 20128 3952 20134 3964
rect 20990 3952 20996 4004
rect 21048 3992 21054 4004
rect 21269 3995 21327 4001
rect 21269 3992 21281 3995
rect 21048 3964 21281 3992
rect 21048 3952 21054 3964
rect 21269 3961 21281 3964
rect 21315 3961 21327 3995
rect 21269 3955 21327 3961
rect 22094 3952 22100 4004
rect 22152 3992 22158 4004
rect 24723 3992 24751 4023
rect 22152 3964 24751 3992
rect 22152 3952 22158 3964
rect 20254 3924 20260 3936
rect 19996 3896 20260 3924
rect 15795 3893 15807 3896
rect 15749 3887 15807 3893
rect 20254 3884 20260 3896
rect 20312 3884 20318 3936
rect 22002 3884 22008 3936
rect 22060 3924 22066 3936
rect 22603 3927 22661 3933
rect 22603 3924 22615 3927
rect 22060 3896 22615 3924
rect 22060 3884 22066 3896
rect 22603 3893 22615 3896
rect 22649 3893 22661 3927
rect 22603 3887 22661 3893
rect 22738 3884 22744 3936
rect 22796 3924 22802 3936
rect 23799 3927 23857 3933
rect 23799 3924 23811 3927
rect 22796 3896 23811 3924
rect 22796 3884 22802 3896
rect 23799 3893 23811 3896
rect 23845 3893 23857 3927
rect 23799 3887 23857 3893
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 4246 3680 4252 3732
rect 4304 3720 4310 3732
rect 4341 3723 4399 3729
rect 4341 3720 4353 3723
rect 4304 3692 4353 3720
rect 4304 3680 4310 3692
rect 4341 3689 4353 3692
rect 4387 3689 4399 3723
rect 7190 3720 7196 3732
rect 7151 3692 7196 3720
rect 4341 3683 4399 3689
rect 7190 3680 7196 3692
rect 7248 3680 7254 3732
rect 10962 3680 10968 3732
rect 11020 3720 11026 3732
rect 12158 3720 12164 3732
rect 11020 3692 12164 3720
rect 11020 3680 11026 3692
rect 12158 3680 12164 3692
rect 12216 3680 12222 3732
rect 12805 3723 12863 3729
rect 12805 3689 12817 3723
rect 12851 3720 12863 3723
rect 12894 3720 12900 3732
rect 12851 3692 12900 3720
rect 12851 3689 12863 3692
rect 12805 3683 12863 3689
rect 12894 3680 12900 3692
rect 12952 3680 12958 3732
rect 14369 3723 14427 3729
rect 14369 3689 14381 3723
rect 14415 3720 14427 3723
rect 14642 3720 14648 3732
rect 14415 3692 14648 3720
rect 14415 3689 14427 3692
rect 14369 3683 14427 3689
rect 14642 3680 14648 3692
rect 14700 3680 14706 3732
rect 15746 3680 15752 3732
rect 15804 3720 15810 3732
rect 15841 3723 15899 3729
rect 15841 3720 15853 3723
rect 15804 3692 15853 3720
rect 15804 3680 15810 3692
rect 15841 3689 15853 3692
rect 15887 3689 15899 3723
rect 15841 3683 15899 3689
rect 15930 3680 15936 3732
rect 15988 3720 15994 3732
rect 16669 3723 16727 3729
rect 16669 3720 16681 3723
rect 15988 3692 16681 3720
rect 15988 3680 15994 3692
rect 16669 3689 16681 3692
rect 16715 3689 16727 3723
rect 16669 3683 16727 3689
rect 16758 3680 16764 3732
rect 16816 3720 16822 3732
rect 19475 3723 19533 3729
rect 19475 3720 19487 3723
rect 16816 3692 19487 3720
rect 16816 3680 16822 3692
rect 19475 3689 19487 3692
rect 19521 3689 19533 3723
rect 19475 3683 19533 3689
rect 19981 3723 20039 3729
rect 19981 3689 19993 3723
rect 20027 3720 20039 3723
rect 20070 3720 20076 3732
rect 20027 3692 20076 3720
rect 20027 3689 20039 3692
rect 19981 3683 20039 3689
rect 20070 3680 20076 3692
rect 20128 3680 20134 3732
rect 20254 3720 20260 3732
rect 20215 3692 20260 3720
rect 20254 3680 20260 3692
rect 20312 3680 20318 3732
rect 22922 3680 22928 3732
rect 22980 3720 22986 3732
rect 24075 3723 24133 3729
rect 24075 3720 24087 3723
rect 22980 3692 24087 3720
rect 22980 3680 22986 3692
rect 24075 3689 24087 3692
rect 24121 3689 24133 3723
rect 25130 3720 25136 3732
rect 25091 3692 25136 3720
rect 24075 3683 24133 3689
rect 25130 3680 25136 3692
rect 25188 3680 25194 3732
rect 4430 3652 4436 3664
rect 1964 3624 4436 3652
rect 1964 3596 1992 3624
rect 4430 3612 4436 3624
rect 4488 3612 4494 3664
rect 6917 3655 6975 3661
rect 6917 3621 6929 3655
rect 6963 3652 6975 3655
rect 7006 3652 7012 3664
rect 6963 3624 7012 3652
rect 6963 3621 6975 3624
rect 6917 3615 6975 3621
rect 7006 3612 7012 3624
rect 7064 3652 7070 3664
rect 7561 3655 7619 3661
rect 7561 3652 7573 3655
rect 7064 3624 7573 3652
rect 7064 3612 7070 3624
rect 7561 3621 7573 3624
rect 7607 3621 7619 3655
rect 7561 3615 7619 3621
rect 8113 3655 8171 3661
rect 8113 3621 8125 3655
rect 8159 3652 8171 3655
rect 8202 3652 8208 3664
rect 8159 3624 8208 3652
rect 8159 3621 8171 3624
rect 8113 3615 8171 3621
rect 8202 3612 8208 3624
rect 8260 3612 8266 3664
rect 8662 3652 8668 3664
rect 8623 3624 8668 3652
rect 8662 3612 8668 3624
rect 8720 3612 8726 3664
rect 11603 3655 11661 3661
rect 11603 3621 11615 3655
rect 11649 3652 11661 3655
rect 11790 3652 11796 3664
rect 11649 3624 11796 3652
rect 11649 3621 11661 3624
rect 11603 3615 11661 3621
rect 11790 3612 11796 3624
rect 11848 3612 11854 3664
rect 12176 3652 12204 3680
rect 13078 3652 13084 3664
rect 12176 3624 13084 3652
rect 13078 3612 13084 3624
rect 13136 3652 13142 3664
rect 13173 3655 13231 3661
rect 13173 3652 13185 3655
rect 13136 3624 13185 3652
rect 13136 3612 13142 3624
rect 13173 3621 13185 3624
rect 13219 3621 13231 3655
rect 13173 3615 13231 3621
rect 15470 3612 15476 3664
rect 15528 3652 15534 3664
rect 15528 3624 15700 3652
rect 15528 3612 15534 3624
rect 1946 3584 1952 3596
rect 1859 3556 1952 3584
rect 1946 3544 1952 3556
rect 2004 3544 2010 3596
rect 2961 3587 3019 3593
rect 2961 3553 2973 3587
rect 3007 3584 3019 3587
rect 3326 3584 3332 3596
rect 3007 3556 3332 3584
rect 3007 3553 3019 3556
rect 2961 3547 3019 3553
rect 3326 3544 3332 3556
rect 3384 3544 3390 3596
rect 3418 3544 3424 3596
rect 3476 3584 3482 3596
rect 4154 3584 4160 3596
rect 3476 3556 4160 3584
rect 3476 3544 3482 3556
rect 4154 3544 4160 3556
rect 4212 3584 4218 3596
rect 4212 3556 4305 3584
rect 4212 3544 4218 3556
rect 4338 3544 4344 3596
rect 4396 3584 4402 3596
rect 4525 3587 4583 3593
rect 4525 3584 4537 3587
rect 4396 3556 4537 3584
rect 4396 3544 4402 3556
rect 4525 3553 4537 3556
rect 4571 3553 4583 3587
rect 4525 3547 4583 3553
rect 6181 3587 6239 3593
rect 6181 3553 6193 3587
rect 6227 3553 6239 3587
rect 6181 3547 6239 3553
rect 6641 3587 6699 3593
rect 6641 3553 6653 3587
rect 6687 3584 6699 3587
rect 7466 3584 7472 3596
rect 6687 3556 7472 3584
rect 6687 3553 6699 3556
rect 6641 3547 6699 3553
rect 4172 3516 4200 3544
rect 6196 3516 6224 3547
rect 6546 3516 6552 3528
rect 4172 3488 6552 3516
rect 6546 3476 6552 3488
rect 6604 3476 6610 3528
rect 3145 3451 3203 3457
rect 3145 3417 3157 3451
rect 3191 3448 3203 3451
rect 4522 3448 4528 3460
rect 3191 3420 4528 3448
rect 3191 3417 3203 3420
rect 3145 3411 3203 3417
rect 4522 3408 4528 3420
rect 4580 3408 4586 3460
rect 5350 3408 5356 3460
rect 5408 3448 5414 3460
rect 6656 3448 6684 3547
rect 7466 3544 7472 3556
rect 7524 3544 7530 3596
rect 9677 3587 9735 3593
rect 9677 3553 9689 3587
rect 9723 3553 9735 3587
rect 10134 3584 10140 3596
rect 10047 3556 10140 3584
rect 9677 3547 9735 3553
rect 8018 3516 8024 3528
rect 7979 3488 8024 3516
rect 8018 3476 8024 3488
rect 8076 3476 8082 3528
rect 8386 3476 8392 3528
rect 8444 3516 8450 3528
rect 9692 3516 9720 3547
rect 10134 3544 10140 3556
rect 10192 3544 10198 3596
rect 10042 3516 10048 3528
rect 8444 3488 10048 3516
rect 8444 3476 8450 3488
rect 10042 3476 10048 3488
rect 10100 3476 10106 3528
rect 5408 3420 6684 3448
rect 5408 3408 5414 3420
rect 9490 3408 9496 3460
rect 9548 3448 9554 3460
rect 10152 3448 10180 3544
rect 10413 3519 10471 3525
rect 10413 3485 10425 3519
rect 10459 3516 10471 3519
rect 11241 3519 11299 3525
rect 11241 3516 11253 3519
rect 10459 3488 11253 3516
rect 10459 3485 10471 3488
rect 10413 3479 10471 3485
rect 11241 3485 11253 3488
rect 11287 3516 11299 3519
rect 11974 3516 11980 3528
rect 11287 3488 11980 3516
rect 11287 3485 11299 3488
rect 11241 3479 11299 3485
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 13081 3519 13139 3525
rect 13081 3485 13093 3519
rect 13127 3516 13139 3519
rect 13998 3516 14004 3528
rect 13127 3488 14004 3516
rect 13127 3485 13139 3488
rect 13081 3479 13139 3485
rect 13998 3476 14004 3488
rect 14056 3516 14062 3528
rect 15470 3516 15476 3528
rect 14056 3488 14780 3516
rect 15431 3488 15476 3516
rect 14056 3476 14062 3488
rect 9548 3420 10180 3448
rect 9548 3408 9554 3420
rect 11698 3408 11704 3460
rect 11756 3448 11762 3460
rect 13446 3448 13452 3460
rect 11756 3420 13452 3448
rect 11756 3408 11762 3420
rect 13446 3408 13452 3420
rect 13504 3448 13510 3460
rect 13633 3451 13691 3457
rect 13633 3448 13645 3451
rect 13504 3420 13645 3448
rect 13504 3408 13510 3420
rect 13633 3417 13645 3420
rect 13679 3448 13691 3451
rect 14645 3451 14703 3457
rect 14645 3448 14657 3451
rect 13679 3420 14657 3448
rect 13679 3417 13691 3420
rect 13633 3411 13691 3417
rect 14645 3417 14657 3420
rect 14691 3417 14703 3451
rect 14752 3448 14780 3488
rect 15470 3476 15476 3488
rect 15528 3476 15534 3528
rect 15672 3516 15700 3624
rect 17862 3612 17868 3664
rect 17920 3652 17926 3664
rect 17957 3655 18015 3661
rect 17957 3652 17969 3655
rect 17920 3624 17969 3652
rect 17920 3612 17926 3624
rect 17957 3621 17969 3624
rect 18003 3652 18015 3655
rect 18230 3652 18236 3664
rect 18003 3624 18236 3652
rect 18003 3621 18015 3624
rect 17957 3615 18015 3621
rect 18230 3612 18236 3624
rect 18288 3612 18294 3664
rect 18690 3612 18696 3664
rect 18748 3652 18754 3664
rect 21818 3652 21824 3664
rect 18748 3624 21824 3652
rect 18748 3612 18754 3624
rect 21818 3612 21824 3624
rect 21876 3612 21882 3664
rect 16206 3544 16212 3596
rect 16264 3584 16270 3596
rect 17681 3587 17739 3593
rect 17681 3584 17693 3587
rect 16264 3556 17693 3584
rect 16264 3544 16270 3556
rect 17681 3553 17693 3556
rect 17727 3553 17739 3587
rect 17681 3547 17739 3553
rect 19404 3587 19462 3593
rect 19404 3553 19416 3587
rect 19450 3584 19462 3587
rect 19610 3584 19616 3596
rect 19450 3556 19616 3584
rect 19450 3553 19462 3556
rect 19404 3547 19462 3553
rect 19610 3544 19616 3556
rect 19668 3584 19674 3596
rect 20346 3584 20352 3596
rect 19668 3556 20352 3584
rect 19668 3544 19674 3556
rect 20346 3544 20352 3556
rect 20404 3544 20410 3596
rect 20968 3587 21026 3593
rect 20968 3553 20980 3587
rect 21014 3584 21026 3587
rect 21174 3584 21180 3596
rect 21014 3556 21180 3584
rect 21014 3553 21026 3556
rect 20968 3547 21026 3553
rect 21174 3544 21180 3556
rect 21232 3544 21238 3596
rect 21980 3587 22038 3593
rect 21980 3553 21992 3587
rect 22026 3584 22038 3587
rect 22094 3584 22100 3596
rect 22026 3556 22100 3584
rect 22026 3553 22038 3556
rect 21980 3547 22038 3553
rect 22094 3544 22100 3556
rect 22152 3544 22158 3596
rect 22992 3587 23050 3593
rect 22992 3553 23004 3587
rect 23038 3584 23050 3587
rect 24004 3587 24062 3593
rect 24004 3584 24016 3587
rect 23038 3556 24016 3584
rect 23038 3553 23050 3556
rect 22992 3547 23050 3553
rect 24004 3553 24016 3556
rect 24050 3584 24062 3587
rect 24210 3584 24216 3596
rect 24050 3556 24216 3584
rect 24050 3553 24062 3556
rect 24004 3547 24062 3553
rect 24210 3544 24216 3556
rect 24268 3544 24274 3596
rect 24946 3584 24952 3596
rect 24907 3556 24952 3584
rect 24946 3544 24952 3556
rect 25004 3544 25010 3596
rect 17865 3519 17923 3525
rect 17865 3516 17877 3519
rect 15672 3488 17877 3516
rect 17865 3485 17877 3488
rect 17911 3516 17923 3519
rect 18230 3516 18236 3528
rect 17911 3488 18236 3516
rect 17911 3485 17923 3488
rect 17865 3479 17923 3485
rect 18230 3476 18236 3488
rect 18288 3476 18294 3528
rect 20806 3516 20812 3528
rect 18432 3488 20812 3516
rect 18432 3457 18460 3488
rect 20806 3476 20812 3488
rect 20864 3476 20870 3528
rect 17681 3451 17739 3457
rect 14752 3420 16620 3448
rect 14645 3411 14703 3417
rect 2133 3383 2191 3389
rect 2133 3349 2145 3383
rect 2179 3380 2191 3383
rect 3878 3380 3884 3392
rect 2179 3352 3884 3380
rect 2179 3349 2191 3352
rect 2133 3343 2191 3349
rect 3878 3340 3884 3352
rect 3936 3340 3942 3392
rect 5074 3380 5080 3392
rect 5035 3352 5080 3380
rect 5074 3340 5080 3352
rect 5132 3340 5138 3392
rect 5442 3340 5448 3392
rect 5500 3380 5506 3392
rect 10134 3380 10140 3392
rect 5500 3352 10140 3380
rect 5500 3340 5506 3352
rect 10134 3340 10140 3352
rect 10192 3340 10198 3392
rect 10686 3380 10692 3392
rect 10647 3352 10692 3380
rect 10686 3340 10692 3352
rect 10744 3340 10750 3392
rect 10962 3340 10968 3392
rect 11020 3380 11026 3392
rect 11057 3383 11115 3389
rect 11057 3380 11069 3383
rect 11020 3352 11069 3380
rect 11020 3340 11026 3352
rect 11057 3349 11069 3352
rect 11103 3349 11115 3383
rect 11057 3343 11115 3349
rect 16022 3340 16028 3392
rect 16080 3380 16086 3392
rect 16393 3383 16451 3389
rect 16393 3380 16405 3383
rect 16080 3352 16405 3380
rect 16080 3340 16086 3352
rect 16393 3349 16405 3352
rect 16439 3349 16451 3383
rect 16592 3380 16620 3420
rect 17681 3417 17693 3451
rect 17727 3448 17739 3451
rect 18417 3451 18475 3457
rect 18417 3448 18429 3451
rect 17727 3420 18429 3448
rect 17727 3417 17739 3420
rect 17681 3411 17739 3417
rect 18417 3417 18429 3420
rect 18463 3417 18475 3451
rect 22051 3451 22109 3457
rect 22051 3448 22063 3451
rect 18417 3411 18475 3417
rect 18524 3420 22063 3448
rect 18524 3380 18552 3420
rect 22051 3417 22063 3420
rect 22097 3417 22109 3451
rect 22051 3411 22109 3417
rect 22186 3408 22192 3460
rect 22244 3448 22250 3460
rect 23063 3451 23121 3457
rect 23063 3448 23075 3451
rect 22244 3420 23075 3448
rect 22244 3408 22250 3420
rect 23063 3417 23075 3420
rect 23109 3417 23121 3451
rect 23063 3411 23121 3417
rect 16592 3352 18552 3380
rect 16393 3343 16451 3349
rect 20346 3340 20352 3392
rect 20404 3380 20410 3392
rect 21039 3383 21097 3389
rect 21039 3380 21051 3383
rect 20404 3352 21051 3380
rect 20404 3340 20410 3352
rect 21039 3349 21051 3352
rect 21085 3349 21097 3383
rect 22462 3380 22468 3392
rect 22375 3352 22468 3380
rect 21039 3343 21097 3349
rect 22462 3340 22468 3352
rect 22520 3380 22526 3392
rect 22646 3380 22652 3392
rect 22520 3352 22652 3380
rect 22520 3340 22526 3352
rect 22646 3340 22652 3352
rect 22704 3340 22710 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1946 3176 1952 3188
rect 1907 3148 1952 3176
rect 1946 3136 1952 3148
rect 2004 3136 2010 3188
rect 3053 3179 3111 3185
rect 3053 3145 3065 3179
rect 3099 3176 3111 3179
rect 3326 3176 3332 3188
rect 3099 3148 3332 3176
rect 3099 3145 3111 3148
rect 3053 3139 3111 3145
rect 3326 3136 3332 3148
rect 3384 3136 3390 3188
rect 4154 3136 4160 3188
rect 4212 3176 4218 3188
rect 4479 3179 4537 3185
rect 4212 3148 4257 3176
rect 4212 3136 4218 3148
rect 4479 3145 4491 3179
rect 4525 3176 4537 3179
rect 4798 3176 4804 3188
rect 4525 3148 4804 3176
rect 4525 3145 4537 3148
rect 4479 3139 4537 3145
rect 4798 3136 4804 3148
rect 4856 3176 4862 3188
rect 5074 3176 5080 3188
rect 4856 3148 5080 3176
rect 4856 3136 4862 3148
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 6546 3176 6552 3188
rect 6507 3148 6552 3176
rect 6546 3136 6552 3148
rect 6604 3136 6610 3188
rect 7926 3176 7932 3188
rect 7887 3148 7932 3176
rect 7926 3136 7932 3148
rect 7984 3136 7990 3188
rect 8202 3176 8208 3188
rect 8163 3148 8208 3176
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 10042 3176 10048 3188
rect 10003 3148 10048 3176
rect 10042 3136 10048 3148
rect 10100 3136 10106 3188
rect 12158 3176 12164 3188
rect 12119 3148 12164 3176
rect 12158 3136 12164 3148
rect 12216 3136 12222 3188
rect 12710 3176 12716 3188
rect 12671 3148 12716 3176
rect 12710 3136 12716 3148
rect 12768 3136 12774 3188
rect 13998 3176 14004 3188
rect 13959 3148 14004 3176
rect 13998 3136 14004 3148
rect 14056 3136 14062 3188
rect 15105 3179 15163 3185
rect 15105 3145 15117 3179
rect 15151 3176 15163 3179
rect 15286 3176 15292 3188
rect 15151 3148 15292 3176
rect 15151 3145 15163 3148
rect 15105 3139 15163 3145
rect 3467 3111 3525 3117
rect 3467 3077 3479 3111
rect 3513 3108 3525 3111
rect 10962 3108 10968 3120
rect 3513 3080 10968 3108
rect 3513 3077 3525 3080
rect 3467 3071 3525 3077
rect 10962 3068 10968 3080
rect 11020 3068 11026 3120
rect 3881 3043 3939 3049
rect 3881 3040 3893 3043
rect 3411 3012 3893 3040
rect 3411 2981 3439 3012
rect 3881 3009 3893 3012
rect 3927 3040 3939 3043
rect 3970 3040 3976 3052
rect 3927 3012 3976 3040
rect 3927 3009 3939 3012
rect 3881 3003 3939 3009
rect 3970 3000 3976 3012
rect 4028 3000 4034 3052
rect 9769 3043 9827 3049
rect 4126 3012 5799 3040
rect 3396 2975 3454 2981
rect 3396 2941 3408 2975
rect 3442 2941 3454 2975
rect 3396 2935 3454 2941
rect 3510 2932 3516 2984
rect 3568 2972 3574 2984
rect 4126 2972 4154 3012
rect 3568 2944 4154 2972
rect 4408 2975 4466 2981
rect 3568 2932 3574 2944
rect 4408 2941 4420 2975
rect 4454 2972 4466 2975
rect 4454 2944 4936 2972
rect 4454 2941 4466 2944
rect 4408 2935 4466 2941
rect 2317 2907 2375 2913
rect 2317 2873 2329 2907
rect 2363 2904 2375 2907
rect 4706 2904 4712 2916
rect 2363 2876 4712 2904
rect 2363 2873 2375 2876
rect 2317 2867 2375 2873
rect 4706 2864 4712 2876
rect 4764 2864 4770 2916
rect 4908 2848 4936 2944
rect 5442 2932 5448 2984
rect 5500 2972 5506 2984
rect 5771 2981 5799 3012
rect 9769 3009 9781 3043
rect 9815 3040 9827 3043
rect 10597 3043 10655 3049
rect 10597 3040 10609 3043
rect 9815 3012 10609 3040
rect 9815 3009 9827 3012
rect 9769 3003 9827 3009
rect 10597 3009 10609 3012
rect 10643 3040 10655 3043
rect 10686 3040 10692 3052
rect 10643 3012 10692 3040
rect 10643 3009 10655 3012
rect 10597 3003 10655 3009
rect 10686 3000 10692 3012
rect 10744 3000 10750 3052
rect 12728 3040 12756 3136
rect 15120 3108 15148 3139
rect 15286 3136 15292 3148
rect 15344 3136 15350 3188
rect 15470 3136 15476 3188
rect 15528 3176 15534 3188
rect 16853 3179 16911 3185
rect 16853 3176 16865 3179
rect 15528 3148 16865 3176
rect 15528 3136 15534 3148
rect 16853 3145 16865 3148
rect 16899 3145 16911 3179
rect 17862 3176 17868 3188
rect 17823 3148 17868 3176
rect 16853 3139 16911 3145
rect 17862 3136 17868 3148
rect 17920 3136 17926 3188
rect 18230 3176 18236 3188
rect 18191 3148 18236 3176
rect 18230 3136 18236 3148
rect 18288 3136 18294 3188
rect 18877 3179 18935 3185
rect 18877 3145 18889 3179
rect 18923 3176 18935 3179
rect 20346 3176 20352 3188
rect 18923 3148 20352 3176
rect 18923 3145 18935 3148
rect 18877 3139 18935 3145
rect 17221 3111 17279 3117
rect 17221 3108 17233 3111
rect 14476 3080 15148 3108
rect 15948 3080 17233 3108
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12728 3012 13001 3040
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 13630 3040 13636 3052
rect 13591 3012 13636 3040
rect 12989 3003 13047 3009
rect 13630 3000 13636 3012
rect 13688 3000 13694 3052
rect 14476 2984 14504 3080
rect 14734 3000 14740 3052
rect 14792 3040 14798 3052
rect 15948 3049 15976 3080
rect 17221 3077 17233 3080
rect 17267 3077 17279 3111
rect 17221 3071 17279 3077
rect 15933 3043 15991 3049
rect 15933 3040 15945 3043
rect 14792 3012 15945 3040
rect 14792 3000 14798 3012
rect 15933 3009 15945 3012
rect 15979 3009 15991 3043
rect 16574 3040 16580 3052
rect 16535 3012 16580 3040
rect 15933 3003 15991 3009
rect 16574 3000 16580 3012
rect 16632 3000 16638 3052
rect 5537 2975 5595 2981
rect 5537 2972 5549 2975
rect 5500 2944 5549 2972
rect 5500 2932 5506 2944
rect 5537 2941 5549 2944
rect 5583 2941 5595 2975
rect 5537 2935 5595 2941
rect 5756 2975 5814 2981
rect 5756 2941 5768 2975
rect 5802 2972 5814 2975
rect 6181 2975 6239 2981
rect 6181 2972 6193 2975
rect 5802 2944 6193 2972
rect 5802 2941 5814 2944
rect 5756 2935 5814 2941
rect 6181 2941 6193 2944
rect 6227 2941 6239 2975
rect 6181 2935 6239 2941
rect 6546 2932 6552 2984
rect 6604 2972 6610 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6604 2944 6837 2972
rect 6604 2932 6610 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 7377 2975 7435 2981
rect 7377 2941 7389 2975
rect 7423 2972 7435 2975
rect 7926 2972 7932 2984
rect 7423 2944 7932 2972
rect 7423 2941 7435 2944
rect 7377 2935 7435 2941
rect 7926 2932 7932 2944
rect 7984 2972 7990 2984
rect 8849 2975 8907 2981
rect 8849 2972 8861 2975
rect 7984 2944 8861 2972
rect 7984 2932 7990 2944
rect 8849 2941 8861 2944
rect 8895 2972 8907 2975
rect 9033 2975 9091 2981
rect 9033 2972 9045 2975
rect 8895 2944 9045 2972
rect 8895 2941 8907 2944
rect 8849 2935 8907 2941
rect 9033 2941 9045 2944
rect 9079 2941 9091 2975
rect 9490 2972 9496 2984
rect 9451 2944 9496 2972
rect 9033 2935 9091 2941
rect 9490 2932 9496 2944
rect 9548 2932 9554 2984
rect 14458 2972 14464 2984
rect 14371 2944 14464 2972
rect 14458 2932 14464 2944
rect 14516 2932 14522 2984
rect 18984 2981 19012 3148
rect 20346 3136 20352 3148
rect 20404 3136 20410 3188
rect 20901 3179 20959 3185
rect 20901 3145 20913 3179
rect 20947 3176 20959 3179
rect 22005 3179 22063 3185
rect 22005 3176 22017 3179
rect 20947 3148 22017 3176
rect 20947 3145 20959 3148
rect 20901 3139 20959 3145
rect 22005 3145 22017 3148
rect 22051 3176 22063 3179
rect 22094 3176 22100 3188
rect 22051 3148 22100 3176
rect 22051 3145 22063 3148
rect 22005 3139 22063 3145
rect 22094 3136 22100 3148
rect 22152 3136 22158 3188
rect 23658 3136 23664 3188
rect 23716 3176 23722 3188
rect 23799 3179 23857 3185
rect 23799 3176 23811 3179
rect 23716 3148 23811 3176
rect 23716 3136 23722 3148
rect 23799 3145 23811 3148
rect 23845 3145 23857 3179
rect 23799 3139 23857 3145
rect 24946 3136 24952 3188
rect 25004 3176 25010 3188
rect 25133 3179 25191 3185
rect 25133 3176 25145 3179
rect 25004 3148 25145 3176
rect 25004 3136 25010 3148
rect 25133 3145 25145 3148
rect 25179 3145 25191 3179
rect 25133 3139 25191 3145
rect 19610 3108 19616 3120
rect 19571 3080 19616 3108
rect 19610 3068 19616 3080
rect 19668 3068 19674 3120
rect 20257 3111 20315 3117
rect 20257 3077 20269 3111
rect 20303 3108 20315 3111
rect 21910 3108 21916 3120
rect 20303 3080 21916 3108
rect 20303 3077 20315 3080
rect 20257 3071 20315 3077
rect 21910 3068 21916 3080
rect 21968 3068 21974 3120
rect 23017 3111 23075 3117
rect 23017 3077 23029 3111
rect 23063 3108 23075 3111
rect 24210 3108 24216 3120
rect 23063 3080 24216 3108
rect 23063 3077 23075 3080
rect 23017 3071 23075 3077
rect 24210 3068 24216 3080
rect 24268 3108 24274 3120
rect 27522 3108 27528 3120
rect 24268 3080 27528 3108
rect 24268 3068 24274 3080
rect 27522 3068 27528 3080
rect 27580 3068 27586 3120
rect 19426 3000 19432 3052
rect 19484 3040 19490 3052
rect 20901 3043 20959 3049
rect 20901 3040 20913 3043
rect 19484 3012 20913 3040
rect 19484 3000 19490 3012
rect 20901 3009 20913 3012
rect 20947 3009 20959 3043
rect 20901 3003 20959 3009
rect 21227 3012 23474 3040
rect 18969 2975 19027 2981
rect 18969 2941 18981 2975
rect 19015 2941 19027 2975
rect 18969 2935 19027 2941
rect 20073 2975 20131 2981
rect 20073 2941 20085 2975
rect 20119 2941 20131 2975
rect 20073 2935 20131 2941
rect 7190 2864 7196 2916
rect 7248 2904 7254 2916
rect 10505 2907 10563 2913
rect 10505 2904 10517 2907
rect 7248 2876 10517 2904
rect 7248 2864 7254 2876
rect 10505 2873 10517 2876
rect 10551 2904 10563 2907
rect 10959 2907 11017 2913
rect 10959 2904 10971 2907
rect 10551 2876 10971 2904
rect 10551 2873 10563 2876
rect 10505 2867 10563 2873
rect 10959 2873 10971 2876
rect 11005 2904 11017 2907
rect 11790 2904 11796 2916
rect 11005 2876 11796 2904
rect 11005 2873 11017 2876
rect 10959 2867 11017 2873
rect 11790 2864 11796 2876
rect 11848 2904 11854 2916
rect 13078 2904 13084 2916
rect 11848 2876 11928 2904
rect 13039 2876 13084 2904
rect 11848 2864 11854 2876
rect 4890 2836 4896 2848
rect 4851 2808 4896 2836
rect 4890 2796 4896 2808
rect 4948 2796 4954 2848
rect 5859 2839 5917 2845
rect 5859 2805 5871 2839
rect 5905 2836 5917 2839
rect 6454 2836 6460 2848
rect 5905 2808 6460 2836
rect 5905 2805 5917 2808
rect 5859 2799 5917 2805
rect 6454 2796 6460 2808
rect 6512 2796 6518 2848
rect 6914 2836 6920 2848
rect 6875 2808 6920 2836
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 11514 2836 11520 2848
rect 11475 2808 11520 2836
rect 11514 2796 11520 2808
rect 11572 2796 11578 2848
rect 11900 2845 11928 2876
rect 13078 2864 13084 2876
rect 13136 2864 13142 2916
rect 15473 2907 15531 2913
rect 15473 2904 15485 2907
rect 13786 2876 15485 2904
rect 11885 2839 11943 2845
rect 11885 2805 11897 2839
rect 11931 2836 11943 2839
rect 13786 2836 13814 2876
rect 15473 2873 15485 2876
rect 15519 2904 15531 2907
rect 15746 2904 15752 2916
rect 15519 2876 15752 2904
rect 15519 2873 15531 2876
rect 15473 2867 15531 2873
rect 15746 2864 15752 2876
rect 15804 2864 15810 2916
rect 16022 2864 16028 2916
rect 16080 2904 16086 2916
rect 16080 2876 16125 2904
rect 16080 2864 16086 2876
rect 16206 2864 16212 2916
rect 16264 2904 16270 2916
rect 20088 2904 20116 2935
rect 20990 2932 20996 2984
rect 21048 2972 21054 2984
rect 21227 2981 21255 3012
rect 21212 2975 21270 2981
rect 21212 2972 21224 2975
rect 21048 2944 21224 2972
rect 21048 2932 21054 2944
rect 21212 2941 21224 2944
rect 21258 2941 21270 2975
rect 21212 2935 21270 2941
rect 22256 2975 22314 2981
rect 22256 2941 22268 2975
rect 22302 2972 22314 2975
rect 22646 2972 22652 2984
rect 22302 2944 22652 2972
rect 22302 2941 22314 2944
rect 22256 2935 22314 2941
rect 22646 2932 22652 2944
rect 22704 2932 22710 2984
rect 23446 2972 23474 3012
rect 23934 3000 23940 3052
rect 23992 3040 23998 3052
rect 25501 3043 25559 3049
rect 25501 3040 25513 3043
rect 23992 3012 25513 3040
rect 23992 3000 23998 3012
rect 24723 2981 24751 3012
rect 25501 3009 25513 3012
rect 25547 3009 25559 3043
rect 25501 3003 25559 3009
rect 23728 2975 23786 2981
rect 23728 2972 23740 2975
rect 23446 2944 23740 2972
rect 23728 2941 23740 2944
rect 23774 2972 23786 2975
rect 24489 2975 24547 2981
rect 24489 2972 24501 2975
rect 23774 2944 24501 2972
rect 23774 2941 23786 2944
rect 23728 2935 23786 2941
rect 24489 2941 24501 2944
rect 24535 2941 24547 2975
rect 24489 2935 24547 2941
rect 24708 2975 24766 2981
rect 24708 2941 24720 2975
rect 24754 2941 24766 2975
rect 24708 2935 24766 2941
rect 20717 2907 20775 2913
rect 20717 2904 20729 2907
rect 16264 2876 18552 2904
rect 20088 2876 20729 2904
rect 16264 2864 16270 2876
rect 14642 2836 14648 2848
rect 11931 2808 13814 2836
rect 14603 2808 14648 2836
rect 11931 2805 11943 2808
rect 11885 2799 11943 2805
rect 14642 2796 14648 2808
rect 14700 2796 14706 2848
rect 18524 2836 18552 2876
rect 20717 2873 20729 2876
rect 20763 2904 20775 2907
rect 24811 2907 24869 2913
rect 24811 2904 24823 2907
rect 20763 2876 24823 2904
rect 20763 2873 20775 2876
rect 20717 2867 20775 2873
rect 24811 2873 24823 2876
rect 24857 2873 24869 2907
rect 24811 2867 24869 2873
rect 19153 2839 19211 2845
rect 19153 2836 19165 2839
rect 18524 2808 19165 2836
rect 19153 2805 19165 2808
rect 19199 2805 19211 2839
rect 20990 2836 20996 2848
rect 20951 2808 20996 2836
rect 19153 2799 19211 2805
rect 20990 2796 20996 2808
rect 21048 2796 21054 2848
rect 21082 2796 21088 2848
rect 21140 2836 21146 2848
rect 21315 2839 21373 2845
rect 21315 2836 21327 2839
rect 21140 2808 21327 2836
rect 21140 2796 21146 2808
rect 21315 2805 21327 2808
rect 21361 2805 21373 2839
rect 21315 2799 21373 2805
rect 22002 2796 22008 2848
rect 22060 2836 22066 2848
rect 22327 2839 22385 2845
rect 22327 2836 22339 2839
rect 22060 2808 22339 2836
rect 22060 2796 22066 2808
rect 22327 2805 22339 2808
rect 22373 2805 22385 2839
rect 22327 2799 22385 2805
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 2087 2635 2145 2641
rect 2087 2601 2099 2635
rect 2133 2632 2145 2635
rect 2774 2632 2780 2644
rect 2133 2604 2780 2632
rect 2133 2601 2145 2604
rect 2087 2595 2145 2601
rect 2774 2592 2780 2604
rect 2832 2592 2838 2644
rect 3513 2635 3571 2641
rect 3513 2601 3525 2635
rect 3559 2632 3571 2635
rect 3694 2632 3700 2644
rect 3559 2604 3700 2632
rect 3559 2601 3571 2604
rect 3513 2595 3571 2601
rect 2016 2499 2074 2505
rect 2016 2465 2028 2499
rect 2062 2496 2074 2499
rect 2498 2496 2504 2508
rect 2062 2468 2504 2496
rect 2062 2465 2074 2468
rect 2016 2459 2074 2465
rect 2498 2456 2504 2468
rect 2556 2456 2562 2508
rect 3012 2499 3070 2505
rect 3012 2465 3024 2499
rect 3058 2496 3070 2499
rect 3528 2496 3556 2595
rect 3694 2592 3700 2604
rect 3752 2592 3758 2644
rect 4338 2632 4344 2644
rect 4299 2604 4344 2632
rect 4338 2592 4344 2604
rect 4396 2592 4402 2644
rect 4939 2635 4997 2641
rect 4939 2601 4951 2635
rect 4985 2632 4997 2635
rect 6270 2632 6276 2644
rect 4985 2604 6276 2632
rect 4985 2601 4997 2604
rect 4939 2595 4997 2601
rect 6270 2592 6276 2604
rect 6328 2592 6334 2644
rect 6454 2592 6460 2644
rect 6512 2632 6518 2644
rect 7837 2635 7895 2641
rect 7837 2632 7849 2635
rect 6512 2604 7849 2632
rect 6512 2592 6518 2604
rect 7837 2601 7849 2604
rect 7883 2632 7895 2635
rect 8018 2632 8024 2644
rect 7883 2604 8024 2632
rect 7883 2601 7895 2604
rect 7837 2595 7895 2601
rect 8018 2592 8024 2604
rect 8076 2592 8082 2644
rect 9582 2592 9588 2644
rect 9640 2632 9646 2644
rect 9907 2635 9965 2641
rect 9907 2632 9919 2635
rect 9640 2604 9919 2632
rect 9640 2592 9646 2604
rect 9907 2601 9919 2604
rect 9953 2601 9965 2635
rect 11974 2632 11980 2644
rect 11935 2604 11980 2632
rect 9907 2595 9965 2601
rect 11974 2592 11980 2604
rect 12032 2592 12038 2644
rect 12989 2635 13047 2641
rect 12989 2601 13001 2635
rect 13035 2632 13047 2635
rect 13078 2632 13084 2644
rect 13035 2604 13084 2632
rect 13035 2601 13047 2604
rect 12989 2595 13047 2601
rect 13078 2592 13084 2604
rect 13136 2592 13142 2644
rect 18049 2635 18107 2641
rect 18049 2632 18061 2635
rect 13648 2604 18061 2632
rect 3878 2524 3884 2576
rect 3936 2564 3942 2576
rect 6178 2564 6184 2576
rect 3936 2536 6184 2564
rect 3936 2524 3942 2536
rect 6178 2524 6184 2536
rect 6236 2524 6242 2576
rect 6365 2567 6423 2573
rect 6365 2533 6377 2567
rect 6411 2564 6423 2567
rect 6546 2564 6552 2576
rect 6411 2536 6552 2564
rect 6411 2533 6423 2536
rect 6365 2527 6423 2533
rect 6546 2524 6552 2536
rect 6604 2524 6610 2576
rect 6733 2567 6791 2573
rect 6733 2533 6745 2567
rect 6779 2564 6791 2567
rect 9030 2564 9036 2576
rect 6779 2536 9036 2564
rect 6779 2533 6791 2536
rect 6733 2527 6791 2533
rect 3058 2468 3556 2496
rect 4868 2499 4926 2505
rect 3058 2465 3070 2468
rect 3012 2459 3070 2465
rect 4868 2465 4880 2499
rect 4914 2496 4926 2499
rect 5077 2499 5135 2505
rect 5077 2496 5089 2499
rect 4914 2468 5089 2496
rect 4914 2465 4926 2468
rect 4868 2459 4926 2465
rect 5077 2465 5089 2468
rect 5123 2465 5135 2499
rect 5077 2459 5135 2465
rect 5813 2499 5871 2505
rect 5813 2465 5825 2499
rect 5859 2496 5871 2499
rect 6748 2496 6776 2527
rect 9030 2524 9036 2536
rect 9088 2524 9094 2576
rect 10873 2567 10931 2573
rect 10873 2533 10885 2567
rect 10919 2564 10931 2567
rect 11149 2567 11207 2573
rect 11149 2564 11161 2567
rect 10919 2536 11161 2564
rect 10919 2533 10931 2536
rect 10873 2527 10931 2533
rect 11149 2533 11161 2536
rect 11195 2564 11207 2567
rect 11514 2564 11520 2576
rect 11195 2536 11520 2564
rect 11195 2533 11207 2536
rect 11149 2527 11207 2533
rect 11514 2524 11520 2536
rect 11572 2564 11578 2576
rect 13648 2573 13676 2604
rect 18049 2601 18061 2604
rect 18095 2632 18107 2635
rect 20993 2635 21051 2641
rect 18095 2604 18552 2632
rect 18095 2601 18107 2604
rect 18049 2595 18107 2601
rect 13265 2567 13323 2573
rect 13265 2564 13277 2567
rect 11572 2536 13277 2564
rect 11572 2524 11578 2536
rect 13265 2533 13277 2536
rect 13311 2564 13323 2567
rect 13633 2567 13691 2573
rect 13633 2564 13645 2567
rect 13311 2536 13645 2564
rect 13311 2533 13323 2536
rect 13265 2527 13323 2533
rect 13633 2533 13645 2536
rect 13679 2533 13691 2567
rect 13633 2527 13691 2533
rect 15933 2567 15991 2573
rect 15933 2533 15945 2567
rect 15979 2564 15991 2567
rect 16022 2564 16028 2576
rect 15979 2536 16028 2564
rect 15979 2533 15991 2536
rect 15933 2527 15991 2533
rect 16022 2524 16028 2536
rect 16080 2564 16086 2576
rect 18524 2573 18552 2604
rect 20993 2601 21005 2635
rect 21039 2632 21051 2635
rect 21174 2632 21180 2644
rect 21039 2604 21180 2632
rect 21039 2601 21051 2604
rect 20993 2595 21051 2601
rect 21174 2592 21180 2604
rect 21232 2592 21238 2644
rect 16393 2567 16451 2573
rect 16393 2564 16405 2567
rect 16080 2536 16405 2564
rect 16080 2524 16086 2536
rect 16393 2533 16405 2536
rect 16439 2564 16451 2567
rect 17221 2567 17279 2573
rect 17221 2564 17233 2567
rect 16439 2536 17233 2564
rect 16439 2533 16451 2536
rect 16393 2527 16451 2533
rect 17221 2533 17233 2536
rect 17267 2533 17279 2567
rect 17221 2527 17279 2533
rect 18509 2567 18567 2573
rect 18509 2533 18521 2567
rect 18555 2533 18567 2567
rect 18509 2527 18567 2533
rect 19429 2567 19487 2573
rect 19429 2533 19441 2567
rect 19475 2564 19487 2567
rect 21082 2564 21088 2576
rect 19475 2536 21088 2564
rect 19475 2533 19487 2536
rect 19429 2527 19487 2533
rect 5859 2468 6776 2496
rect 6917 2499 6975 2505
rect 5859 2465 5871 2468
rect 5813 2459 5871 2465
rect 6917 2465 6929 2499
rect 6963 2465 6975 2499
rect 6917 2459 6975 2465
rect 8021 2499 8079 2505
rect 8021 2465 8033 2499
rect 8067 2496 8079 2499
rect 8570 2496 8576 2508
rect 8067 2468 8576 2496
rect 8067 2465 8079 2468
rect 8021 2459 8079 2465
rect 3099 2431 3157 2437
rect 3099 2397 3111 2431
rect 3145 2428 3157 2431
rect 6932 2428 6960 2459
rect 8570 2456 8576 2468
rect 8628 2496 8634 2508
rect 9836 2499 9894 2505
rect 8628 2468 8708 2496
rect 8628 2456 8634 2468
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 3145 2400 7481 2428
rect 3145 2397 3157 2400
rect 3099 2391 3157 2397
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 5077 2363 5135 2369
rect 5077 2329 5089 2363
rect 5123 2360 5135 2363
rect 5353 2363 5411 2369
rect 5353 2360 5365 2363
rect 5123 2332 5365 2360
rect 5123 2329 5135 2332
rect 5077 2323 5135 2329
rect 5353 2329 5365 2332
rect 5399 2360 5411 2363
rect 6086 2360 6092 2372
rect 5399 2332 6092 2360
rect 5399 2329 5411 2332
rect 5353 2323 5411 2329
rect 6086 2320 6092 2332
rect 6144 2320 6150 2372
rect 8386 2360 8392 2372
rect 7024 2332 8392 2360
rect 2498 2292 2504 2304
rect 2459 2264 2504 2292
rect 2498 2252 2504 2264
rect 2556 2252 2562 2304
rect 4338 2252 4344 2304
rect 4396 2292 4402 2304
rect 5997 2295 6055 2301
rect 5997 2292 6009 2295
rect 4396 2264 6009 2292
rect 4396 2252 4402 2264
rect 5997 2261 6009 2264
rect 6043 2292 6055 2295
rect 7024 2292 7052 2332
rect 8386 2320 8392 2332
rect 8444 2320 8450 2372
rect 8680 2369 8708 2468
rect 9836 2465 9848 2499
rect 9882 2496 9894 2499
rect 10134 2496 10140 2508
rect 9882 2468 10140 2496
rect 9882 2465 9894 2468
rect 9836 2459 9894 2465
rect 10134 2456 10140 2468
rect 10192 2496 10198 2508
rect 10229 2499 10287 2505
rect 10229 2496 10241 2499
rect 10192 2468 10241 2496
rect 10192 2456 10198 2468
rect 10229 2465 10241 2468
rect 10275 2465 10287 2499
rect 10229 2459 10287 2465
rect 11698 2456 11704 2508
rect 11756 2496 11762 2508
rect 11756 2468 11801 2496
rect 11756 2456 11762 2468
rect 17126 2456 17132 2508
rect 17184 2496 17190 2508
rect 17589 2499 17647 2505
rect 17589 2496 17601 2499
rect 17184 2468 17601 2496
rect 17184 2456 17190 2468
rect 17589 2465 17601 2468
rect 17635 2465 17647 2499
rect 17589 2459 17647 2465
rect 11057 2431 11115 2437
rect 11057 2397 11069 2431
rect 11103 2428 11115 2431
rect 13541 2431 13599 2437
rect 11103 2400 12480 2428
rect 11103 2397 11115 2400
rect 11057 2391 11115 2397
rect 8665 2363 8723 2369
rect 8665 2329 8677 2363
rect 8711 2360 8723 2363
rect 9398 2360 9404 2372
rect 8711 2332 9404 2360
rect 8711 2329 8723 2332
rect 8665 2323 8723 2329
rect 9398 2320 9404 2332
rect 9456 2320 9462 2372
rect 12452 2304 12480 2400
rect 13541 2397 13553 2431
rect 13587 2428 13599 2431
rect 16301 2431 16359 2437
rect 13587 2400 14596 2428
rect 13587 2397 13599 2400
rect 13541 2391 13599 2397
rect 13630 2320 13636 2372
rect 13688 2360 13694 2372
rect 14093 2363 14151 2369
rect 14093 2360 14105 2363
rect 13688 2332 14105 2360
rect 13688 2320 13694 2332
rect 14093 2329 14105 2332
rect 14139 2329 14151 2363
rect 14093 2323 14151 2329
rect 6043 2264 7052 2292
rect 7101 2295 7159 2301
rect 6043 2261 6055 2264
rect 5997 2255 6055 2261
rect 7101 2261 7113 2295
rect 7147 2292 7159 2295
rect 7374 2292 7380 2304
rect 7147 2264 7380 2292
rect 7147 2261 7159 2264
rect 7101 2255 7159 2261
rect 7374 2252 7380 2264
rect 7432 2252 7438 2304
rect 8205 2295 8263 2301
rect 8205 2261 8217 2295
rect 8251 2292 8263 2295
rect 8478 2292 8484 2304
rect 8251 2264 8484 2292
rect 8251 2261 8263 2264
rect 8205 2255 8263 2261
rect 8478 2252 8484 2264
rect 8536 2252 8542 2304
rect 9030 2292 9036 2304
rect 8991 2264 9036 2292
rect 9030 2252 9036 2264
rect 9088 2292 9094 2304
rect 9490 2292 9496 2304
rect 9088 2264 9496 2292
rect 9088 2252 9094 2264
rect 9490 2252 9496 2264
rect 9548 2252 9554 2304
rect 12434 2292 12440 2304
rect 12395 2264 12440 2292
rect 12434 2252 12440 2264
rect 12492 2252 12498 2304
rect 14568 2301 14596 2400
rect 16301 2397 16313 2431
rect 16347 2428 16359 2431
rect 17144 2428 17172 2456
rect 16347 2400 17172 2428
rect 18417 2431 18475 2437
rect 16347 2397 16359 2400
rect 16301 2391 16359 2397
rect 18417 2397 18429 2431
rect 18463 2397 18475 2431
rect 18874 2428 18880 2440
rect 18835 2400 18880 2428
rect 18417 2391 18475 2397
rect 16114 2320 16120 2372
rect 16172 2360 16178 2372
rect 16853 2363 16911 2369
rect 16853 2360 16865 2363
rect 16172 2332 16865 2360
rect 16172 2320 16178 2332
rect 16853 2329 16865 2332
rect 16899 2329 16911 2363
rect 18432 2360 18460 2391
rect 18874 2388 18880 2400
rect 18932 2388 18938 2440
rect 19444 2360 19472 2527
rect 21082 2524 21088 2536
rect 21140 2524 21146 2576
rect 22646 2524 22652 2576
rect 22704 2564 22710 2576
rect 22704 2536 24624 2564
rect 22704 2524 22710 2536
rect 19518 2456 19524 2508
rect 19576 2496 19582 2508
rect 24596 2505 24624 2536
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 19576 2468 19901 2496
rect 19576 2456 19582 2468
rect 19889 2465 19901 2468
rect 19935 2496 19947 2499
rect 20441 2499 20499 2505
rect 20441 2496 20453 2499
rect 19935 2468 20453 2496
rect 19935 2465 19947 2468
rect 19889 2459 19947 2465
rect 20441 2465 20453 2468
rect 20487 2465 20499 2499
rect 20441 2459 20499 2465
rect 22097 2499 22155 2505
rect 22097 2465 22109 2499
rect 22143 2465 22155 2499
rect 22097 2459 22155 2465
rect 24581 2499 24639 2505
rect 24581 2465 24593 2499
rect 24627 2496 24639 2499
rect 25133 2499 25191 2505
rect 25133 2496 25145 2499
rect 24627 2468 25145 2496
rect 24627 2465 24639 2468
rect 24581 2459 24639 2465
rect 25133 2465 25145 2468
rect 25179 2465 25191 2499
rect 25133 2459 25191 2465
rect 19610 2388 19616 2440
rect 19668 2428 19674 2440
rect 22112 2428 22140 2459
rect 22649 2431 22707 2437
rect 22649 2428 22661 2431
rect 19668 2400 22661 2428
rect 19668 2388 19674 2400
rect 22649 2397 22661 2400
rect 22695 2397 22707 2431
rect 22649 2391 22707 2397
rect 18432 2332 19472 2360
rect 20073 2363 20131 2369
rect 16853 2323 16911 2329
rect 20073 2329 20085 2363
rect 20119 2360 20131 2363
rect 21266 2360 21272 2372
rect 20119 2332 21272 2360
rect 20119 2329 20131 2332
rect 20073 2323 20131 2329
rect 21266 2320 21272 2332
rect 21324 2320 21330 2372
rect 22281 2363 22339 2369
rect 22281 2329 22293 2363
rect 22327 2360 22339 2363
rect 23934 2360 23940 2372
rect 22327 2332 23940 2360
rect 22327 2329 22339 2332
rect 22281 2323 22339 2329
rect 23934 2320 23940 2332
rect 23992 2320 23998 2372
rect 24765 2363 24823 2369
rect 24765 2329 24777 2363
rect 24811 2360 24823 2363
rect 26418 2360 26424 2372
rect 24811 2332 26424 2360
rect 24811 2329 24823 2332
rect 24765 2323 24823 2329
rect 26418 2320 26424 2332
rect 26476 2320 26482 2372
rect 14553 2295 14611 2301
rect 14553 2261 14565 2295
rect 14599 2292 14611 2295
rect 22186 2292 22192 2304
rect 14599 2264 22192 2292
rect 14599 2261 14611 2264
rect 14553 2255 14611 2261
rect 22186 2252 22192 2264
rect 22244 2252 22250 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 10134 2048 10140 2100
rect 10192 2088 10198 2100
rect 16942 2088 16948 2100
rect 10192 2060 16948 2088
rect 10192 2048 10198 2060
rect 16942 2048 16948 2060
rect 17000 2088 17006 2100
rect 19610 2088 19616 2100
rect 17000 2060 19616 2088
rect 17000 2048 17006 2060
rect 19610 2048 19616 2060
rect 19668 2048 19674 2100
rect 4890 1980 4896 2032
rect 4948 2020 4954 2032
rect 14458 2020 14464 2032
rect 4948 1992 14464 2020
rect 4948 1980 4954 1992
rect 14458 1980 14464 1992
rect 14516 1980 14522 2032
rect 21726 76 21732 128
rect 21784 116 21790 128
rect 23198 116 23204 128
rect 21784 88 23204 116
rect 21784 76 21790 88
rect 23198 76 23204 88
rect 23256 76 23262 128
<< via1 >>
rect 20 27480 72 27532
rect 756 27480 808 27532
rect 2872 27480 2924 27532
rect 3700 27480 3752 27532
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 25136 24939 25188 24948
rect 25136 24905 25145 24939
rect 25145 24905 25179 24939
rect 25179 24905 25188 24939
rect 25136 24896 25188 24905
rect 25136 24692 25188 24744
rect 11428 24556 11480 24608
rect 21272 24556 21324 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 25780 24352 25832 24404
rect 13360 24216 13412 24268
rect 14096 24216 14148 24268
rect 24032 24216 24084 24268
rect 11704 24148 11756 24200
rect 14004 24148 14056 24200
rect 13084 24012 13136 24064
rect 14004 24012 14056 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 5356 23851 5408 23860
rect 5356 23817 5365 23851
rect 5365 23817 5399 23851
rect 5399 23817 5408 23851
rect 5356 23808 5408 23817
rect 6644 23808 6696 23860
rect 1860 23647 1912 23656
rect 1860 23613 1869 23647
rect 1869 23613 1903 23647
rect 1903 23613 1912 23647
rect 1860 23604 1912 23613
rect 5356 23604 5408 23656
rect 6184 23604 6236 23656
rect 9588 23808 9640 23860
rect 12624 23851 12676 23860
rect 12624 23817 12633 23851
rect 12633 23817 12667 23851
rect 12667 23817 12676 23851
rect 12624 23808 12676 23817
rect 13360 23851 13412 23860
rect 13360 23817 13369 23851
rect 13369 23817 13403 23851
rect 13403 23817 13412 23851
rect 13360 23808 13412 23817
rect 16948 23808 17000 23860
rect 24768 23851 24820 23860
rect 24768 23817 24777 23851
rect 24777 23817 24811 23851
rect 24811 23817 24820 23851
rect 24768 23808 24820 23817
rect 13544 23740 13596 23792
rect 12072 23672 12124 23724
rect 12992 23647 13044 23656
rect 12992 23613 13001 23647
rect 13001 23613 13035 23647
rect 13035 23613 13044 23647
rect 12992 23604 13044 23613
rect 13176 23604 13228 23656
rect 2780 23536 2832 23588
rect 13912 23604 13964 23656
rect 15660 23604 15712 23656
rect 16396 23604 16448 23656
rect 16488 23536 16540 23588
rect 7196 23468 7248 23520
rect 13452 23468 13504 23520
rect 14096 23511 14148 23520
rect 14096 23477 14105 23511
rect 14105 23477 14139 23511
rect 14139 23477 14148 23511
rect 18512 23536 18564 23588
rect 18236 23511 18288 23520
rect 14096 23468 14148 23477
rect 18236 23477 18245 23511
rect 18245 23477 18279 23511
rect 18279 23477 18288 23511
rect 18236 23468 18288 23477
rect 24032 23468 24084 23520
rect 25320 23468 25372 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 9588 23264 9640 23316
rect 13176 23264 13228 23316
rect 16488 23264 16540 23316
rect 18052 23264 18104 23316
rect 27252 23264 27304 23316
rect 1584 23128 1636 23180
rect 9680 23128 9732 23180
rect 11336 23128 11388 23180
rect 13912 23128 13964 23180
rect 15476 23128 15528 23180
rect 16764 23128 16816 23180
rect 24676 23128 24728 23180
rect 12164 23103 12216 23112
rect 12164 23069 12173 23103
rect 12173 23069 12207 23103
rect 12207 23069 12216 23103
rect 12164 23060 12216 23069
rect 12716 23060 12768 23112
rect 12808 22992 12860 23044
rect 2596 22924 2648 22976
rect 12900 22924 12952 22976
rect 13176 22924 13228 22976
rect 14740 22924 14792 22976
rect 16028 22924 16080 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 1584 22763 1636 22772
rect 1584 22729 1593 22763
rect 1593 22729 1627 22763
rect 1627 22729 1636 22763
rect 1584 22720 1636 22729
rect 8116 22720 8168 22772
rect 11060 22720 11112 22772
rect 13728 22720 13780 22772
rect 15476 22720 15528 22772
rect 18604 22720 18656 22772
rect 21364 22720 21416 22772
rect 24676 22763 24728 22772
rect 24676 22729 24685 22763
rect 24685 22729 24719 22763
rect 24719 22729 24728 22763
rect 24676 22720 24728 22729
rect 8024 22652 8076 22704
rect 9680 22652 9732 22704
rect 7472 22559 7524 22568
rect 7472 22525 7481 22559
rect 7481 22525 7515 22559
rect 7515 22525 7524 22559
rect 7472 22516 7524 22525
rect 7840 22448 7892 22500
rect 9220 22516 9272 22568
rect 11060 22584 11112 22636
rect 13360 22584 13412 22636
rect 20904 22652 20956 22704
rect 14464 22584 14516 22636
rect 15844 22584 15896 22636
rect 10784 22516 10836 22568
rect 12992 22516 13044 22568
rect 9312 22448 9364 22500
rect 13912 22516 13964 22568
rect 9496 22380 9548 22432
rect 11336 22423 11388 22432
rect 11336 22389 11345 22423
rect 11345 22389 11379 22423
rect 11379 22389 11388 22423
rect 11336 22380 11388 22389
rect 12440 22380 12492 22432
rect 13176 22380 13228 22432
rect 13360 22423 13412 22432
rect 13360 22389 13369 22423
rect 13369 22389 13403 22423
rect 13403 22389 13412 22423
rect 13360 22380 13412 22389
rect 13912 22380 13964 22432
rect 16120 22516 16172 22568
rect 14556 22448 14608 22500
rect 14832 22380 14884 22432
rect 16120 22423 16172 22432
rect 16120 22389 16129 22423
rect 16129 22389 16163 22423
rect 16163 22389 16172 22423
rect 16120 22380 16172 22389
rect 16764 22380 16816 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 7472 22176 7524 22228
rect 12992 22176 13044 22228
rect 14004 22219 14056 22228
rect 13084 22151 13136 22160
rect 13084 22117 13093 22151
rect 13093 22117 13127 22151
rect 13127 22117 13136 22151
rect 13084 22108 13136 22117
rect 14004 22185 14013 22219
rect 14013 22185 14047 22219
rect 14047 22185 14056 22219
rect 14004 22176 14056 22185
rect 14832 22176 14884 22228
rect 15292 22108 15344 22160
rect 7104 22040 7156 22092
rect 8576 22040 8628 22092
rect 10784 22083 10836 22092
rect 10784 22049 10793 22083
rect 10793 22049 10827 22083
rect 10827 22049 10836 22083
rect 10784 22040 10836 22049
rect 12532 22040 12584 22092
rect 15384 22083 15436 22092
rect 15384 22049 15393 22083
rect 15393 22049 15427 22083
rect 15427 22049 15436 22083
rect 15384 22040 15436 22049
rect 16488 22040 16540 22092
rect 17224 22040 17276 22092
rect 18604 22040 18656 22092
rect 21272 22040 21324 22092
rect 14832 21972 14884 22024
rect 17592 21972 17644 22024
rect 9680 21904 9732 21956
rect 10876 21947 10928 21956
rect 10876 21913 10885 21947
rect 10885 21913 10919 21947
rect 10919 21913 10928 21947
rect 10876 21904 10928 21913
rect 12256 21904 12308 21956
rect 17132 21904 17184 21956
rect 8208 21836 8260 21888
rect 8668 21879 8720 21888
rect 8668 21845 8677 21879
rect 8677 21845 8711 21879
rect 8711 21845 8720 21879
rect 8668 21836 8720 21845
rect 9036 21879 9088 21888
rect 9036 21845 9045 21879
rect 9045 21845 9079 21879
rect 9079 21845 9088 21879
rect 9036 21836 9088 21845
rect 9128 21836 9180 21888
rect 11980 21836 12032 21888
rect 12348 21836 12400 21888
rect 15476 21836 15528 21888
rect 16304 21836 16356 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 9036 21632 9088 21684
rect 13084 21632 13136 21684
rect 16488 21632 16540 21684
rect 8576 21564 8628 21616
rect 9680 21607 9732 21616
rect 9680 21573 9689 21607
rect 9689 21573 9723 21607
rect 9723 21573 9732 21607
rect 9680 21564 9732 21573
rect 10876 21564 10928 21616
rect 13636 21564 13688 21616
rect 14004 21564 14056 21616
rect 14096 21564 14148 21616
rect 20904 21675 20956 21684
rect 20904 21641 20913 21675
rect 20913 21641 20947 21675
rect 20947 21641 20956 21675
rect 20904 21632 20956 21641
rect 21272 21675 21324 21684
rect 21272 21641 21281 21675
rect 21281 21641 21315 21675
rect 21315 21641 21324 21675
rect 21272 21632 21324 21641
rect 22008 21632 22060 21684
rect 14648 21496 14700 21548
rect 15384 21496 15436 21548
rect 18328 21564 18380 21616
rect 2136 21428 2188 21480
rect 11060 21428 11112 21480
rect 11704 21428 11756 21480
rect 14832 21428 14884 21480
rect 16120 21428 16172 21480
rect 18420 21428 18472 21480
rect 8668 21360 8720 21412
rect 6920 21292 6972 21344
rect 7104 21335 7156 21344
rect 7104 21301 7113 21335
rect 7113 21301 7147 21335
rect 7147 21301 7156 21335
rect 7104 21292 7156 21301
rect 7932 21292 7984 21344
rect 8116 21335 8168 21344
rect 8116 21301 8125 21335
rect 8125 21301 8159 21335
rect 8159 21301 8168 21335
rect 8116 21292 8168 21301
rect 8484 21292 8536 21344
rect 10048 21292 10100 21344
rect 11060 21292 11112 21344
rect 11796 21292 11848 21344
rect 12532 21292 12584 21344
rect 12992 21292 13044 21344
rect 13084 21292 13136 21344
rect 14372 21360 14424 21412
rect 17960 21360 18012 21412
rect 18604 21539 18656 21548
rect 18604 21505 18613 21539
rect 18613 21505 18647 21539
rect 18647 21505 18656 21539
rect 18604 21496 18656 21505
rect 20904 21428 20956 21480
rect 22836 21360 22888 21412
rect 15568 21292 15620 21344
rect 17224 21292 17276 21344
rect 18052 21292 18104 21344
rect 18604 21292 18656 21344
rect 21548 21292 21600 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 13084 21088 13136 21140
rect 2412 20952 2464 21004
rect 4712 20952 4764 21004
rect 6092 21020 6144 21072
rect 7932 21020 7984 21072
rect 8300 21020 8352 21072
rect 9864 21063 9916 21072
rect 9864 21029 9873 21063
rect 9873 21029 9907 21063
rect 9907 21029 9916 21063
rect 9864 21020 9916 21029
rect 11704 21063 11756 21072
rect 11704 21029 11713 21063
rect 11713 21029 11747 21063
rect 11747 21029 11756 21063
rect 11704 21020 11756 21029
rect 12256 21063 12308 21072
rect 12256 21029 12265 21063
rect 12265 21029 12299 21063
rect 12299 21029 12308 21063
rect 12256 21020 12308 21029
rect 13176 21063 13228 21072
rect 13176 21029 13185 21063
rect 13185 21029 13219 21063
rect 13219 21029 13228 21063
rect 13176 21020 13228 21029
rect 15660 21088 15712 21140
rect 22652 21088 22704 21140
rect 14096 21020 14148 21072
rect 16396 21020 16448 21072
rect 5448 20884 5500 20936
rect 15384 20995 15436 21004
rect 15384 20961 15393 20995
rect 15393 20961 15427 20995
rect 15427 20961 15436 20995
rect 15384 20952 15436 20961
rect 15660 20952 15712 21004
rect 17316 20952 17368 21004
rect 18144 20952 18196 21004
rect 18696 20952 18748 21004
rect 21640 20952 21692 21004
rect 6828 20927 6880 20936
rect 6828 20893 6837 20927
rect 6837 20893 6871 20927
rect 6871 20893 6880 20927
rect 6828 20884 6880 20893
rect 8392 20927 8444 20936
rect 8392 20893 8401 20927
rect 8401 20893 8435 20927
rect 8435 20893 8444 20927
rect 8392 20884 8444 20893
rect 9772 20927 9824 20936
rect 9772 20893 9781 20927
rect 9781 20893 9815 20927
rect 9815 20893 9824 20927
rect 9772 20884 9824 20893
rect 10048 20927 10100 20936
rect 10048 20893 10057 20927
rect 10057 20893 10091 20927
rect 10091 20893 10100 20927
rect 10048 20884 10100 20893
rect 13452 20884 13504 20936
rect 15752 20884 15804 20936
rect 13728 20859 13780 20868
rect 13728 20825 13737 20859
rect 13737 20825 13771 20859
rect 13771 20825 13780 20859
rect 13728 20816 13780 20825
rect 1124 20748 1176 20800
rect 5080 20748 5132 20800
rect 11796 20748 11848 20800
rect 16396 20816 16448 20868
rect 19524 20884 19576 20936
rect 20352 20816 20404 20868
rect 20444 20816 20496 20868
rect 16488 20791 16540 20800
rect 16488 20757 16497 20791
rect 16497 20757 16531 20791
rect 16531 20757 16540 20791
rect 16488 20748 16540 20757
rect 16856 20748 16908 20800
rect 18236 20748 18288 20800
rect 20628 20748 20680 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1584 20587 1636 20596
rect 1584 20553 1593 20587
rect 1593 20553 1627 20587
rect 1627 20553 1636 20587
rect 1584 20544 1636 20553
rect 4712 20587 4764 20596
rect 1308 20340 1360 20392
rect 4712 20553 4721 20587
rect 4721 20553 4755 20587
rect 4755 20553 4764 20587
rect 4712 20544 4764 20553
rect 8300 20544 8352 20596
rect 9036 20544 9088 20596
rect 9864 20544 9916 20596
rect 12164 20544 12216 20596
rect 4160 20476 4212 20528
rect 5448 20476 5500 20528
rect 6828 20451 6880 20460
rect 6828 20417 6837 20451
rect 6837 20417 6871 20451
rect 6871 20417 6880 20451
rect 6828 20408 6880 20417
rect 8944 20451 8996 20460
rect 8944 20417 8953 20451
rect 8953 20417 8987 20451
rect 8987 20417 8996 20451
rect 8944 20408 8996 20417
rect 11060 20408 11112 20460
rect 11704 20408 11756 20460
rect 14372 20544 14424 20596
rect 15660 20587 15712 20596
rect 12992 20476 13044 20528
rect 14832 20476 14884 20528
rect 14740 20451 14792 20460
rect 14740 20417 14749 20451
rect 14749 20417 14783 20451
rect 14783 20417 14792 20451
rect 14740 20408 14792 20417
rect 15660 20553 15669 20587
rect 15669 20553 15703 20587
rect 15703 20553 15712 20587
rect 15660 20544 15712 20553
rect 16672 20544 16724 20596
rect 17316 20587 17368 20596
rect 17316 20553 17325 20587
rect 17325 20553 17359 20587
rect 17359 20553 17368 20587
rect 21640 20587 21692 20596
rect 17316 20544 17368 20553
rect 15384 20476 15436 20528
rect 18972 20476 19024 20528
rect 21640 20553 21649 20587
rect 21649 20553 21683 20587
rect 21683 20553 21692 20587
rect 21640 20544 21692 20553
rect 20352 20476 20404 20528
rect 20812 20476 20864 20528
rect 2412 20247 2464 20256
rect 2412 20213 2421 20247
rect 2421 20213 2455 20247
rect 2455 20213 2464 20247
rect 2412 20204 2464 20213
rect 2688 20204 2740 20256
rect 5448 20383 5500 20392
rect 5448 20349 5457 20383
rect 5457 20349 5491 20383
rect 5491 20349 5500 20383
rect 5448 20340 5500 20349
rect 5632 20315 5684 20324
rect 5632 20281 5641 20315
rect 5641 20281 5675 20315
rect 5675 20281 5684 20315
rect 5632 20272 5684 20281
rect 6644 20315 6696 20324
rect 6644 20281 6653 20315
rect 6653 20281 6687 20315
rect 6687 20281 6696 20315
rect 6644 20272 6696 20281
rect 7656 20272 7708 20324
rect 9036 20315 9088 20324
rect 9036 20281 9045 20315
rect 9045 20281 9079 20315
rect 9079 20281 9088 20315
rect 9036 20272 9088 20281
rect 9404 20272 9456 20324
rect 17868 20340 17920 20392
rect 18604 20383 18656 20392
rect 18604 20349 18613 20383
rect 18613 20349 18647 20383
rect 18647 20349 18656 20383
rect 18604 20340 18656 20349
rect 27620 20476 27672 20528
rect 24676 20408 24728 20460
rect 11152 20315 11204 20324
rect 11152 20281 11161 20315
rect 11161 20281 11195 20315
rect 11195 20281 11204 20315
rect 11152 20272 11204 20281
rect 12992 20272 13044 20324
rect 4896 20204 4948 20256
rect 6092 20204 6144 20256
rect 7748 20247 7800 20256
rect 7748 20213 7757 20247
rect 7757 20213 7791 20247
rect 7791 20213 7800 20247
rect 7748 20204 7800 20213
rect 9956 20247 10008 20256
rect 9956 20213 9965 20247
rect 9965 20213 9999 20247
rect 9999 20213 10008 20247
rect 9956 20204 10008 20213
rect 13728 20204 13780 20256
rect 14832 20315 14884 20324
rect 14832 20281 14841 20315
rect 14841 20281 14875 20315
rect 14875 20281 14884 20315
rect 16396 20315 16448 20324
rect 14832 20272 14884 20281
rect 16396 20281 16405 20315
rect 16405 20281 16439 20315
rect 16439 20281 16448 20315
rect 16396 20272 16448 20281
rect 16488 20315 16540 20324
rect 16488 20281 16497 20315
rect 16497 20281 16531 20315
rect 16531 20281 16540 20315
rect 17040 20315 17092 20324
rect 16488 20272 16540 20281
rect 17040 20281 17049 20315
rect 17049 20281 17083 20315
rect 17083 20281 17092 20315
rect 17040 20272 17092 20281
rect 18788 20315 18840 20324
rect 18788 20281 18797 20315
rect 18797 20281 18831 20315
rect 18831 20281 18840 20315
rect 18788 20272 18840 20281
rect 18144 20204 18196 20256
rect 18696 20204 18748 20256
rect 20168 20204 20220 20256
rect 22284 20383 22336 20392
rect 22284 20349 22293 20383
rect 22293 20349 22327 20383
rect 22327 20349 22336 20383
rect 22284 20340 22336 20349
rect 24216 20340 24268 20392
rect 25044 20340 25096 20392
rect 20536 20272 20588 20324
rect 20720 20204 20772 20256
rect 21088 20204 21140 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 5448 20000 5500 20052
rect 7288 20000 7340 20052
rect 7748 20000 7800 20052
rect 7932 20000 7984 20052
rect 8944 20043 8996 20052
rect 8944 20009 8953 20043
rect 8953 20009 8987 20043
rect 8987 20009 8996 20043
rect 8944 20000 8996 20009
rect 9772 20000 9824 20052
rect 11704 20000 11756 20052
rect 12992 20000 13044 20052
rect 13176 20000 13228 20052
rect 13636 20000 13688 20052
rect 14096 20043 14148 20052
rect 14096 20009 14105 20043
rect 14105 20009 14139 20043
rect 14139 20009 14148 20043
rect 14096 20000 14148 20009
rect 14740 20043 14792 20052
rect 14740 20009 14749 20043
rect 14749 20009 14783 20043
rect 14783 20009 14792 20043
rect 14740 20000 14792 20009
rect 16856 20000 16908 20052
rect 17868 20000 17920 20052
rect 5816 19932 5868 19984
rect 6644 19932 6696 19984
rect 6920 19932 6972 19984
rect 7472 19975 7524 19984
rect 7472 19941 7481 19975
rect 7481 19941 7515 19975
rect 7515 19941 7524 19975
rect 7472 19932 7524 19941
rect 7564 19975 7616 19984
rect 7564 19941 7573 19975
rect 7573 19941 7607 19975
rect 7607 19941 7616 19975
rect 7564 19932 7616 19941
rect 8484 19932 8536 19984
rect 8668 19932 8720 19984
rect 15936 19932 15988 19984
rect 1216 19864 1268 19916
rect 4068 19864 4120 19916
rect 5632 19907 5684 19916
rect 5632 19873 5641 19907
rect 5641 19873 5675 19907
rect 5675 19873 5684 19907
rect 5632 19864 5684 19873
rect 9588 19907 9640 19916
rect 9588 19873 9597 19907
rect 9597 19873 9631 19907
rect 9631 19873 9640 19907
rect 9588 19864 9640 19873
rect 11152 19864 11204 19916
rect 14740 19864 14792 19916
rect 5264 19796 5316 19848
rect 9404 19796 9456 19848
rect 12072 19796 12124 19848
rect 12532 19796 12584 19848
rect 13176 19839 13228 19848
rect 13176 19805 13185 19839
rect 13185 19805 13219 19839
rect 13219 19805 13228 19839
rect 13176 19796 13228 19805
rect 16948 19796 17000 19848
rect 7564 19728 7616 19780
rect 13360 19728 13412 19780
rect 16580 19728 16632 19780
rect 17040 19771 17092 19780
rect 17040 19737 17049 19771
rect 17049 19737 17083 19771
rect 17083 19737 17092 19771
rect 17040 19728 17092 19737
rect 18880 19864 18932 19916
rect 20260 19864 20312 19916
rect 19340 19839 19392 19848
rect 19340 19805 19349 19839
rect 19349 19805 19383 19839
rect 19383 19805 19392 19839
rect 19340 19796 19392 19805
rect 22560 19796 22612 19848
rect 23664 19839 23716 19848
rect 23664 19805 23673 19839
rect 23673 19805 23707 19839
rect 23707 19805 23716 19839
rect 23664 19796 23716 19805
rect 24124 19796 24176 19848
rect 19064 19728 19116 19780
rect 2964 19660 3016 19712
rect 3792 19660 3844 19712
rect 3884 19660 3936 19712
rect 9956 19660 10008 19712
rect 10508 19703 10560 19712
rect 10508 19669 10517 19703
rect 10517 19669 10551 19703
rect 10551 19669 10560 19703
rect 10508 19660 10560 19669
rect 12624 19703 12676 19712
rect 12624 19669 12633 19703
rect 12633 19669 12667 19703
rect 12667 19669 12676 19703
rect 12624 19660 12676 19669
rect 18604 19660 18656 19712
rect 19984 19660 20036 19712
rect 20352 19660 20404 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 1216 19456 1268 19508
rect 5540 19456 5592 19508
rect 7472 19456 7524 19508
rect 8300 19456 8352 19508
rect 8852 19456 8904 19508
rect 11152 19456 11204 19508
rect 7104 19388 7156 19440
rect 10048 19388 10100 19440
rect 11704 19388 11756 19440
rect 12164 19388 12216 19440
rect 12992 19456 13044 19508
rect 13636 19499 13688 19508
rect 13636 19465 13645 19499
rect 13645 19465 13679 19499
rect 13679 19465 13688 19499
rect 13636 19456 13688 19465
rect 15936 19499 15988 19508
rect 15936 19465 15945 19499
rect 15945 19465 15979 19499
rect 15979 19465 15988 19499
rect 15936 19456 15988 19465
rect 16488 19456 16540 19508
rect 16580 19456 16632 19508
rect 18604 19456 18656 19508
rect 19064 19499 19116 19508
rect 19064 19465 19073 19499
rect 19073 19465 19107 19499
rect 19107 19465 19116 19499
rect 19064 19456 19116 19465
rect 24032 19456 24084 19508
rect 17040 19388 17092 19440
rect 18512 19388 18564 19440
rect 5264 19363 5316 19372
rect 5264 19329 5273 19363
rect 5273 19329 5307 19363
rect 5307 19329 5316 19363
rect 5264 19320 5316 19329
rect 8392 19320 8444 19372
rect 9036 19320 9088 19372
rect 9404 19363 9456 19372
rect 9404 19329 9413 19363
rect 9413 19329 9447 19363
rect 9447 19329 9456 19363
rect 9404 19320 9456 19329
rect 13176 19320 13228 19372
rect 14648 19363 14700 19372
rect 14648 19329 14657 19363
rect 14657 19329 14691 19363
rect 14691 19329 14700 19363
rect 14648 19320 14700 19329
rect 16856 19320 16908 19372
rect 18420 19363 18472 19372
rect 18420 19329 18429 19363
rect 18429 19329 18463 19363
rect 18463 19329 18472 19363
rect 18420 19320 18472 19329
rect 18604 19320 18656 19372
rect 1860 19295 1912 19304
rect 1860 19261 1869 19295
rect 1869 19261 1903 19295
rect 1903 19261 1912 19295
rect 1860 19252 1912 19261
rect 4068 19184 4120 19236
rect 2320 19116 2372 19168
rect 2964 19159 3016 19168
rect 2964 19125 2973 19159
rect 2973 19125 3007 19159
rect 3007 19125 3016 19159
rect 2964 19116 3016 19125
rect 3424 19116 3476 19168
rect 4436 19116 4488 19168
rect 4712 19159 4764 19168
rect 4712 19125 4721 19159
rect 4721 19125 4755 19159
rect 4755 19125 4764 19159
rect 4712 19116 4764 19125
rect 6000 19252 6052 19304
rect 5356 19227 5408 19236
rect 5356 19193 5365 19227
rect 5365 19193 5399 19227
rect 5399 19193 5408 19227
rect 5356 19184 5408 19193
rect 6828 19184 6880 19236
rect 7288 19227 7340 19236
rect 7288 19193 7297 19227
rect 7297 19193 7331 19227
rect 7331 19193 7340 19227
rect 7288 19184 7340 19193
rect 8852 19227 8904 19236
rect 8852 19193 8861 19227
rect 8861 19193 8895 19227
rect 8895 19193 8904 19227
rect 8852 19184 8904 19193
rect 8392 19116 8444 19168
rect 9588 19116 9640 19168
rect 10140 19116 10192 19168
rect 10508 19252 10560 19304
rect 11520 19252 11572 19304
rect 12624 19252 12676 19304
rect 17868 19252 17920 19304
rect 11152 19184 11204 19236
rect 12992 19184 13044 19236
rect 14280 19227 14332 19236
rect 14280 19193 14289 19227
rect 14289 19193 14323 19227
rect 14323 19193 14332 19227
rect 14280 19184 14332 19193
rect 14372 19227 14424 19236
rect 14372 19193 14381 19227
rect 14381 19193 14415 19227
rect 14415 19193 14424 19227
rect 14372 19184 14424 19193
rect 16580 19227 16632 19236
rect 16580 19193 16589 19227
rect 16589 19193 16623 19227
rect 16623 19193 16632 19227
rect 16580 19184 16632 19193
rect 14096 19116 14148 19168
rect 14740 19116 14792 19168
rect 17316 19116 17368 19168
rect 17500 19116 17552 19168
rect 18972 19184 19024 19236
rect 19984 19252 20036 19304
rect 21732 19252 21784 19304
rect 19524 19116 19576 19168
rect 20260 19116 20312 19168
rect 21180 19116 21232 19168
rect 24952 19184 25004 19236
rect 22192 19116 22244 19168
rect 24860 19159 24912 19168
rect 24860 19125 24869 19159
rect 24869 19125 24903 19159
rect 24903 19125 24912 19159
rect 24860 19116 24912 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1584 18955 1636 18964
rect 1584 18921 1593 18955
rect 1593 18921 1627 18955
rect 1627 18921 1636 18955
rect 1584 18912 1636 18921
rect 6000 18912 6052 18964
rect 7564 18912 7616 18964
rect 6184 18844 6236 18896
rect 9128 18912 9180 18964
rect 12256 18912 12308 18964
rect 8484 18844 8536 18896
rect 9864 18887 9916 18896
rect 9864 18853 9873 18887
rect 9873 18853 9907 18887
rect 9907 18853 9916 18887
rect 9864 18844 9916 18853
rect 11888 18887 11940 18896
rect 11888 18853 11897 18887
rect 11897 18853 11931 18887
rect 11931 18853 11940 18887
rect 11888 18844 11940 18853
rect 13636 18844 13688 18896
rect 14096 18912 14148 18964
rect 14372 18955 14424 18964
rect 14372 18921 14381 18955
rect 14381 18921 14415 18955
rect 14415 18921 14424 18955
rect 14372 18912 14424 18921
rect 16580 18912 16632 18964
rect 16948 18955 17000 18964
rect 16948 18921 16957 18955
rect 16957 18921 16991 18955
rect 16991 18921 17000 18955
rect 16948 18912 17000 18921
rect 18880 18912 18932 18964
rect 19156 18955 19208 18964
rect 19156 18921 19165 18955
rect 19165 18921 19199 18955
rect 19199 18921 19208 18955
rect 19156 18912 19208 18921
rect 14280 18844 14332 18896
rect 15384 18844 15436 18896
rect 17408 18844 17460 18896
rect 1216 18776 1268 18828
rect 4528 18819 4580 18828
rect 4528 18785 4546 18819
rect 4546 18785 4580 18819
rect 4528 18776 4580 18785
rect 5356 18819 5408 18828
rect 5356 18785 5365 18819
rect 5365 18785 5399 18819
rect 5399 18785 5408 18819
rect 5356 18776 5408 18785
rect 3056 18708 3108 18760
rect 5448 18751 5500 18760
rect 5448 18717 5457 18751
rect 5457 18717 5491 18751
rect 5491 18717 5500 18751
rect 5448 18708 5500 18717
rect 9772 18751 9824 18760
rect 9772 18717 9781 18751
rect 9781 18717 9815 18751
rect 9815 18717 9824 18751
rect 9772 18708 9824 18717
rect 10048 18751 10100 18760
rect 10048 18717 10057 18751
rect 10057 18717 10091 18751
rect 10091 18717 10100 18751
rect 10048 18708 10100 18717
rect 11796 18751 11848 18760
rect 11796 18717 11805 18751
rect 11805 18717 11839 18751
rect 11839 18717 11848 18751
rect 11796 18708 11848 18717
rect 9220 18640 9272 18692
rect 12256 18640 12308 18692
rect 12900 18708 12952 18760
rect 13360 18751 13412 18760
rect 13360 18717 13369 18751
rect 13369 18717 13403 18751
rect 13403 18717 13412 18751
rect 13360 18708 13412 18717
rect 13728 18751 13780 18760
rect 13728 18717 13737 18751
rect 13737 18717 13771 18751
rect 13771 18717 13780 18751
rect 13728 18708 13780 18717
rect 16120 18708 16172 18760
rect 17592 18751 17644 18760
rect 17592 18717 17601 18751
rect 17601 18717 17635 18751
rect 17635 18717 17644 18751
rect 17592 18708 17644 18717
rect 17868 18751 17920 18760
rect 17868 18717 17877 18751
rect 17877 18717 17911 18751
rect 17911 18717 17920 18751
rect 17868 18708 17920 18717
rect 14464 18640 14516 18692
rect 16396 18640 16448 18692
rect 19432 18776 19484 18828
rect 22100 18844 22152 18896
rect 21640 18776 21692 18828
rect 22836 18819 22888 18828
rect 22836 18785 22845 18819
rect 22845 18785 22879 18819
rect 22879 18785 22888 18819
rect 22836 18776 22888 18785
rect 25044 18776 25096 18828
rect 25504 18776 25556 18828
rect 21824 18751 21876 18760
rect 21824 18717 21833 18751
rect 21833 18717 21867 18751
rect 21867 18717 21876 18751
rect 21824 18708 21876 18717
rect 20720 18640 20772 18692
rect 4344 18572 4396 18624
rect 4988 18615 5040 18624
rect 4988 18581 4997 18615
rect 4997 18581 5031 18615
rect 5031 18581 5040 18615
rect 4988 18572 5040 18581
rect 8576 18572 8628 18624
rect 9128 18615 9180 18624
rect 9128 18581 9137 18615
rect 9137 18581 9171 18615
rect 9171 18581 9180 18615
rect 9128 18572 9180 18581
rect 11152 18572 11204 18624
rect 12624 18572 12676 18624
rect 16212 18572 16264 18624
rect 20076 18615 20128 18624
rect 20076 18581 20085 18615
rect 20085 18581 20119 18615
rect 20119 18581 20128 18615
rect 20076 18572 20128 18581
rect 21272 18572 21324 18624
rect 22284 18572 22336 18624
rect 24676 18572 24728 18624
rect 25136 18572 25188 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 1584 18411 1636 18420
rect 1584 18377 1593 18411
rect 1593 18377 1627 18411
rect 1627 18377 1636 18411
rect 1584 18368 1636 18377
rect 2044 18411 2096 18420
rect 2044 18377 2053 18411
rect 2053 18377 2087 18411
rect 2087 18377 2096 18411
rect 2044 18368 2096 18377
rect 3056 18343 3108 18352
rect 3056 18309 3065 18343
rect 3065 18309 3099 18343
rect 3099 18309 3108 18343
rect 8024 18368 8076 18420
rect 8484 18368 8536 18420
rect 8852 18368 8904 18420
rect 4528 18343 4580 18352
rect 3056 18300 3108 18309
rect 4528 18309 4537 18343
rect 4537 18309 4571 18343
rect 4571 18309 4580 18343
rect 4528 18300 4580 18309
rect 6092 18300 6144 18352
rect 11888 18411 11940 18420
rect 9772 18343 9824 18352
rect 9772 18309 9781 18343
rect 9781 18309 9815 18343
rect 9815 18309 9824 18343
rect 9772 18300 9824 18309
rect 5448 18232 5500 18284
rect 6736 18232 6788 18284
rect 9864 18232 9916 18284
rect 2044 18164 2096 18216
rect 3240 18207 3292 18216
rect 1492 18028 1544 18080
rect 3240 18173 3249 18207
rect 3249 18173 3283 18207
rect 3283 18173 3292 18207
rect 3240 18164 3292 18173
rect 4160 18164 4212 18216
rect 4988 18207 5040 18216
rect 4988 18173 4997 18207
rect 4997 18173 5031 18207
rect 5031 18173 5040 18207
rect 4988 18164 5040 18173
rect 5264 18207 5316 18216
rect 5264 18173 5273 18207
rect 5273 18173 5307 18207
rect 5307 18173 5316 18207
rect 5264 18164 5316 18173
rect 7104 18164 7156 18216
rect 8944 18164 8996 18216
rect 11888 18377 11897 18411
rect 11897 18377 11931 18411
rect 11931 18377 11940 18411
rect 11888 18368 11940 18377
rect 13636 18411 13688 18420
rect 13636 18377 13645 18411
rect 13645 18377 13679 18411
rect 13679 18377 13688 18411
rect 13636 18368 13688 18377
rect 15936 18368 15988 18420
rect 17408 18368 17460 18420
rect 17592 18368 17644 18420
rect 18604 18411 18656 18420
rect 18604 18377 18613 18411
rect 18613 18377 18647 18411
rect 18647 18377 18656 18411
rect 18604 18368 18656 18377
rect 18880 18368 18932 18420
rect 21640 18368 21692 18420
rect 24768 18411 24820 18420
rect 24768 18377 24777 18411
rect 24777 18377 24811 18411
rect 24811 18377 24820 18411
rect 24768 18368 24820 18377
rect 18420 18300 18472 18352
rect 11520 18275 11572 18284
rect 11520 18241 11529 18275
rect 11529 18241 11563 18275
rect 11563 18241 11572 18275
rect 11520 18232 11572 18241
rect 13728 18232 13780 18284
rect 11152 18164 11204 18216
rect 11336 18164 11388 18216
rect 12624 18164 12676 18216
rect 7656 18096 7708 18148
rect 9220 18139 9272 18148
rect 9220 18105 9229 18139
rect 9229 18105 9263 18139
rect 9263 18105 9272 18139
rect 9220 18096 9272 18105
rect 6000 18028 6052 18080
rect 6184 18028 6236 18080
rect 8852 18028 8904 18080
rect 12256 18071 12308 18080
rect 12256 18037 12265 18071
rect 12265 18037 12299 18071
rect 12299 18037 12308 18071
rect 12256 18028 12308 18037
rect 13636 18028 13688 18080
rect 13820 18028 13872 18080
rect 14372 18232 14424 18284
rect 14648 18232 14700 18284
rect 17684 18232 17736 18284
rect 24952 18232 25004 18284
rect 16212 18164 16264 18216
rect 18604 18164 18656 18216
rect 20720 18164 20772 18216
rect 24676 18164 24728 18216
rect 14280 18139 14332 18148
rect 14280 18105 14289 18139
rect 14289 18105 14323 18139
rect 14323 18105 14332 18139
rect 14280 18096 14332 18105
rect 15384 18028 15436 18080
rect 17868 18096 17920 18148
rect 18604 18028 18656 18080
rect 19432 18028 19484 18080
rect 20076 18096 20128 18148
rect 20260 18028 20312 18080
rect 21272 18139 21324 18148
rect 21272 18105 21281 18139
rect 21281 18105 21315 18139
rect 21315 18105 21324 18139
rect 21272 18096 21324 18105
rect 21364 18028 21416 18080
rect 22100 18071 22152 18080
rect 22100 18037 22109 18071
rect 22109 18037 22143 18071
rect 22143 18037 22152 18071
rect 22100 18028 22152 18037
rect 22836 18071 22888 18080
rect 22836 18037 22845 18071
rect 22845 18037 22879 18071
rect 22879 18037 22888 18071
rect 22836 18028 22888 18037
rect 25044 18028 25096 18080
rect 25504 18071 25556 18080
rect 25504 18037 25513 18071
rect 25513 18037 25547 18071
rect 25547 18037 25556 18071
rect 25504 18028 25556 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 3884 17867 3936 17876
rect 3884 17833 3893 17867
rect 3893 17833 3927 17867
rect 3927 17833 3936 17867
rect 3884 17824 3936 17833
rect 5264 17867 5316 17876
rect 5264 17833 5273 17867
rect 5273 17833 5307 17867
rect 5307 17833 5316 17867
rect 5264 17824 5316 17833
rect 6184 17867 6236 17876
rect 6184 17833 6193 17867
rect 6193 17833 6227 17867
rect 6227 17833 6236 17867
rect 6184 17824 6236 17833
rect 6736 17867 6788 17876
rect 6736 17833 6745 17867
rect 6745 17833 6779 17867
rect 6779 17833 6788 17867
rect 6736 17824 6788 17833
rect 7104 17824 7156 17876
rect 8852 17824 8904 17876
rect 9220 17867 9272 17876
rect 9220 17833 9229 17867
rect 9229 17833 9263 17867
rect 9263 17833 9272 17867
rect 9220 17824 9272 17833
rect 9772 17824 9824 17876
rect 11796 17867 11848 17876
rect 11796 17833 11805 17867
rect 11805 17833 11839 17867
rect 11839 17833 11848 17867
rect 11796 17824 11848 17833
rect 13360 17867 13412 17876
rect 13360 17833 13369 17867
rect 13369 17833 13403 17867
rect 13403 17833 13412 17867
rect 13360 17824 13412 17833
rect 13636 17824 13688 17876
rect 14188 17824 14240 17876
rect 14280 17824 14332 17876
rect 17316 17824 17368 17876
rect 17592 17824 17644 17876
rect 3516 17799 3568 17808
rect 3516 17765 3525 17799
rect 3525 17765 3559 17799
rect 3559 17765 3568 17799
rect 3516 17756 3568 17765
rect 4160 17756 4212 17808
rect 3608 17688 3660 17740
rect 4528 17731 4580 17740
rect 4528 17697 4537 17731
rect 4537 17697 4571 17731
rect 4571 17697 4580 17731
rect 4528 17688 4580 17697
rect 8300 17756 8352 17808
rect 11336 17799 11388 17808
rect 11336 17765 11345 17799
rect 11345 17765 11379 17799
rect 11379 17765 11388 17799
rect 11336 17756 11388 17765
rect 11888 17756 11940 17808
rect 12256 17756 12308 17808
rect 17408 17756 17460 17808
rect 7564 17731 7616 17740
rect 7564 17697 7573 17731
rect 7573 17697 7607 17731
rect 7607 17697 7616 17731
rect 7564 17688 7616 17697
rect 8576 17688 8628 17740
rect 10600 17731 10652 17740
rect 10600 17697 10609 17731
rect 10609 17697 10643 17731
rect 10643 17697 10652 17731
rect 10600 17688 10652 17697
rect 11152 17731 11204 17740
rect 11152 17697 11161 17731
rect 11161 17697 11195 17731
rect 11195 17697 11204 17731
rect 11152 17688 11204 17697
rect 14740 17688 14792 17740
rect 15660 17731 15712 17740
rect 15660 17697 15669 17731
rect 15669 17697 15703 17731
rect 15703 17697 15712 17731
rect 15660 17688 15712 17697
rect 19156 17824 19208 17876
rect 20076 17824 20128 17876
rect 20260 17867 20312 17876
rect 20260 17833 20269 17867
rect 20269 17833 20303 17867
rect 20303 17833 20312 17867
rect 20260 17824 20312 17833
rect 20996 17867 21048 17876
rect 20996 17833 21005 17867
rect 21005 17833 21039 17867
rect 21039 17833 21048 17867
rect 20996 17824 21048 17833
rect 21364 17824 21416 17876
rect 19156 17688 19208 17740
rect 20260 17688 20312 17740
rect 20720 17688 20772 17740
rect 21640 17688 21692 17740
rect 23020 17731 23072 17740
rect 23020 17697 23029 17731
rect 23029 17697 23063 17731
rect 23063 17697 23072 17731
rect 23020 17688 23072 17697
rect 23848 17688 23900 17740
rect 24676 17688 24728 17740
rect 2780 17620 2832 17672
rect 6000 17620 6052 17672
rect 12164 17663 12216 17672
rect 12164 17629 12173 17663
rect 12173 17629 12207 17663
rect 12207 17629 12216 17663
rect 12164 17620 12216 17629
rect 16764 17663 16816 17672
rect 16764 17629 16773 17663
rect 16773 17629 16807 17663
rect 16807 17629 16816 17663
rect 16764 17620 16816 17629
rect 17040 17620 17092 17672
rect 17868 17620 17920 17672
rect 18880 17620 18932 17672
rect 20812 17620 20864 17672
rect 23480 17663 23532 17672
rect 23480 17629 23489 17663
rect 23489 17629 23523 17663
rect 23523 17629 23532 17663
rect 23480 17620 23532 17629
rect 10968 17552 11020 17604
rect 15292 17552 15344 17604
rect 16580 17595 16632 17604
rect 16580 17561 16589 17595
rect 16589 17561 16623 17595
rect 16623 17561 16632 17595
rect 16580 17552 16632 17561
rect 17500 17552 17552 17604
rect 1216 17484 1268 17536
rect 3148 17527 3200 17536
rect 3148 17493 3157 17527
rect 3157 17493 3191 17527
rect 3191 17493 3200 17527
rect 3148 17484 3200 17493
rect 4160 17484 4212 17536
rect 8392 17484 8444 17536
rect 8852 17527 8904 17536
rect 8852 17493 8861 17527
rect 8861 17493 8895 17527
rect 8895 17493 8904 17527
rect 8852 17484 8904 17493
rect 13084 17527 13136 17536
rect 13084 17493 13093 17527
rect 13093 17493 13127 17527
rect 13127 17493 13136 17527
rect 13084 17484 13136 17493
rect 14280 17484 14332 17536
rect 16120 17484 16172 17536
rect 16948 17484 17000 17536
rect 17684 17484 17736 17536
rect 22744 17484 22796 17536
rect 27620 17484 27672 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 1584 17323 1636 17332
rect 1584 17289 1593 17323
rect 1593 17289 1627 17323
rect 1627 17289 1636 17323
rect 1584 17280 1636 17289
rect 2136 17280 2188 17332
rect 3516 17280 3568 17332
rect 8944 17280 8996 17332
rect 10600 17323 10652 17332
rect 10600 17289 10609 17323
rect 10609 17289 10643 17323
rect 10643 17289 10652 17323
rect 10600 17280 10652 17289
rect 3148 17076 3200 17128
rect 4988 17212 5040 17264
rect 5540 17212 5592 17264
rect 3976 17076 4028 17128
rect 6000 17144 6052 17196
rect 9772 17144 9824 17196
rect 12164 17280 12216 17332
rect 13084 17280 13136 17332
rect 13728 17280 13780 17332
rect 17408 17323 17460 17332
rect 17408 17289 17417 17323
rect 17417 17289 17451 17323
rect 17451 17289 17460 17323
rect 17408 17280 17460 17289
rect 17500 17280 17552 17332
rect 18512 17280 18564 17332
rect 12440 17212 12492 17264
rect 13636 17187 13688 17196
rect 13636 17153 13645 17187
rect 13645 17153 13679 17187
rect 13679 17153 13688 17187
rect 13636 17144 13688 17153
rect 14372 17212 14424 17264
rect 16764 17212 16816 17264
rect 17040 17255 17092 17264
rect 17040 17221 17049 17255
rect 17049 17221 17083 17255
rect 17083 17221 17092 17255
rect 17040 17212 17092 17221
rect 5264 17076 5316 17128
rect 7288 17076 7340 17128
rect 7472 17119 7524 17128
rect 7472 17085 7481 17119
rect 7481 17085 7515 17119
rect 7515 17085 7524 17119
rect 7472 17076 7524 17085
rect 7656 17119 7708 17128
rect 7656 17085 7665 17119
rect 7665 17085 7699 17119
rect 7699 17085 7708 17119
rect 7656 17076 7708 17085
rect 10784 17119 10836 17128
rect 10784 17085 10793 17119
rect 10793 17085 10827 17119
rect 10827 17085 10836 17119
rect 10784 17076 10836 17085
rect 11152 17076 11204 17128
rect 6460 17008 6512 17060
rect 7932 17051 7984 17060
rect 7932 17017 7941 17051
rect 7941 17017 7975 17051
rect 7975 17017 7984 17051
rect 7932 17008 7984 17017
rect 8852 17051 8904 17060
rect 8852 17017 8861 17051
rect 8861 17017 8895 17051
rect 8895 17017 8904 17051
rect 8852 17008 8904 17017
rect 8944 17051 8996 17060
rect 8944 17017 8953 17051
rect 8953 17017 8987 17051
rect 8987 17017 8996 17051
rect 8944 17008 8996 17017
rect 3240 16983 3292 16992
rect 3240 16949 3249 16983
rect 3249 16949 3283 16983
rect 3283 16949 3292 16983
rect 3240 16940 3292 16949
rect 3608 16983 3660 16992
rect 3608 16949 3617 16983
rect 3617 16949 3651 16983
rect 3651 16949 3660 16983
rect 3608 16940 3660 16949
rect 3976 16940 4028 16992
rect 4528 16940 4580 16992
rect 5172 16940 5224 16992
rect 6092 16983 6144 16992
rect 6092 16949 6101 16983
rect 6101 16949 6135 16983
rect 6135 16949 6144 16983
rect 6092 16940 6144 16949
rect 8300 16983 8352 16992
rect 8300 16949 8309 16983
rect 8309 16949 8343 16983
rect 8343 16949 8352 16983
rect 8300 16940 8352 16949
rect 9956 16983 10008 16992
rect 9956 16949 9965 16983
rect 9965 16949 9999 16983
rect 9999 16949 10008 16983
rect 9956 16940 10008 16949
rect 11888 16940 11940 16992
rect 18880 17280 18932 17332
rect 21272 17280 21324 17332
rect 23020 17323 23072 17332
rect 23020 17289 23029 17323
rect 23029 17289 23063 17323
rect 23063 17289 23072 17323
rect 23020 17280 23072 17289
rect 25412 17323 25464 17332
rect 25412 17289 25421 17323
rect 25421 17289 25455 17323
rect 25455 17289 25464 17323
rect 25412 17280 25464 17289
rect 21640 17212 21692 17264
rect 24676 17255 24728 17264
rect 24676 17221 24685 17255
rect 24685 17221 24719 17255
rect 24719 17221 24728 17255
rect 24676 17212 24728 17221
rect 19432 17144 19484 17196
rect 20260 17144 20312 17196
rect 20720 17144 20772 17196
rect 21088 17144 21140 17196
rect 21272 17144 21324 17196
rect 21548 17144 21600 17196
rect 22744 17076 22796 17128
rect 22928 17076 22980 17128
rect 25228 17119 25280 17128
rect 25228 17085 25237 17119
rect 25237 17085 25271 17119
rect 25271 17085 25280 17119
rect 25228 17076 25280 17085
rect 13728 17051 13780 17060
rect 13728 17017 13737 17051
rect 13737 17017 13771 17051
rect 13771 17017 13780 17051
rect 13728 17008 13780 17017
rect 13084 16940 13136 16992
rect 15660 17008 15712 17060
rect 16580 17051 16632 17060
rect 16580 17017 16589 17051
rect 16589 17017 16623 17051
rect 16623 17017 16632 17051
rect 16580 17008 16632 17017
rect 14740 16940 14792 16992
rect 18880 16983 18932 16992
rect 18880 16949 18889 16983
rect 18889 16949 18923 16983
rect 18923 16949 18932 16983
rect 18880 16940 18932 16949
rect 19156 16940 19208 16992
rect 20812 16940 20864 16992
rect 21640 17008 21692 17060
rect 23848 17008 23900 17060
rect 23572 16940 23624 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1584 16779 1636 16788
rect 1584 16745 1593 16779
rect 1593 16745 1627 16779
rect 1627 16745 1636 16779
rect 1584 16736 1636 16745
rect 2320 16779 2372 16788
rect 2320 16745 2329 16779
rect 2329 16745 2363 16779
rect 2363 16745 2372 16779
rect 2320 16736 2372 16745
rect 3516 16736 3568 16788
rect 5264 16779 5316 16788
rect 5264 16745 5273 16779
rect 5273 16745 5307 16779
rect 5307 16745 5316 16779
rect 5264 16736 5316 16745
rect 7564 16779 7616 16788
rect 7564 16745 7573 16779
rect 7573 16745 7607 16779
rect 7607 16745 7616 16779
rect 7564 16736 7616 16745
rect 10784 16779 10836 16788
rect 10784 16745 10793 16779
rect 10793 16745 10827 16779
rect 10827 16745 10836 16779
rect 10784 16736 10836 16745
rect 11888 16779 11940 16788
rect 11888 16745 11897 16779
rect 11897 16745 11931 16779
rect 11931 16745 11940 16779
rect 11888 16736 11940 16745
rect 13728 16736 13780 16788
rect 15292 16736 15344 16788
rect 17408 16736 17460 16788
rect 17776 16736 17828 16788
rect 20720 16779 20772 16788
rect 2596 16668 2648 16720
rect 6184 16668 6236 16720
rect 7656 16668 7708 16720
rect 9864 16711 9916 16720
rect 9864 16677 9873 16711
rect 9873 16677 9907 16711
rect 9907 16677 9916 16711
rect 9864 16668 9916 16677
rect 11980 16668 12032 16720
rect 12532 16668 12584 16720
rect 13360 16711 13412 16720
rect 13360 16677 13369 16711
rect 13369 16677 13403 16711
rect 13403 16677 13412 16711
rect 13360 16668 13412 16677
rect 13636 16711 13688 16720
rect 13636 16677 13645 16711
rect 13645 16677 13679 16711
rect 13679 16677 13688 16711
rect 13636 16668 13688 16677
rect 15384 16668 15436 16720
rect 16764 16668 16816 16720
rect 20720 16745 20729 16779
rect 20729 16745 20763 16779
rect 20763 16745 20772 16779
rect 20720 16736 20772 16745
rect 19248 16668 19300 16720
rect 22836 16736 22888 16788
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 4804 16600 4856 16652
rect 7840 16600 7892 16652
rect 8484 16643 8536 16652
rect 8484 16609 8493 16643
rect 8493 16609 8527 16643
rect 8527 16609 8536 16643
rect 8484 16600 8536 16609
rect 3700 16532 3752 16584
rect 3884 16532 3936 16584
rect 7380 16532 7432 16584
rect 8760 16575 8812 16584
rect 8760 16541 8769 16575
rect 8769 16541 8803 16575
rect 8803 16541 8812 16575
rect 8760 16532 8812 16541
rect 11520 16575 11572 16584
rect 4620 16464 4672 16516
rect 9956 16464 10008 16516
rect 10140 16464 10192 16516
rect 11520 16541 11529 16575
rect 11529 16541 11563 16575
rect 11563 16541 11572 16575
rect 11520 16532 11572 16541
rect 21364 16668 21416 16720
rect 21640 16711 21692 16720
rect 21640 16677 21649 16711
rect 21649 16677 21683 16711
rect 21683 16677 21692 16711
rect 21640 16668 21692 16677
rect 23664 16668 23716 16720
rect 24768 16736 24820 16788
rect 24676 16668 24728 16720
rect 19984 16600 20036 16652
rect 22836 16643 22888 16652
rect 22836 16609 22845 16643
rect 22845 16609 22879 16643
rect 22879 16609 22888 16643
rect 22836 16600 22888 16609
rect 23112 16643 23164 16652
rect 23112 16609 23121 16643
rect 23121 16609 23155 16643
rect 23155 16609 23164 16643
rect 23112 16600 23164 16609
rect 16120 16575 16172 16584
rect 13176 16464 13228 16516
rect 1584 16396 1636 16448
rect 4068 16396 4120 16448
rect 4988 16396 5040 16448
rect 10784 16396 10836 16448
rect 13544 16396 13596 16448
rect 16120 16541 16129 16575
rect 16129 16541 16163 16575
rect 16163 16541 16172 16575
rect 16120 16532 16172 16541
rect 17684 16532 17736 16584
rect 18420 16575 18472 16584
rect 18420 16541 18429 16575
rect 18429 16541 18463 16575
rect 18463 16541 18472 16575
rect 18420 16532 18472 16541
rect 22284 16532 22336 16584
rect 23388 16575 23440 16584
rect 23388 16541 23397 16575
rect 23397 16541 23431 16575
rect 23431 16541 23440 16575
rect 23388 16532 23440 16541
rect 24952 16575 25004 16584
rect 24952 16541 24961 16575
rect 24961 16541 24995 16575
rect 24995 16541 25004 16575
rect 24952 16532 25004 16541
rect 25228 16532 25280 16584
rect 17408 16464 17460 16516
rect 18972 16464 19024 16516
rect 19432 16464 19484 16516
rect 14648 16396 14700 16448
rect 18328 16396 18380 16448
rect 18880 16396 18932 16448
rect 23664 16439 23716 16448
rect 23664 16405 23673 16439
rect 23673 16405 23707 16439
rect 23707 16405 23716 16439
rect 23664 16396 23716 16405
rect 23848 16396 23900 16448
rect 24032 16439 24084 16448
rect 24032 16405 24041 16439
rect 24041 16405 24075 16439
rect 24075 16405 24084 16439
rect 24032 16396 24084 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 1400 16192 1452 16244
rect 4160 16192 4212 16244
rect 6184 16235 6236 16244
rect 6184 16201 6193 16235
rect 6193 16201 6227 16235
rect 6227 16201 6236 16235
rect 6184 16192 6236 16201
rect 9956 16235 10008 16244
rect 9956 16201 9965 16235
rect 9965 16201 9999 16235
rect 9999 16201 10008 16235
rect 9956 16192 10008 16201
rect 13084 16192 13136 16244
rect 13544 16192 13596 16244
rect 13636 16192 13688 16244
rect 16580 16192 16632 16244
rect 17776 16235 17828 16244
rect 17776 16201 17785 16235
rect 17785 16201 17819 16235
rect 17819 16201 17828 16235
rect 17776 16192 17828 16201
rect 22284 16235 22336 16244
rect 22284 16201 22293 16235
rect 22293 16201 22327 16235
rect 22327 16201 22336 16235
rect 22284 16192 22336 16201
rect 23112 16192 23164 16244
rect 24676 16192 24728 16244
rect 25596 16235 25648 16244
rect 25596 16201 25605 16235
rect 25605 16201 25639 16235
rect 25639 16201 25648 16235
rect 25596 16192 25648 16201
rect 1676 16124 1728 16176
rect 2872 16124 2924 16176
rect 4068 16124 4120 16176
rect 2044 15988 2096 16040
rect 112 15852 164 15904
rect 2044 15895 2096 15904
rect 2044 15861 2053 15895
rect 2053 15861 2087 15895
rect 2087 15861 2096 15895
rect 2044 15852 2096 15861
rect 3516 15988 3568 16040
rect 4160 16056 4212 16108
rect 5172 16056 5224 16108
rect 11888 16124 11940 16176
rect 15384 16124 15436 16176
rect 3332 15920 3384 15972
rect 3700 15920 3752 15972
rect 5356 16031 5408 16040
rect 5356 15997 5365 16031
rect 5365 15997 5399 16031
rect 5399 15997 5408 16031
rect 5356 15988 5408 15997
rect 6368 15988 6420 16040
rect 6276 15920 6328 15972
rect 8668 15988 8720 16040
rect 9588 15988 9640 16040
rect 11152 16056 11204 16108
rect 11520 16056 11572 16108
rect 12532 16099 12584 16108
rect 12532 16065 12541 16099
rect 12541 16065 12575 16099
rect 12575 16065 12584 16099
rect 12532 16056 12584 16065
rect 14188 16031 14240 16040
rect 14188 15997 14197 16031
rect 14197 15997 14231 16031
rect 14231 15997 14240 16031
rect 14188 15988 14240 15997
rect 7472 15920 7524 15972
rect 7564 15920 7616 15972
rect 8392 15920 8444 15972
rect 2964 15852 3016 15904
rect 3884 15852 3936 15904
rect 5264 15895 5316 15904
rect 5264 15861 5273 15895
rect 5273 15861 5307 15895
rect 5307 15861 5316 15895
rect 5264 15852 5316 15861
rect 7840 15852 7892 15904
rect 8300 15895 8352 15904
rect 8300 15861 8309 15895
rect 8309 15861 8343 15895
rect 8343 15861 8352 15895
rect 10048 15920 10100 15972
rect 13176 15963 13228 15972
rect 8300 15852 8352 15861
rect 9772 15852 9824 15904
rect 11888 15852 11940 15904
rect 12256 15895 12308 15904
rect 12256 15861 12265 15895
rect 12265 15861 12299 15895
rect 12299 15861 12308 15895
rect 13176 15929 13185 15963
rect 13185 15929 13219 15963
rect 13219 15929 13228 15963
rect 13176 15920 13228 15929
rect 24768 16124 24820 16176
rect 15752 16056 15804 16108
rect 19340 16056 19392 16108
rect 20904 16056 20956 16108
rect 21548 16056 21600 16108
rect 19064 15988 19116 16040
rect 23296 15988 23348 16040
rect 24032 16056 24084 16108
rect 23940 15988 23992 16040
rect 12256 15852 12308 15861
rect 12900 15852 12952 15904
rect 21364 15963 21416 15972
rect 21364 15929 21373 15963
rect 21373 15929 21407 15963
rect 21407 15929 21416 15963
rect 21916 15963 21968 15972
rect 21364 15920 21416 15929
rect 21916 15929 21925 15963
rect 21925 15929 21959 15963
rect 21959 15929 21968 15963
rect 21916 15920 21968 15929
rect 24032 15963 24084 15972
rect 14096 15895 14148 15904
rect 14096 15861 14105 15895
rect 14105 15861 14139 15895
rect 14139 15861 14148 15895
rect 14096 15852 14148 15861
rect 16028 15852 16080 15904
rect 17224 15852 17276 15904
rect 17868 15852 17920 15904
rect 18880 15895 18932 15904
rect 18880 15861 18889 15895
rect 18889 15861 18923 15895
rect 18923 15861 18932 15895
rect 18880 15852 18932 15861
rect 19984 15852 20036 15904
rect 22836 15852 22888 15904
rect 23204 15852 23256 15904
rect 24032 15929 24035 15963
rect 24035 15929 24069 15963
rect 24069 15929 24084 15963
rect 24032 15920 24084 15929
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2964 15648 3016 15700
rect 1952 15555 2004 15564
rect 1952 15521 1961 15555
rect 1961 15521 1995 15555
rect 1995 15521 2004 15555
rect 1952 15512 2004 15521
rect 2964 15555 3016 15564
rect 2964 15521 2973 15555
rect 2973 15521 3007 15555
rect 3007 15521 3016 15555
rect 2964 15512 3016 15521
rect 3240 15648 3292 15700
rect 5448 15648 5500 15700
rect 4160 15580 4212 15632
rect 4988 15580 5040 15632
rect 6184 15648 6236 15700
rect 6368 15648 6420 15700
rect 7564 15648 7616 15700
rect 8668 15691 8720 15700
rect 8668 15657 8677 15691
rect 8677 15657 8711 15691
rect 8711 15657 8720 15691
rect 8668 15648 8720 15657
rect 9404 15648 9456 15700
rect 9864 15648 9916 15700
rect 11520 15691 11572 15700
rect 11520 15657 11529 15691
rect 11529 15657 11563 15691
rect 11563 15657 11572 15691
rect 11520 15648 11572 15657
rect 13452 15648 13504 15700
rect 3240 15512 3292 15564
rect 3884 15512 3936 15564
rect 4528 15512 4580 15564
rect 5264 15512 5316 15564
rect 6184 15512 6236 15564
rect 10048 15580 10100 15632
rect 11888 15580 11940 15632
rect 13268 15623 13320 15632
rect 13268 15589 13277 15623
rect 13277 15589 13311 15623
rect 13311 15589 13320 15623
rect 13912 15648 13964 15700
rect 16120 15648 16172 15700
rect 19340 15648 19392 15700
rect 21364 15648 21416 15700
rect 21548 15691 21600 15700
rect 21548 15657 21557 15691
rect 21557 15657 21591 15691
rect 21591 15657 21600 15691
rect 21548 15648 21600 15657
rect 24032 15691 24084 15700
rect 24032 15657 24041 15691
rect 24041 15657 24075 15691
rect 24075 15657 24084 15691
rect 24032 15648 24084 15657
rect 13268 15580 13320 15589
rect 17960 15580 18012 15632
rect 18144 15580 18196 15632
rect 18420 15580 18472 15632
rect 18880 15580 18932 15632
rect 8760 15512 8812 15564
rect 9956 15555 10008 15564
rect 9956 15521 9965 15555
rect 9965 15521 9999 15555
rect 9999 15521 10008 15555
rect 9956 15512 10008 15521
rect 11796 15512 11848 15564
rect 12256 15512 12308 15564
rect 14556 15512 14608 15564
rect 15752 15555 15804 15564
rect 15752 15521 15761 15555
rect 15761 15521 15795 15555
rect 15795 15521 15804 15555
rect 15752 15512 15804 15521
rect 16672 15512 16724 15564
rect 17316 15555 17368 15564
rect 17316 15521 17325 15555
rect 17325 15521 17359 15555
rect 17359 15521 17368 15555
rect 17316 15512 17368 15521
rect 20812 15512 20864 15564
rect 21824 15512 21876 15564
rect 2872 15487 2924 15496
rect 2872 15453 2881 15487
rect 2881 15453 2915 15487
rect 2915 15453 2924 15487
rect 2872 15444 2924 15453
rect 3700 15444 3752 15496
rect 7104 15487 7156 15496
rect 7104 15453 7113 15487
rect 7113 15453 7147 15487
rect 7147 15453 7156 15487
rect 7104 15444 7156 15453
rect 11704 15487 11756 15496
rect 11704 15453 11713 15487
rect 11713 15453 11747 15487
rect 11747 15453 11756 15487
rect 11704 15444 11756 15453
rect 7196 15376 7248 15428
rect 8484 15376 8536 15428
rect 12900 15376 12952 15428
rect 13176 15376 13228 15428
rect 19524 15444 19576 15496
rect 21548 15444 21600 15496
rect 23204 15580 23256 15632
rect 23388 15512 23440 15564
rect 24032 15512 24084 15564
rect 24216 15512 24268 15564
rect 25412 15555 25464 15564
rect 25412 15521 25421 15555
rect 25421 15521 25455 15555
rect 25455 15521 25464 15555
rect 25412 15512 25464 15521
rect 13912 15376 13964 15428
rect 16120 15376 16172 15428
rect 17684 15376 17736 15428
rect 1860 15351 1912 15360
rect 1860 15317 1869 15351
rect 1869 15317 1903 15351
rect 1903 15317 1912 15351
rect 1860 15308 1912 15317
rect 2412 15351 2464 15360
rect 2412 15317 2421 15351
rect 2421 15317 2455 15351
rect 2455 15317 2464 15351
rect 2412 15308 2464 15317
rect 2596 15308 2648 15360
rect 4804 15351 4856 15360
rect 4804 15317 4813 15351
rect 4813 15317 4847 15351
rect 4847 15317 4856 15351
rect 4804 15308 4856 15317
rect 6552 15351 6604 15360
rect 6552 15317 6561 15351
rect 6561 15317 6595 15351
rect 6595 15317 6604 15351
rect 6552 15308 6604 15317
rect 7012 15308 7064 15360
rect 16396 15308 16448 15360
rect 18604 15308 18656 15360
rect 19156 15308 19208 15360
rect 22192 15308 22244 15360
rect 24676 15308 24728 15360
rect 24952 15351 25004 15360
rect 24952 15317 24961 15351
rect 24961 15317 24995 15351
rect 24995 15317 25004 15351
rect 24952 15308 25004 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2504 15104 2556 15156
rect 2872 15104 2924 15156
rect 4528 15147 4580 15156
rect 4528 15113 4537 15147
rect 4537 15113 4571 15147
rect 4571 15113 4580 15147
rect 4528 15104 4580 15113
rect 9404 15147 9456 15156
rect 9404 15113 9413 15147
rect 9413 15113 9447 15147
rect 9447 15113 9456 15147
rect 9404 15104 9456 15113
rect 10048 15147 10100 15156
rect 10048 15113 10057 15147
rect 10057 15113 10091 15147
rect 10091 15113 10100 15147
rect 10048 15104 10100 15113
rect 11888 15104 11940 15156
rect 12992 15147 13044 15156
rect 12992 15113 13001 15147
rect 13001 15113 13035 15147
rect 13035 15113 13044 15147
rect 12992 15104 13044 15113
rect 13452 15147 13504 15156
rect 13452 15113 13461 15147
rect 13461 15113 13495 15147
rect 13495 15113 13504 15147
rect 13452 15104 13504 15113
rect 15752 15104 15804 15156
rect 17316 15147 17368 15156
rect 17316 15113 17325 15147
rect 17325 15113 17359 15147
rect 17359 15113 17368 15147
rect 17316 15104 17368 15113
rect 19524 15104 19576 15156
rect 2228 15079 2280 15088
rect 2228 15045 2237 15079
rect 2237 15045 2271 15079
rect 2271 15045 2280 15079
rect 2228 15036 2280 15045
rect 4436 15036 4488 15088
rect 6920 15036 6972 15088
rect 11704 15036 11756 15088
rect 14096 15036 14148 15088
rect 2320 15011 2372 15020
rect 2320 14977 2329 15011
rect 2329 14977 2363 15011
rect 2363 14977 2372 15011
rect 2320 14968 2372 14977
rect 2412 14900 2464 14952
rect 2596 14900 2648 14952
rect 2872 14900 2924 14952
rect 3976 14943 4028 14952
rect 3976 14909 3985 14943
rect 3985 14909 4019 14943
rect 4019 14909 4028 14943
rect 3976 14900 4028 14909
rect 4896 14900 4948 14952
rect 4160 14832 4212 14884
rect 5448 14900 5500 14952
rect 7104 14968 7156 15020
rect 7380 15011 7432 15020
rect 7380 14977 7389 15011
rect 7389 14977 7423 15011
rect 7423 14977 7432 15011
rect 7380 14968 7432 14977
rect 7932 14968 7984 15020
rect 8484 15011 8536 15020
rect 8484 14977 8493 15011
rect 8493 14977 8527 15011
rect 8527 14977 8536 15011
rect 8484 14968 8536 14977
rect 10784 14968 10836 15020
rect 6736 14900 6788 14952
rect 11060 14943 11112 14952
rect 11060 14909 11069 14943
rect 11069 14909 11103 14943
rect 11103 14909 11112 14943
rect 11060 14900 11112 14909
rect 13820 14968 13872 15020
rect 14188 14968 14240 15020
rect 17040 15036 17092 15088
rect 18972 15036 19024 15088
rect 16212 15011 16264 15020
rect 12164 14900 12216 14952
rect 12992 14900 13044 14952
rect 16212 14977 16221 15011
rect 16221 14977 16255 15011
rect 16255 14977 16264 15011
rect 16212 14968 16264 14977
rect 19432 14968 19484 15020
rect 5724 14832 5776 14884
rect 6920 14875 6972 14884
rect 6920 14841 6929 14875
rect 6929 14841 6963 14875
rect 6963 14841 6972 14875
rect 6920 14832 6972 14841
rect 7012 14875 7064 14884
rect 7012 14841 7021 14875
rect 7021 14841 7055 14875
rect 7055 14841 7064 14875
rect 7012 14832 7064 14841
rect 11520 14875 11572 14884
rect 1952 14764 2004 14816
rect 2596 14764 2648 14816
rect 5172 14764 5224 14816
rect 6184 14807 6236 14816
rect 6184 14773 6193 14807
rect 6193 14773 6227 14807
rect 6227 14773 6236 14807
rect 6184 14764 6236 14773
rect 6644 14764 6696 14816
rect 8300 14807 8352 14816
rect 8300 14773 8309 14807
rect 8309 14773 8343 14807
rect 8343 14773 8352 14807
rect 11520 14841 11529 14875
rect 11529 14841 11563 14875
rect 11563 14841 11572 14875
rect 11520 14832 11572 14841
rect 14372 14875 14424 14884
rect 8300 14764 8352 14773
rect 10692 14764 10744 14816
rect 11612 14764 11664 14816
rect 11888 14807 11940 14816
rect 11888 14773 11897 14807
rect 11897 14773 11931 14807
rect 11931 14773 11940 14807
rect 11888 14764 11940 14773
rect 12440 14764 12492 14816
rect 13452 14764 13504 14816
rect 14372 14841 14381 14875
rect 14381 14841 14415 14875
rect 14415 14841 14424 14875
rect 14372 14832 14424 14841
rect 16396 14900 16448 14952
rect 18604 14943 18656 14952
rect 17684 14764 17736 14816
rect 18604 14909 18613 14943
rect 18613 14909 18647 14943
rect 18647 14909 18656 14943
rect 18604 14900 18656 14909
rect 19156 14943 19208 14952
rect 19156 14909 19165 14943
rect 19165 14909 19199 14943
rect 19199 14909 19208 14943
rect 23112 15104 23164 15156
rect 23388 15147 23440 15156
rect 23388 15113 23397 15147
rect 23397 15113 23431 15147
rect 23431 15113 23440 15147
rect 23388 15104 23440 15113
rect 24676 15104 24728 15156
rect 19984 15036 20036 15088
rect 20536 15011 20588 15020
rect 20536 14977 20545 15011
rect 20545 14977 20579 15011
rect 20579 14977 20588 15011
rect 20536 14968 20588 14977
rect 22008 15036 22060 15088
rect 23204 15036 23256 15088
rect 21916 14968 21968 15020
rect 24952 14968 25004 15020
rect 25228 15011 25280 15020
rect 25228 14977 25237 15011
rect 25237 14977 25271 15011
rect 25271 14977 25280 15011
rect 25228 14968 25280 14977
rect 19156 14900 19208 14909
rect 18144 14764 18196 14816
rect 18420 14807 18472 14816
rect 18420 14773 18429 14807
rect 18429 14773 18463 14807
rect 18463 14773 18472 14807
rect 18420 14764 18472 14773
rect 20812 14832 20864 14884
rect 22192 14875 22244 14884
rect 22192 14841 22201 14875
rect 22201 14841 22235 14875
rect 22235 14841 22244 14875
rect 22192 14832 22244 14841
rect 24676 14875 24728 14884
rect 24676 14841 24685 14875
rect 24685 14841 24719 14875
rect 24719 14841 24728 14875
rect 24676 14832 24728 14841
rect 21548 14764 21600 14816
rect 24860 14764 24912 14816
rect 25412 14764 25464 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2320 14560 2372 14612
rect 2964 14603 3016 14612
rect 2964 14569 2973 14603
rect 2973 14569 3007 14603
rect 3007 14569 3016 14603
rect 2964 14560 3016 14569
rect 3884 14560 3936 14612
rect 5264 14560 5316 14612
rect 7012 14560 7064 14612
rect 7104 14560 7156 14612
rect 7380 14560 7432 14612
rect 8484 14603 8536 14612
rect 2044 14535 2096 14544
rect 2044 14501 2053 14535
rect 2053 14501 2087 14535
rect 2087 14501 2096 14535
rect 2044 14492 2096 14501
rect 2780 14492 2832 14544
rect 3976 14492 4028 14544
rect 4528 14492 4580 14544
rect 6552 14492 6604 14544
rect 7656 14535 7708 14544
rect 7656 14501 7665 14535
rect 7665 14501 7699 14535
rect 7699 14501 7708 14535
rect 7656 14492 7708 14501
rect 8484 14569 8493 14603
rect 8493 14569 8527 14603
rect 8527 14569 8536 14603
rect 8484 14560 8536 14569
rect 9496 14603 9548 14612
rect 9496 14569 9505 14603
rect 9505 14569 9539 14603
rect 9539 14569 9548 14603
rect 9496 14560 9548 14569
rect 10140 14560 10192 14612
rect 10784 14603 10836 14612
rect 9772 14492 9824 14544
rect 10784 14569 10793 14603
rect 10793 14569 10827 14603
rect 10827 14569 10836 14603
rect 10784 14560 10836 14569
rect 13452 14560 13504 14612
rect 14280 14560 14332 14612
rect 16948 14603 17000 14612
rect 11796 14535 11848 14544
rect 11796 14501 11805 14535
rect 11805 14501 11839 14535
rect 11839 14501 11848 14535
rect 11796 14492 11848 14501
rect 13636 14492 13688 14544
rect 13912 14535 13964 14544
rect 13912 14501 13921 14535
rect 13921 14501 13955 14535
rect 13955 14501 13964 14535
rect 13912 14492 13964 14501
rect 15384 14492 15436 14544
rect 16948 14569 16957 14603
rect 16957 14569 16991 14603
rect 16991 14569 17000 14603
rect 16948 14560 17000 14569
rect 18788 14560 18840 14612
rect 20536 14603 20588 14612
rect 20536 14569 20545 14603
rect 20545 14569 20579 14603
rect 20579 14569 20588 14603
rect 20536 14560 20588 14569
rect 22192 14560 22244 14612
rect 23480 14560 23532 14612
rect 18236 14492 18288 14544
rect 19156 14492 19208 14544
rect 19432 14535 19484 14544
rect 19432 14501 19441 14535
rect 19441 14501 19475 14535
rect 19475 14501 19484 14535
rect 19432 14492 19484 14501
rect 21088 14535 21140 14544
rect 21088 14501 21097 14535
rect 21097 14501 21131 14535
rect 21131 14501 21140 14535
rect 21088 14492 21140 14501
rect 21640 14535 21692 14544
rect 21640 14501 21649 14535
rect 21649 14501 21683 14535
rect 21683 14501 21692 14535
rect 21640 14492 21692 14501
rect 21824 14492 21876 14544
rect 23296 14535 23348 14544
rect 23296 14501 23305 14535
rect 23305 14501 23339 14535
rect 23339 14501 23348 14535
rect 23296 14492 23348 14501
rect 24768 14560 24820 14612
rect 24676 14492 24728 14544
rect 5540 14424 5592 14476
rect 6092 14467 6144 14476
rect 6092 14433 6101 14467
rect 6101 14433 6135 14467
rect 6135 14433 6144 14467
rect 6092 14424 6144 14433
rect 17316 14467 17368 14476
rect 2136 14356 2188 14408
rect 3056 14356 3108 14408
rect 5724 14356 5776 14408
rect 6368 14399 6420 14408
rect 6368 14365 6377 14399
rect 6377 14365 6411 14399
rect 6411 14365 6420 14399
rect 6368 14356 6420 14365
rect 8576 14356 8628 14408
rect 11704 14399 11756 14408
rect 9220 14288 9272 14340
rect 9680 14288 9732 14340
rect 11704 14365 11713 14399
rect 11713 14365 11747 14399
rect 11747 14365 11756 14399
rect 11704 14356 11756 14365
rect 12532 14356 12584 14408
rect 13268 14399 13320 14408
rect 13268 14365 13277 14399
rect 13277 14365 13311 14399
rect 13311 14365 13320 14399
rect 13268 14356 13320 14365
rect 15660 14399 15712 14408
rect 14832 14288 14884 14340
rect 15660 14365 15669 14399
rect 15669 14365 15703 14399
rect 15703 14365 15712 14399
rect 15660 14356 15712 14365
rect 17316 14433 17325 14467
rect 17325 14433 17359 14467
rect 17359 14433 17368 14467
rect 17316 14424 17368 14433
rect 22928 14424 22980 14476
rect 23112 14467 23164 14476
rect 23112 14433 23121 14467
rect 23121 14433 23155 14467
rect 23155 14433 23164 14467
rect 23112 14424 23164 14433
rect 17592 14356 17644 14408
rect 19984 14399 20036 14408
rect 15568 14288 15620 14340
rect 19984 14365 19993 14399
rect 19993 14365 20027 14399
rect 20027 14365 20036 14399
rect 19984 14356 20036 14365
rect 20168 14356 20220 14408
rect 21916 14356 21968 14408
rect 19524 14288 19576 14340
rect 20444 14288 20496 14340
rect 22008 14288 22060 14340
rect 24952 14356 25004 14408
rect 4344 14220 4396 14272
rect 8392 14220 8444 14272
rect 8852 14263 8904 14272
rect 8852 14229 8861 14263
rect 8861 14229 8895 14263
rect 8895 14229 8904 14263
rect 8852 14220 8904 14229
rect 14464 14220 14516 14272
rect 22836 14220 22888 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 2044 14016 2096 14068
rect 4528 14016 4580 14068
rect 4620 14016 4672 14068
rect 9404 14016 9456 14068
rect 9772 14016 9824 14068
rect 9956 14059 10008 14068
rect 9956 14025 9965 14059
rect 9965 14025 9999 14059
rect 9999 14025 10008 14059
rect 9956 14016 10008 14025
rect 11520 14016 11572 14068
rect 2320 13948 2372 14000
rect 2780 13948 2832 14000
rect 3700 13948 3752 14000
rect 3884 13948 3936 14000
rect 4896 13948 4948 14000
rect 9220 13991 9272 14000
rect 9220 13957 9229 13991
rect 9229 13957 9263 13991
rect 9263 13957 9272 13991
rect 9220 13948 9272 13957
rect 1584 13880 1636 13932
rect 3332 13880 3384 13932
rect 3976 13880 4028 13932
rect 5172 13880 5224 13932
rect 4620 13812 4672 13864
rect 6368 13880 6420 13932
rect 8852 13880 8904 13932
rect 4344 13744 4396 13796
rect 8300 13812 8352 13864
rect 6552 13787 6604 13796
rect 6552 13753 6561 13787
rect 6561 13753 6595 13787
rect 6595 13753 6604 13787
rect 6552 13744 6604 13753
rect 9496 13880 9548 13932
rect 13820 14016 13872 14068
rect 15384 14059 15436 14068
rect 15384 14025 15393 14059
rect 15393 14025 15427 14059
rect 15427 14025 15436 14059
rect 15384 14016 15436 14025
rect 17316 14016 17368 14068
rect 17592 14059 17644 14068
rect 17592 14025 17601 14059
rect 17601 14025 17635 14059
rect 17635 14025 17644 14059
rect 17592 14016 17644 14025
rect 19432 14016 19484 14068
rect 21088 14016 21140 14068
rect 21916 14059 21968 14068
rect 21916 14025 21925 14059
rect 21925 14025 21959 14059
rect 21959 14025 21968 14059
rect 21916 14016 21968 14025
rect 22928 14059 22980 14068
rect 22928 14025 22937 14059
rect 22937 14025 22971 14059
rect 22971 14025 22980 14059
rect 22928 14016 22980 14025
rect 23388 14016 23440 14068
rect 24676 14016 24728 14068
rect 24768 14016 24820 14068
rect 25412 14016 25464 14068
rect 12532 13948 12584 14000
rect 15292 13948 15344 14000
rect 18328 13948 18380 14000
rect 20076 13948 20128 14000
rect 14280 13923 14332 13932
rect 14280 13889 14289 13923
rect 14289 13889 14323 13923
rect 14323 13889 14332 13923
rect 14280 13880 14332 13889
rect 14372 13880 14424 13932
rect 15660 13880 15712 13932
rect 16212 13923 16264 13932
rect 16212 13889 16221 13923
rect 16221 13889 16255 13923
rect 16255 13889 16264 13923
rect 16212 13880 16264 13889
rect 16488 13923 16540 13932
rect 16488 13889 16497 13923
rect 16497 13889 16531 13923
rect 16531 13889 16540 13923
rect 16488 13880 16540 13889
rect 18788 13880 18840 13932
rect 20720 13880 20772 13932
rect 21640 13948 21692 14000
rect 23112 13948 23164 14000
rect 22652 13880 22704 13932
rect 23020 13880 23072 13932
rect 23480 13880 23532 13932
rect 11796 13812 11848 13864
rect 22008 13812 22060 13864
rect 22376 13812 22428 13864
rect 25228 13812 25280 13864
rect 5448 13676 5500 13728
rect 6276 13676 6328 13728
rect 9956 13744 10008 13796
rect 10048 13744 10100 13796
rect 10692 13744 10744 13796
rect 11888 13676 11940 13728
rect 13176 13676 13228 13728
rect 13636 13719 13688 13728
rect 13636 13685 13645 13719
rect 13645 13685 13679 13719
rect 13679 13685 13688 13719
rect 13636 13676 13688 13685
rect 16580 13744 16632 13796
rect 17408 13676 17460 13728
rect 17592 13676 17644 13728
rect 18144 13676 18196 13728
rect 21088 13787 21140 13796
rect 21088 13753 21097 13787
rect 21097 13753 21131 13787
rect 21131 13753 21140 13787
rect 21088 13744 21140 13753
rect 19064 13676 19116 13728
rect 23296 13676 23348 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 2228 13472 2280 13524
rect 2412 13472 2464 13524
rect 2780 13472 2832 13524
rect 3700 13515 3752 13524
rect 3700 13481 3709 13515
rect 3709 13481 3743 13515
rect 3743 13481 3752 13515
rect 3700 13472 3752 13481
rect 4436 13472 4488 13524
rect 6092 13472 6144 13524
rect 7656 13515 7708 13524
rect 7656 13481 7665 13515
rect 7665 13481 7699 13515
rect 7699 13481 7708 13515
rect 7656 13472 7708 13481
rect 8300 13515 8352 13524
rect 8300 13481 8309 13515
rect 8309 13481 8343 13515
rect 8343 13481 8352 13515
rect 8300 13472 8352 13481
rect 8576 13472 8628 13524
rect 9680 13472 9732 13524
rect 10692 13515 10744 13524
rect 10692 13481 10701 13515
rect 10701 13481 10735 13515
rect 10735 13481 10744 13515
rect 10692 13472 10744 13481
rect 11704 13515 11756 13524
rect 11704 13481 11713 13515
rect 11713 13481 11747 13515
rect 11747 13481 11756 13515
rect 11704 13472 11756 13481
rect 11888 13472 11940 13524
rect 13176 13472 13228 13524
rect 13268 13472 13320 13524
rect 14832 13472 14884 13524
rect 16212 13515 16264 13524
rect 16212 13481 16221 13515
rect 16221 13481 16255 13515
rect 16255 13481 16264 13515
rect 16212 13472 16264 13481
rect 16948 13472 17000 13524
rect 18236 13472 18288 13524
rect 19524 13472 19576 13524
rect 21088 13472 21140 13524
rect 24676 13515 24728 13524
rect 24676 13481 24685 13515
rect 24685 13481 24719 13515
rect 24719 13481 24728 13515
rect 24676 13472 24728 13481
rect 25136 13515 25188 13524
rect 25136 13481 25145 13515
rect 25145 13481 25179 13515
rect 25179 13481 25188 13515
rect 25136 13472 25188 13481
rect 1676 13404 1728 13456
rect 1860 13336 1912 13388
rect 2596 13404 2648 13456
rect 2964 13404 3016 13456
rect 6552 13404 6604 13456
rect 7564 13404 7616 13456
rect 9864 13447 9916 13456
rect 2780 13336 2832 13388
rect 4344 13379 4396 13388
rect 4344 13345 4353 13379
rect 4353 13345 4387 13379
rect 4387 13345 4396 13379
rect 4344 13336 4396 13345
rect 4436 13336 4488 13388
rect 4620 13336 4672 13388
rect 9864 13413 9873 13447
rect 9873 13413 9907 13447
rect 9907 13413 9916 13447
rect 9864 13404 9916 13413
rect 9956 13404 10008 13456
rect 13820 13447 13872 13456
rect 13820 13413 13829 13447
rect 13829 13413 13863 13447
rect 13863 13413 13872 13447
rect 13820 13404 13872 13413
rect 16304 13404 16356 13456
rect 16764 13447 16816 13456
rect 16764 13413 16773 13447
rect 16773 13413 16807 13447
rect 16807 13413 16816 13447
rect 16764 13404 16816 13413
rect 16856 13447 16908 13456
rect 16856 13413 16865 13447
rect 16865 13413 16899 13447
rect 16899 13413 16908 13447
rect 16856 13404 16908 13413
rect 17224 13404 17276 13456
rect 17408 13404 17460 13456
rect 17868 13404 17920 13456
rect 18420 13447 18472 13456
rect 18420 13413 18429 13447
rect 18429 13413 18463 13447
rect 18463 13413 18472 13447
rect 18420 13404 18472 13413
rect 18604 13404 18656 13456
rect 15292 13379 15344 13388
rect 15292 13345 15301 13379
rect 15301 13345 15335 13379
rect 15335 13345 15344 13379
rect 15292 13336 15344 13345
rect 21456 13404 21508 13456
rect 23296 13404 23348 13456
rect 23848 13447 23900 13456
rect 23848 13413 23851 13447
rect 23851 13413 23885 13447
rect 23885 13413 23900 13447
rect 23848 13404 23900 13413
rect 3516 13268 3568 13320
rect 3148 13132 3200 13184
rect 3976 13132 4028 13184
rect 6184 13175 6236 13184
rect 6184 13141 6193 13175
rect 6193 13141 6227 13175
rect 6227 13141 6236 13175
rect 6736 13268 6788 13320
rect 8024 13268 8076 13320
rect 9404 13268 9456 13320
rect 10876 13268 10928 13320
rect 11520 13268 11572 13320
rect 12348 13268 12400 13320
rect 13728 13311 13780 13320
rect 13728 13277 13737 13311
rect 13737 13277 13771 13311
rect 13771 13277 13780 13311
rect 13728 13268 13780 13277
rect 13912 13268 13964 13320
rect 16948 13268 17000 13320
rect 14188 13200 14240 13252
rect 15200 13200 15252 13252
rect 17224 13200 17276 13252
rect 18328 13268 18380 13320
rect 20168 13268 20220 13320
rect 20996 13268 21048 13320
rect 21364 13268 21416 13320
rect 23572 13336 23624 13388
rect 23756 13336 23808 13388
rect 25412 13336 25464 13388
rect 27712 13336 27764 13388
rect 21548 13268 21600 13320
rect 22100 13268 22152 13320
rect 6184 13132 6236 13141
rect 7196 13132 7248 13184
rect 12532 13132 12584 13184
rect 15844 13175 15896 13184
rect 15844 13141 15853 13175
rect 15853 13141 15887 13175
rect 15887 13141 15896 13175
rect 15844 13132 15896 13141
rect 23664 13200 23716 13252
rect 24216 13200 24268 13252
rect 20536 13132 20588 13184
rect 20720 13175 20772 13184
rect 20720 13141 20729 13175
rect 20729 13141 20763 13175
rect 20763 13141 20772 13175
rect 20720 13132 20772 13141
rect 21088 13132 21140 13184
rect 22376 13132 22428 13184
rect 24676 13132 24728 13184
rect 25504 13132 25556 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2228 12928 2280 12980
rect 2688 12928 2740 12980
rect 2780 12971 2832 12980
rect 2780 12937 2789 12971
rect 2789 12937 2823 12971
rect 2823 12937 2832 12971
rect 4344 12971 4396 12980
rect 2780 12928 2832 12937
rect 1860 12835 1912 12844
rect 1860 12801 1866 12835
rect 1866 12801 1912 12835
rect 1860 12792 1912 12801
rect 2412 12792 2464 12844
rect 4344 12937 4353 12971
rect 4353 12937 4387 12971
rect 4387 12937 4396 12971
rect 4344 12928 4396 12937
rect 6552 12928 6604 12980
rect 7012 12971 7064 12980
rect 7012 12937 7021 12971
rect 7021 12937 7055 12971
rect 7055 12937 7064 12971
rect 7012 12928 7064 12937
rect 10876 12971 10928 12980
rect 10876 12937 10885 12971
rect 10885 12937 10919 12971
rect 10919 12937 10928 12971
rect 10876 12928 10928 12937
rect 13820 12928 13872 12980
rect 16764 12928 16816 12980
rect 17868 12971 17920 12980
rect 17868 12937 17877 12971
rect 17877 12937 17911 12971
rect 17911 12937 17920 12971
rect 17868 12928 17920 12937
rect 3516 12860 3568 12912
rect 4252 12860 4304 12912
rect 3148 12724 3200 12776
rect 5448 12792 5500 12844
rect 3516 12724 3568 12776
rect 3700 12767 3752 12776
rect 3700 12733 3709 12767
rect 3709 12733 3743 12767
rect 3743 12733 3752 12767
rect 3700 12724 3752 12733
rect 8208 12860 8260 12912
rect 8484 12860 8536 12912
rect 8576 12860 8628 12912
rect 10140 12860 10192 12912
rect 11888 12860 11940 12912
rect 15660 12860 15712 12912
rect 16580 12903 16632 12912
rect 16580 12869 16589 12903
rect 16589 12869 16623 12903
rect 16623 12869 16632 12903
rect 18420 12928 18472 12980
rect 20168 12971 20220 12980
rect 20168 12937 20177 12971
rect 20177 12937 20211 12971
rect 20211 12937 20220 12971
rect 20168 12928 20220 12937
rect 21456 12928 21508 12980
rect 23572 12928 23624 12980
rect 23848 12971 23900 12980
rect 23848 12937 23857 12971
rect 23857 12937 23891 12971
rect 23891 12937 23900 12971
rect 23848 12928 23900 12937
rect 25412 12971 25464 12980
rect 25412 12937 25421 12971
rect 25421 12937 25455 12971
rect 25455 12937 25464 12971
rect 25412 12928 25464 12937
rect 16580 12860 16632 12869
rect 6184 12792 6236 12844
rect 6552 12792 6604 12844
rect 6092 12724 6144 12776
rect 8024 12792 8076 12844
rect 10968 12792 11020 12844
rect 12532 12835 12584 12844
rect 12532 12801 12541 12835
rect 12541 12801 12575 12835
rect 12575 12801 12584 12835
rect 12532 12792 12584 12801
rect 15108 12835 15160 12844
rect 15108 12801 15117 12835
rect 15117 12801 15151 12835
rect 15151 12801 15160 12835
rect 15108 12792 15160 12801
rect 3332 12631 3384 12640
rect 3332 12597 3341 12631
rect 3341 12597 3375 12631
rect 3375 12597 3384 12631
rect 3332 12588 3384 12597
rect 3516 12588 3568 12640
rect 7012 12656 7064 12708
rect 8024 12656 8076 12708
rect 14556 12767 14608 12776
rect 10048 12699 10100 12708
rect 10048 12665 10057 12699
rect 10057 12665 10091 12699
rect 10091 12665 10100 12699
rect 10048 12656 10100 12665
rect 12808 12656 12860 12708
rect 13452 12656 13504 12708
rect 13912 12699 13964 12708
rect 13912 12665 13921 12699
rect 13921 12665 13955 12699
rect 13955 12665 13964 12699
rect 14556 12733 14565 12767
rect 14565 12733 14599 12767
rect 14599 12733 14608 12767
rect 17776 12792 17828 12844
rect 14556 12724 14608 12733
rect 15844 12724 15896 12776
rect 17684 12724 17736 12776
rect 18972 12767 19024 12776
rect 18972 12733 18981 12767
rect 18981 12733 19015 12767
rect 19015 12733 19024 12767
rect 18972 12724 19024 12733
rect 13912 12656 13964 12665
rect 14464 12656 14516 12708
rect 14832 12699 14884 12708
rect 14832 12665 14841 12699
rect 14841 12665 14875 12699
rect 14875 12665 14884 12699
rect 14832 12656 14884 12665
rect 7564 12631 7616 12640
rect 7564 12597 7573 12631
rect 7573 12597 7607 12631
rect 7607 12597 7616 12631
rect 7564 12588 7616 12597
rect 9864 12588 9916 12640
rect 11520 12631 11572 12640
rect 11520 12597 11529 12631
rect 11529 12597 11563 12631
rect 11563 12597 11572 12631
rect 11520 12588 11572 12597
rect 11704 12588 11756 12640
rect 11888 12631 11940 12640
rect 11888 12597 11897 12631
rect 11897 12597 11931 12631
rect 11931 12597 11940 12631
rect 11888 12588 11940 12597
rect 15660 12588 15712 12640
rect 18144 12656 18196 12708
rect 22192 12860 22244 12912
rect 22376 12860 22428 12912
rect 24952 12903 25004 12912
rect 24952 12869 24961 12903
rect 24961 12869 24995 12903
rect 24995 12869 25004 12903
rect 24952 12860 25004 12869
rect 20812 12835 20864 12844
rect 20812 12801 20821 12835
rect 20821 12801 20855 12835
rect 20855 12801 20864 12835
rect 20812 12792 20864 12801
rect 21088 12835 21140 12844
rect 21088 12801 21097 12835
rect 21097 12801 21131 12835
rect 21131 12801 21140 12835
rect 21088 12792 21140 12801
rect 25136 12792 25188 12844
rect 16856 12631 16908 12640
rect 16856 12597 16865 12631
rect 16865 12597 16899 12631
rect 16899 12597 16908 12631
rect 16856 12588 16908 12597
rect 17316 12588 17368 12640
rect 18696 12588 18748 12640
rect 19524 12588 19576 12640
rect 21824 12588 21876 12640
rect 24492 12699 24544 12708
rect 24492 12665 24501 12699
rect 24501 12665 24535 12699
rect 24535 12665 24544 12699
rect 24492 12656 24544 12665
rect 24676 12656 24728 12708
rect 23112 12588 23164 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1952 12384 2004 12436
rect 3332 12384 3384 12436
rect 3608 12384 3660 12436
rect 5080 12384 5132 12436
rect 7012 12427 7064 12436
rect 2228 12359 2280 12368
rect 2228 12325 2237 12359
rect 2237 12325 2271 12359
rect 2271 12325 2280 12359
rect 2228 12316 2280 12325
rect 3792 12316 3844 12368
rect 3976 12316 4028 12368
rect 5540 12316 5592 12368
rect 7012 12393 7021 12427
rect 7021 12393 7055 12427
rect 7055 12393 7064 12427
rect 7012 12384 7064 12393
rect 8024 12427 8076 12436
rect 8024 12393 8033 12427
rect 8033 12393 8067 12427
rect 8067 12393 8076 12427
rect 8024 12384 8076 12393
rect 9312 12384 9364 12436
rect 7748 12316 7800 12368
rect 10968 12384 11020 12436
rect 11520 12427 11572 12436
rect 11520 12393 11529 12427
rect 11529 12393 11563 12427
rect 11563 12393 11572 12427
rect 11520 12384 11572 12393
rect 13728 12384 13780 12436
rect 17684 12427 17736 12436
rect 17684 12393 17693 12427
rect 17693 12393 17727 12427
rect 17727 12393 17736 12427
rect 17684 12384 17736 12393
rect 9864 12359 9916 12368
rect 9864 12325 9873 12359
rect 9873 12325 9907 12359
rect 9907 12325 9916 12359
rect 9864 12316 9916 12325
rect 10232 12316 10284 12368
rect 13636 12316 13688 12368
rect 14556 12316 14608 12368
rect 15660 12316 15712 12368
rect 21364 12427 21416 12436
rect 21364 12393 21373 12427
rect 21373 12393 21407 12427
rect 21407 12393 21416 12427
rect 21364 12384 21416 12393
rect 24492 12384 24544 12436
rect 1768 12248 1820 12300
rect 3700 12248 3752 12300
rect 2504 12180 2556 12232
rect 4988 12248 5040 12300
rect 5356 12291 5408 12300
rect 5356 12257 5365 12291
rect 5365 12257 5399 12291
rect 5399 12257 5408 12291
rect 5356 12248 5408 12257
rect 6000 12291 6052 12300
rect 6000 12257 6009 12291
rect 6009 12257 6043 12291
rect 6043 12257 6052 12291
rect 6000 12248 6052 12257
rect 6092 12248 6144 12300
rect 6828 12248 6880 12300
rect 8760 12248 8812 12300
rect 6644 12223 6696 12232
rect 6644 12189 6653 12223
rect 6653 12189 6687 12223
rect 6687 12189 6696 12223
rect 6644 12180 6696 12189
rect 7380 12180 7432 12232
rect 10140 12223 10192 12232
rect 10140 12189 10149 12223
rect 10149 12189 10183 12223
rect 10183 12189 10192 12223
rect 10140 12180 10192 12189
rect 12164 12248 12216 12300
rect 14372 12248 14424 12300
rect 19524 12316 19576 12368
rect 19984 12359 20036 12368
rect 19984 12325 19993 12359
rect 19993 12325 20027 12359
rect 20027 12325 20036 12359
rect 19984 12316 20036 12325
rect 22468 12359 22520 12368
rect 22468 12325 22477 12359
rect 22477 12325 22511 12359
rect 22511 12325 22520 12359
rect 22468 12316 22520 12325
rect 24768 12316 24820 12368
rect 25044 12316 25096 12368
rect 17592 12291 17644 12300
rect 17592 12257 17601 12291
rect 17601 12257 17635 12291
rect 17635 12257 17644 12291
rect 17592 12248 17644 12257
rect 17684 12248 17736 12300
rect 19064 12248 19116 12300
rect 21456 12248 21508 12300
rect 11888 12180 11940 12232
rect 14096 12180 14148 12232
rect 9864 12112 9916 12164
rect 13452 12155 13504 12164
rect 13452 12121 13461 12155
rect 13461 12121 13495 12155
rect 13495 12121 13504 12155
rect 13452 12112 13504 12121
rect 1860 12044 1912 12096
rect 3884 12087 3936 12096
rect 3884 12053 3893 12087
rect 3893 12053 3927 12087
rect 3927 12053 3936 12087
rect 3884 12044 3936 12053
rect 4344 12087 4396 12096
rect 4344 12053 4353 12087
rect 4353 12053 4387 12087
rect 4387 12053 4396 12087
rect 4344 12044 4396 12053
rect 4528 12044 4580 12096
rect 4896 12044 4948 12096
rect 12808 12044 12860 12096
rect 15292 12044 15344 12096
rect 16304 12044 16356 12096
rect 16856 12044 16908 12096
rect 17040 12087 17092 12096
rect 17040 12053 17049 12087
rect 17049 12053 17083 12087
rect 17083 12053 17092 12087
rect 17040 12044 17092 12053
rect 18420 12044 18472 12096
rect 20536 12180 20588 12232
rect 22376 12223 22428 12232
rect 22376 12189 22385 12223
rect 22385 12189 22419 12223
rect 22419 12189 22428 12223
rect 22376 12180 22428 12189
rect 22652 12223 22704 12232
rect 22652 12189 22661 12223
rect 22661 12189 22695 12223
rect 22695 12189 22704 12223
rect 22652 12180 22704 12189
rect 18972 12112 19024 12164
rect 22928 12112 22980 12164
rect 23296 12112 23348 12164
rect 25412 12180 25464 12232
rect 21916 12087 21968 12096
rect 21916 12053 21925 12087
rect 21925 12053 21959 12087
rect 21959 12053 21968 12087
rect 21916 12044 21968 12053
rect 22652 12044 22704 12096
rect 25044 12044 25096 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1768 11840 1820 11892
rect 2228 11840 2280 11892
rect 2872 11883 2924 11892
rect 2872 11849 2881 11883
rect 2881 11849 2915 11883
rect 2915 11849 2924 11883
rect 2872 11840 2924 11849
rect 4344 11840 4396 11892
rect 4804 11840 4856 11892
rect 5540 11840 5592 11892
rect 6000 11840 6052 11892
rect 8668 11840 8720 11892
rect 10232 11883 10284 11892
rect 10232 11849 10241 11883
rect 10241 11849 10275 11883
rect 10275 11849 10284 11883
rect 10232 11840 10284 11849
rect 12164 11883 12216 11892
rect 12164 11849 12173 11883
rect 12173 11849 12207 11883
rect 12207 11849 12216 11883
rect 12164 11840 12216 11849
rect 14096 11883 14148 11892
rect 14096 11849 14105 11883
rect 14105 11849 14139 11883
rect 14139 11849 14148 11883
rect 19524 11883 19576 11892
rect 14096 11840 14148 11849
rect 3332 11772 3384 11824
rect 3700 11815 3752 11824
rect 3700 11781 3709 11815
rect 3709 11781 3743 11815
rect 3743 11781 3752 11815
rect 3700 11772 3752 11781
rect 2504 11704 2556 11756
rect 5816 11772 5868 11824
rect 7840 11772 7892 11824
rect 9864 11772 9916 11824
rect 10692 11772 10744 11824
rect 13728 11772 13780 11824
rect 14004 11772 14056 11824
rect 7748 11747 7800 11756
rect 7748 11713 7757 11747
rect 7757 11713 7791 11747
rect 7791 11713 7800 11747
rect 7748 11704 7800 11713
rect 8116 11704 8168 11756
rect 9312 11747 9364 11756
rect 9312 11713 9321 11747
rect 9321 11713 9355 11747
rect 9355 11713 9364 11747
rect 9312 11704 9364 11713
rect 9956 11747 10008 11756
rect 9956 11713 9965 11747
rect 9965 11713 9999 11747
rect 9999 11713 10008 11747
rect 9956 11704 10008 11713
rect 12440 11704 12492 11756
rect 15292 11747 15344 11756
rect 15292 11713 15301 11747
rect 15301 11713 15335 11747
rect 15335 11713 15344 11747
rect 15292 11704 15344 11713
rect 15660 11704 15712 11756
rect 17040 11772 17092 11824
rect 16488 11747 16540 11756
rect 16488 11713 16497 11747
rect 16497 11713 16531 11747
rect 16531 11713 16540 11747
rect 16488 11704 16540 11713
rect 2228 11679 2280 11688
rect 2228 11645 2237 11679
rect 2237 11645 2271 11679
rect 2271 11645 2280 11679
rect 2228 11636 2280 11645
rect 3884 11636 3936 11688
rect 5356 11679 5408 11688
rect 5356 11645 5365 11679
rect 5365 11645 5399 11679
rect 5399 11645 5408 11679
rect 5356 11636 5408 11645
rect 5448 11636 5500 11688
rect 8576 11636 8628 11688
rect 9128 11636 9180 11688
rect 3608 11568 3660 11620
rect 4344 11568 4396 11620
rect 7840 11611 7892 11620
rect 7840 11577 7849 11611
rect 7849 11577 7883 11611
rect 7883 11577 7892 11611
rect 7840 11568 7892 11577
rect 2412 11500 2464 11552
rect 2596 11500 2648 11552
rect 4436 11500 4488 11552
rect 7380 11500 7432 11552
rect 8024 11500 8076 11552
rect 8852 11500 8904 11552
rect 9588 11500 9640 11552
rect 10048 11500 10100 11552
rect 11152 11636 11204 11688
rect 14740 11679 14792 11688
rect 14740 11645 14749 11679
rect 14749 11645 14783 11679
rect 14783 11645 14792 11679
rect 14740 11636 14792 11645
rect 15108 11679 15160 11688
rect 15108 11645 15117 11679
rect 15117 11645 15151 11679
rect 15151 11645 15160 11679
rect 15108 11636 15160 11645
rect 11520 11611 11572 11620
rect 11520 11577 11529 11611
rect 11529 11577 11563 11611
rect 11563 11577 11572 11611
rect 11520 11568 11572 11577
rect 12808 11611 12860 11620
rect 12808 11577 12817 11611
rect 12817 11577 12851 11611
rect 12851 11577 12860 11611
rect 12808 11568 12860 11577
rect 13360 11611 13412 11620
rect 13360 11577 13369 11611
rect 13369 11577 13403 11611
rect 13403 11577 13412 11611
rect 13360 11568 13412 11577
rect 11888 11543 11940 11552
rect 11888 11509 11897 11543
rect 11897 11509 11931 11543
rect 11931 11509 11940 11543
rect 11888 11500 11940 11509
rect 13636 11543 13688 11552
rect 13636 11509 13645 11543
rect 13645 11509 13679 11543
rect 13679 11509 13688 11543
rect 13636 11500 13688 11509
rect 16304 11611 16356 11620
rect 16304 11577 16313 11611
rect 16313 11577 16347 11611
rect 16347 11577 16356 11611
rect 16304 11568 16356 11577
rect 17684 11772 17736 11824
rect 19524 11849 19533 11883
rect 19533 11849 19567 11883
rect 19567 11849 19576 11883
rect 19524 11840 19576 11849
rect 22468 11840 22520 11892
rect 22836 11840 22888 11892
rect 24124 11840 24176 11892
rect 25412 11883 25464 11892
rect 20168 11772 20220 11824
rect 20352 11772 20404 11824
rect 17592 11747 17644 11756
rect 17592 11713 17601 11747
rect 17601 11713 17635 11747
rect 17635 11713 17644 11747
rect 17592 11704 17644 11713
rect 22376 11772 22428 11824
rect 20536 11704 20588 11756
rect 22652 11747 22704 11756
rect 22652 11713 22661 11747
rect 22661 11713 22695 11747
rect 22695 11713 22704 11747
rect 22652 11704 22704 11713
rect 25412 11849 25421 11883
rect 25421 11849 25455 11883
rect 25455 11849 25464 11883
rect 25412 11840 25464 11849
rect 25044 11815 25096 11824
rect 25044 11781 25053 11815
rect 25053 11781 25087 11815
rect 25087 11781 25096 11815
rect 25044 11772 25096 11781
rect 18236 11500 18288 11552
rect 18972 11679 19024 11688
rect 18972 11645 18981 11679
rect 18981 11645 19015 11679
rect 19015 11645 19024 11679
rect 18972 11636 19024 11645
rect 22008 11611 22060 11620
rect 22008 11577 22017 11611
rect 22017 11577 22051 11611
rect 22051 11577 22060 11611
rect 22008 11568 22060 11577
rect 18788 11543 18840 11552
rect 18788 11509 18797 11543
rect 18797 11509 18831 11543
rect 18831 11509 18840 11543
rect 18788 11500 18840 11509
rect 20260 11543 20312 11552
rect 20260 11509 20269 11543
rect 20269 11509 20303 11543
rect 20303 11509 20312 11543
rect 20260 11500 20312 11509
rect 21456 11543 21508 11552
rect 21456 11509 21465 11543
rect 21465 11509 21499 11543
rect 21499 11509 21508 11543
rect 21456 11500 21508 11509
rect 21732 11543 21784 11552
rect 21732 11509 21741 11543
rect 21741 11509 21775 11543
rect 21775 11509 21784 11543
rect 24584 11611 24636 11620
rect 24584 11577 24593 11611
rect 24593 11577 24627 11611
rect 24627 11577 24636 11611
rect 24584 11568 24636 11577
rect 21732 11500 21784 11509
rect 24768 11500 24820 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1860 11296 1912 11348
rect 3700 11296 3752 11348
rect 3884 11296 3936 11348
rect 5540 11296 5592 11348
rect 5816 11339 5868 11348
rect 5816 11305 5825 11339
rect 5825 11305 5859 11339
rect 5859 11305 5868 11339
rect 5816 11296 5868 11305
rect 6092 11339 6144 11348
rect 6092 11305 6101 11339
rect 6101 11305 6135 11339
rect 6135 11305 6144 11339
rect 6092 11296 6144 11305
rect 7840 11296 7892 11348
rect 8208 11296 8260 11348
rect 9312 11339 9364 11348
rect 1492 11228 1544 11280
rect 2504 11228 2556 11280
rect 3148 11228 3200 11280
rect 1768 11160 1820 11212
rect 2412 11203 2464 11212
rect 2412 11169 2421 11203
rect 2421 11169 2455 11203
rect 2455 11169 2464 11203
rect 2412 11160 2464 11169
rect 2780 11160 2832 11212
rect 3608 11228 3660 11280
rect 3608 11092 3660 11144
rect 3976 11160 4028 11212
rect 4252 11228 4304 11280
rect 4804 11271 4856 11280
rect 4804 11237 4813 11271
rect 4813 11237 4847 11271
rect 4847 11237 4856 11271
rect 4804 11228 4856 11237
rect 6368 11228 6420 11280
rect 5448 11160 5500 11212
rect 4252 11135 4304 11144
rect 4252 11101 4258 11135
rect 4258 11101 4304 11135
rect 4252 11092 4304 11101
rect 4436 11135 4488 11144
rect 4436 11101 4445 11135
rect 4445 11101 4479 11135
rect 4479 11101 4488 11135
rect 4436 11092 4488 11101
rect 6736 11228 6788 11280
rect 8024 11228 8076 11280
rect 9312 11305 9321 11339
rect 9321 11305 9355 11339
rect 9355 11305 9364 11339
rect 9312 11296 9364 11305
rect 12440 11296 12492 11348
rect 15108 11296 15160 11348
rect 16120 11296 16172 11348
rect 16304 11296 16356 11348
rect 18328 11296 18380 11348
rect 18788 11296 18840 11348
rect 19432 11339 19484 11348
rect 9404 11228 9456 11280
rect 9864 11271 9916 11280
rect 9864 11237 9873 11271
rect 9873 11237 9907 11271
rect 9907 11237 9916 11271
rect 9864 11228 9916 11237
rect 11704 11228 11756 11280
rect 12624 11228 12676 11280
rect 13360 11228 13412 11280
rect 16580 11271 16632 11280
rect 16580 11237 16589 11271
rect 16589 11237 16623 11271
rect 16623 11237 16632 11271
rect 16580 11228 16632 11237
rect 17776 11228 17828 11280
rect 18972 11228 19024 11280
rect 6644 11203 6696 11212
rect 6644 11169 6653 11203
rect 6653 11169 6687 11203
rect 6687 11169 6696 11203
rect 6644 11160 6696 11169
rect 8300 11160 8352 11212
rect 15292 11203 15344 11212
rect 15292 11169 15301 11203
rect 15301 11169 15335 11203
rect 15335 11169 15344 11203
rect 15292 11160 15344 11169
rect 2136 11024 2188 11076
rect 2688 11024 2740 11076
rect 3332 11024 3384 11076
rect 3884 10956 3936 11008
rect 7564 11024 7616 11076
rect 8484 11092 8536 11144
rect 9772 11135 9824 11144
rect 9772 11101 9781 11135
rect 9781 11101 9815 11135
rect 9815 11101 9824 11135
rect 9772 11092 9824 11101
rect 9956 11092 10008 11144
rect 11520 11092 11572 11144
rect 14004 11092 14056 11144
rect 16948 11135 17000 11144
rect 11152 11024 11204 11076
rect 13636 11024 13688 11076
rect 4344 10999 4396 11008
rect 4344 10965 4353 10999
rect 4353 10965 4387 10999
rect 4387 10965 4396 10999
rect 4344 10956 4396 10965
rect 4988 10956 5040 11008
rect 5172 10956 5224 11008
rect 7840 10999 7892 11008
rect 7840 10965 7849 10999
rect 7849 10965 7883 10999
rect 7883 10965 7892 10999
rect 7840 10956 7892 10965
rect 8852 10999 8904 11008
rect 8852 10965 8861 10999
rect 8861 10965 8895 10999
rect 8895 10965 8904 10999
rect 8852 10956 8904 10965
rect 11796 10956 11848 11008
rect 12808 10956 12860 11008
rect 13084 10956 13136 11008
rect 15384 11024 15436 11076
rect 16948 11101 16957 11135
rect 16957 11101 16991 11135
rect 16991 11101 17000 11135
rect 16948 11092 17000 11101
rect 17868 11092 17920 11144
rect 19432 11305 19441 11339
rect 19441 11305 19475 11339
rect 19475 11305 19484 11339
rect 19432 11296 19484 11305
rect 20352 11339 20404 11348
rect 20352 11305 20361 11339
rect 20361 11305 20395 11339
rect 20395 11305 20404 11339
rect 20352 11296 20404 11305
rect 22192 11296 22244 11348
rect 22836 11339 22888 11348
rect 22836 11305 22845 11339
rect 22845 11305 22879 11339
rect 22879 11305 22888 11339
rect 22836 11296 22888 11305
rect 24584 11296 24636 11348
rect 23480 11228 23532 11280
rect 19248 11160 19300 11212
rect 20076 11160 20128 11212
rect 20812 11203 20864 11212
rect 20812 11169 20821 11203
rect 20821 11169 20855 11203
rect 20855 11169 20864 11203
rect 20812 11160 20864 11169
rect 21272 11160 21324 11212
rect 24768 11160 24820 11212
rect 19616 11092 19668 11144
rect 20260 11092 20312 11144
rect 21088 11092 21140 11144
rect 22284 11092 22336 11144
rect 23664 11135 23716 11144
rect 23664 11101 23673 11135
rect 23673 11101 23707 11135
rect 23707 11101 23716 11135
rect 23664 11092 23716 11101
rect 24032 11092 24084 11144
rect 25228 11092 25280 11144
rect 20168 11024 20220 11076
rect 17592 10956 17644 11008
rect 20076 10956 20128 11008
rect 21364 10999 21416 11008
rect 21364 10965 21373 10999
rect 21373 10965 21407 10999
rect 21407 10965 21416 10999
rect 21364 10956 21416 10965
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1768 10752 1820 10804
rect 2136 10752 2188 10804
rect 2320 10752 2372 10804
rect 3056 10752 3108 10804
rect 4344 10752 4396 10804
rect 5356 10752 5408 10804
rect 6736 10752 6788 10804
rect 13636 10752 13688 10804
rect 14464 10752 14516 10804
rect 15660 10752 15712 10804
rect 17868 10795 17920 10804
rect 17868 10761 17877 10795
rect 17877 10761 17911 10795
rect 17911 10761 17920 10795
rect 17868 10752 17920 10761
rect 21732 10752 21784 10804
rect 23480 10795 23532 10804
rect 23480 10761 23489 10795
rect 23489 10761 23523 10795
rect 23523 10761 23532 10795
rect 23480 10752 23532 10761
rect 24676 10752 24728 10804
rect 25228 10795 25280 10804
rect 25228 10761 25237 10795
rect 25237 10761 25271 10795
rect 25271 10761 25280 10795
rect 25228 10752 25280 10761
rect 25596 10795 25648 10804
rect 25596 10761 25605 10795
rect 25605 10761 25639 10795
rect 25639 10761 25648 10795
rect 25596 10752 25648 10761
rect 3332 10684 3384 10736
rect 2412 10616 2464 10668
rect 3056 10616 3108 10668
rect 3700 10684 3752 10736
rect 4068 10727 4120 10736
rect 4068 10693 4077 10727
rect 4077 10693 4111 10727
rect 4111 10693 4120 10727
rect 4068 10684 4120 10693
rect 13360 10684 13412 10736
rect 20 10548 72 10600
rect 2320 10591 2372 10600
rect 2320 10557 2329 10591
rect 2329 10557 2363 10591
rect 2363 10557 2372 10591
rect 2320 10548 2372 10557
rect 3792 10591 3844 10600
rect 3792 10557 3801 10591
rect 3801 10557 3835 10591
rect 3835 10557 3844 10591
rect 3792 10548 3844 10557
rect 4988 10616 5040 10668
rect 5448 10616 5500 10668
rect 7104 10659 7156 10668
rect 7104 10625 7113 10659
rect 7113 10625 7147 10659
rect 7147 10625 7156 10659
rect 7104 10616 7156 10625
rect 7840 10616 7892 10668
rect 9128 10616 9180 10668
rect 12808 10659 12860 10668
rect 12808 10625 12817 10659
rect 12817 10625 12851 10659
rect 12851 10625 12860 10659
rect 12808 10616 12860 10625
rect 12900 10616 12952 10668
rect 14372 10659 14424 10668
rect 14372 10625 14381 10659
rect 14381 10625 14415 10659
rect 14415 10625 14424 10659
rect 14372 10616 14424 10625
rect 14924 10684 14976 10736
rect 14832 10616 14884 10668
rect 16120 10659 16172 10668
rect 16120 10625 16129 10659
rect 16129 10625 16163 10659
rect 16163 10625 16172 10659
rect 16120 10616 16172 10625
rect 5264 10548 5316 10600
rect 10140 10591 10192 10600
rect 4068 10480 4120 10532
rect 5356 10523 5408 10532
rect 5356 10489 5365 10523
rect 5365 10489 5399 10523
rect 5399 10489 5408 10523
rect 5356 10480 5408 10489
rect 6736 10480 6788 10532
rect 7196 10480 7248 10532
rect 2504 10455 2556 10464
rect 2504 10421 2513 10455
rect 2513 10421 2547 10455
rect 2547 10421 2556 10455
rect 2504 10412 2556 10421
rect 3700 10412 3752 10464
rect 3976 10412 4028 10464
rect 5632 10455 5684 10464
rect 5632 10421 5641 10455
rect 5641 10421 5675 10455
rect 5675 10421 5684 10455
rect 5632 10412 5684 10421
rect 8300 10412 8352 10464
rect 10140 10557 10149 10591
rect 10149 10557 10183 10591
rect 10183 10557 10192 10591
rect 10140 10548 10192 10557
rect 8760 10480 8812 10532
rect 8852 10412 8904 10464
rect 11704 10480 11756 10532
rect 15292 10548 15344 10600
rect 17960 10548 18012 10600
rect 19248 10591 19300 10600
rect 19248 10557 19257 10591
rect 19257 10557 19291 10591
rect 19291 10557 19300 10591
rect 19248 10548 19300 10557
rect 19616 10591 19668 10600
rect 19616 10557 19625 10591
rect 19625 10557 19659 10591
rect 19659 10557 19668 10591
rect 19616 10548 19668 10557
rect 21364 10616 21416 10668
rect 21456 10548 21508 10600
rect 22836 10548 22888 10600
rect 24584 10548 24636 10600
rect 25596 10548 25648 10600
rect 12624 10480 12676 10532
rect 13452 10523 13504 10532
rect 12440 10412 12492 10464
rect 13452 10489 13461 10523
rect 13461 10489 13495 10523
rect 13495 10489 13504 10523
rect 13452 10480 13504 10489
rect 14464 10523 14516 10532
rect 14464 10489 14473 10523
rect 14473 10489 14507 10523
rect 14507 10489 14516 10523
rect 14464 10480 14516 10489
rect 15660 10480 15712 10532
rect 17224 10480 17276 10532
rect 19432 10480 19484 10532
rect 22192 10480 22244 10532
rect 23480 10480 23532 10532
rect 23756 10480 23808 10532
rect 14740 10412 14792 10464
rect 16580 10412 16632 10464
rect 18512 10412 18564 10464
rect 20812 10412 20864 10464
rect 21732 10412 21784 10464
rect 22284 10455 22336 10464
rect 22284 10421 22293 10455
rect 22293 10421 22327 10455
rect 22327 10421 22336 10455
rect 22284 10412 22336 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2320 10208 2372 10260
rect 4712 10251 4764 10260
rect 1952 10072 2004 10124
rect 3976 10140 4028 10192
rect 4712 10217 4721 10251
rect 4721 10217 4755 10251
rect 4755 10217 4764 10251
rect 4712 10208 4764 10217
rect 5540 10208 5592 10260
rect 7196 10208 7248 10260
rect 9864 10251 9916 10260
rect 9864 10217 9873 10251
rect 9873 10217 9907 10251
rect 9907 10217 9916 10251
rect 9864 10208 9916 10217
rect 10140 10208 10192 10260
rect 11152 10251 11204 10260
rect 11152 10217 11161 10251
rect 11161 10217 11195 10251
rect 11195 10217 11204 10251
rect 11152 10208 11204 10217
rect 11520 10251 11572 10260
rect 11520 10217 11529 10251
rect 11529 10217 11563 10251
rect 11563 10217 11572 10251
rect 11520 10208 11572 10217
rect 12808 10208 12860 10260
rect 14004 10251 14056 10260
rect 14004 10217 14013 10251
rect 14013 10217 14047 10251
rect 14047 10217 14056 10251
rect 14004 10208 14056 10217
rect 14924 10208 14976 10260
rect 18328 10208 18380 10260
rect 19524 10208 19576 10260
rect 23756 10251 23808 10260
rect 23756 10217 23765 10251
rect 23765 10217 23799 10251
rect 23799 10217 23808 10251
rect 23756 10208 23808 10217
rect 24584 10251 24636 10260
rect 24584 10217 24593 10251
rect 24593 10217 24627 10251
rect 24627 10217 24636 10251
rect 24584 10208 24636 10217
rect 5448 10140 5500 10192
rect 7104 10183 7156 10192
rect 7104 10149 7113 10183
rect 7113 10149 7147 10183
rect 7147 10149 7156 10183
rect 7104 10140 7156 10149
rect 10048 10140 10100 10192
rect 4068 10115 4120 10124
rect 4068 10081 4077 10115
rect 4077 10081 4111 10115
rect 4111 10081 4120 10115
rect 4068 10072 4120 10081
rect 6000 10072 6052 10124
rect 6368 10115 6420 10124
rect 6368 10081 6377 10115
rect 6377 10081 6411 10115
rect 6411 10081 6420 10115
rect 6368 10072 6420 10081
rect 6460 10072 6512 10124
rect 7196 10072 7248 10124
rect 8024 10072 8076 10124
rect 10692 10115 10744 10124
rect 3792 10004 3844 10056
rect 4160 10004 4212 10056
rect 4436 10047 4488 10056
rect 4436 10013 4445 10047
rect 4445 10013 4479 10047
rect 4479 10013 4488 10047
rect 4436 10004 4488 10013
rect 7840 10004 7892 10056
rect 10692 10081 10701 10115
rect 10701 10081 10735 10115
rect 10735 10081 10744 10115
rect 12624 10183 12676 10192
rect 12624 10149 12633 10183
rect 12633 10149 12667 10183
rect 12667 10149 12676 10183
rect 12624 10140 12676 10149
rect 13636 10140 13688 10192
rect 14372 10183 14424 10192
rect 14372 10149 14381 10183
rect 14381 10149 14415 10183
rect 14415 10149 14424 10183
rect 14372 10140 14424 10149
rect 16120 10183 16172 10192
rect 16120 10149 16129 10183
rect 16129 10149 16163 10183
rect 16163 10149 16172 10183
rect 16120 10140 16172 10149
rect 16580 10140 16632 10192
rect 18512 10183 18564 10192
rect 18512 10149 18521 10183
rect 18521 10149 18555 10183
rect 18555 10149 18564 10183
rect 18512 10140 18564 10149
rect 18604 10183 18656 10192
rect 18604 10149 18613 10183
rect 18613 10149 18647 10183
rect 18647 10149 18656 10183
rect 21088 10183 21140 10192
rect 18604 10140 18656 10149
rect 21088 10149 21097 10183
rect 21097 10149 21131 10183
rect 21131 10149 21140 10183
rect 21088 10140 21140 10149
rect 23664 10140 23716 10192
rect 11704 10115 11756 10124
rect 10692 10072 10744 10081
rect 11704 10081 11713 10115
rect 11713 10081 11747 10115
rect 11747 10081 11756 10115
rect 11704 10072 11756 10081
rect 15568 10072 15620 10124
rect 16028 10072 16080 10124
rect 22744 10115 22796 10124
rect 22744 10081 22753 10115
rect 22753 10081 22787 10115
rect 22787 10081 22796 10115
rect 22744 10072 22796 10081
rect 23204 10115 23256 10124
rect 23204 10081 23213 10115
rect 23213 10081 23247 10115
rect 23247 10081 23256 10115
rect 23204 10072 23256 10081
rect 23388 10072 23440 10124
rect 8392 10047 8444 10056
rect 8392 10013 8401 10047
rect 8401 10013 8435 10047
rect 8435 10013 8444 10047
rect 8392 10004 8444 10013
rect 13268 10004 13320 10056
rect 14280 10004 14332 10056
rect 16948 10004 17000 10056
rect 18880 10047 18932 10056
rect 18880 10013 18889 10047
rect 18889 10013 18923 10047
rect 18923 10013 18932 10047
rect 18880 10004 18932 10013
rect 21180 10004 21232 10056
rect 1860 9868 1912 9920
rect 3148 9868 3200 9920
rect 5356 9979 5408 9988
rect 5356 9945 5365 9979
rect 5365 9945 5399 9979
rect 5399 9945 5408 9979
rect 5356 9936 5408 9945
rect 4252 9911 4304 9920
rect 4252 9877 4276 9911
rect 4276 9877 4304 9911
rect 4252 9868 4304 9877
rect 8208 9936 8260 9988
rect 11888 9979 11940 9988
rect 11888 9945 11897 9979
rect 11897 9945 11931 9979
rect 11931 9945 11940 9979
rect 11888 9936 11940 9945
rect 8484 9868 8536 9920
rect 12992 9868 13044 9920
rect 16488 9936 16540 9988
rect 21916 10004 21968 10056
rect 23572 10004 23624 10056
rect 25044 10004 25096 10056
rect 19248 9868 19300 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 1860 9596 1912 9648
rect 2412 9639 2464 9648
rect 2412 9605 2421 9639
rect 2421 9605 2455 9639
rect 2455 9605 2464 9639
rect 2412 9596 2464 9605
rect 112 9528 164 9580
rect 2688 9664 2740 9716
rect 4160 9664 4212 9716
rect 10048 9664 10100 9716
rect 11428 9664 11480 9716
rect 13636 9707 13688 9716
rect 1952 9460 2004 9512
rect 2136 9503 2188 9512
rect 2136 9469 2145 9503
rect 2145 9469 2179 9503
rect 2179 9469 2188 9503
rect 2136 9460 2188 9469
rect 2596 9528 2648 9580
rect 4068 9571 4120 9580
rect 4068 9537 4077 9571
rect 4077 9537 4111 9571
rect 4111 9537 4120 9571
rect 4068 9528 4120 9537
rect 3976 9460 4028 9512
rect 4252 9596 4304 9648
rect 9588 9596 9640 9648
rect 10692 9596 10744 9648
rect 11704 9596 11756 9648
rect 4620 9528 4672 9580
rect 6736 9528 6788 9580
rect 7380 9571 7432 9580
rect 4344 9460 4396 9512
rect 5080 9460 5132 9512
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 7564 9528 7616 9580
rect 8300 9528 8352 9580
rect 13636 9673 13645 9707
rect 13645 9673 13679 9707
rect 13679 9673 13688 9707
rect 13636 9664 13688 9673
rect 15660 9664 15712 9716
rect 18236 9664 18288 9716
rect 19524 9664 19576 9716
rect 13360 9596 13412 9648
rect 12992 9571 13044 9580
rect 12992 9537 13001 9571
rect 13001 9537 13035 9571
rect 13035 9537 13044 9571
rect 12992 9528 13044 9537
rect 18880 9596 18932 9648
rect 21916 9664 21968 9716
rect 22744 9707 22796 9716
rect 22744 9673 22753 9707
rect 22753 9673 22787 9707
rect 22787 9673 22796 9707
rect 22744 9664 22796 9673
rect 25044 9707 25096 9716
rect 25044 9673 25053 9707
rect 25053 9673 25087 9707
rect 25087 9673 25096 9707
rect 25044 9664 25096 9673
rect 25412 9707 25464 9716
rect 25412 9673 25421 9707
rect 25421 9673 25455 9707
rect 25455 9673 25464 9707
rect 25412 9664 25464 9673
rect 23204 9596 23256 9648
rect 14556 9528 14608 9580
rect 14740 9571 14792 9580
rect 14740 9537 14749 9571
rect 14749 9537 14783 9571
rect 14783 9537 14792 9571
rect 14740 9528 14792 9537
rect 15476 9528 15528 9580
rect 18328 9571 18380 9580
rect 18328 9537 18337 9571
rect 18337 9537 18371 9571
rect 18371 9537 18380 9571
rect 18328 9528 18380 9537
rect 20076 9571 20128 9580
rect 20076 9537 20085 9571
rect 20085 9537 20119 9571
rect 20119 9537 20128 9571
rect 20076 9528 20128 9537
rect 20352 9571 20404 9580
rect 20352 9537 20361 9571
rect 20361 9537 20395 9571
rect 20395 9537 20404 9571
rect 20352 9528 20404 9537
rect 22284 9571 22336 9580
rect 22284 9537 22293 9571
rect 22293 9537 22327 9571
rect 22327 9537 22336 9571
rect 22284 9528 22336 9537
rect 22928 9528 22980 9580
rect 7196 9460 7248 9512
rect 8208 9460 8260 9512
rect 8484 9503 8536 9512
rect 8484 9469 8493 9503
rect 8493 9469 8527 9503
rect 8527 9469 8536 9503
rect 8484 9460 8536 9469
rect 11244 9503 11296 9512
rect 2044 9324 2096 9376
rect 3424 9324 3476 9376
rect 3700 9435 3752 9444
rect 3700 9401 3709 9435
rect 3709 9401 3743 9435
rect 3743 9401 3752 9435
rect 3700 9392 3752 9401
rect 8300 9392 8352 9444
rect 11244 9469 11253 9503
rect 11253 9469 11287 9503
rect 11287 9469 11296 9503
rect 11244 9460 11296 9469
rect 15292 9460 15344 9512
rect 16856 9503 16908 9512
rect 16856 9469 16865 9503
rect 16865 9469 16899 9503
rect 16899 9469 16908 9503
rect 16856 9460 16908 9469
rect 21548 9503 21600 9512
rect 11520 9435 11572 9444
rect 11520 9401 11529 9435
rect 11529 9401 11563 9435
rect 11563 9401 11572 9435
rect 11520 9392 11572 9401
rect 15568 9435 15620 9444
rect 6368 9324 6420 9376
rect 7748 9324 7800 9376
rect 8024 9367 8076 9376
rect 8024 9333 8033 9367
rect 8033 9333 8067 9367
rect 8067 9333 8076 9367
rect 8024 9324 8076 9333
rect 10784 9324 10836 9376
rect 12624 9324 12676 9376
rect 14004 9367 14056 9376
rect 14004 9333 14013 9367
rect 14013 9333 14047 9367
rect 14047 9333 14056 9367
rect 15568 9401 15577 9435
rect 15577 9401 15611 9435
rect 15611 9401 15620 9435
rect 15568 9392 15620 9401
rect 16488 9392 16540 9444
rect 17776 9392 17828 9444
rect 17960 9392 18012 9444
rect 18972 9435 19024 9444
rect 18972 9401 18981 9435
rect 18981 9401 19015 9435
rect 19015 9401 19024 9435
rect 18972 9392 19024 9401
rect 21548 9469 21557 9503
rect 21557 9469 21591 9503
rect 21591 9469 21600 9503
rect 21548 9460 21600 9469
rect 22744 9460 22796 9512
rect 22836 9460 22888 9512
rect 24124 9503 24176 9512
rect 24124 9469 24133 9503
rect 24133 9469 24167 9503
rect 24167 9469 24176 9503
rect 24124 9460 24176 9469
rect 25136 9460 25188 9512
rect 23480 9392 23532 9444
rect 14004 9324 14056 9333
rect 18604 9324 18656 9376
rect 19984 9324 20036 9376
rect 21364 9367 21416 9376
rect 21364 9333 21373 9367
rect 21373 9333 21407 9367
rect 21407 9333 21416 9367
rect 21364 9324 21416 9333
rect 23664 9324 23716 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2412 9120 2464 9172
rect 3424 9120 3476 9172
rect 3700 9120 3752 9172
rect 6000 9120 6052 9172
rect 6460 9120 6512 9172
rect 6736 9120 6788 9172
rect 7012 9120 7064 9172
rect 9772 9120 9824 9172
rect 13268 9120 13320 9172
rect 14004 9120 14056 9172
rect 14556 9163 14608 9172
rect 14556 9129 14565 9163
rect 14565 9129 14599 9163
rect 14599 9129 14608 9163
rect 14556 9120 14608 9129
rect 16580 9163 16632 9172
rect 16580 9129 16589 9163
rect 16589 9129 16623 9163
rect 16623 9129 16632 9163
rect 16580 9120 16632 9129
rect 17960 9163 18012 9172
rect 17960 9129 17969 9163
rect 17969 9129 18003 9163
rect 18003 9129 18012 9163
rect 17960 9120 18012 9129
rect 18512 9120 18564 9172
rect 21088 9163 21140 9172
rect 21088 9129 21097 9163
rect 21097 9129 21131 9163
rect 21131 9129 21140 9163
rect 21088 9120 21140 9129
rect 22744 9163 22796 9172
rect 22744 9129 22753 9163
rect 22753 9129 22787 9163
rect 22787 9129 22796 9163
rect 22744 9120 22796 9129
rect 23112 9163 23164 9172
rect 23112 9129 23121 9163
rect 23121 9129 23155 9163
rect 23155 9129 23164 9163
rect 23112 9120 23164 9129
rect 24124 9163 24176 9172
rect 24124 9129 24133 9163
rect 24133 9129 24167 9163
rect 24167 9129 24176 9163
rect 24124 9120 24176 9129
rect 3884 9052 3936 9104
rect 4344 9052 4396 9104
rect 2044 8984 2096 9036
rect 2504 8984 2556 9036
rect 6460 9027 6512 9036
rect 6460 8993 6469 9027
rect 6469 8993 6503 9027
rect 6503 8993 6512 9027
rect 6460 8984 6512 8993
rect 6736 9027 6788 9036
rect 6736 8993 6745 9027
rect 6745 8993 6779 9027
rect 6779 8993 6788 9027
rect 6736 8984 6788 8993
rect 8116 8984 8168 9036
rect 8300 9027 8352 9036
rect 8300 8993 8309 9027
rect 8309 8993 8343 9027
rect 8343 8993 8352 9027
rect 8300 8984 8352 8993
rect 9864 9027 9916 9036
rect 9864 8993 9873 9027
rect 9873 8993 9907 9027
rect 9907 8993 9916 9027
rect 9864 8984 9916 8993
rect 10968 9052 11020 9104
rect 12440 9095 12492 9104
rect 12440 9061 12449 9095
rect 12449 9061 12483 9095
rect 12483 9061 12492 9095
rect 12440 9052 12492 9061
rect 13452 9052 13504 9104
rect 14280 9052 14332 9104
rect 17224 9052 17276 9104
rect 19156 9052 19208 9104
rect 20076 9095 20128 9104
rect 20076 9061 20085 9095
rect 20085 9061 20119 9095
rect 20119 9061 20128 9095
rect 20076 9052 20128 9061
rect 21180 9052 21232 9104
rect 21640 9095 21692 9104
rect 21640 9061 21649 9095
rect 21649 9061 21683 9095
rect 21683 9061 21692 9095
rect 21640 9052 21692 9061
rect 23296 9052 23348 9104
rect 3792 8916 3844 8968
rect 3884 8959 3936 8968
rect 3884 8925 3893 8959
rect 3893 8925 3927 8959
rect 3927 8925 3936 8959
rect 4436 8959 4488 8968
rect 3884 8916 3936 8925
rect 4436 8925 4445 8959
rect 4445 8925 4479 8959
rect 4479 8925 4488 8959
rect 4436 8916 4488 8925
rect 6920 8959 6972 8968
rect 6920 8925 6929 8959
rect 6929 8925 6963 8959
rect 6963 8925 6972 8959
rect 6920 8916 6972 8925
rect 9680 8916 9732 8968
rect 11704 8984 11756 9036
rect 15660 9027 15712 9036
rect 15660 8993 15669 9027
rect 15669 8993 15703 9027
rect 15703 8993 15712 9027
rect 15660 8984 15712 8993
rect 15844 8984 15896 9036
rect 17776 8984 17828 9036
rect 18788 9027 18840 9036
rect 18788 8993 18797 9027
rect 18797 8993 18831 9027
rect 18831 8993 18840 9027
rect 18788 8984 18840 8993
rect 19984 8984 20036 9036
rect 22928 8984 22980 9036
rect 23480 9027 23532 9036
rect 23480 8993 23489 9027
rect 23489 8993 23523 9027
rect 23523 8993 23532 9027
rect 23480 8984 23532 8993
rect 24860 8984 24912 9036
rect 11520 8916 11572 8968
rect 13544 8916 13596 8968
rect 16212 8959 16264 8968
rect 16212 8925 16221 8959
rect 16221 8925 16255 8959
rect 16255 8925 16264 8959
rect 16212 8916 16264 8925
rect 17040 8959 17092 8968
rect 17040 8925 17049 8959
rect 17049 8925 17083 8959
rect 17083 8925 17092 8959
rect 17040 8916 17092 8925
rect 20352 8916 20404 8968
rect 3424 8848 3476 8900
rect 4160 8848 4212 8900
rect 6368 8848 6420 8900
rect 8116 8891 8168 8900
rect 1676 8780 1728 8832
rect 1860 8780 1912 8832
rect 4068 8780 4120 8832
rect 4344 8823 4396 8832
rect 4344 8789 4353 8823
rect 4353 8789 4387 8823
rect 4387 8789 4396 8823
rect 4344 8780 4396 8789
rect 4528 8823 4580 8832
rect 4528 8789 4537 8823
rect 4537 8789 4571 8823
rect 4571 8789 4580 8823
rect 4528 8780 4580 8789
rect 7840 8823 7892 8832
rect 7840 8789 7849 8823
rect 7849 8789 7883 8823
rect 7883 8789 7892 8823
rect 7840 8780 7892 8789
rect 8116 8857 8125 8891
rect 8125 8857 8159 8891
rect 8159 8857 8168 8891
rect 8116 8848 8168 8857
rect 12900 8848 12952 8900
rect 16948 8891 17000 8900
rect 16948 8857 16957 8891
rect 16957 8857 16991 8891
rect 16991 8857 17000 8891
rect 16948 8848 17000 8857
rect 8484 8780 8536 8832
rect 11796 8823 11848 8832
rect 11796 8789 11805 8823
rect 11805 8789 11839 8823
rect 11839 8789 11848 8823
rect 11796 8780 11848 8789
rect 18328 8823 18380 8832
rect 18328 8789 18337 8823
rect 18337 8789 18371 8823
rect 18371 8789 18380 8823
rect 18328 8780 18380 8789
rect 21180 8848 21232 8900
rect 22744 8916 22796 8968
rect 23572 8916 23624 8968
rect 21272 8780 21324 8832
rect 22468 8848 22520 8900
rect 23020 8848 23072 8900
rect 23940 8780 23992 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2136 8576 2188 8628
rect 3148 8619 3200 8628
rect 3148 8585 3157 8619
rect 3157 8585 3191 8619
rect 3191 8585 3200 8619
rect 3148 8576 3200 8585
rect 4344 8576 4396 8628
rect 5448 8576 5500 8628
rect 6736 8576 6788 8628
rect 7196 8576 7248 8628
rect 8300 8576 8352 8628
rect 10968 8576 11020 8628
rect 12440 8576 12492 8628
rect 17224 8619 17276 8628
rect 17224 8585 17233 8619
rect 17233 8585 17267 8619
rect 17267 8585 17276 8619
rect 17224 8576 17276 8585
rect 19156 8619 19208 8628
rect 19156 8585 19165 8619
rect 19165 8585 19199 8619
rect 19199 8585 19208 8619
rect 19156 8576 19208 8585
rect 19984 8576 20036 8628
rect 21640 8576 21692 8628
rect 3884 8508 3936 8560
rect 4160 8508 4212 8560
rect 7656 8508 7708 8560
rect 12992 8508 13044 8560
rect 14464 8508 14516 8560
rect 16120 8551 16172 8560
rect 16120 8517 16129 8551
rect 16129 8517 16163 8551
rect 16163 8517 16172 8551
rect 16120 8508 16172 8517
rect 4712 8440 4764 8492
rect 14280 8483 14332 8492
rect 14280 8449 14289 8483
rect 14289 8449 14323 8483
rect 14323 8449 14332 8483
rect 14280 8440 14332 8449
rect 14556 8483 14608 8492
rect 14556 8449 14565 8483
rect 14565 8449 14599 8483
rect 14599 8449 14608 8483
rect 14556 8440 14608 8449
rect 14740 8440 14792 8492
rect 1492 8415 1544 8424
rect 1492 8381 1501 8415
rect 1501 8381 1535 8415
rect 1535 8381 1544 8415
rect 1492 8372 1544 8381
rect 5724 8415 5776 8424
rect 1952 8236 2004 8288
rect 2596 8236 2648 8288
rect 2872 8279 2924 8288
rect 2872 8245 2881 8279
rect 2881 8245 2915 8279
rect 2915 8245 2924 8279
rect 2872 8236 2924 8245
rect 5724 8381 5733 8415
rect 5733 8381 5767 8415
rect 5767 8381 5776 8415
rect 5724 8372 5776 8381
rect 7380 8415 7432 8424
rect 7380 8381 7389 8415
rect 7389 8381 7423 8415
rect 7423 8381 7432 8415
rect 7380 8372 7432 8381
rect 8116 8372 8168 8424
rect 8668 8372 8720 8424
rect 4344 8347 4396 8356
rect 4344 8313 4353 8347
rect 4353 8313 4387 8347
rect 4387 8313 4396 8347
rect 4896 8347 4948 8356
rect 4344 8304 4396 8313
rect 4896 8313 4905 8347
rect 4905 8313 4939 8347
rect 4939 8313 4948 8347
rect 4896 8304 4948 8313
rect 6368 8304 6420 8356
rect 9588 8372 9640 8424
rect 17684 8508 17736 8560
rect 18972 8508 19024 8560
rect 17040 8440 17092 8492
rect 18880 8483 18932 8492
rect 18880 8449 18889 8483
rect 18889 8449 18923 8483
rect 18923 8449 18932 8483
rect 18880 8440 18932 8449
rect 20076 8440 20128 8492
rect 23112 8576 23164 8628
rect 25412 8619 25464 8628
rect 25412 8585 25421 8619
rect 25421 8585 25455 8619
rect 25455 8585 25464 8619
rect 25412 8576 25464 8585
rect 23388 8551 23440 8560
rect 23388 8517 23397 8551
rect 23397 8517 23431 8551
rect 23431 8517 23440 8551
rect 23388 8508 23440 8517
rect 23940 8440 23992 8492
rect 9864 8304 9916 8356
rect 10692 8304 10744 8356
rect 10876 8347 10928 8356
rect 10876 8313 10885 8347
rect 10885 8313 10919 8347
rect 10919 8313 10928 8347
rect 10876 8304 10928 8313
rect 11796 8347 11848 8356
rect 11796 8313 11805 8347
rect 11805 8313 11839 8347
rect 11839 8313 11848 8347
rect 11796 8304 11848 8313
rect 12440 8304 12492 8356
rect 3884 8236 3936 8288
rect 6460 8236 6512 8288
rect 8024 8236 8076 8288
rect 9220 8236 9272 8288
rect 16580 8372 16632 8424
rect 16856 8372 16908 8424
rect 22376 8372 22428 8424
rect 23112 8372 23164 8424
rect 25228 8415 25280 8424
rect 25228 8381 25237 8415
rect 25237 8381 25271 8415
rect 25271 8381 25280 8415
rect 25228 8372 25280 8381
rect 17408 8304 17460 8356
rect 18328 8347 18380 8356
rect 18328 8313 18337 8347
rect 18337 8313 18371 8347
rect 18371 8313 18380 8347
rect 18328 8304 18380 8313
rect 19984 8304 20036 8356
rect 15660 8236 15712 8288
rect 15936 8236 15988 8288
rect 19156 8236 19208 8288
rect 20996 8236 21048 8288
rect 22744 8304 22796 8356
rect 21364 8236 21416 8288
rect 22928 8236 22980 8288
rect 23388 8236 23440 8288
rect 23480 8236 23532 8288
rect 23848 8347 23900 8356
rect 23848 8313 23857 8347
rect 23857 8313 23891 8347
rect 23891 8313 23900 8347
rect 23848 8304 23900 8313
rect 24124 8236 24176 8288
rect 24860 8236 24912 8288
rect 25412 8236 25464 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1860 8032 1912 8084
rect 2044 8032 2096 8084
rect 3148 8032 3200 8084
rect 3516 8075 3568 8084
rect 3516 8041 3525 8075
rect 3525 8041 3559 8075
rect 3559 8041 3568 8075
rect 3516 8032 3568 8041
rect 4068 8032 4120 8084
rect 5724 8075 5776 8084
rect 3608 7964 3660 8016
rect 5724 8041 5733 8075
rect 5733 8041 5767 8075
rect 5767 8041 5776 8075
rect 5724 8032 5776 8041
rect 4436 7964 4488 8016
rect 6092 7964 6144 8016
rect 8208 8032 8260 8084
rect 9588 8032 9640 8084
rect 13544 8075 13596 8084
rect 13544 8041 13553 8075
rect 13553 8041 13587 8075
rect 13587 8041 13596 8075
rect 13544 8032 13596 8041
rect 15568 8075 15620 8084
rect 15568 8041 15577 8075
rect 15577 8041 15611 8075
rect 15611 8041 15620 8075
rect 15568 8032 15620 8041
rect 17408 8032 17460 8084
rect 18328 8075 18380 8084
rect 18328 8041 18337 8075
rect 18337 8041 18371 8075
rect 18371 8041 18380 8075
rect 18328 8032 18380 8041
rect 1952 7896 2004 7948
rect 2688 7939 2740 7948
rect 2688 7905 2697 7939
rect 2697 7905 2731 7939
rect 2731 7905 2740 7939
rect 2688 7896 2740 7905
rect 2964 7939 3016 7948
rect 2964 7905 2973 7939
rect 2973 7905 3007 7939
rect 3007 7905 3016 7939
rect 2964 7896 3016 7905
rect 3424 7896 3476 7948
rect 6368 7896 6420 7948
rect 9864 7964 9916 8016
rect 10692 7964 10744 8016
rect 6736 7939 6788 7948
rect 6736 7905 6745 7939
rect 6745 7905 6779 7939
rect 6779 7905 6788 7939
rect 6736 7896 6788 7905
rect 7840 7896 7892 7948
rect 8024 7939 8076 7948
rect 8024 7905 8033 7939
rect 8033 7905 8067 7939
rect 8067 7905 8076 7939
rect 8024 7896 8076 7905
rect 8300 7939 8352 7948
rect 8300 7905 8309 7939
rect 8309 7905 8343 7939
rect 8343 7905 8352 7939
rect 8300 7896 8352 7905
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 10600 7896 10652 7948
rect 11244 7939 11296 7948
rect 11244 7905 11253 7939
rect 11253 7905 11287 7939
rect 11287 7905 11296 7939
rect 11244 7896 11296 7905
rect 12440 7964 12492 8016
rect 12992 7964 13044 8016
rect 13452 7964 13504 8016
rect 17224 7964 17276 8016
rect 18788 8007 18840 8016
rect 18788 7973 18797 8007
rect 18797 7973 18831 8007
rect 18831 7973 18840 8007
rect 18788 7964 18840 7973
rect 20352 8032 20404 8084
rect 19432 7964 19484 8016
rect 21088 8007 21140 8016
rect 21088 7973 21097 8007
rect 21097 7973 21131 8007
rect 21131 7973 21140 8007
rect 21088 7964 21140 7973
rect 24032 8032 24084 8084
rect 22744 7964 22796 8016
rect 14096 7939 14148 7948
rect 14096 7905 14105 7939
rect 14105 7905 14139 7939
rect 14139 7905 14148 7939
rect 14096 7896 14148 7905
rect 3516 7828 3568 7880
rect 4160 7828 4212 7880
rect 4436 7828 4488 7880
rect 12164 7828 12216 7880
rect 16396 7896 16448 7948
rect 23848 7896 23900 7948
rect 24676 7896 24728 7948
rect 16120 7828 16172 7880
rect 17408 7871 17460 7880
rect 17408 7837 17417 7871
rect 17417 7837 17451 7871
rect 17451 7837 17460 7871
rect 17408 7828 17460 7837
rect 19340 7828 19392 7880
rect 848 7760 900 7812
rect 1492 7760 1544 7812
rect 3700 7760 3752 7812
rect 6368 7760 6420 7812
rect 7380 7760 7432 7812
rect 8208 7760 8260 7812
rect 9772 7760 9824 7812
rect 10876 7760 10928 7812
rect 12256 7760 12308 7812
rect 15844 7760 15896 7812
rect 16488 7760 16540 7812
rect 18788 7760 18840 7812
rect 18972 7760 19024 7812
rect 20720 7828 20772 7880
rect 3976 7692 4028 7744
rect 4344 7692 4396 7744
rect 7748 7692 7800 7744
rect 9956 7692 10008 7744
rect 13268 7735 13320 7744
rect 13268 7701 13277 7735
rect 13277 7701 13311 7735
rect 13311 7701 13320 7735
rect 13268 7692 13320 7701
rect 13544 7692 13596 7744
rect 16580 7692 16632 7744
rect 20076 7692 20128 7744
rect 22008 7735 22060 7744
rect 22008 7701 22017 7735
rect 22017 7701 22051 7735
rect 22051 7701 22060 7735
rect 22008 7692 22060 7701
rect 23756 7692 23808 7744
rect 24124 7692 24176 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 1584 7531 1636 7540
rect 1584 7497 1593 7531
rect 1593 7497 1627 7531
rect 1627 7497 1636 7531
rect 1584 7488 1636 7497
rect 1952 7531 2004 7540
rect 1952 7497 1961 7531
rect 1961 7497 1995 7531
rect 1995 7497 2004 7531
rect 1952 7488 2004 7497
rect 4068 7488 4120 7540
rect 7196 7531 7248 7540
rect 7196 7497 7205 7531
rect 7205 7497 7239 7531
rect 7239 7497 7248 7531
rect 7196 7488 7248 7497
rect 7288 7488 7340 7540
rect 9680 7531 9732 7540
rect 9680 7497 9689 7531
rect 9689 7497 9723 7531
rect 9723 7497 9732 7531
rect 9680 7488 9732 7497
rect 12164 7531 12216 7540
rect 12164 7497 12173 7531
rect 12173 7497 12207 7531
rect 12207 7497 12216 7531
rect 12164 7488 12216 7497
rect 12440 7488 12492 7540
rect 13268 7531 13320 7540
rect 13268 7497 13277 7531
rect 13277 7497 13311 7531
rect 13311 7497 13320 7531
rect 13268 7488 13320 7497
rect 14096 7488 14148 7540
rect 16120 7488 16172 7540
rect 16396 7531 16448 7540
rect 16396 7497 16405 7531
rect 16405 7497 16439 7531
rect 16439 7497 16448 7531
rect 16396 7488 16448 7497
rect 17500 7488 17552 7540
rect 19432 7531 19484 7540
rect 19432 7497 19441 7531
rect 19441 7497 19475 7531
rect 19475 7497 19484 7531
rect 19432 7488 19484 7497
rect 21088 7488 21140 7540
rect 22744 7488 22796 7540
rect 2688 7420 2740 7472
rect 5356 7420 5408 7472
rect 3700 7352 3752 7404
rect 5448 7352 5500 7404
rect 1124 7284 1176 7336
rect 3148 7327 3200 7336
rect 1768 7216 1820 7268
rect 3148 7293 3157 7327
rect 3157 7293 3191 7327
rect 3191 7293 3200 7327
rect 3148 7284 3200 7293
rect 4252 7327 4304 7336
rect 4252 7293 4261 7327
rect 4261 7293 4295 7327
rect 4295 7293 4304 7327
rect 4252 7284 4304 7293
rect 4804 7284 4856 7336
rect 8392 7420 8444 7472
rect 12900 7420 12952 7472
rect 8208 7352 8260 7404
rect 7564 7284 7616 7336
rect 8024 7284 8076 7336
rect 8300 7327 8352 7336
rect 8300 7293 8309 7327
rect 8309 7293 8343 7327
rect 8343 7293 8352 7327
rect 8300 7284 8352 7293
rect 9404 7352 9456 7404
rect 9956 7352 10008 7404
rect 10600 7395 10652 7404
rect 10600 7361 10609 7395
rect 10609 7361 10643 7395
rect 10643 7361 10652 7395
rect 10600 7352 10652 7361
rect 13452 7395 13504 7404
rect 13452 7361 13461 7395
rect 13461 7361 13495 7395
rect 13495 7361 13504 7395
rect 13452 7352 13504 7361
rect 10784 7327 10836 7336
rect 3332 7216 3384 7268
rect 2136 7148 2188 7200
rect 2964 7148 3016 7200
rect 6276 7216 6328 7268
rect 7840 7216 7892 7268
rect 9036 7259 9088 7268
rect 9036 7225 9045 7259
rect 9045 7225 9079 7259
rect 9079 7225 9088 7259
rect 9036 7216 9088 7225
rect 4068 7191 4120 7200
rect 4068 7157 4077 7191
rect 4077 7157 4111 7191
rect 4111 7157 4120 7191
rect 4068 7148 4120 7157
rect 4436 7191 4488 7200
rect 4436 7157 4445 7191
rect 4445 7157 4479 7191
rect 4479 7157 4488 7191
rect 4436 7148 4488 7157
rect 4712 7148 4764 7200
rect 6368 7148 6420 7200
rect 8024 7148 8076 7200
rect 10784 7293 10793 7327
rect 10793 7293 10827 7327
rect 10827 7293 10836 7327
rect 10784 7284 10836 7293
rect 11060 7284 11112 7336
rect 15016 7352 15068 7404
rect 18236 7420 18288 7472
rect 21272 7420 21324 7472
rect 15292 7284 15344 7336
rect 17224 7352 17276 7404
rect 18972 7352 19024 7404
rect 20260 7352 20312 7404
rect 11520 7259 11572 7268
rect 11520 7225 11529 7259
rect 11529 7225 11563 7259
rect 11563 7225 11572 7259
rect 11520 7216 11572 7225
rect 14096 7259 14148 7268
rect 13268 7148 13320 7200
rect 14096 7225 14105 7259
rect 14105 7225 14139 7259
rect 14139 7225 14148 7259
rect 14096 7216 14148 7225
rect 14556 7216 14608 7268
rect 13728 7148 13780 7200
rect 21824 7284 21876 7336
rect 23572 7352 23624 7404
rect 22100 7284 22152 7336
rect 23848 7284 23900 7336
rect 25044 7284 25096 7336
rect 15660 7259 15712 7268
rect 15660 7225 15669 7259
rect 15669 7225 15703 7259
rect 15703 7225 15712 7259
rect 15660 7216 15712 7225
rect 18144 7259 18196 7268
rect 18144 7225 18153 7259
rect 18153 7225 18187 7259
rect 18187 7225 18196 7259
rect 18144 7216 18196 7225
rect 18236 7259 18288 7268
rect 18236 7225 18245 7259
rect 18245 7225 18279 7259
rect 18279 7225 18288 7259
rect 18236 7216 18288 7225
rect 20628 7259 20680 7268
rect 20628 7225 20637 7259
rect 20637 7225 20671 7259
rect 20671 7225 20680 7259
rect 21180 7259 21232 7268
rect 20628 7216 20680 7225
rect 21180 7225 21189 7259
rect 21189 7225 21223 7259
rect 21223 7225 21232 7259
rect 21180 7216 21232 7225
rect 22652 7216 22704 7268
rect 23388 7216 23440 7268
rect 19432 7148 19484 7200
rect 21824 7191 21876 7200
rect 21824 7157 21833 7191
rect 21833 7157 21867 7191
rect 21867 7157 21876 7191
rect 21824 7148 21876 7157
rect 23756 7191 23808 7200
rect 23756 7157 23765 7191
rect 23765 7157 23799 7191
rect 23799 7157 23808 7191
rect 23756 7148 23808 7157
rect 24676 7191 24728 7200
rect 24676 7157 24685 7191
rect 24685 7157 24719 7191
rect 24719 7157 24728 7191
rect 24676 7148 24728 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 1676 6987 1728 6996
rect 1676 6953 1685 6987
rect 1685 6953 1719 6987
rect 1719 6953 1728 6987
rect 1676 6944 1728 6953
rect 2964 6944 3016 6996
rect 3424 6944 3476 6996
rect 4252 6987 4304 6996
rect 4252 6953 4261 6987
rect 4261 6953 4295 6987
rect 4295 6953 4304 6987
rect 4252 6944 4304 6953
rect 6092 6987 6144 6996
rect 2412 6919 2464 6928
rect 2412 6885 2421 6919
rect 2421 6885 2455 6919
rect 2455 6885 2464 6919
rect 2412 6876 2464 6885
rect 2504 6876 2556 6928
rect 5172 6919 5224 6928
rect 5172 6885 5181 6919
rect 5181 6885 5215 6919
rect 5215 6885 5224 6919
rect 5172 6876 5224 6885
rect 6092 6953 6101 6987
rect 6101 6953 6135 6987
rect 6135 6953 6144 6987
rect 6092 6944 6144 6953
rect 7472 6944 7524 6996
rect 11244 6944 11296 6996
rect 11520 6944 11572 6996
rect 12440 6944 12492 6996
rect 15016 6987 15068 6996
rect 6736 6876 6788 6928
rect 7564 6919 7616 6928
rect 2136 6851 2188 6860
rect 2136 6817 2145 6851
rect 2145 6817 2179 6851
rect 2179 6817 2188 6851
rect 2136 6808 2188 6817
rect 6276 6808 6328 6860
rect 6828 6808 6880 6860
rect 7012 6851 7064 6860
rect 7012 6817 7021 6851
rect 7021 6817 7055 6851
rect 7055 6817 7064 6851
rect 7012 6808 7064 6817
rect 7564 6885 7573 6919
rect 7573 6885 7607 6919
rect 7607 6885 7616 6919
rect 7564 6876 7616 6885
rect 8208 6876 8260 6928
rect 13360 6919 13412 6928
rect 13360 6885 13369 6919
rect 13369 6885 13403 6919
rect 13403 6885 13412 6919
rect 13360 6876 13412 6885
rect 15016 6953 15025 6987
rect 15025 6953 15059 6987
rect 15059 6953 15068 6987
rect 15016 6944 15068 6953
rect 17224 6944 17276 6996
rect 18144 6944 18196 6996
rect 20076 6944 20128 6996
rect 20628 6944 20680 6996
rect 22560 6944 22612 6996
rect 13912 6876 13964 6928
rect 8116 6851 8168 6860
rect 8116 6817 8125 6851
rect 8125 6817 8159 6851
rect 8159 6817 8168 6851
rect 8116 6808 8168 6817
rect 9956 6808 10008 6860
rect 11060 6808 11112 6860
rect 11888 6851 11940 6860
rect 11888 6817 11897 6851
rect 11897 6817 11931 6851
rect 11931 6817 11940 6851
rect 11888 6808 11940 6817
rect 12256 6808 12308 6860
rect 16396 6876 16448 6928
rect 16120 6808 16172 6860
rect 16212 6808 16264 6860
rect 17592 6851 17644 6860
rect 17592 6817 17601 6851
rect 17601 6817 17635 6851
rect 17635 6817 17644 6851
rect 17592 6808 17644 6817
rect 2504 6740 2556 6792
rect 3424 6740 3476 6792
rect 4252 6740 4304 6792
rect 5540 6740 5592 6792
rect 7104 6783 7156 6792
rect 7104 6749 7113 6783
rect 7113 6749 7147 6783
rect 7147 6749 7156 6783
rect 7104 6740 7156 6749
rect 10784 6783 10836 6792
rect 10784 6749 10793 6783
rect 10793 6749 10827 6783
rect 10827 6749 10836 6783
rect 10784 6740 10836 6749
rect 3792 6672 3844 6724
rect 4896 6672 4948 6724
rect 6460 6672 6512 6724
rect 3056 6647 3108 6656
rect 3056 6613 3065 6647
rect 3065 6613 3099 6647
rect 3099 6613 3108 6647
rect 3056 6604 3108 6613
rect 3424 6647 3476 6656
rect 3424 6613 3433 6647
rect 3433 6613 3467 6647
rect 3467 6613 3476 6647
rect 3424 6604 3476 6613
rect 4804 6604 4856 6656
rect 6184 6604 6236 6656
rect 8024 6604 8076 6656
rect 8300 6604 8352 6656
rect 9312 6604 9364 6656
rect 11060 6647 11112 6656
rect 11060 6613 11069 6647
rect 11069 6613 11103 6647
rect 11103 6613 11112 6647
rect 11060 6604 11112 6613
rect 13452 6740 13504 6792
rect 15844 6783 15896 6792
rect 15844 6749 15853 6783
rect 15853 6749 15887 6783
rect 15887 6749 15896 6783
rect 15844 6740 15896 6749
rect 18052 6876 18104 6928
rect 20260 6919 20312 6928
rect 20260 6885 20269 6919
rect 20269 6885 20303 6919
rect 20303 6885 20312 6919
rect 20260 6876 20312 6885
rect 20996 6876 21048 6928
rect 22744 6876 22796 6928
rect 24216 6876 24268 6928
rect 24952 6876 25004 6928
rect 18236 6808 18288 6860
rect 19524 6808 19576 6860
rect 19616 6808 19668 6860
rect 22836 6808 22888 6860
rect 20812 6740 20864 6792
rect 22652 6783 22704 6792
rect 22652 6749 22661 6783
rect 22661 6749 22695 6783
rect 22695 6749 22704 6783
rect 22652 6740 22704 6749
rect 24032 6740 24084 6792
rect 24676 6740 24728 6792
rect 14004 6672 14056 6724
rect 17408 6715 17460 6724
rect 17408 6681 17417 6715
rect 17417 6681 17451 6715
rect 17451 6681 17460 6715
rect 17408 6672 17460 6681
rect 20628 6647 20680 6656
rect 20628 6613 20637 6647
rect 20637 6613 20671 6647
rect 20671 6613 20680 6647
rect 20628 6604 20680 6613
rect 23848 6647 23900 6656
rect 23848 6613 23857 6647
rect 23857 6613 23891 6647
rect 23891 6613 23900 6647
rect 23848 6604 23900 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 1768 6400 1820 6452
rect 3056 6400 3108 6452
rect 5172 6400 5224 6452
rect 6276 6443 6328 6452
rect 6276 6409 6285 6443
rect 6285 6409 6319 6443
rect 6319 6409 6328 6443
rect 6276 6400 6328 6409
rect 6828 6400 6880 6452
rect 11888 6443 11940 6452
rect 5540 6332 5592 6384
rect 1492 6264 1544 6316
rect 3792 6264 3844 6316
rect 4436 6264 4488 6316
rect 6828 6264 6880 6316
rect 7104 6264 7156 6316
rect 8944 6264 8996 6316
rect 9864 6264 9916 6316
rect 11888 6409 11897 6443
rect 11897 6409 11931 6443
rect 11931 6409 11940 6443
rect 11888 6400 11940 6409
rect 12348 6400 12400 6452
rect 13360 6400 13412 6452
rect 16120 6400 16172 6452
rect 18052 6400 18104 6452
rect 19432 6400 19484 6452
rect 20996 6443 21048 6452
rect 20996 6409 21005 6443
rect 21005 6409 21039 6443
rect 21039 6409 21048 6443
rect 20996 6400 21048 6409
rect 22652 6400 22704 6452
rect 24216 6400 24268 6452
rect 24952 6400 25004 6452
rect 25320 6400 25372 6452
rect 13544 6332 13596 6384
rect 15200 6332 15252 6384
rect 17224 6332 17276 6384
rect 22744 6375 22796 6384
rect 22744 6341 22753 6375
rect 22753 6341 22787 6375
rect 22787 6341 22796 6375
rect 22744 6332 22796 6341
rect 12440 6307 12492 6316
rect 1676 6196 1728 6248
rect 3332 6196 3384 6248
rect 6920 6196 6972 6248
rect 8116 6196 8168 6248
rect 12440 6273 12449 6307
rect 12449 6273 12483 6307
rect 12483 6273 12492 6307
rect 12440 6264 12492 6273
rect 15660 6264 15712 6316
rect 19248 6264 19300 6316
rect 2504 6171 2556 6180
rect 2504 6137 2513 6171
rect 2513 6137 2547 6171
rect 2547 6137 2556 6171
rect 2504 6128 2556 6137
rect 2964 6128 3016 6180
rect 2412 6060 2464 6112
rect 4068 6060 4120 6112
rect 7840 6060 7892 6112
rect 10140 6128 10192 6180
rect 11060 6196 11112 6248
rect 13728 6196 13780 6248
rect 11152 6171 11204 6180
rect 11152 6137 11161 6171
rect 11161 6137 11195 6171
rect 11195 6137 11204 6171
rect 11152 6128 11204 6137
rect 12348 6128 12400 6180
rect 14004 6171 14056 6180
rect 14004 6137 14013 6171
rect 14013 6137 14047 6171
rect 14047 6137 14056 6171
rect 14004 6128 14056 6137
rect 18972 6196 19024 6248
rect 19616 6239 19668 6248
rect 19616 6205 19625 6239
rect 19625 6205 19659 6239
rect 19659 6205 19668 6239
rect 19616 6196 19668 6205
rect 19984 6196 20036 6248
rect 21916 6196 21968 6248
rect 22008 6239 22060 6248
rect 22008 6205 22017 6239
rect 22017 6205 22051 6239
rect 22051 6205 22060 6239
rect 22008 6196 22060 6205
rect 23848 6196 23900 6248
rect 24308 6196 24360 6248
rect 25136 6196 25188 6248
rect 9956 6060 10008 6112
rect 13544 6060 13596 6112
rect 14096 6060 14148 6112
rect 15200 6060 15252 6112
rect 19432 6128 19484 6180
rect 20076 6128 20128 6180
rect 20812 6128 20864 6180
rect 16304 6103 16356 6112
rect 16304 6069 16313 6103
rect 16313 6069 16347 6103
rect 16347 6069 16356 6103
rect 16304 6060 16356 6069
rect 19524 6060 19576 6112
rect 21824 6103 21876 6112
rect 21824 6069 21833 6103
rect 21833 6069 21867 6103
rect 21867 6069 21876 6103
rect 21824 6060 21876 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1216 5856 1268 5908
rect 2136 5899 2188 5908
rect 2136 5865 2145 5899
rect 2145 5865 2179 5899
rect 2179 5865 2188 5899
rect 2136 5856 2188 5865
rect 2872 5899 2924 5908
rect 2872 5865 2881 5899
rect 2881 5865 2915 5899
rect 2915 5865 2924 5899
rect 2872 5856 2924 5865
rect 3516 5899 3568 5908
rect 3516 5865 3525 5899
rect 3525 5865 3559 5899
rect 3559 5865 3568 5899
rect 3516 5856 3568 5865
rect 4344 5856 4396 5908
rect 5172 5856 5224 5908
rect 5540 5856 5592 5908
rect 7104 5899 7156 5908
rect 7104 5865 7113 5899
rect 7113 5865 7147 5899
rect 7147 5865 7156 5899
rect 7104 5856 7156 5865
rect 8944 5856 8996 5908
rect 12256 5856 12308 5908
rect 16396 5856 16448 5908
rect 17500 5899 17552 5908
rect 17500 5865 17509 5899
rect 17509 5865 17543 5899
rect 17543 5865 17552 5899
rect 17500 5856 17552 5865
rect 17592 5856 17644 5908
rect 19248 5899 19300 5908
rect 19248 5865 19257 5899
rect 19257 5865 19291 5899
rect 19291 5865 19300 5899
rect 19248 5856 19300 5865
rect 20076 5856 20128 5908
rect 4068 5788 4120 5840
rect 1492 5720 1544 5772
rect 3056 5763 3108 5772
rect 3056 5729 3065 5763
rect 3065 5729 3099 5763
rect 3099 5729 3108 5763
rect 3056 5720 3108 5729
rect 4988 5720 5040 5772
rect 6000 5788 6052 5840
rect 7840 5788 7892 5840
rect 10692 5788 10744 5840
rect 12348 5788 12400 5840
rect 13728 5831 13780 5840
rect 13728 5797 13737 5831
rect 13737 5797 13771 5831
rect 13771 5797 13780 5831
rect 13728 5788 13780 5797
rect 15200 5788 15252 5840
rect 15476 5788 15528 5840
rect 14280 5763 14332 5772
rect 14280 5729 14289 5763
rect 14289 5729 14323 5763
rect 14323 5729 14332 5763
rect 14280 5720 14332 5729
rect 15292 5720 15344 5772
rect 15844 5720 15896 5772
rect 17408 5763 17460 5772
rect 17408 5729 17417 5763
rect 17417 5729 17451 5763
rect 17451 5729 17460 5763
rect 17408 5720 17460 5729
rect 18052 5720 18104 5772
rect 18328 5720 18380 5772
rect 21364 5788 21416 5840
rect 22744 5788 22796 5840
rect 24308 5788 24360 5840
rect 19984 5720 20036 5772
rect 21272 5763 21324 5772
rect 21272 5729 21281 5763
rect 21281 5729 21315 5763
rect 21315 5729 21324 5763
rect 21272 5720 21324 5729
rect 4160 5695 4212 5704
rect 4160 5661 4169 5695
rect 4169 5661 4203 5695
rect 4203 5661 4212 5695
rect 4160 5652 4212 5661
rect 6092 5652 6144 5704
rect 6460 5695 6512 5704
rect 6460 5661 6469 5695
rect 6469 5661 6503 5695
rect 6503 5661 6512 5695
rect 6460 5652 6512 5661
rect 9588 5652 9640 5704
rect 10968 5652 11020 5704
rect 11888 5652 11940 5704
rect 2964 5584 3016 5636
rect 5080 5584 5132 5636
rect 8024 5584 8076 5636
rect 8668 5627 8720 5636
rect 8668 5593 8677 5627
rect 8677 5593 8711 5627
rect 8711 5593 8720 5627
rect 8668 5584 8720 5593
rect 11520 5584 11572 5636
rect 18880 5652 18932 5704
rect 22008 5720 22060 5772
rect 22284 5763 22336 5772
rect 22284 5729 22293 5763
rect 22293 5729 22327 5763
rect 22327 5729 22336 5763
rect 22284 5720 22336 5729
rect 24216 5763 24268 5772
rect 21916 5652 21968 5704
rect 24216 5729 24225 5763
rect 24225 5729 24259 5763
rect 24259 5729 24268 5763
rect 24216 5720 24268 5729
rect 25136 5720 25188 5772
rect 23756 5584 23808 5636
rect 3700 5516 3752 5568
rect 9956 5516 10008 5568
rect 10140 5559 10192 5568
rect 10140 5525 10149 5559
rect 10149 5525 10183 5559
rect 10183 5525 10192 5559
rect 10140 5516 10192 5525
rect 14556 5559 14608 5568
rect 14556 5525 14565 5559
rect 14565 5525 14599 5559
rect 14599 5525 14608 5559
rect 14556 5516 14608 5525
rect 16580 5559 16632 5568
rect 16580 5525 16589 5559
rect 16589 5525 16623 5559
rect 16623 5525 16632 5559
rect 16580 5516 16632 5525
rect 23204 5559 23256 5568
rect 23204 5525 23213 5559
rect 23213 5525 23247 5559
rect 23247 5525 23256 5559
rect 23204 5516 23256 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 1584 5355 1636 5364
rect 1584 5321 1593 5355
rect 1593 5321 1627 5355
rect 1627 5321 1636 5355
rect 1584 5312 1636 5321
rect 2412 5312 2464 5364
rect 3056 5312 3108 5364
rect 4896 5312 4948 5364
rect 6000 5355 6052 5364
rect 6000 5321 6009 5355
rect 6009 5321 6043 5355
rect 6043 5321 6052 5355
rect 6000 5312 6052 5321
rect 7840 5355 7892 5364
rect 7840 5321 7849 5355
rect 7849 5321 7883 5355
rect 7883 5321 7892 5355
rect 7840 5312 7892 5321
rect 9036 5312 9088 5364
rect 5540 5244 5592 5296
rect 4160 5176 4212 5228
rect 4620 5176 4672 5228
rect 1400 5151 1452 5160
rect 1400 5117 1409 5151
rect 1409 5117 1443 5151
rect 1443 5117 1452 5151
rect 1400 5108 1452 5117
rect 3424 5151 3476 5160
rect 3424 5117 3433 5151
rect 3433 5117 3467 5151
rect 3467 5117 3476 5151
rect 3424 5108 3476 5117
rect 3700 5151 3752 5160
rect 3700 5117 3709 5151
rect 3709 5117 3743 5151
rect 3743 5117 3752 5151
rect 3700 5108 3752 5117
rect 7932 5244 7984 5296
rect 8576 5244 8628 5296
rect 9128 5244 9180 5296
rect 9864 5219 9916 5228
rect 9864 5185 9873 5219
rect 9873 5185 9907 5219
rect 9907 5185 9916 5219
rect 9864 5176 9916 5185
rect 12348 5312 12400 5364
rect 13728 5355 13780 5364
rect 13728 5321 13737 5355
rect 13737 5321 13771 5355
rect 13771 5321 13780 5355
rect 13728 5312 13780 5321
rect 15844 5312 15896 5364
rect 17408 5355 17460 5364
rect 15936 5244 15988 5296
rect 17408 5321 17417 5355
rect 17417 5321 17451 5355
rect 17451 5321 17460 5355
rect 17408 5312 17460 5321
rect 18052 5312 18104 5364
rect 18328 5355 18380 5364
rect 18328 5321 18337 5355
rect 18337 5321 18371 5355
rect 18371 5321 18380 5355
rect 18328 5312 18380 5321
rect 20628 5312 20680 5364
rect 22744 5312 22796 5364
rect 23204 5312 23256 5364
rect 23848 5312 23900 5364
rect 24216 5312 24268 5364
rect 16672 5244 16724 5296
rect 10784 5176 10836 5228
rect 12992 5176 13044 5228
rect 14556 5176 14608 5228
rect 15292 5176 15344 5228
rect 15476 5176 15528 5228
rect 16764 5176 16816 5228
rect 19984 5244 20036 5296
rect 21180 5244 21232 5296
rect 20076 5176 20128 5228
rect 21824 5219 21876 5228
rect 21824 5185 21833 5219
rect 21833 5185 21867 5219
rect 21867 5185 21876 5219
rect 21824 5176 21876 5185
rect 24124 5176 24176 5228
rect 4528 5040 4580 5092
rect 4804 5040 4856 5092
rect 4896 5083 4948 5092
rect 4896 5049 4905 5083
rect 4905 5049 4939 5083
rect 4939 5049 4948 5083
rect 8024 5083 8076 5092
rect 4896 5040 4948 5049
rect 8024 5049 8033 5083
rect 8033 5049 8067 5083
rect 8067 5049 8076 5083
rect 8024 5040 8076 5049
rect 8668 5083 8720 5092
rect 4068 4972 4120 5024
rect 8668 5049 8677 5083
rect 8677 5049 8711 5083
rect 8711 5049 8720 5083
rect 8668 5040 8720 5049
rect 8300 4972 8352 5024
rect 12348 5040 12400 5092
rect 10692 4972 10744 5024
rect 19156 5108 19208 5160
rect 19340 5108 19392 5160
rect 15936 5040 15988 5092
rect 16580 5040 16632 5092
rect 16672 5040 16724 5092
rect 20996 5108 21048 5160
rect 23756 5083 23808 5092
rect 23756 5049 23765 5083
rect 23765 5049 23799 5083
rect 23799 5049 23808 5083
rect 23756 5040 23808 5049
rect 23848 5083 23900 5092
rect 23848 5049 23857 5083
rect 23857 5049 23891 5083
rect 23891 5049 23900 5083
rect 23848 5040 23900 5049
rect 20444 5015 20496 5024
rect 20444 4981 20453 5015
rect 20453 4981 20487 5015
rect 20487 4981 20496 5015
rect 20444 4972 20496 4981
rect 21272 5015 21324 5024
rect 21272 4981 21281 5015
rect 21281 4981 21315 5015
rect 21315 4981 21324 5015
rect 21272 4972 21324 4981
rect 22744 5015 22796 5024
rect 22744 4981 22753 5015
rect 22753 4981 22787 5015
rect 22787 4981 22796 5015
rect 22744 4972 22796 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1124 4768 1176 4820
rect 2504 4811 2556 4820
rect 2504 4777 2513 4811
rect 2513 4777 2547 4811
rect 2547 4777 2556 4811
rect 2504 4768 2556 4777
rect 3700 4768 3752 4820
rect 4160 4768 4212 4820
rect 7196 4768 7248 4820
rect 8300 4811 8352 4820
rect 8300 4777 8309 4811
rect 8309 4777 8343 4811
rect 8343 4777 8352 4811
rect 8300 4768 8352 4777
rect 12992 4811 13044 4820
rect 12992 4777 13001 4811
rect 13001 4777 13035 4811
rect 13035 4777 13044 4811
rect 12992 4768 13044 4777
rect 4620 4700 4672 4752
rect 4896 4743 4948 4752
rect 4896 4709 4905 4743
rect 4905 4709 4939 4743
rect 4939 4709 4948 4743
rect 4896 4700 4948 4709
rect 6092 4700 6144 4752
rect 8668 4700 8720 4752
rect 11796 4743 11848 4752
rect 11796 4709 11799 4743
rect 11799 4709 11833 4743
rect 11833 4709 11848 4743
rect 11796 4700 11848 4709
rect 12348 4700 12400 4752
rect 13452 4743 13504 4752
rect 13452 4709 13461 4743
rect 13461 4709 13495 4743
rect 13495 4709 13504 4743
rect 13452 4700 13504 4709
rect 13544 4743 13596 4752
rect 13544 4709 13553 4743
rect 13553 4709 13587 4743
rect 13587 4709 13596 4743
rect 13544 4700 13596 4709
rect 14280 4700 14332 4752
rect 1952 4632 2004 4684
rect 2964 4675 3016 4684
rect 2964 4641 2973 4675
rect 2973 4641 3007 4675
rect 3007 4641 3016 4675
rect 2964 4632 3016 4641
rect 7472 4632 7524 4684
rect 9220 4632 9272 4684
rect 9864 4675 9916 4684
rect 9864 4641 9873 4675
rect 9873 4641 9907 4675
rect 9907 4641 9916 4675
rect 9864 4632 9916 4641
rect 10140 4632 10192 4684
rect 11888 4632 11940 4684
rect 4804 4607 4856 4616
rect 4804 4573 4813 4607
rect 4813 4573 4847 4607
rect 4847 4573 4856 4607
rect 4804 4564 4856 4573
rect 6920 4564 6972 4616
rect 11152 4564 11204 4616
rect 15752 4768 15804 4820
rect 16764 4811 16816 4820
rect 16764 4777 16773 4811
rect 16773 4777 16807 4811
rect 16807 4777 16816 4811
rect 16764 4768 16816 4777
rect 19340 4768 19392 4820
rect 20904 4768 20956 4820
rect 15936 4743 15988 4752
rect 15936 4709 15945 4743
rect 15945 4709 15979 4743
rect 15979 4709 15988 4743
rect 15936 4700 15988 4709
rect 17224 4700 17276 4752
rect 17408 4700 17460 4752
rect 21824 4768 21876 4820
rect 22284 4811 22336 4820
rect 22284 4777 22293 4811
rect 22293 4777 22327 4811
rect 22327 4777 22336 4811
rect 22284 4768 22336 4777
rect 23756 4768 23808 4820
rect 24768 4811 24820 4820
rect 24768 4777 24777 4811
rect 24777 4777 24811 4811
rect 24811 4777 24820 4811
rect 24768 4768 24820 4777
rect 22744 4700 22796 4752
rect 17500 4632 17552 4684
rect 19248 4632 19300 4684
rect 24584 4675 24636 4684
rect 24584 4641 24593 4675
rect 24593 4641 24627 4675
rect 24627 4641 24636 4675
rect 24584 4632 24636 4641
rect 10968 4539 11020 4548
rect 10968 4505 10977 4539
rect 10977 4505 11011 4539
rect 11011 4505 11020 4539
rect 10968 4496 11020 4505
rect 4252 4471 4304 4480
rect 4252 4437 4261 4471
rect 4261 4437 4295 4471
rect 4295 4437 4304 4471
rect 4252 4428 4304 4437
rect 8852 4471 8904 4480
rect 8852 4437 8861 4471
rect 8861 4437 8895 4471
rect 8895 4437 8904 4471
rect 8852 4428 8904 4437
rect 10692 4428 10744 4480
rect 12900 4428 12952 4480
rect 13360 4428 13412 4480
rect 14464 4471 14516 4480
rect 14464 4437 14473 4471
rect 14473 4437 14507 4471
rect 14507 4437 14516 4471
rect 14464 4428 14516 4437
rect 16212 4607 16264 4616
rect 16212 4573 16221 4607
rect 16221 4573 16255 4607
rect 16255 4573 16264 4607
rect 16212 4564 16264 4573
rect 20996 4607 21048 4616
rect 20996 4573 21005 4607
rect 21005 4573 21039 4607
rect 21039 4573 21048 4607
rect 20996 4564 21048 4573
rect 21272 4607 21324 4616
rect 21272 4573 21281 4607
rect 21281 4573 21315 4607
rect 21315 4573 21324 4607
rect 21272 4564 21324 4573
rect 22928 4607 22980 4616
rect 22928 4573 22937 4607
rect 22937 4573 22971 4607
rect 22971 4573 22980 4607
rect 22928 4564 22980 4573
rect 24032 4564 24084 4616
rect 24216 4496 24268 4548
rect 25596 4496 25648 4548
rect 16764 4428 16816 4480
rect 18236 4471 18288 4480
rect 18236 4437 18245 4471
rect 18245 4437 18279 4471
rect 18279 4437 18288 4471
rect 18236 4428 18288 4437
rect 18604 4471 18656 4480
rect 18604 4437 18613 4471
rect 18613 4437 18647 4471
rect 18647 4437 18656 4471
rect 18604 4428 18656 4437
rect 25136 4428 25188 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 1492 4224 1544 4276
rect 1952 4267 2004 4276
rect 1952 4233 1961 4267
rect 1961 4233 1995 4267
rect 1995 4233 2004 4267
rect 1952 4224 2004 4233
rect 2964 4199 3016 4208
rect 2964 4165 2973 4199
rect 2973 4165 3007 4199
rect 3007 4165 3016 4199
rect 2964 4156 3016 4165
rect 4896 4224 4948 4276
rect 11152 4224 11204 4276
rect 13544 4267 13596 4276
rect 13544 4233 13553 4267
rect 13553 4233 13587 4267
rect 13587 4233 13596 4267
rect 13544 4224 13596 4233
rect 14556 4224 14608 4276
rect 15936 4224 15988 4276
rect 17500 4224 17552 4276
rect 18236 4224 18288 4276
rect 19248 4224 19300 4276
rect 20904 4267 20956 4276
rect 20904 4233 20913 4267
rect 20913 4233 20947 4267
rect 20947 4233 20956 4267
rect 20904 4224 20956 4233
rect 22744 4224 22796 4276
rect 24032 4224 24084 4276
rect 25228 4267 25280 4276
rect 25228 4233 25237 4267
rect 25237 4233 25271 4267
rect 25271 4233 25280 4267
rect 25228 4224 25280 4233
rect 9772 4156 9824 4208
rect 9864 4199 9916 4208
rect 9864 4165 9873 4199
rect 9873 4165 9907 4199
rect 9907 4165 9916 4199
rect 9864 4156 9916 4165
rect 13636 4156 13688 4208
rect 16672 4156 16724 4208
rect 19340 4199 19392 4208
rect 2596 4088 2648 4140
rect 3516 4088 3568 4140
rect 3608 4063 3660 4072
rect 3608 4029 3617 4063
rect 3617 4029 3651 4063
rect 3651 4029 3660 4063
rect 3608 4020 3660 4029
rect 1768 3952 1820 4004
rect 4068 4088 4120 4140
rect 4252 4088 4304 4140
rect 6276 4088 6328 4140
rect 8852 4131 8904 4140
rect 8852 4097 8861 4131
rect 8861 4097 8895 4131
rect 8895 4097 8904 4131
rect 8852 4088 8904 4097
rect 9128 4131 9180 4140
rect 9128 4097 9137 4131
rect 9137 4097 9171 4131
rect 9171 4097 9180 4131
rect 9128 4088 9180 4097
rect 10968 4088 11020 4140
rect 11520 4131 11572 4140
rect 11520 4097 11529 4131
rect 11529 4097 11563 4131
rect 11563 4097 11572 4131
rect 11520 4088 11572 4097
rect 7012 4063 7064 4072
rect 7012 4029 7021 4063
rect 7021 4029 7055 4063
rect 7055 4029 7064 4063
rect 7012 4020 7064 4029
rect 3792 3884 3844 3936
rect 4160 3884 4212 3936
rect 6920 3952 6972 4004
rect 10876 3995 10928 4004
rect 7196 3884 7248 3936
rect 8208 3884 8260 3936
rect 10876 3961 10885 3995
rect 10885 3961 10919 3995
rect 10919 3961 10928 3995
rect 10876 3952 10928 3961
rect 10968 3995 11020 4004
rect 10968 3961 10977 3995
rect 10977 3961 11011 3995
rect 11011 3961 11020 3995
rect 12900 3995 12952 4004
rect 10968 3952 11020 3961
rect 12900 3961 12909 3995
rect 12909 3961 12943 3995
rect 12943 3961 12952 3995
rect 12900 3952 12952 3961
rect 10140 3884 10192 3936
rect 11796 3927 11848 3936
rect 11796 3893 11805 3927
rect 11805 3893 11839 3927
rect 11839 3893 11848 3927
rect 11796 3884 11848 3893
rect 14648 4088 14700 4140
rect 16212 4088 16264 4140
rect 17408 4088 17460 4140
rect 18604 4088 18656 4140
rect 19340 4165 19349 4199
rect 19349 4165 19383 4199
rect 19383 4165 19392 4199
rect 19340 4156 19392 4165
rect 19432 4156 19484 4208
rect 24216 4199 24268 4208
rect 24216 4165 24225 4199
rect 24225 4165 24259 4199
rect 24259 4165 24268 4199
rect 24216 4156 24268 4165
rect 24676 4156 24728 4208
rect 15936 3995 15988 4004
rect 14372 3884 14424 3936
rect 15936 3961 15945 3995
rect 15945 3961 15979 3995
rect 15979 3961 15988 3995
rect 15936 3952 15988 3961
rect 16304 3952 16356 4004
rect 16580 3995 16632 4004
rect 16580 3961 16589 3995
rect 16589 3961 16623 3995
rect 16623 3961 16632 3995
rect 16580 3952 16632 3961
rect 18236 3952 18288 4004
rect 20076 4088 20128 4140
rect 20444 4088 20496 4140
rect 21272 4088 21324 4140
rect 22836 4088 22888 4140
rect 21824 4020 21876 4072
rect 22008 4020 22060 4072
rect 20076 3995 20128 4004
rect 20076 3961 20085 3995
rect 20085 3961 20119 3995
rect 20119 3961 20128 3995
rect 20076 3952 20128 3961
rect 20996 3952 21048 4004
rect 22100 3952 22152 4004
rect 20260 3884 20312 3936
rect 22008 3884 22060 3936
rect 22744 3884 22796 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 4252 3680 4304 3732
rect 7196 3723 7248 3732
rect 7196 3689 7205 3723
rect 7205 3689 7239 3723
rect 7239 3689 7248 3723
rect 7196 3680 7248 3689
rect 10968 3680 11020 3732
rect 12164 3723 12216 3732
rect 12164 3689 12173 3723
rect 12173 3689 12207 3723
rect 12207 3689 12216 3723
rect 12164 3680 12216 3689
rect 12900 3680 12952 3732
rect 14648 3680 14700 3732
rect 15752 3680 15804 3732
rect 15936 3680 15988 3732
rect 16764 3680 16816 3732
rect 20076 3680 20128 3732
rect 20260 3723 20312 3732
rect 20260 3689 20269 3723
rect 20269 3689 20303 3723
rect 20303 3689 20312 3723
rect 20260 3680 20312 3689
rect 22928 3680 22980 3732
rect 25136 3723 25188 3732
rect 25136 3689 25145 3723
rect 25145 3689 25179 3723
rect 25179 3689 25188 3723
rect 25136 3680 25188 3689
rect 4436 3612 4488 3664
rect 7012 3612 7064 3664
rect 8208 3612 8260 3664
rect 8668 3655 8720 3664
rect 8668 3621 8677 3655
rect 8677 3621 8711 3655
rect 8711 3621 8720 3655
rect 8668 3612 8720 3621
rect 11796 3612 11848 3664
rect 13084 3612 13136 3664
rect 15476 3612 15528 3664
rect 1952 3587 2004 3596
rect 1952 3553 1961 3587
rect 1961 3553 1995 3587
rect 1995 3553 2004 3587
rect 1952 3544 2004 3553
rect 3332 3544 3384 3596
rect 3424 3544 3476 3596
rect 4160 3587 4212 3596
rect 4160 3553 4169 3587
rect 4169 3553 4203 3587
rect 4203 3553 4212 3587
rect 4160 3544 4212 3553
rect 4344 3544 4396 3596
rect 6552 3476 6604 3528
rect 4528 3408 4580 3460
rect 5356 3408 5408 3460
rect 7472 3544 7524 3596
rect 10140 3587 10192 3596
rect 8024 3519 8076 3528
rect 8024 3485 8033 3519
rect 8033 3485 8067 3519
rect 8067 3485 8076 3519
rect 8024 3476 8076 3485
rect 8392 3476 8444 3528
rect 10140 3553 10149 3587
rect 10149 3553 10183 3587
rect 10183 3553 10192 3587
rect 10140 3544 10192 3553
rect 10048 3476 10100 3528
rect 9496 3408 9548 3460
rect 11980 3476 12032 3528
rect 14004 3476 14056 3528
rect 15476 3519 15528 3528
rect 11704 3408 11756 3460
rect 13452 3408 13504 3460
rect 15476 3485 15485 3519
rect 15485 3485 15519 3519
rect 15519 3485 15528 3519
rect 15476 3476 15528 3485
rect 17868 3612 17920 3664
rect 18236 3612 18288 3664
rect 18696 3612 18748 3664
rect 21824 3612 21876 3664
rect 16212 3544 16264 3596
rect 19616 3544 19668 3596
rect 20352 3544 20404 3596
rect 21180 3544 21232 3596
rect 22100 3544 22152 3596
rect 24216 3544 24268 3596
rect 24952 3587 25004 3596
rect 24952 3553 24961 3587
rect 24961 3553 24995 3587
rect 24995 3553 25004 3587
rect 24952 3544 25004 3553
rect 18236 3476 18288 3528
rect 20812 3476 20864 3528
rect 3884 3340 3936 3392
rect 5080 3383 5132 3392
rect 5080 3349 5089 3383
rect 5089 3349 5123 3383
rect 5123 3349 5132 3383
rect 5080 3340 5132 3349
rect 5448 3340 5500 3392
rect 10140 3340 10192 3392
rect 10692 3383 10744 3392
rect 10692 3349 10701 3383
rect 10701 3349 10735 3383
rect 10735 3349 10744 3383
rect 10692 3340 10744 3349
rect 10968 3340 11020 3392
rect 16028 3340 16080 3392
rect 22192 3408 22244 3460
rect 20352 3340 20404 3392
rect 22468 3383 22520 3392
rect 22468 3349 22477 3383
rect 22477 3349 22511 3383
rect 22511 3349 22520 3383
rect 22468 3340 22520 3349
rect 22652 3340 22704 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1952 3179 2004 3188
rect 1952 3145 1961 3179
rect 1961 3145 1995 3179
rect 1995 3145 2004 3179
rect 1952 3136 2004 3145
rect 3332 3136 3384 3188
rect 4160 3179 4212 3188
rect 4160 3145 4169 3179
rect 4169 3145 4203 3179
rect 4203 3145 4212 3179
rect 4160 3136 4212 3145
rect 4804 3136 4856 3188
rect 5080 3136 5132 3188
rect 6552 3179 6604 3188
rect 6552 3145 6561 3179
rect 6561 3145 6595 3179
rect 6595 3145 6604 3179
rect 6552 3136 6604 3145
rect 7932 3179 7984 3188
rect 7932 3145 7941 3179
rect 7941 3145 7975 3179
rect 7975 3145 7984 3179
rect 7932 3136 7984 3145
rect 8208 3179 8260 3188
rect 8208 3145 8217 3179
rect 8217 3145 8251 3179
rect 8251 3145 8260 3179
rect 8208 3136 8260 3145
rect 10048 3179 10100 3188
rect 10048 3145 10057 3179
rect 10057 3145 10091 3179
rect 10091 3145 10100 3179
rect 10048 3136 10100 3145
rect 12164 3179 12216 3188
rect 12164 3145 12173 3179
rect 12173 3145 12207 3179
rect 12207 3145 12216 3179
rect 12164 3136 12216 3145
rect 12716 3179 12768 3188
rect 12716 3145 12725 3179
rect 12725 3145 12759 3179
rect 12759 3145 12768 3179
rect 12716 3136 12768 3145
rect 14004 3179 14056 3188
rect 14004 3145 14013 3179
rect 14013 3145 14047 3179
rect 14047 3145 14056 3179
rect 14004 3136 14056 3145
rect 10968 3068 11020 3120
rect 3976 3000 4028 3052
rect 3516 2932 3568 2984
rect 4712 2864 4764 2916
rect 5448 2932 5500 2984
rect 10692 3000 10744 3052
rect 15292 3136 15344 3188
rect 15476 3136 15528 3188
rect 17868 3179 17920 3188
rect 17868 3145 17877 3179
rect 17877 3145 17911 3179
rect 17911 3145 17920 3179
rect 17868 3136 17920 3145
rect 18236 3179 18288 3188
rect 18236 3145 18245 3179
rect 18245 3145 18279 3179
rect 18279 3145 18288 3179
rect 18236 3136 18288 3145
rect 13636 3043 13688 3052
rect 13636 3009 13645 3043
rect 13645 3009 13679 3043
rect 13679 3009 13688 3043
rect 13636 3000 13688 3009
rect 14740 3000 14792 3052
rect 16580 3043 16632 3052
rect 16580 3009 16589 3043
rect 16589 3009 16623 3043
rect 16623 3009 16632 3043
rect 16580 3000 16632 3009
rect 6552 2932 6604 2984
rect 7932 2932 7984 2984
rect 9496 2975 9548 2984
rect 9496 2941 9505 2975
rect 9505 2941 9539 2975
rect 9539 2941 9548 2975
rect 9496 2932 9548 2941
rect 14464 2975 14516 2984
rect 14464 2941 14473 2975
rect 14473 2941 14507 2975
rect 14507 2941 14516 2975
rect 14464 2932 14516 2941
rect 20352 3136 20404 3188
rect 22100 3136 22152 3188
rect 23664 3136 23716 3188
rect 24952 3136 25004 3188
rect 19616 3111 19668 3120
rect 19616 3077 19625 3111
rect 19625 3077 19659 3111
rect 19659 3077 19668 3111
rect 19616 3068 19668 3077
rect 21916 3068 21968 3120
rect 24216 3111 24268 3120
rect 24216 3077 24225 3111
rect 24225 3077 24259 3111
rect 24259 3077 24268 3111
rect 24216 3068 24268 3077
rect 27528 3068 27580 3120
rect 19432 3000 19484 3052
rect 7196 2864 7248 2916
rect 11796 2864 11848 2916
rect 13084 2907 13136 2916
rect 4896 2839 4948 2848
rect 4896 2805 4905 2839
rect 4905 2805 4939 2839
rect 4939 2805 4948 2839
rect 4896 2796 4948 2805
rect 6460 2796 6512 2848
rect 6920 2839 6972 2848
rect 6920 2805 6929 2839
rect 6929 2805 6963 2839
rect 6963 2805 6972 2839
rect 6920 2796 6972 2805
rect 11520 2839 11572 2848
rect 11520 2805 11529 2839
rect 11529 2805 11563 2839
rect 11563 2805 11572 2839
rect 11520 2796 11572 2805
rect 13084 2873 13093 2907
rect 13093 2873 13127 2907
rect 13127 2873 13136 2907
rect 13084 2864 13136 2873
rect 15752 2864 15804 2916
rect 16028 2907 16080 2916
rect 16028 2873 16037 2907
rect 16037 2873 16071 2907
rect 16071 2873 16080 2907
rect 16028 2864 16080 2873
rect 16212 2864 16264 2916
rect 20996 2932 21048 2984
rect 22652 2932 22704 2984
rect 23940 3000 23992 3052
rect 14648 2839 14700 2848
rect 14648 2805 14657 2839
rect 14657 2805 14691 2839
rect 14691 2805 14700 2839
rect 14648 2796 14700 2805
rect 20996 2839 21048 2848
rect 20996 2805 21005 2839
rect 21005 2805 21039 2839
rect 21039 2805 21048 2839
rect 20996 2796 21048 2805
rect 21088 2796 21140 2848
rect 22008 2796 22060 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 2780 2592 2832 2644
rect 2504 2456 2556 2508
rect 3700 2592 3752 2644
rect 4344 2635 4396 2644
rect 4344 2601 4353 2635
rect 4353 2601 4387 2635
rect 4387 2601 4396 2635
rect 4344 2592 4396 2601
rect 6276 2592 6328 2644
rect 6460 2592 6512 2644
rect 8024 2592 8076 2644
rect 9588 2592 9640 2644
rect 11980 2635 12032 2644
rect 11980 2601 11989 2635
rect 11989 2601 12023 2635
rect 12023 2601 12032 2635
rect 11980 2592 12032 2601
rect 13084 2592 13136 2644
rect 3884 2524 3936 2576
rect 6184 2524 6236 2576
rect 6552 2524 6604 2576
rect 9036 2524 9088 2576
rect 11520 2524 11572 2576
rect 16028 2524 16080 2576
rect 21180 2592 21232 2644
rect 8576 2456 8628 2508
rect 6092 2320 6144 2372
rect 2504 2295 2556 2304
rect 2504 2261 2513 2295
rect 2513 2261 2547 2295
rect 2547 2261 2556 2295
rect 2504 2252 2556 2261
rect 4344 2252 4396 2304
rect 8392 2320 8444 2372
rect 10140 2456 10192 2508
rect 11704 2499 11756 2508
rect 11704 2465 11713 2499
rect 11713 2465 11747 2499
rect 11747 2465 11756 2499
rect 11704 2456 11756 2465
rect 17132 2456 17184 2508
rect 9404 2320 9456 2372
rect 13636 2320 13688 2372
rect 7380 2252 7432 2304
rect 8484 2252 8536 2304
rect 9036 2295 9088 2304
rect 9036 2261 9045 2295
rect 9045 2261 9079 2295
rect 9079 2261 9088 2295
rect 9496 2295 9548 2304
rect 9036 2252 9088 2261
rect 9496 2261 9505 2295
rect 9505 2261 9539 2295
rect 9539 2261 9548 2295
rect 9496 2252 9548 2261
rect 12440 2295 12492 2304
rect 12440 2261 12449 2295
rect 12449 2261 12483 2295
rect 12483 2261 12492 2295
rect 12440 2252 12492 2261
rect 18880 2431 18932 2440
rect 16120 2320 16172 2372
rect 18880 2397 18889 2431
rect 18889 2397 18923 2431
rect 18923 2397 18932 2431
rect 18880 2388 18932 2397
rect 21088 2524 21140 2576
rect 22652 2524 22704 2576
rect 19524 2456 19576 2508
rect 19616 2388 19668 2440
rect 21272 2320 21324 2372
rect 23940 2320 23992 2372
rect 26424 2320 26476 2372
rect 22192 2252 22244 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 10140 2048 10192 2100
rect 16948 2048 17000 2100
rect 19616 2048 19668 2100
rect 4896 1980 4948 2032
rect 14464 1980 14516 2032
rect 21732 76 21784 128
rect 23204 76 23256 128
<< metal2 >>
rect 20 27532 72 27538
rect 754 27532 810 28000
rect 754 27520 756 27532
rect 20 27474 72 27480
rect 808 27520 810 27532
rect 1780 27526 2176 27554
rect 756 27474 808 27480
rect 32 10606 60 27474
rect 768 27443 796 27474
rect 1214 26888 1270 26897
rect 1214 26823 1270 26832
rect 1124 20800 1176 20806
rect 1124 20742 1176 20748
rect 112 15904 164 15910
rect 112 15846 164 15852
rect 124 13977 152 15846
rect 110 13968 166 13977
rect 110 13903 166 13912
rect 110 11248 166 11257
rect 110 11183 166 11192
rect 20 10600 72 10606
rect 20 10542 72 10548
rect 124 9586 152 11183
rect 112 9580 164 9586
rect 112 9522 164 9528
rect 848 7812 900 7818
rect 848 7754 900 7760
rect 478 82 534 480
rect 860 82 888 7754
rect 1136 7342 1164 20742
rect 1228 19922 1256 26823
rect 1582 24168 1638 24177
rect 1582 24103 1638 24112
rect 1596 23186 1624 24103
rect 1584 23180 1636 23186
rect 1584 23122 1636 23128
rect 1596 22778 1624 23122
rect 1584 22772 1636 22778
rect 1584 22714 1636 22720
rect 1582 21312 1638 21321
rect 1582 21247 1638 21256
rect 1596 20602 1624 21247
rect 1584 20596 1636 20602
rect 1584 20538 1636 20544
rect 1308 20392 1360 20398
rect 1308 20334 1360 20340
rect 1216 19916 1268 19922
rect 1216 19858 1268 19864
rect 1228 19514 1256 19858
rect 1216 19508 1268 19514
rect 1216 19450 1268 19456
rect 1216 18828 1268 18834
rect 1216 18770 1268 18776
rect 1228 17542 1256 18770
rect 1216 17536 1268 17542
rect 1216 17478 1268 17484
rect 1124 7336 1176 7342
rect 1124 7278 1176 7284
rect 1136 4826 1164 7278
rect 1228 5914 1256 17478
rect 1320 15745 1348 20334
rect 1582 20088 1638 20097
rect 1582 20023 1638 20032
rect 1596 18970 1624 20023
rect 1584 18964 1636 18970
rect 1584 18906 1636 18912
rect 1582 18728 1638 18737
rect 1582 18663 1638 18672
rect 1596 18426 1624 18663
rect 1584 18420 1636 18426
rect 1584 18362 1636 18368
rect 1492 18080 1544 18086
rect 1492 18022 1544 18028
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1412 16250 1440 16594
rect 1400 16244 1452 16250
rect 1400 16186 1452 16192
rect 1306 15736 1362 15745
rect 1306 15671 1362 15680
rect 1504 11286 1532 18022
rect 1582 17504 1638 17513
rect 1582 17439 1638 17448
rect 1596 17338 1624 17439
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 1582 16960 1638 16969
rect 1582 16895 1638 16904
rect 1596 16794 1624 16895
rect 1584 16788 1636 16794
rect 1584 16730 1636 16736
rect 1584 16448 1636 16454
rect 1584 16390 1636 16396
rect 1596 13938 1624 16390
rect 1676 16176 1728 16182
rect 1676 16118 1728 16124
rect 1584 13932 1636 13938
rect 1584 13874 1636 13880
rect 1582 13832 1638 13841
rect 1582 13767 1638 13776
rect 1492 11280 1544 11286
rect 1492 11222 1544 11228
rect 1596 8514 1624 13767
rect 1688 13462 1716 16118
rect 1676 13456 1728 13462
rect 1676 13398 1728 13404
rect 1780 12306 1808 27526
rect 2148 27520 2176 27526
rect 2226 27520 2282 28000
rect 2872 27532 2924 27538
rect 2148 27492 2268 27520
rect 3698 27532 3754 28000
rect 3698 27520 3700 27532
rect 2872 27474 2924 27480
rect 3752 27520 3754 27532
rect 5170 27554 5226 28000
rect 5170 27526 5396 27554
rect 5170 27520 5226 27526
rect 3700 27474 3752 27480
rect 1858 25392 1914 25401
rect 1858 25327 1914 25336
rect 1872 23662 1900 25327
rect 1860 23656 1912 23662
rect 1860 23598 1912 23604
rect 2780 23588 2832 23594
rect 2780 23530 2832 23536
rect 2596 22976 2648 22982
rect 2596 22918 2648 22924
rect 1858 22672 1914 22681
rect 1858 22607 1914 22616
rect 1872 19310 1900 22607
rect 2136 21480 2188 21486
rect 2136 21422 2188 21428
rect 2042 20360 2098 20369
rect 2042 20295 2098 20304
rect 1860 19304 1912 19310
rect 1860 19246 1912 19252
rect 2056 18426 2084 20295
rect 2044 18420 2096 18426
rect 2044 18362 2096 18368
rect 2056 18222 2084 18362
rect 2044 18216 2096 18222
rect 2044 18158 2096 18164
rect 2148 17338 2176 21422
rect 2412 21004 2464 21010
rect 2412 20946 2464 20952
rect 2424 20262 2452 20946
rect 2412 20256 2464 20262
rect 2412 20198 2464 20204
rect 2320 19168 2372 19174
rect 2320 19110 2372 19116
rect 2136 17332 2188 17338
rect 2136 17274 2188 17280
rect 2332 16794 2360 19110
rect 2320 16788 2372 16794
rect 2148 16748 2320 16776
rect 2044 16040 2096 16046
rect 2042 16008 2044 16017
rect 2096 16008 2098 16017
rect 2042 15943 2098 15952
rect 2056 15910 2084 15943
rect 2044 15904 2096 15910
rect 2044 15846 2096 15852
rect 1952 15564 2004 15570
rect 1952 15506 2004 15512
rect 1860 15360 1912 15366
rect 1860 15302 1912 15308
rect 1872 13394 1900 15302
rect 1964 14822 1992 15506
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 2044 14544 2096 14550
rect 2044 14486 2096 14492
rect 2056 14074 2084 14486
rect 2148 14414 2176 16748
rect 2320 16730 2372 16736
rect 2424 16674 2452 20198
rect 2608 16726 2636 22918
rect 2792 22409 2820 23530
rect 2778 22400 2834 22409
rect 2778 22335 2834 22344
rect 2688 20256 2740 20262
rect 2688 20198 2740 20204
rect 2332 16646 2452 16674
rect 2596 16720 2648 16726
rect 2596 16662 2648 16668
rect 2332 15201 2360 16646
rect 2412 15360 2464 15366
rect 2412 15302 2464 15308
rect 2596 15360 2648 15366
rect 2596 15302 2648 15308
rect 2318 15192 2374 15201
rect 2318 15127 2374 15136
rect 2228 15088 2280 15094
rect 2228 15030 2280 15036
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2044 14068 2096 14074
rect 2044 14010 2096 14016
rect 2240 13530 2268 15030
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2332 14618 2360 14962
rect 2424 14958 2452 15302
rect 2504 15156 2556 15162
rect 2504 15098 2556 15104
rect 2412 14952 2464 14958
rect 2412 14894 2464 14900
rect 2320 14612 2372 14618
rect 2320 14554 2372 14560
rect 2332 14006 2360 14554
rect 2320 14000 2372 14006
rect 2320 13942 2372 13948
rect 2424 13814 2452 14894
rect 2332 13786 2452 13814
rect 2228 13524 2280 13530
rect 2228 13466 2280 13472
rect 1860 13388 1912 13394
rect 1912 13348 1992 13376
rect 1860 13330 1912 13336
rect 1860 12844 1912 12850
rect 1860 12786 1912 12792
rect 1768 12300 1820 12306
rect 1768 12242 1820 12248
rect 1780 11898 1808 12242
rect 1872 12102 1900 12786
rect 1964 12442 1992 13348
rect 2240 12986 2268 13466
rect 2228 12980 2280 12986
rect 2228 12922 2280 12928
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 2240 12374 2268 12922
rect 2228 12368 2280 12374
rect 2228 12310 2280 12316
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1768 11892 1820 11898
rect 1768 11834 1820 11840
rect 1780 11218 1808 11834
rect 1872 11354 1900 12038
rect 2240 11898 2268 12310
rect 2228 11892 2280 11898
rect 2228 11834 2280 11840
rect 2228 11688 2280 11694
rect 2332 11676 2360 13786
rect 2412 13524 2464 13530
rect 2412 13466 2464 13472
rect 2424 12850 2452 13466
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 2280 11648 2360 11676
rect 2228 11630 2280 11636
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1780 10810 1808 11154
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1872 9926 1900 11290
rect 2136 11076 2188 11082
rect 2188 11036 2268 11064
rect 2136 11018 2188 11024
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 1952 10124 2004 10130
rect 1952 10066 2004 10072
rect 1860 9920 1912 9926
rect 1766 9888 1822 9897
rect 1860 9862 1912 9868
rect 1766 9823 1822 9832
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1412 8486 1624 8514
rect 1216 5908 1268 5914
rect 1216 5850 1268 5856
rect 1412 5166 1440 8486
rect 1492 8424 1544 8430
rect 1492 8366 1544 8372
rect 1504 7818 1532 8366
rect 1582 7984 1638 7993
rect 1582 7919 1638 7928
rect 1492 7812 1544 7818
rect 1492 7754 1544 7760
rect 1596 7546 1624 7919
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1688 7002 1716 8774
rect 1780 7970 1808 9823
rect 1872 9654 1900 9862
rect 1860 9648 1912 9654
rect 1860 9590 1912 9596
rect 1872 8838 1900 9590
rect 1964 9518 1992 10066
rect 2148 10033 2176 10746
rect 2134 10024 2190 10033
rect 2134 9959 2190 9968
rect 2148 9518 2176 9959
rect 2240 9674 2268 11036
rect 2332 10810 2360 11648
rect 2424 11558 2452 12786
rect 2516 12238 2544 15098
rect 2608 14958 2636 15302
rect 2596 14952 2648 14958
rect 2596 14894 2648 14900
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2608 13462 2636 14758
rect 2596 13456 2648 13462
rect 2596 13398 2648 13404
rect 2700 12986 2728 20198
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 2792 14550 2820 17614
rect 2884 16182 2912 27474
rect 3712 27443 3740 27474
rect 5368 23866 5396 27526
rect 6642 27520 6698 28000
rect 8114 27520 8170 28000
rect 9586 27520 9642 28000
rect 11058 27520 11114 28000
rect 12530 27554 12586 28000
rect 12530 27526 12664 27554
rect 12530 27520 12586 27526
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 6656 23866 6684 27520
rect 5356 23860 5408 23866
rect 5356 23802 5408 23808
rect 6644 23860 6696 23866
rect 6644 23802 6696 23808
rect 5368 23662 5396 23802
rect 5356 23656 5408 23662
rect 5356 23598 5408 23604
rect 6184 23656 6236 23662
rect 6184 23598 6236 23604
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 6092 21072 6144 21078
rect 6092 21014 6144 21020
rect 4712 21004 4764 21010
rect 4712 20946 4764 20952
rect 4724 20602 4752 20946
rect 5448 20936 5500 20942
rect 5448 20878 5500 20884
rect 5080 20800 5132 20806
rect 5080 20742 5132 20748
rect 4712 20596 4764 20602
rect 4712 20538 4764 20544
rect 4160 20528 4212 20534
rect 4160 20470 4212 20476
rect 3698 19952 3754 19961
rect 3698 19887 3754 19896
rect 4068 19916 4120 19922
rect 2964 19712 3016 19718
rect 2964 19654 3016 19660
rect 2976 19174 3004 19654
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 3424 19168 3476 19174
rect 3424 19110 3476 19116
rect 2976 16980 3004 19110
rect 3056 18760 3108 18766
rect 3056 18702 3108 18708
rect 3238 18728 3294 18737
rect 3068 18358 3096 18702
rect 3238 18663 3294 18672
rect 3056 18352 3108 18358
rect 3056 18294 3108 18300
rect 3252 18222 3280 18663
rect 3240 18216 3292 18222
rect 3240 18158 3292 18164
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 3160 17134 3188 17478
rect 3148 17128 3200 17134
rect 3148 17070 3200 17076
rect 3240 16992 3292 16998
rect 2976 16952 3188 16980
rect 2872 16176 2924 16182
rect 2872 16118 2924 16124
rect 2964 15904 3016 15910
rect 2964 15846 3016 15852
rect 2976 15706 3004 15846
rect 2964 15700 3016 15706
rect 2964 15642 3016 15648
rect 2964 15564 3016 15570
rect 2964 15506 3016 15512
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 2884 15162 2912 15438
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 2872 14952 2924 14958
rect 2872 14894 2924 14900
rect 2780 14544 2832 14550
rect 2780 14486 2832 14492
rect 2780 14000 2832 14006
rect 2780 13942 2832 13948
rect 2792 13530 2820 13942
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2792 12986 2820 13330
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 2780 12980 2832 12986
rect 2780 12922 2832 12928
rect 2884 12832 2912 14894
rect 2976 14618 3004 15506
rect 3054 15192 3110 15201
rect 3054 15127 3110 15136
rect 2964 14612 3016 14618
rect 2964 14554 3016 14560
rect 2976 13814 3004 14554
rect 3068 14414 3096 15127
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 3160 13814 3188 16952
rect 3240 16934 3292 16940
rect 3252 15706 3280 16934
rect 3332 15972 3384 15978
rect 3332 15914 3384 15920
rect 3240 15700 3292 15706
rect 3240 15642 3292 15648
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 3252 13977 3280 15506
rect 3344 14521 3372 15914
rect 3330 14512 3386 14521
rect 3330 14447 3386 14456
rect 3238 13968 3294 13977
rect 3238 13903 3294 13912
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 2976 13786 3096 13814
rect 3160 13786 3280 13814
rect 2964 13456 3016 13462
rect 2964 13398 3016 13404
rect 2792 12804 2912 12832
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2516 11762 2544 12174
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2412 11552 2464 11558
rect 2412 11494 2464 11500
rect 2516 11286 2544 11698
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2504 11280 2556 11286
rect 2504 11222 2556 11228
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 2424 10674 2452 11154
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2320 10600 2372 10606
rect 2320 10542 2372 10548
rect 2332 10266 2360 10542
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2240 9654 2452 9674
rect 2240 9648 2464 9654
rect 2240 9646 2412 9648
rect 2412 9590 2464 9596
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 2136 9512 2188 9518
rect 2136 9454 2188 9460
rect 1860 8832 1912 8838
rect 1860 8774 1912 8780
rect 1872 8090 1900 8774
rect 1964 8294 1992 9454
rect 2044 9376 2096 9382
rect 2044 9318 2096 9324
rect 2056 9042 2084 9318
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 1952 8288 2004 8294
rect 1952 8230 2004 8236
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 1780 7942 1900 7970
rect 1964 7954 1992 8230
rect 2056 8090 2084 8978
rect 2148 8634 2176 9454
rect 2424 9178 2452 9590
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2516 9042 2544 10406
rect 2608 9586 2636 11494
rect 2792 11393 2820 12804
rect 2870 12744 2926 12753
rect 2870 12679 2926 12688
rect 2884 11898 2912 12679
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2976 11778 3004 13398
rect 2884 11750 3004 11778
rect 2778 11384 2834 11393
rect 2778 11319 2834 11328
rect 2792 11218 2820 11319
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2688 11076 2740 11082
rect 2688 11018 2740 11024
rect 2700 9722 2728 11018
rect 2884 9897 2912 11750
rect 3068 10810 3096 13786
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3160 12782 3188 13126
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 2870 9888 2926 9897
rect 2870 9823 2926 9832
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2504 9036 2556 9042
rect 2504 8978 2556 8984
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 1768 7268 1820 7274
rect 1768 7210 1820 7216
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1582 6760 1638 6769
rect 1582 6695 1638 6704
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 1504 5778 1532 6258
rect 1492 5772 1544 5778
rect 1492 5714 1544 5720
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 1124 4820 1176 4826
rect 1124 4762 1176 4768
rect 1504 4282 1532 5714
rect 1596 5370 1624 6695
rect 1688 6254 1716 6938
rect 1780 6458 1808 7210
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1584 5364 1636 5370
rect 1584 5306 1636 5312
rect 1492 4276 1544 4282
rect 1492 4218 1544 4224
rect 1768 4004 1820 4010
rect 1768 3946 1820 3952
rect 478 54 888 82
rect 1490 82 1546 480
rect 1780 82 1808 3946
rect 1872 2417 1900 7942
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 1964 7546 1992 7890
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 2136 7200 2188 7206
rect 2136 7142 2188 7148
rect 2148 6866 2176 7142
rect 2516 6934 2544 8978
rect 2608 8809 2636 9522
rect 3068 9489 3096 10610
rect 3160 9926 3188 11222
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3054 9480 3110 9489
rect 3054 9415 3110 9424
rect 3146 9344 3202 9353
rect 3146 9279 3202 9288
rect 2594 8800 2650 8809
rect 2594 8735 2650 8744
rect 2608 8294 2636 8735
rect 3160 8634 3188 9279
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 2872 8288 2924 8294
rect 2872 8230 2924 8236
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2700 7478 2728 7890
rect 2688 7472 2740 7478
rect 2688 7414 2740 7420
rect 2412 6928 2464 6934
rect 2412 6870 2464 6876
rect 2504 6928 2556 6934
rect 2504 6870 2556 6876
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 2148 5914 2176 6802
rect 2424 6118 2452 6870
rect 2516 6798 2544 6870
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2504 6180 2556 6186
rect 2504 6122 2556 6128
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 1950 5400 2006 5409
rect 1950 5335 2006 5344
rect 2412 5364 2464 5370
rect 1964 4690 1992 5335
rect 2412 5306 2464 5312
rect 1952 4684 2004 4690
rect 1952 4626 2004 4632
rect 1964 4282 1992 4626
rect 1952 4276 2004 4282
rect 1952 4218 2004 4224
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 1964 3194 1992 3538
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 1858 2408 1914 2417
rect 1858 2343 1914 2352
rect 1490 54 1808 82
rect 2424 82 2452 5306
rect 2516 4826 2544 6122
rect 2884 5914 2912 8230
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2976 7206 3004 7890
rect 3160 7342 3188 8026
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2976 7002 3004 7142
rect 2964 6996 3016 7002
rect 2964 6938 3016 6944
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 3068 6458 3096 6598
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 2964 6180 3016 6186
rect 3068 6168 3096 6394
rect 3016 6140 3096 6168
rect 2964 6122 3016 6128
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 2964 5636 3016 5642
rect 2964 5578 3016 5584
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2976 4690 3004 5578
rect 3068 5370 3096 5714
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 2594 4312 2650 4321
rect 2594 4247 2650 4256
rect 2608 4146 2636 4247
rect 2976 4214 3004 4626
rect 2964 4208 3016 4214
rect 2778 4176 2834 4185
rect 2596 4140 2648 4146
rect 2964 4150 3016 4156
rect 2778 4111 2834 4120
rect 2596 4082 2648 4088
rect 2792 2650 2820 4111
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 2516 2310 2544 2450
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 2516 1737 2544 2246
rect 2502 1728 2558 1737
rect 2502 1663 2558 1672
rect 2502 82 2558 480
rect 2424 54 2558 82
rect 3252 82 3280 13786
rect 3344 12646 3372 13874
rect 3332 12640 3384 12646
rect 3332 12582 3384 12588
rect 3332 12436 3384 12442
rect 3332 12378 3384 12384
rect 3344 12209 3372 12378
rect 3330 12200 3386 12209
rect 3330 12135 3386 12144
rect 3332 11824 3384 11830
rect 3332 11766 3384 11772
rect 3344 11082 3372 11766
rect 3332 11076 3384 11082
rect 3332 11018 3384 11024
rect 3344 10742 3372 11018
rect 3332 10736 3384 10742
rect 3332 10678 3384 10684
rect 3436 10554 3464 19110
rect 3516 17808 3568 17814
rect 3516 17750 3568 17756
rect 3528 17338 3556 17750
rect 3608 17740 3660 17746
rect 3608 17682 3660 17688
rect 3516 17332 3568 17338
rect 3516 17274 3568 17280
rect 3620 16998 3648 17682
rect 3608 16992 3660 16998
rect 3608 16934 3660 16940
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 3528 16046 3556 16730
rect 3516 16040 3568 16046
rect 3516 15982 3568 15988
rect 3528 13326 3556 15982
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 3528 12918 3556 13262
rect 3516 12912 3568 12918
rect 3516 12854 3568 12860
rect 3516 12776 3568 12782
rect 3516 12718 3568 12724
rect 3528 12646 3556 12718
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3344 10526 3464 10554
rect 3344 7721 3372 10526
rect 3422 9752 3478 9761
rect 3422 9687 3478 9696
rect 3436 9382 3464 9687
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3436 9178 3464 9318
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3424 8900 3476 8906
rect 3424 8842 3476 8848
rect 3436 7954 3464 8842
rect 3528 8090 3556 12582
rect 3620 12442 3648 16934
rect 3712 16590 3740 19887
rect 4068 19858 4120 19864
rect 3792 19712 3844 19718
rect 3792 19654 3844 19660
rect 3884 19712 3936 19718
rect 3884 19654 3936 19660
rect 3700 16584 3752 16590
rect 3700 16526 3752 16532
rect 3700 15972 3752 15978
rect 3700 15914 3752 15920
rect 3712 15502 3740 15914
rect 3700 15496 3752 15502
rect 3700 15438 3752 15444
rect 3700 14000 3752 14006
rect 3700 13942 3752 13948
rect 3712 13530 3740 13942
rect 3804 13814 3832 19654
rect 3896 17882 3924 19654
rect 4080 19242 4108 19858
rect 4068 19236 4120 19242
rect 4068 19178 4120 19184
rect 4172 18222 4200 20470
rect 4896 20256 4948 20262
rect 4896 20198 4948 20204
rect 4436 19168 4488 19174
rect 4436 19110 4488 19116
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 4344 18624 4396 18630
rect 4344 18566 4396 18572
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 3884 17876 3936 17882
rect 3884 17818 3936 17824
rect 3896 17116 3924 17818
rect 4172 17814 4200 18158
rect 4160 17808 4212 17814
rect 4160 17750 4212 17756
rect 4160 17536 4212 17542
rect 4160 17478 4212 17484
rect 3976 17128 4028 17134
rect 3896 17088 3976 17116
rect 3976 17070 4028 17076
rect 3976 16992 4028 16998
rect 3976 16934 4028 16940
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3896 15910 3924 16526
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3896 15570 3924 15846
rect 3884 15564 3936 15570
rect 3884 15506 3936 15512
rect 3988 14958 4016 16934
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 4080 16182 4108 16390
rect 4172 16250 4200 17478
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 3976 14952 4028 14958
rect 3896 14912 3976 14940
rect 3896 14618 3924 14912
rect 3976 14894 4028 14900
rect 3884 14612 3936 14618
rect 3884 14554 3936 14560
rect 3896 14006 3924 14554
rect 3976 14544 4028 14550
rect 3976 14486 4028 14492
rect 3884 14000 3936 14006
rect 3884 13942 3936 13948
rect 3988 13938 4016 14486
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 3804 13786 3924 13814
rect 3700 13524 3752 13530
rect 3700 13466 3752 13472
rect 3712 12782 3740 13466
rect 3896 12889 3924 13786
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 3882 12880 3938 12889
rect 3882 12815 3938 12824
rect 3700 12776 3752 12782
rect 3700 12718 3752 12724
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3988 12374 4016 13126
rect 3792 12368 3844 12374
rect 3792 12310 3844 12316
rect 3976 12368 4028 12374
rect 3976 12310 4028 12316
rect 3700 12300 3752 12306
rect 3700 12242 3752 12248
rect 3712 11830 3740 12242
rect 3700 11824 3752 11830
rect 3700 11766 3752 11772
rect 3608 11620 3660 11626
rect 3608 11562 3660 11568
rect 3620 11286 3648 11562
rect 3700 11348 3752 11354
rect 3700 11290 3752 11296
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3620 9353 3648 11086
rect 3712 10742 3740 11290
rect 3700 10736 3752 10742
rect 3700 10678 3752 10684
rect 3804 10606 3832 12310
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3896 11694 3924 12038
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 3896 11354 3924 11630
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 3884 11008 3936 11014
rect 3884 10950 3936 10956
rect 3792 10600 3844 10606
rect 3792 10542 3844 10548
rect 3700 10464 3752 10470
rect 3700 10406 3752 10412
rect 3712 9625 3740 10406
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3698 9616 3754 9625
rect 3698 9551 3754 9560
rect 3700 9444 3752 9450
rect 3700 9386 3752 9392
rect 3606 9344 3662 9353
rect 3606 9279 3662 9288
rect 3712 9178 3740 9386
rect 3700 9172 3752 9178
rect 3700 9114 3752 9120
rect 3804 8974 3832 9998
rect 3896 9110 3924 10950
rect 3988 10470 4016 11154
rect 4080 10826 4108 16118
rect 4160 16108 4212 16114
rect 4160 16050 4212 16056
rect 4172 15638 4200 16050
rect 4160 15632 4212 15638
rect 4160 15574 4212 15580
rect 4160 14884 4212 14890
rect 4160 14826 4212 14832
rect 4172 11257 4200 14826
rect 4356 14278 4384 18566
rect 4448 15094 4476 19110
rect 4528 18828 4580 18834
rect 4528 18770 4580 18776
rect 4540 18358 4568 18770
rect 4528 18352 4580 18358
rect 4528 18294 4580 18300
rect 4528 17740 4580 17746
rect 4528 17682 4580 17688
rect 4540 16998 4568 17682
rect 4528 16992 4580 16998
rect 4528 16934 4580 16940
rect 4620 16516 4672 16522
rect 4620 16458 4672 16464
rect 4528 15564 4580 15570
rect 4528 15506 4580 15512
rect 4540 15162 4568 15506
rect 4528 15156 4580 15162
rect 4528 15098 4580 15104
rect 4436 15088 4488 15094
rect 4436 15030 4488 15036
rect 4528 14544 4580 14550
rect 4528 14486 4580 14492
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 4540 14074 4568 14486
rect 4632 14074 4660 16458
rect 4528 14068 4580 14074
rect 4528 14010 4580 14016
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4620 13864 4672 13870
rect 4526 13832 4582 13841
rect 4344 13796 4396 13802
rect 4620 13806 4672 13812
rect 4526 13767 4582 13776
rect 4344 13738 4396 13744
rect 4356 13394 4384 13738
rect 4436 13524 4488 13530
rect 4436 13466 4488 13472
rect 4448 13394 4476 13466
rect 4344 13388 4396 13394
rect 4344 13330 4396 13336
rect 4436 13388 4488 13394
rect 4436 13330 4488 13336
rect 4356 12986 4384 13330
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 4252 12912 4304 12918
rect 4252 12854 4304 12860
rect 4264 11286 4292 12854
rect 4540 12102 4568 13767
rect 4632 13394 4660 13806
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4528 12096 4580 12102
rect 4528 12038 4580 12044
rect 4356 11898 4384 12038
rect 4344 11892 4396 11898
rect 4344 11834 4396 11840
rect 4356 11626 4384 11834
rect 4344 11620 4396 11626
rect 4344 11562 4396 11568
rect 4252 11280 4304 11286
rect 4158 11248 4214 11257
rect 4252 11222 4304 11228
rect 4158 11183 4214 11192
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4080 10798 4200 10826
rect 4080 10742 4108 10798
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 4068 10532 4120 10538
rect 4068 10474 4120 10480
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3976 10192 4028 10198
rect 3976 10134 4028 10140
rect 3988 9518 4016 10134
rect 4080 10130 4108 10474
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 4172 10062 4200 10798
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4172 9761 4200 9998
rect 4264 9926 4292 11086
rect 4356 11014 4384 11562
rect 4436 11552 4488 11558
rect 4436 11494 4488 11500
rect 4448 11150 4476 11494
rect 4436 11144 4488 11150
rect 4436 11086 4488 11092
rect 4344 11008 4396 11014
rect 4344 10950 4396 10956
rect 4356 10810 4384 10950
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4448 10062 4476 11086
rect 4724 10266 4752 19110
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 4816 15366 4844 16594
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 4816 11898 4844 15302
rect 4908 14958 4936 20198
rect 4988 18624 5040 18630
rect 4988 18566 5040 18572
rect 5000 18222 5028 18566
rect 4988 18216 5040 18222
rect 4988 18158 5040 18164
rect 4988 17264 5040 17270
rect 4988 17206 5040 17212
rect 5000 16454 5028 17206
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 4988 15632 5040 15638
rect 4988 15574 5040 15580
rect 4896 14952 4948 14958
rect 4896 14894 4948 14900
rect 4908 14793 4936 14894
rect 4894 14784 4950 14793
rect 4894 14719 4950 14728
rect 4896 14000 4948 14006
rect 4896 13942 4948 13948
rect 4908 12186 4936 13942
rect 5000 12306 5028 15574
rect 5092 12442 5120 20742
rect 5460 20534 5488 20878
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5448 20528 5500 20534
rect 5448 20470 5500 20476
rect 5460 20398 5488 20470
rect 5448 20392 5500 20398
rect 5448 20334 5500 20340
rect 5460 20058 5488 20334
rect 5632 20324 5684 20330
rect 5632 20266 5684 20272
rect 5448 20052 5500 20058
rect 5448 19994 5500 20000
rect 5644 19922 5672 20266
rect 6104 20262 6132 21014
rect 6092 20256 6144 20262
rect 6092 20198 6144 20204
rect 5816 19984 5868 19990
rect 5816 19926 5868 19932
rect 5632 19916 5684 19922
rect 5552 19876 5632 19904
rect 5264 19848 5316 19854
rect 5264 19790 5316 19796
rect 5276 19378 5304 19790
rect 5552 19514 5580 19876
rect 5632 19858 5684 19864
rect 5828 19825 5856 19926
rect 5814 19816 5870 19825
rect 5814 19751 5870 19760
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5540 19508 5592 19514
rect 5540 19450 5592 19456
rect 5264 19372 5316 19378
rect 5264 19314 5316 19320
rect 6000 19304 6052 19310
rect 6000 19246 6052 19252
rect 5356 19236 5408 19242
rect 5356 19178 5408 19184
rect 5368 18834 5396 19178
rect 6012 18970 6040 19246
rect 6000 18964 6052 18970
rect 6000 18906 6052 18912
rect 5356 18828 5408 18834
rect 5356 18770 5408 18776
rect 5448 18760 5500 18766
rect 5448 18702 5500 18708
rect 5460 18290 5488 18702
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5448 18284 5500 18290
rect 5448 18226 5500 18232
rect 5264 18216 5316 18222
rect 5264 18158 5316 18164
rect 5276 17882 5304 18158
rect 6012 18086 6040 18906
rect 6104 18358 6132 20198
rect 6196 18902 6224 23598
rect 7196 23520 7248 23526
rect 7196 23462 7248 23468
rect 7104 22092 7156 22098
rect 7104 22034 7156 22040
rect 7116 21350 7144 22034
rect 6920 21344 6972 21350
rect 6920 21286 6972 21292
rect 7104 21344 7156 21350
rect 7104 21286 7156 21292
rect 6828 20936 6880 20942
rect 6828 20878 6880 20884
rect 6840 20466 6868 20878
rect 6828 20460 6880 20466
rect 6828 20402 6880 20408
rect 6644 20324 6696 20330
rect 6644 20266 6696 20272
rect 6656 19990 6684 20266
rect 6932 19990 6960 21286
rect 6644 19984 6696 19990
rect 6644 19926 6696 19932
rect 6920 19984 6972 19990
rect 6920 19926 6972 19932
rect 6274 19680 6330 19689
rect 6274 19615 6330 19624
rect 6184 18896 6236 18902
rect 6184 18838 6236 18844
rect 6196 18601 6224 18838
rect 6182 18592 6238 18601
rect 6182 18527 6238 18536
rect 6092 18352 6144 18358
rect 6092 18294 6144 18300
rect 6000 18080 6052 18086
rect 6000 18022 6052 18028
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 5276 17134 5304 17818
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5540 17264 5592 17270
rect 5540 17206 5592 17212
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 5172 16992 5224 16998
rect 5172 16934 5224 16940
rect 5184 16114 5212 16934
rect 5276 16794 5304 17070
rect 5264 16788 5316 16794
rect 5264 16730 5316 16736
rect 5172 16108 5224 16114
rect 5172 16050 5224 16056
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 5276 15570 5304 15846
rect 5264 15564 5316 15570
rect 5264 15506 5316 15512
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5184 13938 5212 14758
rect 5276 14618 5304 15506
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5368 13977 5396 15982
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5460 14958 5488 15642
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 5552 14482 5580 17206
rect 6012 17202 6040 17614
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 6104 17082 6132 18294
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 6196 17882 6224 18022
rect 6184 17876 6236 17882
rect 6184 17818 6236 17824
rect 6012 17054 6132 17082
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5724 14884 5776 14890
rect 5724 14826 5776 14832
rect 5540 14476 5592 14482
rect 5460 14436 5540 14464
rect 5354 13968 5410 13977
rect 5172 13932 5224 13938
rect 5354 13903 5410 13912
rect 5172 13874 5224 13880
rect 5460 13734 5488 14436
rect 5540 14418 5592 14424
rect 5736 14414 5764 14826
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5448 13728 5500 13734
rect 5170 13696 5226 13705
rect 5448 13670 5500 13676
rect 5170 13631 5226 13640
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 5078 12336 5134 12345
rect 4988 12300 5040 12306
rect 5184 12322 5212 13631
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5134 12294 5212 12322
rect 5356 12300 5408 12306
rect 5078 12271 5134 12280
rect 4988 12242 5040 12248
rect 4908 12158 5028 12186
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4802 11792 4858 11801
rect 4802 11727 4858 11736
rect 4816 11286 4844 11727
rect 4804 11280 4856 11286
rect 4804 11222 4856 11228
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4618 10160 4674 10169
rect 4618 10095 4674 10104
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 4158 9752 4214 9761
rect 4158 9687 4160 9696
rect 4212 9687 4214 9696
rect 4160 9658 4212 9664
rect 4264 9654 4292 9862
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 4342 9616 4398 9625
rect 4068 9580 4120 9586
rect 4632 9586 4660 10095
rect 4908 9674 4936 12038
rect 5000 11014 5028 12158
rect 4988 11008 5040 11014
rect 4988 10950 5040 10956
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 4724 9646 4936 9674
rect 4342 9551 4398 9560
rect 4620 9580 4672 9586
rect 4068 9522 4120 9528
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3884 9104 3936 9110
rect 3988 9081 4016 9454
rect 3884 9046 3936 9052
rect 3974 9072 4030 9081
rect 3974 9007 4030 9016
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3608 8016 3660 8022
rect 3608 7958 3660 7964
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 3330 7712 3386 7721
rect 3330 7647 3386 7656
rect 3332 7268 3384 7274
rect 3332 7210 3384 7216
rect 3344 6780 3372 7210
rect 3436 7002 3464 7890
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 3424 6792 3476 6798
rect 3344 6752 3424 6780
rect 3424 6734 3476 6740
rect 3436 6662 3464 6734
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3332 6248 3384 6254
rect 3332 6190 3384 6196
rect 3344 3602 3372 6190
rect 3436 5166 3464 6598
rect 3528 5914 3556 7822
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3424 5160 3476 5166
rect 3424 5102 3476 5108
rect 3436 3602 3464 5102
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 3344 3194 3372 3538
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3528 2990 3556 4082
rect 3620 4078 3648 7958
rect 3700 7812 3752 7818
rect 3804 7800 3832 8910
rect 3896 8566 3924 8910
rect 4080 8838 4108 9522
rect 4356 9518 4384 9551
rect 4620 9522 4672 9528
rect 4344 9512 4396 9518
rect 4344 9454 4396 9460
rect 4342 9344 4398 9353
rect 4342 9279 4398 9288
rect 4356 9110 4384 9279
rect 4344 9104 4396 9110
rect 4344 9046 4396 9052
rect 4436 8968 4488 8974
rect 4342 8936 4398 8945
rect 4160 8900 4212 8906
rect 4436 8910 4488 8916
rect 4342 8871 4398 8880
rect 4160 8842 4212 8848
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 3884 8560 3936 8566
rect 4080 8548 4108 8774
rect 4172 8566 4200 8842
rect 4356 8838 4384 8871
rect 4344 8832 4396 8838
rect 4448 8809 4476 8910
rect 4528 8832 4580 8838
rect 4344 8774 4396 8780
rect 4434 8800 4490 8809
rect 4356 8634 4384 8774
rect 4528 8774 4580 8780
rect 4434 8735 4490 8744
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4160 8560 4212 8566
rect 3936 8520 4016 8548
rect 4080 8520 4160 8548
rect 3884 8502 3936 8508
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3752 7772 3832 7800
rect 3700 7754 3752 7760
rect 3698 7712 3754 7721
rect 3698 7647 3754 7656
rect 3712 7410 3740 7647
rect 3700 7404 3752 7410
rect 3700 7346 3752 7352
rect 3792 6724 3844 6730
rect 3792 6666 3844 6672
rect 3804 6322 3832 6666
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3712 5166 3740 5510
rect 3790 5400 3846 5409
rect 3790 5335 3846 5344
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3712 4826 3740 5102
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3608 4072 3660 4078
rect 3804 4026 3832 5335
rect 3896 4154 3924 8230
rect 3988 7750 4016 8520
rect 4160 8502 4212 8508
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 4080 7546 4108 8026
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4068 7200 4120 7206
rect 4172 7188 4200 7822
rect 4356 7750 4384 8298
rect 4436 8016 4488 8022
rect 4436 7958 4488 7964
rect 4448 7886 4476 7958
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 4120 7160 4200 7188
rect 4068 7142 4120 7148
rect 4080 6118 4108 7142
rect 4264 7002 4292 7278
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4264 6798 4292 6938
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4080 5846 4108 6054
rect 4356 5914 4384 7686
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4448 6322 4476 7142
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 4080 5030 4108 5782
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 4172 5234 4200 5646
rect 4160 5228 4212 5234
rect 4540 5216 4568 8774
rect 4724 8616 4752 9646
rect 4632 8588 4752 8616
rect 4632 5409 4660 8588
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4724 7206 4752 8434
rect 4896 8356 4948 8362
rect 4896 8298 4948 8304
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4618 5400 4674 5409
rect 4618 5335 4674 5344
rect 4160 5170 4212 5176
rect 4448 5188 4568 5216
rect 4620 5228 4672 5234
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 3896 4126 4016 4154
rect 4080 4146 4108 4966
rect 4172 4826 4200 5170
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4264 4146 4292 4422
rect 3608 4014 3660 4020
rect 3712 3998 3832 4026
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3712 2650 3740 3998
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3804 3233 3832 3878
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3790 3224 3846 3233
rect 3790 3159 3846 3168
rect 3700 2644 3752 2650
rect 3700 2586 3752 2592
rect 3896 2582 3924 3334
rect 3988 3058 4016 4126
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4080 3924 4108 4082
rect 4160 3936 4212 3942
rect 4080 3896 4160 3924
rect 4160 3878 4212 3884
rect 4264 3738 4292 4082
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4448 3670 4476 5188
rect 4620 5170 4672 5176
rect 4528 5092 4580 5098
rect 4528 5034 4580 5040
rect 4436 3664 4488 3670
rect 4436 3606 4488 3612
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4172 3194 4200 3538
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 3988 2961 4016 2994
rect 3974 2952 4030 2961
rect 3974 2887 4030 2896
rect 4356 2650 4384 3538
rect 4540 3466 4568 5034
rect 4632 4758 4660 5170
rect 4620 4752 4672 4758
rect 4620 4694 4672 4700
rect 4528 3460 4580 3466
rect 4528 3402 4580 3408
rect 4724 2922 4752 7142
rect 4816 6662 4844 7278
rect 4908 6730 4936 8298
rect 4896 6724 4948 6730
rect 4896 6666 4948 6672
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 4816 5098 4844 6598
rect 5000 5778 5028 10610
rect 5092 9518 5120 12271
rect 5356 12242 5408 12248
rect 5368 12209 5396 12242
rect 5354 12200 5410 12209
rect 5354 12135 5410 12144
rect 5368 11694 5396 12135
rect 5460 11694 5488 12786
rect 5540 12368 5592 12374
rect 5540 12310 5592 12316
rect 5552 11898 5580 12310
rect 6012 12306 6040 17054
rect 6092 16992 6144 16998
rect 6196 16980 6224 17818
rect 6144 16952 6224 16980
rect 6092 16934 6144 16940
rect 6104 15552 6132 16934
rect 6184 16720 6236 16726
rect 6184 16662 6236 16668
rect 6196 16250 6224 16662
rect 6184 16244 6236 16250
rect 6184 16186 6236 16192
rect 6196 15706 6224 16186
rect 6288 15978 6316 19615
rect 7116 19446 7144 21286
rect 7104 19440 7156 19446
rect 7104 19382 7156 19388
rect 6828 19236 6880 19242
rect 6828 19178 6880 19184
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 6748 17882 6776 18226
rect 6736 17876 6788 17882
rect 6736 17818 6788 17824
rect 6460 17060 6512 17066
rect 6460 17002 6512 17008
rect 6368 16040 6420 16046
rect 6368 15982 6420 15988
rect 6276 15972 6328 15978
rect 6276 15914 6328 15920
rect 6380 15706 6408 15982
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6368 15700 6420 15706
rect 6368 15642 6420 15648
rect 6184 15564 6236 15570
rect 6104 15524 6184 15552
rect 6184 15506 6236 15512
rect 6196 14822 6224 15506
rect 6184 14816 6236 14822
rect 6184 14758 6236 14764
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 6104 13530 6132 14418
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 6380 13938 6408 14350
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6276 13728 6328 13734
rect 6276 13670 6328 13676
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6104 12782 6132 13466
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 6196 12850 6224 13126
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 6092 12776 6144 12782
rect 6092 12718 6144 12724
rect 6104 12306 6132 12718
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6012 11898 6040 12242
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 5816 11824 5868 11830
rect 5816 11766 5868 11772
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5460 11336 5488 11630
rect 5828 11354 5856 11766
rect 6104 11354 6132 12242
rect 5368 11308 5488 11336
rect 5540 11348 5592 11354
rect 5172 11008 5224 11014
rect 5172 10950 5224 10956
rect 5184 9674 5212 10950
rect 5368 10810 5396 11308
rect 5540 11290 5592 11296
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5356 10804 5408 10810
rect 5276 10764 5356 10792
rect 5276 10606 5304 10764
rect 5356 10746 5408 10752
rect 5460 10674 5488 11154
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 5368 9994 5396 10474
rect 5552 10266 5580 11290
rect 6288 11234 6316 13670
rect 6366 11384 6422 11393
rect 6366 11319 6422 11328
rect 6380 11286 6408 11319
rect 6196 11206 6316 11234
rect 6368 11280 6420 11286
rect 6368 11222 6420 11228
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5356 9988 5408 9994
rect 5356 9930 5408 9936
rect 5368 9897 5396 9930
rect 5354 9888 5410 9897
rect 5354 9823 5410 9832
rect 5184 9646 5396 9674
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 5092 5642 5120 9454
rect 5368 7478 5396 9646
rect 5460 8634 5488 10134
rect 5644 10033 5672 10406
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 5630 10024 5686 10033
rect 5630 9959 5686 9968
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6012 9178 6040 10066
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5736 8090 5764 8366
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 6092 8016 6144 8022
rect 6092 7958 6144 7964
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5356 7472 5408 7478
rect 5356 7414 5408 7420
rect 5368 7313 5396 7414
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5354 7304 5410 7313
rect 5354 7239 5410 7248
rect 5172 6928 5224 6934
rect 5172 6870 5224 6876
rect 5184 6458 5212 6870
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5184 5914 5212 6394
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5080 5636 5132 5642
rect 5080 5578 5132 5584
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 4908 5098 4936 5306
rect 4804 5092 4856 5098
rect 4804 5034 4856 5040
rect 4896 5092 4948 5098
rect 4896 5034 4948 5040
rect 4908 4758 4936 5034
rect 4896 4752 4948 4758
rect 4896 4694 4948 4700
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4816 3194 4844 4558
rect 4908 4282 4936 4694
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 5356 3460 5408 3466
rect 5356 3402 5408 3408
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 5092 3194 5120 3334
rect 5368 3210 5396 3402
rect 5460 3398 5488 7346
rect 6104 7002 6132 7958
rect 6092 6996 6144 7002
rect 6092 6938 6144 6944
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5552 6390 5580 6734
rect 6196 6662 6224 11206
rect 6472 10130 6500 17002
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6564 14550 6592 15302
rect 6736 14952 6788 14958
rect 6736 14894 6788 14900
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 6552 14544 6604 14550
rect 6552 14486 6604 14492
rect 6552 13796 6604 13802
rect 6656 13784 6684 14758
rect 6604 13756 6684 13784
rect 6552 13738 6604 13744
rect 6564 13462 6592 13738
rect 6552 13456 6604 13462
rect 6552 13398 6604 13404
rect 6564 12986 6592 13398
rect 6748 13326 6776 14894
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6564 12850 6592 12922
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6840 12306 6868 19178
rect 7104 18216 7156 18222
rect 7104 18158 7156 18164
rect 7116 17882 7144 18158
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 7208 16697 7236 23462
rect 8128 22778 8156 27520
rect 9600 23866 9628 27520
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 9588 23860 9640 23866
rect 9588 23802 9640 23808
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 9588 23316 9640 23322
rect 9588 23258 9640 23264
rect 8116 22772 8168 22778
rect 8116 22714 8168 22720
rect 8024 22704 8076 22710
rect 8024 22646 8076 22652
rect 8758 22672 8814 22681
rect 7472 22568 7524 22574
rect 7472 22510 7524 22516
rect 7484 22234 7512 22510
rect 7840 22500 7892 22506
rect 7840 22442 7892 22448
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 7656 20324 7708 20330
rect 7656 20266 7708 20272
rect 7288 20052 7340 20058
rect 7288 19994 7340 20000
rect 7300 19242 7328 19994
rect 7472 19984 7524 19990
rect 7472 19926 7524 19932
rect 7564 19984 7616 19990
rect 7564 19926 7616 19932
rect 7484 19514 7512 19926
rect 7576 19786 7604 19926
rect 7564 19780 7616 19786
rect 7564 19722 7616 19728
rect 7472 19508 7524 19514
rect 7472 19450 7524 19456
rect 7288 19236 7340 19242
rect 7288 19178 7340 19184
rect 7576 18970 7604 19722
rect 7564 18964 7616 18970
rect 7564 18906 7616 18912
rect 7668 18154 7696 20266
rect 7748 20256 7800 20262
rect 7748 20198 7800 20204
rect 7760 20058 7788 20198
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 7852 19334 7880 22442
rect 7932 21344 7984 21350
rect 7932 21286 7984 21292
rect 7944 21078 7972 21286
rect 7932 21072 7984 21078
rect 7932 21014 7984 21020
rect 7944 20058 7972 21014
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 7760 19306 7880 19334
rect 7656 18148 7708 18154
rect 7656 18090 7708 18096
rect 7564 17740 7616 17746
rect 7564 17682 7616 17688
rect 7470 17232 7526 17241
rect 7470 17167 7526 17176
rect 7484 17134 7512 17167
rect 7288 17128 7340 17134
rect 7288 17070 7340 17076
rect 7472 17128 7524 17134
rect 7472 17070 7524 17076
rect 7194 16688 7250 16697
rect 7194 16623 7250 16632
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 6920 15088 6972 15094
rect 6920 15030 6972 15036
rect 6932 14890 6960 15030
rect 7024 14890 7052 15302
rect 7116 15026 7144 15438
rect 7196 15428 7248 15434
rect 7196 15370 7248 15376
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 6920 14884 6972 14890
rect 6920 14826 6972 14832
rect 7012 14884 7064 14890
rect 7012 14826 7064 14832
rect 7024 14618 7052 14826
rect 7116 14618 7144 14962
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7010 13968 7066 13977
rect 7010 13903 7066 13912
rect 7024 12986 7052 13903
rect 7208 13190 7236 15370
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 7024 12442 7052 12650
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6656 11218 6684 12174
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6748 10810 6776 11222
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 6748 10538 6776 10746
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 7116 10198 7144 10610
rect 7196 10532 7248 10538
rect 7196 10474 7248 10480
rect 7208 10266 7236 10474
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 6380 9382 6408 10066
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6472 9178 6500 10066
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6748 9489 6776 9522
rect 7208 9518 7236 10066
rect 7196 9512 7248 9518
rect 6734 9480 6790 9489
rect 7196 9454 7248 9460
rect 6734 9415 6790 9424
rect 6748 9178 6776 9415
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 6458 9072 6514 9081
rect 6458 9007 6460 9016
rect 6512 9007 6514 9016
rect 6736 9036 6788 9042
rect 6460 8978 6512 8984
rect 6736 8978 6788 8984
rect 6368 8900 6420 8906
rect 6368 8842 6420 8848
rect 6380 8362 6408 8842
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 6380 7954 6408 8298
rect 6472 8294 6500 8978
rect 6748 8634 6776 8978
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6460 8288 6512 8294
rect 6460 8230 6512 8236
rect 6642 7984 6698 7993
rect 6368 7948 6420 7954
rect 6642 7919 6698 7928
rect 6736 7948 6788 7954
rect 6368 7890 6420 7896
rect 6368 7812 6420 7818
rect 6368 7754 6420 7760
rect 6276 7268 6328 7274
rect 6276 7210 6328 7216
rect 6288 6866 6316 7210
rect 6380 7206 6408 7754
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6288 6458 6316 6802
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 5552 5914 5580 6326
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5552 5302 5580 5850
rect 6000 5840 6052 5846
rect 6000 5782 6052 5788
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6012 5370 6040 5782
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6000 5364 6052 5370
rect 6000 5306 6052 5312
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 6104 4758 6132 5646
rect 6092 4752 6144 4758
rect 5538 4720 5594 4729
rect 6092 4694 6144 4700
rect 5538 4655 5594 4664
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5446 3224 5502 3233
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 5080 3188 5132 3194
rect 5368 3182 5446 3210
rect 5446 3159 5502 3168
rect 5080 3130 5132 3136
rect 5460 2990 5488 3159
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 4712 2916 4764 2922
rect 4712 2858 4764 2864
rect 4896 2848 4948 2854
rect 4896 2790 4948 2796
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 3884 2576 3936 2582
rect 3884 2518 3936 2524
rect 4356 2310 4384 2586
rect 4344 2304 4396 2310
rect 4344 2246 4396 2252
rect 4908 2038 4936 2790
rect 4896 2032 4948 2038
rect 4896 1974 4948 1980
rect 3514 82 3570 480
rect 3252 54 3570 82
rect 478 0 534 54
rect 1490 0 1546 54
rect 2502 0 2558 54
rect 3514 0 3570 54
rect 4618 82 4674 480
rect 4908 82 4936 1974
rect 4618 54 4936 82
rect 5552 82 5580 4655
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6288 2650 6316 4082
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 6184 2576 6236 2582
rect 6184 2518 6236 2524
rect 6196 2417 6224 2518
rect 6182 2408 6238 2417
rect 6092 2372 6144 2378
rect 6182 2343 6238 2352
rect 6092 2314 6144 2320
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6104 2145 6132 2314
rect 6090 2136 6146 2145
rect 6090 2071 6146 2080
rect 6380 1193 6408 7142
rect 6460 6724 6512 6730
rect 6460 6666 6512 6672
rect 6472 5710 6500 6666
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6656 4154 6684 7919
rect 6736 7890 6788 7896
rect 6748 6934 6776 7890
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6840 6458 6868 6802
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6840 6322 6868 6394
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6932 6254 6960 8910
rect 7024 6866 7052 9114
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7208 7546 7236 8570
rect 7300 7546 7328 17070
rect 7576 16794 7604 17682
rect 7656 17128 7708 17134
rect 7656 17070 7708 17076
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7668 16726 7696 17070
rect 7656 16720 7708 16726
rect 7656 16662 7708 16668
rect 7380 16584 7432 16590
rect 7380 16526 7432 16532
rect 7392 15026 7420 16526
rect 7472 15972 7524 15978
rect 7472 15914 7524 15920
rect 7564 15972 7616 15978
rect 7564 15914 7616 15920
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7392 14618 7420 14962
rect 7484 14929 7512 15914
rect 7576 15706 7604 15914
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7470 14920 7526 14929
rect 7470 14855 7526 14864
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7392 13841 7420 14554
rect 7378 13832 7434 13841
rect 7378 13767 7434 13776
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7392 11558 7420 12174
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7392 9586 7420 11494
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7392 7818 7420 8366
rect 7380 7812 7432 7818
rect 7380 7754 7432 7760
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7484 7002 7512 14855
rect 7656 14544 7708 14550
rect 7656 14486 7708 14492
rect 7668 13530 7696 14486
rect 7760 13705 7788 19306
rect 8036 18426 8064 22646
rect 8758 22607 8814 22616
rect 8576 22092 8628 22098
rect 8576 22034 8628 22040
rect 8208 21888 8260 21894
rect 8208 21830 8260 21836
rect 8116 21344 8168 21350
rect 8116 21286 8168 21292
rect 8128 20369 8156 21286
rect 8114 20360 8170 20369
rect 8114 20295 8170 20304
rect 8024 18420 8076 18426
rect 8024 18362 8076 18368
rect 7932 17060 7984 17066
rect 7932 17002 7984 17008
rect 7840 16652 7892 16658
rect 7840 16594 7892 16600
rect 7852 15910 7880 16594
rect 7840 15904 7892 15910
rect 7840 15846 7892 15852
rect 7746 13696 7802 13705
rect 7746 13631 7802 13640
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 7564 13456 7616 13462
rect 7564 13398 7616 13404
rect 7576 12646 7604 13398
rect 7564 12640 7616 12646
rect 7564 12582 7616 12588
rect 7576 11082 7604 12582
rect 7852 12458 7880 15846
rect 7944 15026 7972 17002
rect 7932 15020 7984 15026
rect 7932 14962 7984 14968
rect 8036 13814 8064 18362
rect 8220 13814 8248 21830
rect 8588 21622 8616 22034
rect 8668 21888 8720 21894
rect 8668 21830 8720 21836
rect 8576 21616 8628 21622
rect 8576 21558 8628 21564
rect 8484 21344 8536 21350
rect 8484 21286 8536 21292
rect 8300 21072 8352 21078
rect 8300 21014 8352 21020
rect 8312 20602 8340 21014
rect 8392 20936 8444 20942
rect 8496 20924 8524 21286
rect 8444 20896 8524 20924
rect 8392 20878 8444 20884
rect 8300 20596 8352 20602
rect 8300 20538 8352 20544
rect 8312 19514 8340 20538
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 8404 19378 8432 20878
rect 8588 20233 8616 21558
rect 8680 21418 8708 21830
rect 8668 21412 8720 21418
rect 8668 21354 8720 21360
rect 8574 20224 8630 20233
rect 8574 20159 8630 20168
rect 8484 19984 8536 19990
rect 8484 19926 8536 19932
rect 8392 19372 8444 19378
rect 8392 19314 8444 19320
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8300 17808 8352 17814
rect 8300 17750 8352 17756
rect 8312 16998 8340 17750
rect 8404 17542 8432 19110
rect 8496 18902 8524 19926
rect 8588 19553 8616 20159
rect 8680 19990 8708 21354
rect 8668 19984 8720 19990
rect 8668 19926 8720 19932
rect 8574 19544 8630 19553
rect 8574 19479 8630 19488
rect 8484 18896 8536 18902
rect 8484 18838 8536 18844
rect 8496 18426 8524 18838
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8484 18420 8536 18426
rect 8484 18362 8536 18368
rect 8588 17746 8616 18566
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8312 15910 8340 16934
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8392 15972 8444 15978
rect 8496 15960 8524 16594
rect 8444 15932 8524 15960
rect 8392 15914 8444 15920
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 8312 14822 8340 15846
rect 8496 15434 8524 15932
rect 8484 15428 8536 15434
rect 8484 15370 8536 15376
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 8496 14618 8524 14962
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8588 14498 8616 17682
rect 8772 16674 8800 22607
rect 9220 22568 9272 22574
rect 9220 22510 9272 22516
rect 9036 21888 9088 21894
rect 9036 21830 9088 21836
rect 9128 21888 9180 21894
rect 9128 21830 9180 21836
rect 9048 21690 9076 21830
rect 9036 21684 9088 21690
rect 9036 21626 9088 21632
rect 9036 20596 9088 20602
rect 9036 20538 9088 20544
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 8956 20058 8984 20402
rect 9048 20330 9076 20538
rect 9036 20324 9088 20330
rect 9036 20266 9088 20272
rect 8944 20052 8996 20058
rect 8944 19994 8996 20000
rect 8852 19508 8904 19514
rect 9048 19496 9076 20266
rect 8852 19450 8904 19456
rect 8956 19468 9076 19496
rect 8864 19242 8892 19450
rect 8852 19236 8904 19242
rect 8852 19178 8904 19184
rect 8864 18426 8892 19178
rect 8852 18420 8904 18426
rect 8852 18362 8904 18368
rect 8864 18086 8892 18362
rect 8956 18222 8984 19468
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 9048 18612 9076 19314
rect 9140 18970 9168 21830
rect 9232 21729 9260 22510
rect 9312 22500 9364 22506
rect 9312 22442 9364 22448
rect 9218 21720 9274 21729
rect 9218 21655 9274 21664
rect 9128 18964 9180 18970
rect 9128 18906 9180 18912
rect 9220 18692 9272 18698
rect 9220 18634 9272 18640
rect 9128 18624 9180 18630
rect 9048 18584 9128 18612
rect 9128 18566 9180 18572
rect 8944 18216 8996 18222
rect 8944 18158 8996 18164
rect 8852 18080 8904 18086
rect 8852 18022 8904 18028
rect 8864 17882 8892 18022
rect 8852 17876 8904 17882
rect 8852 17818 8904 17824
rect 8852 17536 8904 17542
rect 8852 17478 8904 17484
rect 8864 17066 8892 17478
rect 8956 17338 8984 18158
rect 8944 17332 8996 17338
rect 8944 17274 8996 17280
rect 8956 17066 8984 17274
rect 9140 17105 9168 18566
rect 9232 18154 9260 18634
rect 9220 18148 9272 18154
rect 9220 18090 9272 18096
rect 9232 17882 9260 18090
rect 9220 17876 9272 17882
rect 9220 17818 9272 17824
rect 9126 17096 9182 17105
rect 8852 17060 8904 17066
rect 8852 17002 8904 17008
rect 8944 17060 8996 17066
rect 9126 17031 9182 17040
rect 8944 17002 8996 17008
rect 8772 16646 8984 16674
rect 8760 16584 8812 16590
rect 8760 16526 8812 16532
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8680 15706 8708 15982
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 8772 15570 8800 16526
rect 8760 15564 8812 15570
rect 8760 15506 8812 15512
rect 8496 14470 8616 14498
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 7668 12430 7880 12458
rect 7944 13786 8064 13814
rect 8128 13786 8248 13814
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 7668 12209 7696 12430
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7654 12200 7710 12209
rect 7654 12135 7710 12144
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7576 7342 7604 9522
rect 7668 8566 7696 12135
rect 7760 11762 7788 12310
rect 7840 11824 7892 11830
rect 7840 11766 7892 11772
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7852 11626 7880 11766
rect 7840 11620 7892 11626
rect 7840 11562 7892 11568
rect 7852 11354 7880 11562
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 7840 11008 7892 11014
rect 7840 10950 7892 10956
rect 7852 10674 7880 10950
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 7760 7750 7788 9318
rect 7852 8838 7880 9998
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7852 7954 7880 8774
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7576 6934 7604 7278
rect 7564 6928 7616 6934
rect 7564 6870 7616 6876
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7116 6322 7144 6734
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 7116 5914 7144 6258
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6656 4126 6868 4154
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6564 3194 6592 3470
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6564 2990 6592 3130
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6472 2650 6500 2790
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 6564 2582 6592 2926
rect 6552 2576 6604 2582
rect 6552 2518 6604 2524
rect 6366 1184 6422 1193
rect 6366 1119 6422 1128
rect 5630 82 5686 480
rect 5552 54 5686 82
rect 4618 0 4674 54
rect 5630 0 5686 54
rect 6642 82 6698 480
rect 6840 82 6868 4126
rect 6932 4010 6960 4558
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 6920 4004 6972 4010
rect 6920 3946 6972 3952
rect 6932 2854 6960 3946
rect 7024 3670 7052 4014
rect 7208 3942 7236 4762
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7208 3738 7236 3878
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 7012 3664 7064 3670
rect 7012 3606 7064 3612
rect 7208 2922 7236 3674
rect 7484 3602 7512 4626
rect 7760 4154 7788 7686
rect 7852 7274 7880 7890
rect 7840 7268 7892 7274
rect 7840 7210 7892 7216
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7852 5846 7880 6054
rect 7840 5840 7892 5846
rect 7840 5782 7892 5788
rect 7852 5370 7880 5782
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7944 5302 7972 13786
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 8036 12850 8064 13262
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 8024 12708 8076 12714
rect 8024 12650 8076 12656
rect 8036 12442 8064 12650
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 8036 11558 8064 12378
rect 8128 11762 8156 13786
rect 8312 13530 8340 13806
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8208 12912 8260 12918
rect 8208 12854 8260 12860
rect 8116 11756 8168 11762
rect 8116 11698 8168 11704
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 8036 11286 8064 11494
rect 8220 11354 8248 12854
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8024 11280 8076 11286
rect 8024 11222 8076 11228
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 8312 10470 8340 11154
rect 8404 11132 8432 14214
rect 8496 12918 8524 14470
rect 8576 14408 8628 14414
rect 8576 14350 8628 14356
rect 8588 13530 8616 14350
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8864 13938 8892 14214
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8588 12918 8616 13466
rect 8484 12912 8536 12918
rect 8484 12854 8536 12860
rect 8576 12912 8628 12918
rect 8576 12854 8628 12860
rect 8588 11694 8616 12854
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8484 11144 8536 11150
rect 8404 11104 8484 11132
rect 8484 11086 8536 11092
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 8036 9382 8064 10066
rect 8208 9988 8260 9994
rect 8208 9930 8260 9936
rect 8220 9518 8248 9930
rect 8312 9586 8340 10406
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 8036 8294 8064 9318
rect 8116 9036 8168 9042
rect 8220 9024 8248 9454
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 8312 9042 8340 9386
rect 8168 8996 8248 9024
rect 8116 8978 8168 8984
rect 8116 8900 8168 8906
rect 8116 8842 8168 8848
rect 8128 8430 8156 8842
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 8036 7954 8064 8230
rect 8220 8090 8248 8996
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8312 8634 8340 8978
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 8312 7954 8340 8570
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8036 7342 8064 7890
rect 8208 7812 8260 7818
rect 8208 7754 8260 7760
rect 8220 7410 8248 7754
rect 8404 7478 8432 9998
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8496 9518 8524 9862
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8496 8838 8524 9454
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8680 8430 8708 11834
rect 8772 10538 8800 12242
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8864 11014 8892 11494
rect 8852 11008 8904 11014
rect 8852 10950 8904 10956
rect 8760 10532 8812 10538
rect 8760 10474 8812 10480
rect 8864 10470 8892 10950
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 8036 6662 8064 7142
rect 8220 6934 8248 7346
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 8128 6254 8156 6802
rect 8312 6662 8340 7278
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8956 6322 8984 16646
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 9232 14006 9260 14282
rect 9220 14000 9272 14006
rect 9220 13942 9272 13948
rect 9034 13424 9090 13433
rect 9034 13359 9090 13368
rect 9048 10577 9076 13359
rect 9324 12442 9352 22442
rect 9496 22432 9548 22438
rect 9496 22374 9548 22380
rect 9404 20324 9456 20330
rect 9404 20266 9456 20272
rect 9416 19854 9444 20266
rect 9404 19848 9456 19854
rect 9404 19790 9456 19796
rect 9416 19378 9444 19790
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 9416 15162 9444 15642
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9508 14618 9536 22374
rect 9600 19922 9628 23258
rect 9680 23180 9732 23186
rect 9680 23122 9732 23128
rect 9692 22710 9720 23122
rect 11072 22778 11100 27520
rect 11428 24608 11480 24614
rect 11428 24550 11480 24556
rect 11336 23180 11388 23186
rect 11336 23122 11388 23128
rect 11060 22772 11112 22778
rect 11060 22714 11112 22720
rect 9680 22704 9732 22710
rect 9680 22646 9732 22652
rect 11060 22636 11112 22642
rect 11060 22578 11112 22584
rect 10784 22568 10836 22574
rect 10784 22510 10836 22516
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10796 22098 10824 22510
rect 10784 22092 10836 22098
rect 10784 22034 10836 22040
rect 10796 22001 10824 22034
rect 10782 21992 10838 22001
rect 9680 21956 9732 21962
rect 10782 21927 10838 21936
rect 10876 21956 10928 21962
rect 9680 21898 9732 21904
rect 10876 21898 10928 21904
rect 9692 21622 9720 21898
rect 10888 21622 10916 21898
rect 9680 21616 9732 21622
rect 9680 21558 9732 21564
rect 10876 21616 10928 21622
rect 10876 21558 10928 21564
rect 9692 20913 9720 21558
rect 11072 21486 11100 22578
rect 11348 22438 11376 23122
rect 11336 22432 11388 22438
rect 11336 22374 11388 22380
rect 11060 21480 11112 21486
rect 11060 21422 11112 21428
rect 10048 21344 10100 21350
rect 10048 21286 10100 21292
rect 11060 21344 11112 21350
rect 11060 21286 11112 21292
rect 9864 21072 9916 21078
rect 9864 21014 9916 21020
rect 9772 20936 9824 20942
rect 9678 20904 9734 20913
rect 9772 20878 9824 20884
rect 9678 20839 9734 20848
rect 9784 20058 9812 20878
rect 9876 20602 9904 21014
rect 10060 20942 10088 21286
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10048 20936 10100 20942
rect 10048 20878 10100 20884
rect 9864 20596 9916 20602
rect 9864 20538 9916 20544
rect 11072 20466 11100 21286
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 11152 20324 11204 20330
rect 11152 20266 11204 20272
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 9772 20052 9824 20058
rect 9772 19994 9824 20000
rect 9588 19916 9640 19922
rect 9588 19858 9640 19864
rect 9600 19174 9628 19858
rect 9968 19718 9996 20198
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 11164 19922 11192 20266
rect 11152 19916 11204 19922
rect 11152 19858 11204 19864
rect 9956 19712 10008 19718
rect 9956 19654 10008 19660
rect 10508 19712 10560 19718
rect 10508 19654 10560 19660
rect 10048 19440 10100 19446
rect 10048 19382 10100 19388
rect 9588 19168 9640 19174
rect 9588 19110 9640 19116
rect 9864 18896 9916 18902
rect 9864 18838 9916 18844
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9784 18358 9812 18702
rect 9772 18352 9824 18358
rect 9772 18294 9824 18300
rect 9784 17882 9812 18294
rect 9876 18290 9904 18838
rect 10060 18766 10088 19382
rect 10520 19310 10548 19654
rect 11164 19514 11192 19858
rect 11152 19508 11204 19514
rect 11152 19450 11204 19456
rect 10508 19304 10560 19310
rect 10508 19246 10560 19252
rect 11152 19236 11204 19242
rect 11152 19178 11204 19184
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 10048 18760 10100 18766
rect 10152 18737 10180 19110
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10048 18702 10100 18708
rect 10138 18728 10194 18737
rect 10138 18663 10194 18672
rect 11164 18630 11192 19178
rect 11152 18624 11204 18630
rect 11152 18566 11204 18572
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 11164 18222 11192 18566
rect 11152 18216 11204 18222
rect 11152 18158 11204 18164
rect 11336 18216 11388 18222
rect 11336 18158 11388 18164
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9784 17202 9812 17818
rect 11164 17746 11192 18158
rect 11348 17814 11376 18158
rect 11336 17808 11388 17814
rect 11336 17750 11388 17756
rect 10600 17740 10652 17746
rect 10600 17682 10652 17688
rect 11152 17740 11204 17746
rect 11152 17682 11204 17688
rect 10612 17338 10640 17682
rect 10968 17604 11020 17610
rect 10968 17546 11020 17552
rect 10600 17332 10652 17338
rect 10600 17274 10652 17280
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 9864 16720 9916 16726
rect 9864 16662 9916 16668
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9416 13326 9444 14010
rect 9508 13938 9536 14554
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9140 10674 9168 11630
rect 9324 11354 9352 11698
rect 9600 11558 9628 15982
rect 9772 15904 9824 15910
rect 9772 15846 9824 15852
rect 9784 14550 9812 15846
rect 9876 15706 9904 16662
rect 9968 16522 9996 16934
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10796 16794 10824 17070
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 9956 16516 10008 16522
rect 9956 16458 10008 16464
rect 10140 16516 10192 16522
rect 10140 16458 10192 16464
rect 9968 16250 9996 16458
rect 9956 16244 10008 16250
rect 9956 16186 10008 16192
rect 10048 15972 10100 15978
rect 10048 15914 10100 15920
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 10060 15638 10088 15914
rect 10048 15632 10100 15638
rect 10048 15574 10100 15580
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9772 14544 9824 14550
rect 9772 14486 9824 14492
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 9692 13530 9720 14282
rect 9784 14074 9812 14486
rect 9968 14074 9996 15506
rect 10060 15162 10088 15574
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 10152 14618 10180 16458
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 10690 16008 10746 16017
rect 10690 15943 10746 15952
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10704 14822 10732 15943
rect 10796 15026 10824 16390
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10796 14618 10824 14962
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9956 13796 10008 13802
rect 9956 13738 10008 13744
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 10692 13796 10744 13802
rect 10692 13738 10744 13744
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9968 13462 9996 13738
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9956 13456 10008 13462
rect 9956 13398 10008 13404
rect 9876 12646 9904 13398
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 9876 12374 9904 12582
rect 9864 12368 9916 12374
rect 9864 12310 9916 12316
rect 9876 12170 9904 12310
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9864 11824 9916 11830
rect 9864 11766 9916 11772
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9876 11286 9904 11766
rect 9968 11762 9996 13398
rect 10060 12714 10088 13738
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10704 13530 10732 13738
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10876 13320 10928 13326
rect 10690 13288 10746 13297
rect 10876 13262 10928 13268
rect 10690 13223 10746 13232
rect 10140 12912 10192 12918
rect 10140 12854 10192 12860
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 10152 12238 10180 12854
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10232 12368 10284 12374
rect 10232 12310 10284 12316
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 10244 11898 10272 12310
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10704 11830 10732 13223
rect 10888 12986 10916 13262
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10980 12850 11008 17546
rect 11164 17134 11192 17682
rect 11152 17128 11204 17134
rect 11152 17070 11204 17076
rect 11164 16114 11192 17070
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 11072 13977 11100 14894
rect 11058 13968 11114 13977
rect 11058 13903 11114 13912
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 10980 12442 11008 12786
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 9404 11280 9456 11286
rect 9404 11222 9456 11228
rect 9864 11280 9916 11286
rect 9864 11222 9916 11228
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9034 10568 9090 10577
rect 9034 10503 9090 10512
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9036 7268 9088 7274
rect 9036 7210 9088 7216
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 8956 5914 8984 6258
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 8024 5636 8076 5642
rect 8024 5578 8076 5584
rect 8668 5636 8720 5642
rect 8668 5578 8720 5584
rect 8036 5409 8064 5578
rect 8022 5400 8078 5409
rect 8022 5335 8078 5344
rect 7932 5296 7984 5302
rect 7932 5238 7984 5244
rect 8036 5098 8064 5335
rect 8576 5296 8628 5302
rect 8576 5238 8628 5244
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8312 4826 8340 4966
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 7760 4126 7972 4154
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7944 3194 7972 4126
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8220 3670 8248 3878
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 7944 2990 7972 3130
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 7196 2916 7248 2922
rect 7196 2858 7248 2864
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 8036 2650 8064 3470
rect 8220 3194 8248 3606
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 8404 2378 8432 3470
rect 8588 2514 8616 5238
rect 8680 5098 8708 5578
rect 9048 5370 9076 7210
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 8668 5092 8720 5098
rect 8668 5034 8720 5040
rect 8680 4758 8708 5034
rect 8668 4752 8720 4758
rect 8668 4694 8720 4700
rect 8680 3670 8708 4694
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 8864 4146 8892 4422
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 9048 2582 9076 5306
rect 9128 5296 9180 5302
rect 9128 5238 9180 5244
rect 9140 4146 9168 5238
rect 9232 4690 9260 8230
rect 9416 7410 9444 11222
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9600 8430 9628 9590
rect 9784 9178 9812 11086
rect 9876 10266 9904 11222
rect 9968 11150 9996 11698
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 10060 10962 10088 11494
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 11164 11082 11192 11630
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 9968 10934 10088 10962
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9600 8090 9628 8366
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9692 7954 9720 8910
rect 9876 8362 9904 8978
rect 9864 8356 9916 8362
rect 9864 8298 9916 8304
rect 9876 8022 9904 8298
rect 9864 8016 9916 8022
rect 9864 7958 9916 7964
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9692 7546 9720 7890
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9036 2576 9088 2582
rect 9036 2518 9088 2524
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 9034 2408 9090 2417
rect 8392 2372 8444 2378
rect 9034 2343 9090 2352
rect 8392 2314 8444 2320
rect 9048 2310 9076 2343
rect 7380 2304 7432 2310
rect 7380 2246 7432 2252
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 6642 54 6868 82
rect 7392 82 7420 2246
rect 7654 82 7710 480
rect 7392 54 7710 82
rect 8496 82 8524 2246
rect 8758 82 8814 480
rect 9324 105 9352 6598
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9496 3460 9548 3466
rect 9496 3402 9548 3408
rect 9508 2990 9536 3402
rect 9496 2984 9548 2990
rect 9496 2926 9548 2932
rect 9404 2372 9456 2378
rect 9404 2314 9456 2320
rect 8496 54 8814 82
rect 6642 0 6698 54
rect 7654 0 7710 54
rect 8758 0 8814 54
rect 9310 96 9366 105
rect 9416 82 9444 2314
rect 9508 2310 9536 2926
rect 9600 2650 9628 5646
rect 9784 4214 9812 7754
rect 9968 7750 9996 10934
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 10046 10296 10102 10305
rect 10152 10266 10180 10542
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 11164 10266 11192 11018
rect 10046 10231 10102 10240
rect 10140 10260 10192 10266
rect 10060 10198 10088 10231
rect 10140 10202 10192 10208
rect 11152 10260 11204 10266
rect 11152 10202 11204 10208
rect 10048 10192 10100 10198
rect 10048 10134 10100 10140
rect 10060 9722 10088 10134
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 9968 6866 9996 7346
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9876 5234 9904 6258
rect 9968 6118 9996 6802
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 9968 5574 9996 6054
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 9876 4214 9904 4626
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9864 4208 9916 4214
rect 9864 4150 9916 4156
rect 10060 3534 10088 9658
rect 10704 9654 10732 10066
rect 11440 9722 11468 24550
rect 11704 24200 11756 24206
rect 11704 24142 11756 24148
rect 11716 21486 11744 24142
rect 12636 23866 12664 27526
rect 14002 27520 14058 28000
rect 15474 27520 15530 28000
rect 16946 27520 17002 28000
rect 18064 27526 18368 27554
rect 13360 24268 13412 24274
rect 13360 24210 13412 24216
rect 13084 24064 13136 24070
rect 13084 24006 13136 24012
rect 12624 23860 12676 23866
rect 12624 23802 12676 23808
rect 12072 23724 12124 23730
rect 12072 23666 12124 23672
rect 11980 21888 12032 21894
rect 11980 21830 12032 21836
rect 11704 21480 11756 21486
rect 11704 21422 11756 21428
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 11704 21072 11756 21078
rect 11704 21014 11756 21020
rect 11716 20466 11744 21014
rect 11808 20806 11836 21286
rect 11796 20800 11848 20806
rect 11796 20742 11848 20748
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 11716 19446 11744 19994
rect 11704 19440 11756 19446
rect 11704 19382 11756 19388
rect 11520 19304 11572 19310
rect 11520 19246 11572 19252
rect 11532 18290 11560 19246
rect 11888 18896 11940 18902
rect 11888 18838 11940 18844
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11520 18284 11572 18290
rect 11520 18226 11572 18232
rect 11808 17882 11836 18702
rect 11900 18426 11928 18838
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11796 17876 11848 17882
rect 11796 17818 11848 17824
rect 11888 17808 11940 17814
rect 11888 17750 11940 17756
rect 11900 16998 11928 17750
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11900 16794 11928 16934
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 11532 16114 11560 16526
rect 11900 16182 11928 16730
rect 11992 16726 12020 21830
rect 12084 19961 12112 23666
rect 12992 23656 13044 23662
rect 12992 23598 13044 23604
rect 12164 23112 12216 23118
rect 12164 23054 12216 23060
rect 12716 23112 12768 23118
rect 12716 23054 12768 23060
rect 12176 20602 12204 23054
rect 12440 22432 12492 22438
rect 12440 22374 12492 22380
rect 12256 21956 12308 21962
rect 12256 21898 12308 21904
rect 12268 21078 12296 21898
rect 12348 21888 12400 21894
rect 12348 21830 12400 21836
rect 12256 21072 12308 21078
rect 12256 21014 12308 21020
rect 12164 20596 12216 20602
rect 12164 20538 12216 20544
rect 12070 19952 12126 19961
rect 12070 19887 12126 19896
rect 12072 19848 12124 19854
rect 12072 19790 12124 19796
rect 11980 16720 12032 16726
rect 11980 16662 12032 16668
rect 11888 16176 11940 16182
rect 11888 16118 11940 16124
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11532 15706 11560 16050
rect 11900 15910 11928 16118
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 11520 15700 11572 15706
rect 11520 15642 11572 15648
rect 11900 15638 11928 15846
rect 11888 15632 11940 15638
rect 11888 15574 11940 15580
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11716 15094 11744 15438
rect 11704 15088 11756 15094
rect 11704 15030 11756 15036
rect 11520 14884 11572 14890
rect 11520 14826 11572 14832
rect 11532 14074 11560 14826
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11532 12646 11560 13262
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11532 12442 11560 12582
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11532 11150 11560 11562
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11532 10266 11560 11086
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11428 9716 11480 9722
rect 11428 9658 11480 9664
rect 10692 9648 10744 9654
rect 10692 9590 10744 9596
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10704 8022 10732 8298
rect 10692 8016 10744 8022
rect 10692 7958 10744 7964
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 10612 7410 10640 7890
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10796 7342 10824 9318
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 10980 8634 11008 9046
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 10888 7818 10916 8298
rect 11256 7954 11284 9454
rect 11520 9444 11572 9450
rect 11520 9386 11572 9392
rect 11532 8974 11560 9386
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11624 7993 11652 14758
rect 11808 14550 11836 15506
rect 11900 15162 11928 15574
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11900 14822 11928 15098
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 11796 14544 11848 14550
rect 11702 14512 11758 14521
rect 11796 14486 11848 14492
rect 11702 14447 11758 14456
rect 11716 14414 11744 14447
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 11716 13530 11744 14350
rect 11808 13870 11836 14486
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11900 13734 11928 14758
rect 12084 13814 12112 19790
rect 12164 19440 12216 19446
rect 12164 19382 12216 19388
rect 12176 18068 12204 19382
rect 12268 18970 12296 21014
rect 12256 18964 12308 18970
rect 12256 18906 12308 18912
rect 12268 18698 12296 18906
rect 12256 18692 12308 18698
rect 12256 18634 12308 18640
rect 12256 18080 12308 18086
rect 12176 18040 12256 18068
rect 12256 18022 12308 18028
rect 12268 17814 12296 18022
rect 12256 17808 12308 17814
rect 12256 17750 12308 17756
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 12176 17338 12204 17614
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 12268 15570 12296 15846
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 12164 14952 12216 14958
rect 12164 14894 12216 14900
rect 11992 13786 12112 13814
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 11900 13530 11928 13670
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11900 12918 11928 13466
rect 11888 12912 11940 12918
rect 11888 12854 11940 12860
rect 11900 12646 11928 12854
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11716 11286 11744 12582
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11900 11558 11928 12174
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 11704 11280 11756 11286
rect 11704 11222 11756 11228
rect 11716 10538 11744 11222
rect 11796 11008 11848 11014
rect 11796 10950 11848 10956
rect 11704 10532 11756 10538
rect 11704 10474 11756 10480
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11716 9654 11744 10066
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 11716 9042 11744 9590
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11808 8838 11836 10950
rect 11900 9994 11928 11494
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 11900 9897 11928 9930
rect 11886 9888 11942 9897
rect 11886 9823 11942 9832
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11808 8362 11836 8774
rect 11796 8356 11848 8362
rect 11796 8298 11848 8304
rect 11610 7984 11666 7993
rect 11244 7948 11296 7954
rect 11610 7919 11666 7928
rect 11244 7890 11296 7896
rect 10876 7812 10928 7818
rect 10876 7754 10928 7760
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 11072 6866 11100 7278
rect 11256 7002 11284 7890
rect 11520 7268 11572 7274
rect 11520 7210 11572 7216
rect 11532 7002 11560 7210
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11520 6996 11572 7002
rect 11520 6938 11572 6944
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10140 6180 10192 6186
rect 10140 6122 10192 6128
rect 10152 5574 10180 6122
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10152 4690 10180 5510
rect 10704 5030 10732 5782
rect 10796 5234 10824 6734
rect 11072 6662 11100 6802
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11072 6254 11100 6598
rect 11900 6458 11928 6802
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 11152 6180 11204 6186
rect 11152 6122 11204 6128
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10152 3942 10180 4626
rect 10704 4486 10732 4966
rect 10980 4554 11008 5646
rect 11058 5128 11114 5137
rect 11058 5063 11114 5072
rect 10968 4548 11020 4554
rect 10968 4490 11020 4496
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 10980 4010 11008 4082
rect 10876 4004 10928 4010
rect 10876 3946 10928 3952
rect 10968 4004 11020 4010
rect 10968 3946 11020 3952
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10152 3602 10180 3878
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10060 3194 10088 3470
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 10692 3392 10744 3398
rect 10888 3380 10916 3946
rect 10980 3738 11008 3946
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 10968 3392 11020 3398
rect 10888 3352 10968 3380
rect 10692 3334 10744 3340
rect 10968 3334 11020 3340
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 10152 2514 10180 3334
rect 10704 3058 10732 3334
rect 10980 3126 11008 3334
rect 10968 3120 11020 3126
rect 10968 3062 11020 3068
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 9496 2304 9548 2310
rect 9496 2246 9548 2252
rect 10152 2106 10180 2450
rect 10140 2100 10192 2106
rect 10140 2042 10192 2048
rect 9770 82 9826 480
rect 9416 54 9826 82
rect 9310 31 9366 40
rect 9770 0 9826 54
rect 10782 82 10838 480
rect 11072 82 11100 5063
rect 11164 4622 11192 6122
rect 11888 5704 11940 5710
rect 11888 5646 11940 5652
rect 11520 5636 11572 5642
rect 11520 5578 11572 5584
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11164 4282 11192 4558
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11532 4146 11560 5578
rect 11796 4752 11848 4758
rect 11796 4694 11848 4700
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11808 3942 11836 4694
rect 11900 4690 11928 5646
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11992 4154 12020 13786
rect 12070 12880 12126 12889
rect 12070 12815 12126 12824
rect 12084 4321 12112 12815
rect 12176 12306 12204 14894
rect 12360 13326 12388 21830
rect 12452 17270 12480 22374
rect 12532 22092 12584 22098
rect 12532 22034 12584 22040
rect 12544 21350 12572 22034
rect 12532 21344 12584 21350
rect 12532 21286 12584 21292
rect 12544 19854 12572 21286
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12624 19712 12676 19718
rect 12624 19654 12676 19660
rect 12636 19310 12664 19654
rect 12624 19304 12676 19310
rect 12624 19246 12676 19252
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12636 18222 12664 18566
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12440 17264 12492 17270
rect 12440 17206 12492 17212
rect 12452 16017 12480 17206
rect 12532 16720 12584 16726
rect 12532 16662 12584 16668
rect 12544 16114 12572 16662
rect 12532 16108 12584 16114
rect 12532 16050 12584 16056
rect 12438 16008 12494 16017
rect 12438 15943 12494 15952
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12176 11898 12204 12242
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12452 11762 12480 14758
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 12544 14006 12572 14350
rect 12532 14000 12584 14006
rect 12532 13942 12584 13948
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12544 12850 12572 13126
rect 12532 12844 12584 12850
rect 12532 12786 12584 12792
rect 12440 11756 12492 11762
rect 12440 11698 12492 11704
rect 12452 11354 12480 11698
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12636 10538 12664 11222
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 9110 12480 10406
rect 12636 10198 12664 10474
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12636 9382 12664 10134
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 12452 8634 12480 9046
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12452 8362 12480 8570
rect 12440 8356 12492 8362
rect 12440 8298 12492 8304
rect 12452 8022 12480 8298
rect 12440 8016 12492 8022
rect 12440 7958 12492 7964
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12176 7546 12204 7822
rect 12256 7812 12308 7818
rect 12256 7754 12308 7760
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 12268 6866 12296 7754
rect 12452 7546 12480 7958
rect 12440 7540 12492 7546
rect 12360 7500 12440 7528
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 12268 5914 12296 6802
rect 12360 6458 12388 7500
rect 12440 7482 12492 7488
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12360 6186 12388 6394
rect 12452 6322 12480 6938
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12348 6180 12400 6186
rect 12348 6122 12400 6128
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 12360 5846 12388 6122
rect 12348 5840 12400 5846
rect 12348 5782 12400 5788
rect 12360 5370 12388 5782
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12360 5098 12388 5306
rect 12348 5092 12400 5098
rect 12348 5034 12400 5040
rect 12360 4758 12388 5034
rect 12348 4752 12400 4758
rect 12348 4694 12400 4700
rect 12070 4312 12126 4321
rect 12070 4247 12126 4256
rect 11900 4126 12020 4154
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11808 3670 11836 3878
rect 11796 3664 11848 3670
rect 11796 3606 11848 3612
rect 11704 3460 11756 3466
rect 11704 3402 11756 3408
rect 11520 2848 11572 2854
rect 11520 2790 11572 2796
rect 11532 2582 11560 2790
rect 11520 2576 11572 2582
rect 11520 2518 11572 2524
rect 11716 2514 11744 3402
rect 11808 2922 11836 3606
rect 11900 2961 11928 4126
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11886 2952 11942 2961
rect 11796 2916 11848 2922
rect 11886 2887 11942 2896
rect 11796 2858 11848 2864
rect 11992 2650 12020 3470
rect 12176 3194 12204 3674
rect 12728 3194 12756 23054
rect 12808 23044 12860 23050
rect 12808 22986 12860 22992
rect 12820 13814 12848 22986
rect 12900 22976 12952 22982
rect 12900 22918 12952 22924
rect 12912 18766 12940 22918
rect 13004 22574 13032 23598
rect 12992 22568 13044 22574
rect 12992 22510 13044 22516
rect 12992 22228 13044 22234
rect 12992 22170 13044 22176
rect 13004 21350 13032 22170
rect 13096 22166 13124 24006
rect 13372 23866 13400 24210
rect 14016 24206 14044 27520
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14096 24268 14148 24274
rect 14096 24210 14148 24216
rect 14004 24200 14056 24206
rect 14004 24142 14056 24148
rect 14004 24064 14056 24070
rect 14004 24006 14056 24012
rect 13360 23860 13412 23866
rect 13360 23802 13412 23808
rect 13176 23656 13228 23662
rect 13176 23598 13228 23604
rect 13188 23322 13216 23598
rect 13176 23316 13228 23322
rect 13176 23258 13228 23264
rect 13176 22976 13228 22982
rect 13228 22936 13308 22964
rect 13176 22918 13228 22924
rect 13176 22432 13228 22438
rect 13176 22374 13228 22380
rect 13084 22160 13136 22166
rect 13084 22102 13136 22108
rect 13096 21690 13124 22102
rect 13084 21684 13136 21690
rect 13084 21626 13136 21632
rect 12992 21344 13044 21350
rect 12992 21286 13044 21292
rect 13084 21344 13136 21350
rect 13084 21286 13136 21292
rect 13004 20534 13032 21286
rect 13096 21146 13124 21286
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 13188 21078 13216 22374
rect 13176 21072 13228 21078
rect 13176 21014 13228 21020
rect 12992 20528 13044 20534
rect 12992 20470 13044 20476
rect 13004 20330 13032 20470
rect 12992 20324 13044 20330
rect 12992 20266 13044 20272
rect 13004 20058 13032 20266
rect 13188 20058 13216 21014
rect 12992 20052 13044 20058
rect 12992 19994 13044 20000
rect 13176 20052 13228 20058
rect 13176 19994 13228 20000
rect 13176 19848 13228 19854
rect 13176 19790 13228 19796
rect 12992 19508 13044 19514
rect 12992 19450 13044 19456
rect 13004 19242 13032 19450
rect 13188 19378 13216 19790
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 12992 19236 13044 19242
rect 12992 19178 13044 19184
rect 12900 18760 12952 18766
rect 12900 18702 12952 18708
rect 12990 18592 13046 18601
rect 12990 18527 13046 18536
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 12912 15434 12940 15846
rect 12900 15428 12952 15434
rect 12900 15370 12952 15376
rect 13004 15162 13032 18527
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 13096 17338 13124 17478
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 13084 16992 13136 16998
rect 13084 16934 13136 16940
rect 13096 16250 13124 16934
rect 13176 16516 13228 16522
rect 13176 16458 13228 16464
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 13188 15978 13216 16458
rect 13176 15972 13228 15978
rect 13176 15914 13228 15920
rect 13188 15434 13216 15914
rect 13280 15638 13308 22936
rect 13372 22642 13400 23802
rect 13544 23792 13596 23798
rect 13544 23734 13596 23740
rect 13452 23520 13504 23526
rect 13452 23462 13504 23468
rect 13360 22636 13412 22642
rect 13360 22578 13412 22584
rect 13372 22545 13400 22578
rect 13358 22536 13414 22545
rect 13358 22471 13414 22480
rect 13360 22432 13412 22438
rect 13360 22374 13412 22380
rect 13372 19786 13400 22374
rect 13464 20942 13492 23462
rect 13452 20936 13504 20942
rect 13452 20878 13504 20884
rect 13360 19780 13412 19786
rect 13360 19722 13412 19728
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13372 17882 13400 18702
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 13556 17320 13584 23734
rect 13912 23656 13964 23662
rect 13912 23598 13964 23604
rect 13924 23186 13952 23598
rect 13912 23180 13964 23186
rect 13912 23122 13964 23128
rect 13728 22772 13780 22778
rect 13728 22714 13780 22720
rect 13636 21616 13688 21622
rect 13740 21604 13768 22714
rect 13924 22574 13952 23122
rect 13912 22568 13964 22574
rect 13912 22510 13964 22516
rect 13912 22432 13964 22438
rect 13912 22374 13964 22380
rect 13688 21576 13768 21604
rect 13636 21558 13688 21564
rect 13728 20868 13780 20874
rect 13728 20810 13780 20816
rect 13740 20262 13768 20810
rect 13728 20256 13780 20262
rect 13728 20198 13780 20204
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 13648 19514 13676 19994
rect 13636 19508 13688 19514
rect 13636 19450 13688 19456
rect 13636 18896 13688 18902
rect 13636 18838 13688 18844
rect 13648 18426 13676 18838
rect 13740 18766 13768 20198
rect 13728 18760 13780 18766
rect 13728 18702 13780 18708
rect 13636 18420 13688 18426
rect 13636 18362 13688 18368
rect 13648 18086 13676 18362
rect 13740 18290 13768 18702
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13636 18080 13688 18086
rect 13636 18022 13688 18028
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13636 17876 13688 17882
rect 13636 17818 13688 17824
rect 13372 17292 13584 17320
rect 13372 16726 13400 17292
rect 13648 17202 13676 17818
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 13636 17196 13688 17202
rect 13556 17156 13636 17184
rect 13360 16720 13412 16726
rect 13360 16662 13412 16668
rect 13556 16454 13584 17156
rect 13636 17138 13688 17144
rect 13740 17066 13768 17274
rect 13728 17060 13780 17066
rect 13728 17002 13780 17008
rect 13832 16946 13860 18022
rect 13648 16918 13860 16946
rect 13648 16726 13676 16918
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13636 16720 13688 16726
rect 13740 16697 13768 16730
rect 13636 16662 13688 16668
rect 13726 16688 13782 16697
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13648 16250 13676 16662
rect 13726 16623 13782 16632
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 13636 16244 13688 16250
rect 13636 16186 13688 16192
rect 13452 15700 13504 15706
rect 13452 15642 13504 15648
rect 13268 15632 13320 15638
rect 13268 15574 13320 15580
rect 13176 15428 13228 15434
rect 13176 15370 13228 15376
rect 13464 15162 13492 15642
rect 12992 15156 13044 15162
rect 12992 15098 13044 15104
rect 13452 15156 13504 15162
rect 13452 15098 13504 15104
rect 13004 14958 13032 15098
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 13464 14822 13492 15098
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13464 14618 13492 14758
rect 13452 14612 13504 14618
rect 13452 14554 13504 14560
rect 13266 14512 13322 14521
rect 13266 14447 13322 14456
rect 13280 14414 13308 14447
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 12820 13786 13124 13814
rect 12808 12708 12860 12714
rect 12808 12650 12860 12656
rect 12820 12102 12848 12650
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12820 11626 12848 12038
rect 12808 11620 12860 11626
rect 12808 11562 12860 11568
rect 12820 11014 12848 11562
rect 13096 11014 13124 13786
rect 13176 13728 13228 13734
rect 13176 13670 13228 13676
rect 13188 13530 13216 13670
rect 13280 13530 13308 14350
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13452 12708 13504 12714
rect 13452 12650 13504 12656
rect 13464 12170 13492 12650
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13360 11620 13412 11626
rect 13360 11562 13412 11568
rect 13372 11286 13400 11562
rect 13360 11280 13412 11286
rect 13360 11222 13412 11228
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 13084 11008 13136 11014
rect 13084 10950 13136 10956
rect 13372 10742 13400 11222
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12820 10577 12848 10610
rect 12806 10568 12862 10577
rect 12806 10503 12862 10512
rect 12820 10266 12848 10503
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 12912 8906 12940 10610
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 13004 9586 13032 9862
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 12900 8900 12952 8906
rect 12900 8842 12952 8848
rect 12912 7478 12940 8842
rect 13004 8566 13032 9522
rect 13280 9178 13308 9998
rect 13372 9654 13400 10678
rect 13464 10538 13492 12106
rect 13452 10532 13504 10538
rect 13452 10474 13504 10480
rect 13360 9648 13412 9654
rect 13360 9590 13412 9596
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 13464 9110 13492 10474
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13556 9058 13584 16186
rect 13924 15706 13952 22374
rect 14016 22234 14044 24006
rect 14108 23526 14136 24210
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 14096 23520 14148 23526
rect 14096 23462 14148 23468
rect 15488 23186 15516 27520
rect 16960 23866 16988 27520
rect 16948 23860 17000 23866
rect 16948 23802 17000 23808
rect 15660 23656 15712 23662
rect 15660 23598 15712 23604
rect 16396 23656 16448 23662
rect 16396 23598 16448 23604
rect 15476 23180 15528 23186
rect 15476 23122 15528 23128
rect 14740 22976 14792 22982
rect 14740 22918 14792 22924
rect 14464 22636 14516 22642
rect 14464 22578 14516 22584
rect 14004 22228 14056 22234
rect 14004 22170 14056 22176
rect 14016 21622 14044 22170
rect 14004 21616 14056 21622
rect 14004 21558 14056 21564
rect 14096 21616 14148 21622
rect 14096 21558 14148 21564
rect 14108 21162 14136 21558
rect 14372 21412 14424 21418
rect 14372 21354 14424 21360
rect 14016 21134 14136 21162
rect 13912 15700 13964 15706
rect 13832 15660 13912 15688
rect 13832 15026 13860 15660
rect 13912 15642 13964 15648
rect 13912 15428 13964 15434
rect 13912 15370 13964 15376
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13924 14550 13952 15370
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13912 14544 13964 14550
rect 13912 14486 13964 14492
rect 13648 13734 13676 14486
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13832 13462 13860 14010
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13740 12442 13768 13262
rect 13832 12986 13860 13398
rect 13924 13326 13952 14486
rect 13912 13320 13964 13326
rect 13912 13262 13964 13268
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13912 12708 13964 12714
rect 13912 12650 13964 12656
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13636 12368 13688 12374
rect 13636 12310 13688 12316
rect 13648 11558 13676 12310
rect 13924 12209 13952 12650
rect 13910 12200 13966 12209
rect 13910 12135 13966 12144
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13648 11082 13676 11494
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 13648 10810 13676 11018
rect 13636 10804 13688 10810
rect 13636 10746 13688 10752
rect 13648 10198 13676 10746
rect 13636 10192 13688 10198
rect 13636 10134 13688 10140
rect 13648 9722 13676 10134
rect 13636 9716 13688 9722
rect 13636 9658 13688 9664
rect 13556 9030 13676 9058
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 12992 8560 13044 8566
rect 12992 8502 13044 8508
rect 13004 8022 13032 8502
rect 13556 8090 13584 8910
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 12992 8016 13044 8022
rect 12992 7958 13044 7964
rect 13452 8016 13504 8022
rect 13452 7958 13504 7964
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 13280 7546 13308 7686
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 13280 7206 13308 7482
rect 13464 7410 13492 7958
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 13360 6928 13412 6934
rect 13360 6870 13412 6876
rect 13372 6458 13400 6870
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 13004 4826 13032 5170
rect 12992 4820 13044 4826
rect 12992 4762 13044 4768
rect 13372 4486 13400 6394
rect 13464 4758 13492 6734
rect 13556 6390 13584 7686
rect 13544 6384 13596 6390
rect 13544 6326 13596 6332
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13556 4758 13584 6054
rect 13648 5137 13676 9030
rect 13740 7206 13768 11766
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13740 6254 13768 7142
rect 13924 6934 13952 12135
rect 14016 11830 14044 21134
rect 14096 21072 14148 21078
rect 14096 21014 14148 21020
rect 14108 20058 14136 21014
rect 14384 20602 14412 21354
rect 14372 20596 14424 20602
rect 14200 20556 14372 20584
rect 14096 20052 14148 20058
rect 14096 19994 14148 20000
rect 14096 19168 14148 19174
rect 14096 19110 14148 19116
rect 14108 18970 14136 19110
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 14200 17882 14228 20556
rect 14372 20538 14424 20544
rect 14280 19236 14332 19242
rect 14280 19178 14332 19184
rect 14372 19236 14424 19242
rect 14372 19178 14424 19184
rect 14292 18902 14320 19178
rect 14384 18970 14412 19178
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14280 18896 14332 18902
rect 14280 18838 14332 18844
rect 14476 18698 14504 22578
rect 14556 22500 14608 22506
rect 14556 22442 14608 22448
rect 14568 21729 14596 22442
rect 14554 21720 14610 21729
rect 14554 21655 14610 21664
rect 14648 21548 14700 21554
rect 14648 21490 14700 21496
rect 14660 19689 14688 21490
rect 14752 20466 14780 22918
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15488 22778 15516 23122
rect 15476 22772 15528 22778
rect 15476 22714 15528 22720
rect 14832 22432 14884 22438
rect 14832 22374 14884 22380
rect 14844 22234 14872 22374
rect 14832 22228 14884 22234
rect 14832 22170 14884 22176
rect 15292 22160 15344 22166
rect 15292 22102 15344 22108
rect 14832 22024 14884 22030
rect 14832 21966 14884 21972
rect 14844 21486 14872 21966
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14832 21480 14884 21486
rect 14832 21422 14884 21428
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14832 20528 14884 20534
rect 14832 20470 14884 20476
rect 14740 20460 14792 20466
rect 14740 20402 14792 20408
rect 14752 20058 14780 20402
rect 14844 20330 14872 20470
rect 14832 20324 14884 20330
rect 14832 20266 14884 20272
rect 14740 20052 14792 20058
rect 14740 19994 14792 20000
rect 14740 19916 14792 19922
rect 14740 19858 14792 19864
rect 14646 19680 14702 19689
rect 14646 19615 14702 19624
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 14464 18692 14516 18698
rect 14464 18634 14516 18640
rect 14660 18290 14688 19314
rect 14752 19174 14780 19858
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14740 19168 14792 19174
rect 14740 19110 14792 19116
rect 14752 18601 14780 19110
rect 14738 18592 14794 18601
rect 14738 18527 14794 18536
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14648 18284 14700 18290
rect 14648 18226 14700 18232
rect 14280 18148 14332 18154
rect 14280 18090 14332 18096
rect 14292 17882 14320 18090
rect 14188 17876 14240 17882
rect 14188 17818 14240 17824
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14188 16040 14240 16046
rect 14188 15982 14240 15988
rect 14096 15904 14148 15910
rect 14096 15846 14148 15852
rect 14108 15094 14136 15846
rect 14096 15088 14148 15094
rect 14096 15030 14148 15036
rect 14200 15026 14228 15982
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 14292 14770 14320 17478
rect 14384 17270 14412 18226
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 14372 17264 14424 17270
rect 14372 17206 14424 17212
rect 14752 16998 14780 17682
rect 15304 17610 15332 22102
rect 15384 22092 15436 22098
rect 15384 22034 15436 22040
rect 15396 21554 15424 22034
rect 15476 21888 15528 21894
rect 15476 21830 15528 21836
rect 15384 21548 15436 21554
rect 15384 21490 15436 21496
rect 15384 21004 15436 21010
rect 15384 20946 15436 20952
rect 15396 20534 15424 20946
rect 15384 20528 15436 20534
rect 15384 20470 15436 20476
rect 15384 18896 15436 18902
rect 15384 18838 15436 18844
rect 15396 18086 15424 18838
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 15292 17604 15344 17610
rect 15292 17546 15344 17552
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14740 16992 14792 16998
rect 14740 16934 14792 16940
rect 14648 16448 14700 16454
rect 14648 16390 14700 16396
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14372 14884 14424 14890
rect 14372 14826 14424 14832
rect 14200 14742 14320 14770
rect 14200 13376 14228 14742
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14292 13938 14320 14554
rect 14384 13938 14412 14826
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14372 13932 14424 13938
rect 14372 13874 14424 13880
rect 14476 13841 14504 14214
rect 14462 13832 14518 13841
rect 14462 13767 14518 13776
rect 14568 13716 14596 15506
rect 14476 13688 14596 13716
rect 14200 13348 14320 13376
rect 14188 13252 14240 13258
rect 14188 13194 14240 13200
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 14108 11898 14136 12174
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14004 11824 14056 11830
rect 14004 11766 14056 11772
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 14016 10266 14044 11086
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 14016 9178 14044 9318
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 14108 7546 14136 7890
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 14096 7268 14148 7274
rect 14096 7210 14148 7216
rect 13912 6928 13964 6934
rect 13912 6870 13964 6876
rect 14004 6724 14056 6730
rect 14004 6666 14056 6672
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 14016 6186 14044 6666
rect 14108 6361 14136 7210
rect 14094 6352 14150 6361
rect 14094 6287 14150 6296
rect 14004 6180 14056 6186
rect 14004 6122 14056 6128
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 13728 5840 13780 5846
rect 13728 5782 13780 5788
rect 13740 5370 13768 5782
rect 14108 5409 14136 6054
rect 14094 5400 14150 5409
rect 13728 5364 13780 5370
rect 14094 5335 14150 5344
rect 13728 5306 13780 5312
rect 13634 5128 13690 5137
rect 13634 5063 13690 5072
rect 13452 4752 13504 4758
rect 13452 4694 13504 4700
rect 13544 4752 13596 4758
rect 13544 4694 13596 4700
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 13360 4480 13412 4486
rect 13360 4422 13412 4428
rect 12912 4010 12940 4422
rect 12900 4004 12952 4010
rect 12900 3946 12952 3952
rect 12912 3738 12940 3946
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 13084 3664 13136 3670
rect 13084 3606 13136 3612
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 12990 2952 13046 2961
rect 13096 2922 13124 3606
rect 13464 3466 13492 4694
rect 13556 4282 13584 4694
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 13636 4208 13688 4214
rect 13636 4150 13688 4156
rect 13452 3460 13504 3466
rect 13452 3402 13504 3408
rect 13648 3058 13676 4150
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 14016 3194 14044 3470
rect 14004 3188 14056 3194
rect 14004 3130 14056 3136
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 12990 2887 13046 2896
rect 13084 2916 13136 2922
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12070 2000 12126 2009
rect 12070 1935 12126 1944
rect 10782 54 11100 82
rect 11794 82 11850 480
rect 12084 82 12112 1935
rect 12452 1873 12480 2246
rect 12438 1864 12494 1873
rect 12438 1799 12494 1808
rect 11794 54 12112 82
rect 12898 82 12954 480
rect 13004 82 13032 2887
rect 13084 2858 13136 2864
rect 13096 2650 13124 2858
rect 13084 2644 13136 2650
rect 13084 2586 13136 2592
rect 13648 2378 13676 2994
rect 13636 2372 13688 2378
rect 13636 2314 13688 2320
rect 14200 2145 14228 13194
rect 14292 10062 14320 13348
rect 14476 12714 14504 13688
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14464 12708 14516 12714
rect 14464 12650 14516 12656
rect 14568 12374 14596 12718
rect 14556 12368 14608 12374
rect 14556 12310 14608 12316
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 14384 10674 14412 12242
rect 14464 10804 14516 10810
rect 14464 10746 14516 10752
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14384 10198 14412 10610
rect 14476 10538 14504 10746
rect 14464 10532 14516 10538
rect 14464 10474 14516 10480
rect 14372 10192 14424 10198
rect 14372 10134 14424 10140
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14462 9888 14518 9897
rect 14462 9823 14518 9832
rect 14280 9104 14332 9110
rect 14280 9046 14332 9052
rect 14292 8498 14320 9046
rect 14476 8566 14504 9823
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14568 9178 14596 9522
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14464 8560 14516 8566
rect 14464 8502 14516 8508
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14568 7274 14596 8434
rect 14556 7268 14608 7274
rect 14556 7210 14608 7216
rect 14280 5772 14332 5778
rect 14280 5714 14332 5720
rect 14292 4758 14320 5714
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14568 5234 14596 5510
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14280 4752 14332 4758
rect 14280 4694 14332 4700
rect 14464 4480 14516 4486
rect 14464 4422 14516 4428
rect 14372 3936 14424 3942
rect 14476 3924 14504 4422
rect 14568 4282 14596 5170
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 14660 4146 14688 16390
rect 14752 13433 14780 16934
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14832 14340 14884 14346
rect 14832 14282 14884 14288
rect 14844 13530 14872 14282
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15304 14006 15332 16730
rect 15396 16726 15424 18022
rect 15384 16720 15436 16726
rect 15384 16662 15436 16668
rect 15396 16182 15424 16662
rect 15384 16176 15436 16182
rect 15384 16118 15436 16124
rect 15384 14544 15436 14550
rect 15384 14486 15436 14492
rect 15396 14074 15424 14486
rect 15384 14068 15436 14074
rect 15384 14010 15436 14016
rect 15292 14000 15344 14006
rect 15198 13968 15254 13977
rect 15292 13942 15344 13948
rect 15198 13903 15254 13912
rect 14922 13832 14978 13841
rect 14922 13767 14978 13776
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 14738 13424 14794 13433
rect 14738 13359 14794 13368
rect 14936 13172 14964 13767
rect 15212 13258 15240 13903
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15200 13252 15252 13258
rect 15200 13194 15252 13200
rect 14752 13144 14964 13172
rect 14752 11694 14780 13144
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15108 12844 15160 12850
rect 15304 12832 15332 13330
rect 15160 12804 15332 12832
rect 15108 12786 15160 12792
rect 15120 12753 15148 12786
rect 15106 12744 15162 12753
rect 14832 12708 14884 12714
rect 15106 12679 15162 12688
rect 14832 12650 14884 12656
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14752 10470 14780 11630
rect 14844 10674 14872 12650
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15304 11762 15332 12038
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15108 11688 15160 11694
rect 15108 11630 15160 11636
rect 15120 11354 15148 11630
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14924 10736 14976 10742
rect 14924 10678 14976 10684
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14936 10266 14964 10678
rect 15304 10606 15332 11154
rect 15384 11076 15436 11082
rect 15384 11018 15436 11024
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14752 8498 14780 9522
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 15028 7002 15056 7346
rect 15304 7342 15332 9454
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15016 6996 15068 7002
rect 15016 6938 15068 6944
rect 15290 6760 15346 6769
rect 15290 6695 15346 6704
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15200 6384 15252 6390
rect 15200 6326 15252 6332
rect 15212 6118 15240 6326
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15212 5846 15240 6054
rect 15200 5840 15252 5846
rect 15200 5782 15252 5788
rect 15304 5778 15332 6695
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15304 5234 15332 5714
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 15290 4992 15346 5001
rect 15290 4927 15346 4936
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14738 4312 14794 4321
rect 14956 4304 15252 4324
rect 14738 4247 14794 4256
rect 14648 4140 14700 4146
rect 14648 4082 14700 4088
rect 14424 3896 14504 3924
rect 14372 3878 14424 3884
rect 14476 3641 14504 3896
rect 14660 3738 14688 4082
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14462 3632 14518 3641
rect 14462 3567 14518 3576
rect 14752 3058 14780 4247
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15304 3194 15332 4927
rect 15396 4154 15424 11018
rect 15488 9586 15516 21830
rect 15568 21344 15620 21350
rect 15568 21286 15620 21292
rect 15580 14346 15608 21286
rect 15672 21146 15700 23598
rect 16028 22976 16080 22982
rect 16028 22918 16080 22924
rect 15844 22636 15896 22642
rect 15844 22578 15896 22584
rect 15660 21140 15712 21146
rect 15660 21082 15712 21088
rect 15660 21004 15712 21010
rect 15660 20946 15712 20952
rect 15672 20602 15700 20946
rect 15752 20936 15804 20942
rect 15752 20878 15804 20884
rect 15660 20596 15712 20602
rect 15660 20538 15712 20544
rect 15660 17740 15712 17746
rect 15660 17682 15712 17688
rect 15672 17066 15700 17682
rect 15660 17060 15712 17066
rect 15660 17002 15712 17008
rect 15764 16114 15792 20878
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15752 15564 15804 15570
rect 15752 15506 15804 15512
rect 15764 15162 15792 15506
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15568 14340 15620 14346
rect 15568 14282 15620 14288
rect 15672 13938 15700 14350
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15856 13814 15884 22578
rect 15936 19984 15988 19990
rect 15936 19926 15988 19932
rect 15948 19514 15976 19926
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 15948 18426 15976 19450
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 16040 16266 16068 22918
rect 16120 22568 16172 22574
rect 16120 22510 16172 22516
rect 16132 22438 16160 22510
rect 16120 22432 16172 22438
rect 16120 22374 16172 22380
rect 16132 21486 16160 22374
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 16120 21480 16172 21486
rect 16120 21422 16172 21428
rect 16132 20369 16160 21422
rect 16118 20360 16174 20369
rect 16118 20295 16174 20304
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 16132 17542 16160 18702
rect 16212 18624 16264 18630
rect 16212 18566 16264 18572
rect 16224 18222 16252 18566
rect 16212 18216 16264 18222
rect 16212 18158 16264 18164
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 15764 13786 15884 13814
rect 15948 16238 16068 16266
rect 15660 12912 15712 12918
rect 15660 12854 15712 12860
rect 15672 12646 15700 12854
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15672 12374 15700 12582
rect 15660 12368 15712 12374
rect 15660 12310 15712 12316
rect 15672 11762 15700 12310
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15672 10810 15700 11698
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15672 10538 15700 10746
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15580 9450 15608 10066
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15568 9444 15620 9450
rect 15568 9386 15620 9392
rect 15672 9042 15700 9658
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15672 8294 15700 8978
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15568 8084 15620 8090
rect 15568 8026 15620 8032
rect 15476 5840 15528 5846
rect 15476 5782 15528 5788
rect 15488 5234 15516 5782
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15396 4126 15516 4154
rect 15488 3670 15516 4126
rect 15476 3664 15528 3670
rect 15476 3606 15528 3612
rect 15476 3528 15528 3534
rect 15580 3516 15608 8026
rect 15660 7268 15712 7274
rect 15660 7210 15712 7216
rect 15672 6322 15700 7210
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15764 4826 15792 13786
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15856 12782 15884 13126
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 15844 9036 15896 9042
rect 15844 8978 15896 8984
rect 15856 8673 15884 8978
rect 15948 8956 15976 16238
rect 16028 15904 16080 15910
rect 16028 15846 16080 15852
rect 16040 10130 16068 15846
rect 16132 15706 16160 16526
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 16120 15428 16172 15434
rect 16120 15370 16172 15376
rect 16132 11354 16160 15370
rect 16224 15026 16252 18158
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 16212 13932 16264 13938
rect 16212 13874 16264 13880
rect 16224 13530 16252 13874
rect 16212 13524 16264 13530
rect 16212 13466 16264 13472
rect 16316 13462 16344 21830
rect 16408 21078 16436 23598
rect 16488 23588 16540 23594
rect 16488 23530 16540 23536
rect 16500 23322 16528 23530
rect 18064 23322 18092 27526
rect 18340 27418 18368 27526
rect 18418 27520 18474 28000
rect 19536 27526 19840 27554
rect 18432 27418 18460 27520
rect 18340 27390 18460 27418
rect 18234 23624 18290 23633
rect 18234 23559 18290 23568
rect 18512 23588 18564 23594
rect 18248 23526 18276 23559
rect 18512 23530 18564 23536
rect 18236 23520 18288 23526
rect 18524 23497 18552 23530
rect 18236 23462 18288 23468
rect 18510 23488 18566 23497
rect 18510 23423 18566 23432
rect 16488 23316 16540 23322
rect 16488 23258 16540 23264
rect 18052 23316 18104 23322
rect 18052 23258 18104 23264
rect 16500 22098 16528 23258
rect 16764 23180 16816 23186
rect 16764 23122 16816 23128
rect 16776 22438 16804 23122
rect 18604 22772 18656 22778
rect 18604 22714 18656 22720
rect 16764 22432 16816 22438
rect 16764 22374 16816 22380
rect 16488 22092 16540 22098
rect 16488 22034 16540 22040
rect 16500 21690 16528 22034
rect 16488 21684 16540 21690
rect 16488 21626 16540 21632
rect 16396 21072 16448 21078
rect 16396 21014 16448 21020
rect 16396 20868 16448 20874
rect 16396 20810 16448 20816
rect 16408 20330 16436 20810
rect 16488 20800 16540 20806
rect 16488 20742 16540 20748
rect 16500 20330 16528 20742
rect 16672 20596 16724 20602
rect 16672 20538 16724 20544
rect 16396 20324 16448 20330
rect 16396 20266 16448 20272
rect 16488 20324 16540 20330
rect 16488 20266 16540 20272
rect 16408 19825 16436 20266
rect 16394 19816 16450 19825
rect 16394 19751 16450 19760
rect 16500 19514 16528 20266
rect 16580 19780 16632 19786
rect 16580 19722 16632 19728
rect 16592 19514 16620 19722
rect 16488 19508 16540 19514
rect 16488 19450 16540 19456
rect 16580 19508 16632 19514
rect 16580 19450 16632 19456
rect 16500 19224 16528 19450
rect 16580 19236 16632 19242
rect 16500 19196 16580 19224
rect 16580 19178 16632 19184
rect 16592 18970 16620 19178
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 16396 18692 16448 18698
rect 16396 18634 16448 18640
rect 16408 17241 16436 18634
rect 16580 17604 16632 17610
rect 16580 17546 16632 17552
rect 16394 17232 16450 17241
rect 16394 17167 16450 17176
rect 16592 17066 16620 17546
rect 16580 17060 16632 17066
rect 16580 17002 16632 17008
rect 16592 16250 16620 17002
rect 16580 16244 16632 16250
rect 16580 16186 16632 16192
rect 16684 15570 16712 20538
rect 16776 19258 16804 22374
rect 18616 22098 18644 22714
rect 17224 22092 17276 22098
rect 17224 22034 17276 22040
rect 18604 22092 18656 22098
rect 18604 22034 18656 22040
rect 17132 21956 17184 21962
rect 17132 21898 17184 21904
rect 16856 20800 16908 20806
rect 16856 20742 16908 20748
rect 16868 20058 16896 20742
rect 17040 20324 17092 20330
rect 17040 20266 17092 20272
rect 16856 20052 16908 20058
rect 16856 19994 16908 20000
rect 16868 19378 16896 19994
rect 16948 19848 17000 19854
rect 16948 19790 17000 19796
rect 16856 19372 16908 19378
rect 16856 19314 16908 19320
rect 16776 19230 16896 19258
rect 16764 17672 16816 17678
rect 16764 17614 16816 17620
rect 16776 17270 16804 17614
rect 16764 17264 16816 17270
rect 16764 17206 16816 17212
rect 16776 16726 16804 17206
rect 16764 16720 16816 16726
rect 16764 16662 16816 16668
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16670 15464 16726 15473
rect 16670 15399 16726 15408
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 16408 14958 16436 15302
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 16488 13932 16540 13938
rect 16488 13874 16540 13880
rect 16304 13456 16356 13462
rect 16304 13398 16356 13404
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 16316 11626 16344 12038
rect 16500 11762 16528 13874
rect 16580 13796 16632 13802
rect 16580 13738 16632 13744
rect 16592 12918 16620 13738
rect 16580 12912 16632 12918
rect 16580 12854 16632 12860
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 16304 11620 16356 11626
rect 16304 11562 16356 11568
rect 16316 11354 16344 11562
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 16132 10198 16160 10610
rect 16120 10192 16172 10198
rect 16120 10134 16172 10140
rect 16028 10124 16080 10130
rect 16028 10066 16080 10072
rect 16500 9994 16528 11698
rect 16580 11280 16632 11286
rect 16580 11222 16632 11228
rect 16592 10470 16620 11222
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16592 10198 16620 10406
rect 16580 10192 16632 10198
rect 16580 10134 16632 10140
rect 16488 9988 16540 9994
rect 16488 9930 16540 9936
rect 16488 9444 16540 9450
rect 16488 9386 16540 9392
rect 16212 8968 16264 8974
rect 15948 8928 16068 8956
rect 15842 8664 15898 8673
rect 15842 8599 15898 8608
rect 15856 7818 15884 8599
rect 15936 8288 15988 8294
rect 15936 8230 15988 8236
rect 15844 7812 15896 7818
rect 15844 7754 15896 7760
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 15856 5778 15884 6734
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15856 5370 15884 5714
rect 15844 5364 15896 5370
rect 15844 5306 15896 5312
rect 15948 5302 15976 8230
rect 15936 5296 15988 5302
rect 15936 5238 15988 5244
rect 15936 5092 15988 5098
rect 15936 5034 15988 5040
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 15948 4758 15976 5034
rect 15936 4752 15988 4758
rect 15936 4694 15988 4700
rect 15948 4282 15976 4694
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 16040 4154 16068 8928
rect 16212 8910 16264 8916
rect 16120 8560 16172 8566
rect 16120 8502 16172 8508
rect 16132 7886 16160 8502
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 16132 7546 16160 7822
rect 16120 7540 16172 7546
rect 16120 7482 16172 7488
rect 16224 6866 16252 8910
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16408 7546 16436 7890
rect 16500 7818 16528 9386
rect 16592 9178 16620 10134
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16488 7812 16540 7818
rect 16488 7754 16540 7760
rect 16592 7750 16620 8366
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16396 6928 16448 6934
rect 16396 6870 16448 6876
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16132 6458 16160 6802
rect 16120 6452 16172 6458
rect 16120 6394 16172 6400
rect 16304 6112 16356 6118
rect 16304 6054 16356 6060
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 16040 4126 16160 4154
rect 16224 4146 16252 4558
rect 15936 4004 15988 4010
rect 16132 3992 16160 4126
rect 16212 4140 16264 4146
rect 16212 4082 16264 4088
rect 15988 3964 16160 3992
rect 15936 3946 15988 3952
rect 15948 3738 15976 3946
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 15528 3488 15608 3516
rect 15476 3470 15528 3476
rect 15488 3194 15516 3470
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 13818 2136 13874 2145
rect 13818 2071 13874 2080
rect 14186 2136 14242 2145
rect 14186 2071 14242 2080
rect 12898 54 13032 82
rect 13832 82 13860 2071
rect 14476 2038 14504 2926
rect 15764 2922 15792 3674
rect 16224 3602 16252 4082
rect 16316 4010 16344 6054
rect 16408 5914 16436 6870
rect 16592 6225 16620 7686
rect 16578 6216 16634 6225
rect 16578 6151 16634 6160
rect 16396 5908 16448 5914
rect 16396 5850 16448 5856
rect 16580 5568 16632 5574
rect 16580 5510 16632 5516
rect 16592 5098 16620 5510
rect 16684 5302 16712 15399
rect 16868 13977 16896 19230
rect 16960 18970 16988 19790
rect 17052 19786 17080 20266
rect 17040 19780 17092 19786
rect 17040 19722 17092 19728
rect 17052 19446 17080 19722
rect 17040 19440 17092 19446
rect 17040 19382 17092 19388
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 17040 17672 17092 17678
rect 17040 17614 17092 17620
rect 16948 17536 17000 17542
rect 16948 17478 17000 17484
rect 16960 14618 16988 17478
rect 17052 17270 17080 17614
rect 17040 17264 17092 17270
rect 17040 17206 17092 17212
rect 17040 15088 17092 15094
rect 17040 15030 17092 15036
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 16854 13968 16910 13977
rect 16854 13903 16910 13912
rect 17052 13814 17080 15030
rect 16960 13786 17080 13814
rect 16960 13530 16988 13786
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 16764 13456 16816 13462
rect 16764 13398 16816 13404
rect 16856 13456 16908 13462
rect 16856 13398 16908 13404
rect 16776 12986 16804 13398
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 16868 12646 16896 13398
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16868 12102 16896 12582
rect 16856 12096 16908 12102
rect 16856 12038 16908 12044
rect 16960 11150 16988 13262
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 17052 11830 17080 12038
rect 17040 11824 17092 11830
rect 17040 11766 17092 11772
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16868 8430 16896 9454
rect 16960 8906 16988 9998
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 16948 8900 17000 8906
rect 16948 8842 17000 8848
rect 17052 8498 17080 8910
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 16672 5296 16724 5302
rect 16672 5238 16724 5244
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16672 5092 16724 5098
rect 16672 5034 16724 5040
rect 16684 4214 16712 5034
rect 16776 4826 16804 5170
rect 16764 4820 16816 4826
rect 16816 4780 16896 4808
rect 16764 4762 16816 4768
rect 16764 4480 16816 4486
rect 16764 4422 16816 4428
rect 16672 4208 16724 4214
rect 16672 4154 16724 4156
rect 16592 4150 16724 4154
rect 16592 4126 16712 4150
rect 16592 4010 16620 4126
rect 16304 4004 16356 4010
rect 16304 3946 16356 3952
rect 16580 4004 16632 4010
rect 16580 3946 16632 3952
rect 16212 3596 16264 3602
rect 16212 3538 16264 3544
rect 16028 3392 16080 3398
rect 16028 3334 16080 3340
rect 16040 2922 16068 3334
rect 16224 3040 16252 3538
rect 16592 3058 16620 3946
rect 16776 3738 16804 4422
rect 16868 4049 16896 4780
rect 16854 4040 16910 4049
rect 16854 3975 16910 3984
rect 16764 3732 16816 3738
rect 16764 3674 16816 3680
rect 16132 3012 16252 3040
rect 16580 3052 16632 3058
rect 15752 2916 15804 2922
rect 15752 2858 15804 2864
rect 16028 2916 16080 2922
rect 16028 2858 16080 2864
rect 14648 2848 14700 2854
rect 14648 2790 14700 2796
rect 14464 2032 14516 2038
rect 14464 1974 14516 1980
rect 13910 82 13966 480
rect 13832 54 13966 82
rect 14660 82 14688 2790
rect 16040 2582 16068 2858
rect 16028 2576 16080 2582
rect 16028 2518 16080 2524
rect 16132 2378 16160 3012
rect 16580 2994 16632 3000
rect 16212 2916 16264 2922
rect 16212 2858 16264 2864
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14922 82 14978 480
rect 14660 54 14978 82
rect 10782 0 10838 54
rect 11794 0 11850 54
rect 12898 0 12954 54
rect 13910 0 13966 54
rect 14922 0 14978 54
rect 15934 82 15990 480
rect 16224 82 16252 2858
rect 17144 2514 17172 21898
rect 17236 21350 17264 22034
rect 17592 22024 17644 22030
rect 17512 22001 17592 22012
rect 17498 21992 17592 22001
rect 17554 21984 17592 21992
rect 17592 21966 17644 21972
rect 17498 21927 17554 21936
rect 18328 21616 18380 21622
rect 18328 21558 18380 21564
rect 17960 21412 18012 21418
rect 17960 21354 18012 21360
rect 17224 21344 17276 21350
rect 17224 21286 17276 21292
rect 17236 15910 17264 21286
rect 17316 21004 17368 21010
rect 17316 20946 17368 20952
rect 17328 20913 17356 20946
rect 17314 20904 17370 20913
rect 17314 20839 17370 20848
rect 17328 20602 17356 20839
rect 17316 20596 17368 20602
rect 17316 20538 17368 20544
rect 17868 20392 17920 20398
rect 17868 20334 17920 20340
rect 17880 20058 17908 20334
rect 17868 20052 17920 20058
rect 17788 20012 17868 20040
rect 17316 19168 17368 19174
rect 17316 19110 17368 19116
rect 17500 19168 17552 19174
rect 17500 19110 17552 19116
rect 17328 17882 17356 19110
rect 17408 18896 17460 18902
rect 17408 18838 17460 18844
rect 17420 18426 17448 18838
rect 17408 18420 17460 18426
rect 17408 18362 17460 18368
rect 17316 17876 17368 17882
rect 17316 17818 17368 17824
rect 17408 17808 17460 17814
rect 17408 17750 17460 17756
rect 17420 17338 17448 17750
rect 17512 17610 17540 19110
rect 17592 18760 17644 18766
rect 17592 18702 17644 18708
rect 17604 18426 17632 18702
rect 17592 18420 17644 18426
rect 17592 18362 17644 18368
rect 17604 17882 17632 18362
rect 17684 18284 17736 18290
rect 17684 18226 17736 18232
rect 17592 17876 17644 17882
rect 17592 17818 17644 17824
rect 17500 17604 17552 17610
rect 17500 17546 17552 17552
rect 17696 17542 17724 18226
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 17408 17332 17460 17338
rect 17408 17274 17460 17280
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17420 16794 17448 17274
rect 17408 16788 17460 16794
rect 17408 16730 17460 16736
rect 17408 16516 17460 16522
rect 17408 16458 17460 16464
rect 17224 15904 17276 15910
rect 17224 15846 17276 15852
rect 17222 15736 17278 15745
rect 17222 15671 17278 15680
rect 17236 13462 17264 15671
rect 17316 15564 17368 15570
rect 17316 15506 17368 15512
rect 17328 15162 17356 15506
rect 17316 15156 17368 15162
rect 17316 15098 17368 15104
rect 17328 14482 17356 15098
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 17328 14074 17356 14418
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17224 13456 17276 13462
rect 17224 13398 17276 13404
rect 17224 13252 17276 13258
rect 17328 13240 17356 14010
rect 17420 13734 17448 16458
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 17408 13456 17460 13462
rect 17408 13398 17460 13404
rect 17276 13212 17356 13240
rect 17224 13194 17276 13200
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17328 10713 17356 12582
rect 17314 10704 17370 10713
rect 17314 10639 17370 10648
rect 17224 10532 17276 10538
rect 17224 10474 17276 10480
rect 17236 9110 17264 10474
rect 17224 9104 17276 9110
rect 17224 9046 17276 9052
rect 17236 8634 17264 9046
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17236 8022 17264 8570
rect 17224 8016 17276 8022
rect 17224 7958 17276 7964
rect 17236 7410 17264 7958
rect 17224 7404 17276 7410
rect 17224 7346 17276 7352
rect 17236 7002 17264 7346
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17236 6390 17264 6938
rect 17224 6384 17276 6390
rect 17224 6326 17276 6332
rect 17236 4758 17264 6326
rect 17328 5001 17356 10639
rect 17420 8362 17448 13398
rect 17408 8356 17460 8362
rect 17408 8298 17460 8304
rect 17420 8090 17448 8298
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17420 6730 17448 7822
rect 17512 7546 17540 17274
rect 17788 16946 17816 20012
rect 17868 19994 17920 20000
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17880 18766 17908 19246
rect 17868 18760 17920 18766
rect 17868 18702 17920 18708
rect 17880 18154 17908 18702
rect 17868 18148 17920 18154
rect 17868 18090 17920 18096
rect 17880 17678 17908 18090
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 17604 16918 17816 16946
rect 17604 14414 17632 16918
rect 17776 16788 17828 16794
rect 17776 16730 17828 16736
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17696 15434 17724 16526
rect 17788 16250 17816 16730
rect 17776 16244 17828 16250
rect 17776 16186 17828 16192
rect 17868 15904 17920 15910
rect 17788 15864 17868 15892
rect 17684 15428 17736 15434
rect 17684 15370 17736 15376
rect 17682 14920 17738 14929
rect 17682 14855 17738 14864
rect 17696 14822 17724 14855
rect 17684 14816 17736 14822
rect 17684 14758 17736 14764
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17604 14074 17632 14350
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17604 13841 17632 14010
rect 17590 13832 17646 13841
rect 17590 13767 17646 13776
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 17604 12306 17632 13670
rect 17788 12850 17816 15864
rect 17868 15846 17920 15852
rect 17972 15722 18000 21354
rect 18052 21344 18104 21350
rect 18052 21286 18104 21292
rect 17880 15694 18000 15722
rect 17880 13462 17908 15694
rect 17960 15632 18012 15638
rect 17960 15574 18012 15580
rect 17868 13456 17920 13462
rect 17868 13398 17920 13404
rect 17880 12986 17908 13398
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17684 12776 17736 12782
rect 17684 12718 17736 12724
rect 17696 12442 17724 12718
rect 17684 12436 17736 12442
rect 17684 12378 17736 12384
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17604 11762 17632 12242
rect 17696 11830 17724 12242
rect 17684 11824 17736 11830
rect 17684 11766 17736 11772
rect 17592 11756 17644 11762
rect 17592 11698 17644 11704
rect 17604 11098 17632 11698
rect 17788 11286 17816 12786
rect 17776 11280 17828 11286
rect 17776 11222 17828 11228
rect 17866 11248 17922 11257
rect 17866 11183 17922 11192
rect 17880 11150 17908 11183
rect 17868 11144 17920 11150
rect 17604 11070 17724 11098
rect 17868 11086 17920 11092
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17604 7721 17632 10950
rect 17696 8566 17724 11070
rect 17880 10810 17908 11086
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 17972 10606 18000 15574
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 17776 9444 17828 9450
rect 17776 9386 17828 9392
rect 17960 9444 18012 9450
rect 17960 9386 18012 9392
rect 17788 9042 17816 9386
rect 17972 9178 18000 9386
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 17776 9036 17828 9042
rect 17776 8978 17828 8984
rect 17684 8560 17736 8566
rect 17684 8502 17736 8508
rect 17590 7712 17646 7721
rect 17590 7647 17646 7656
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 18064 6934 18092 21286
rect 18144 21004 18196 21010
rect 18144 20946 18196 20952
rect 18156 20262 18184 20946
rect 18236 20800 18288 20806
rect 18236 20742 18288 20748
rect 18144 20256 18196 20262
rect 18144 20198 18196 20204
rect 18156 15638 18184 20198
rect 18144 15632 18196 15638
rect 18144 15574 18196 15580
rect 18144 14816 18196 14822
rect 18144 14758 18196 14764
rect 18156 13734 18184 14758
rect 18248 14550 18276 20742
rect 18340 16454 18368 21558
rect 18616 21554 18644 22034
rect 18604 21548 18656 21554
rect 18604 21490 18656 21496
rect 18420 21480 18472 21486
rect 18472 21440 18552 21468
rect 18616 21457 18644 21490
rect 18420 21422 18472 21428
rect 18524 21332 18552 21440
rect 18602 21448 18658 21457
rect 18602 21383 18658 21392
rect 18604 21344 18656 21350
rect 18524 21304 18604 21332
rect 18524 19446 18552 21304
rect 18604 21286 18656 21292
rect 18696 21004 18748 21010
rect 18696 20946 18748 20952
rect 18604 20392 18656 20398
rect 18604 20334 18656 20340
rect 18616 19718 18644 20334
rect 18708 20262 18736 20946
rect 19536 20942 19564 27526
rect 19812 27418 19840 27526
rect 19890 27520 19946 28000
rect 21362 27520 21418 28000
rect 22834 27520 22890 28000
rect 24306 27520 24362 28000
rect 25778 27520 25834 28000
rect 27250 27520 27306 28000
rect 19904 27418 19932 27520
rect 19812 27390 19932 27418
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 21272 24608 21324 24614
rect 21272 24550 21324 24556
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20902 24168 20958 24177
rect 20902 24103 20958 24112
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 20916 22710 20944 24103
rect 20904 22704 20956 22710
rect 21284 22681 21312 24550
rect 21376 22778 21404 27520
rect 21364 22772 21416 22778
rect 21364 22714 21416 22720
rect 20904 22646 20956 22652
rect 21270 22672 21326 22681
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 20916 21690 20944 22646
rect 21270 22607 21326 22616
rect 21272 22092 21324 22098
rect 21272 22034 21324 22040
rect 21284 21690 21312 22034
rect 20904 21684 20956 21690
rect 20904 21626 20956 21632
rect 21272 21684 21324 21690
rect 21272 21626 21324 21632
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 20904 21480 20956 21486
rect 20904 21422 20956 21428
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19524 20936 19576 20942
rect 19524 20878 19576 20884
rect 20352 20868 20404 20874
rect 20352 20810 20404 20816
rect 20444 20868 20496 20874
rect 20444 20810 20496 20816
rect 20364 20534 20392 20810
rect 18972 20528 19024 20534
rect 18972 20470 19024 20476
rect 20352 20528 20404 20534
rect 20352 20470 20404 20476
rect 18788 20324 18840 20330
rect 18788 20266 18840 20272
rect 18696 20256 18748 20262
rect 18696 20198 18748 20204
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18604 19508 18656 19514
rect 18604 19450 18656 19456
rect 18512 19440 18564 19446
rect 18512 19382 18564 19388
rect 18420 19372 18472 19378
rect 18420 19314 18472 19320
rect 18432 18358 18460 19314
rect 18420 18352 18472 18358
rect 18420 18294 18472 18300
rect 18432 16590 18460 18294
rect 18524 17338 18552 19382
rect 18616 19378 18644 19450
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 18616 18426 18644 19314
rect 18604 18420 18656 18426
rect 18604 18362 18656 18368
rect 18616 18222 18644 18362
rect 18604 18216 18656 18222
rect 18604 18158 18656 18164
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18512 17332 18564 17338
rect 18512 17274 18564 17280
rect 18510 17232 18566 17241
rect 18510 17167 18566 17176
rect 18420 16584 18472 16590
rect 18420 16526 18472 16532
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 18420 15632 18472 15638
rect 18420 15574 18472 15580
rect 18432 14822 18460 15574
rect 18524 14929 18552 17167
rect 18616 15366 18644 18022
rect 18604 15360 18656 15366
rect 18604 15302 18656 15308
rect 18604 14952 18656 14958
rect 18510 14920 18566 14929
rect 18604 14894 18656 14900
rect 18510 14855 18566 14864
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18236 14544 18288 14550
rect 18236 14486 18288 14492
rect 18328 14000 18380 14006
rect 18328 13942 18380 13948
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 18156 12714 18184 13670
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18144 12708 18196 12714
rect 18144 12650 18196 12656
rect 18248 11558 18276 13466
rect 18340 13326 18368 13942
rect 18420 13456 18472 13462
rect 18420 13398 18472 13404
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 18248 9722 18276 11494
rect 18340 11354 18368 13262
rect 18432 12986 18460 13398
rect 18420 12980 18472 12986
rect 18420 12922 18472 12928
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18328 11348 18380 11354
rect 18328 11290 18380 11296
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18340 9586 18368 10202
rect 18328 9580 18380 9586
rect 18328 9522 18380 9528
rect 18328 8832 18380 8838
rect 18328 8774 18380 8780
rect 18340 8362 18368 8774
rect 18328 8356 18380 8362
rect 18328 8298 18380 8304
rect 18340 8090 18368 8298
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18236 7472 18288 7478
rect 18236 7414 18288 7420
rect 18248 7274 18276 7414
rect 18144 7268 18196 7274
rect 18144 7210 18196 7216
rect 18236 7268 18288 7274
rect 18236 7210 18288 7216
rect 18156 7002 18184 7210
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 18052 6928 18104 6934
rect 18052 6870 18104 6876
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17408 6724 17460 6730
rect 17408 6666 17460 6672
rect 17604 5914 17632 6802
rect 18064 6458 18092 6870
rect 18248 6866 18276 7210
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 18052 6452 18104 6458
rect 18052 6394 18104 6400
rect 17500 5908 17552 5914
rect 17500 5850 17552 5856
rect 17592 5908 17644 5914
rect 17592 5850 17644 5856
rect 17408 5772 17460 5778
rect 17408 5714 17460 5720
rect 17420 5370 17448 5714
rect 17408 5364 17460 5370
rect 17408 5306 17460 5312
rect 17314 4992 17370 5001
rect 17314 4927 17370 4936
rect 17224 4752 17276 4758
rect 17224 4694 17276 4700
rect 17408 4752 17460 4758
rect 17408 4694 17460 4700
rect 17420 4146 17448 4694
rect 17512 4690 17540 5850
rect 18064 5778 18092 6394
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 18328 5772 18380 5778
rect 18328 5714 18380 5720
rect 18064 5370 18092 5714
rect 18340 5370 18368 5714
rect 18052 5364 18104 5370
rect 18052 5306 18104 5312
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 17500 4684 17552 4690
rect 17500 4626 17552 4632
rect 17512 4282 17540 4626
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 18248 4282 18276 4422
rect 17500 4276 17552 4282
rect 17500 4218 17552 4224
rect 18236 4276 18288 4282
rect 18236 4218 18288 4224
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 18248 4010 18276 4218
rect 18432 4185 18460 12038
rect 18524 10554 18552 14855
rect 18616 13462 18644 14894
rect 18604 13456 18656 13462
rect 18604 13398 18656 13404
rect 18708 12646 18736 20198
rect 18800 14618 18828 20266
rect 18880 19916 18932 19922
rect 18880 19858 18932 19864
rect 18892 18970 18920 19858
rect 18984 19242 19012 20470
rect 20168 20256 20220 20262
rect 20168 20198 20220 20204
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 19064 19780 19116 19786
rect 19064 19722 19116 19728
rect 19076 19514 19104 19722
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 18972 19236 19024 19242
rect 18972 19178 19024 19184
rect 18880 18964 18932 18970
rect 18880 18906 18932 18912
rect 18892 18426 18920 18906
rect 18880 18420 18932 18426
rect 18880 18362 18932 18368
rect 18880 17672 18932 17678
rect 18880 17614 18932 17620
rect 18892 17338 18920 17614
rect 18880 17332 18932 17338
rect 18880 17274 18932 17280
rect 18880 16992 18932 16998
rect 18880 16934 18932 16940
rect 18892 16454 18920 16934
rect 18984 16522 19012 19178
rect 18972 16516 19024 16522
rect 18972 16458 19024 16464
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18892 15910 18920 16390
rect 19076 16130 19104 19450
rect 19156 18964 19208 18970
rect 19156 18906 19208 18912
rect 19168 17882 19196 18906
rect 19156 17876 19208 17882
rect 19156 17818 19208 17824
rect 19156 17740 19208 17746
rect 19156 17682 19208 17688
rect 19168 16998 19196 17682
rect 19246 17096 19302 17105
rect 19246 17031 19302 17040
rect 19156 16992 19208 16998
rect 19156 16934 19208 16940
rect 19260 16726 19288 17031
rect 19248 16720 19300 16726
rect 19248 16662 19300 16668
rect 18984 16102 19104 16130
rect 19352 16114 19380 19790
rect 19984 19712 20036 19718
rect 19984 19654 20036 19660
rect 19996 19310 20024 19654
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 19524 19168 19576 19174
rect 19524 19110 19576 19116
rect 19432 18828 19484 18834
rect 19432 18770 19484 18776
rect 19444 18086 19472 18770
rect 19432 18080 19484 18086
rect 19432 18022 19484 18028
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19444 16522 19472 17138
rect 19432 16516 19484 16522
rect 19432 16458 19484 16464
rect 19340 16108 19392 16114
rect 18880 15904 18932 15910
rect 18880 15846 18932 15852
rect 18892 15638 18920 15846
rect 18880 15632 18932 15638
rect 18880 15574 18932 15580
rect 18984 15094 19012 16102
rect 19340 16050 19392 16056
rect 19064 16040 19116 16046
rect 19064 15982 19116 15988
rect 18972 15088 19024 15094
rect 18972 15030 19024 15036
rect 18788 14612 18840 14618
rect 18788 14554 18840 14560
rect 18800 13938 18828 14554
rect 18788 13932 18840 13938
rect 18788 13874 18840 13880
rect 19076 13734 19104 15982
rect 19352 15706 19380 16050
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19156 15360 19208 15366
rect 19156 15302 19208 15308
rect 19168 14958 19196 15302
rect 19444 15026 19472 16458
rect 19536 15502 19564 19110
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19996 17762 20024 19246
rect 20076 18624 20128 18630
rect 20076 18566 20128 18572
rect 20088 18154 20116 18566
rect 20076 18148 20128 18154
rect 20076 18090 20128 18096
rect 20088 17882 20116 18090
rect 20076 17876 20128 17882
rect 20076 17818 20128 17824
rect 19996 17734 20116 17762
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 19996 15910 20024 16594
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19996 15609 20024 15846
rect 19982 15600 20038 15609
rect 19982 15535 20038 15544
rect 19524 15496 19576 15502
rect 19524 15438 19576 15444
rect 19536 15162 19564 15438
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19984 15088 20036 15094
rect 19984 15030 20036 15036
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19156 14952 19208 14958
rect 19156 14894 19208 14900
rect 19168 14550 19196 14894
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19156 14544 19208 14550
rect 19156 14486 19208 14492
rect 19432 14544 19484 14550
rect 19432 14486 19484 14492
rect 19444 14074 19472 14486
rect 19996 14414 20024 15030
rect 19984 14408 20036 14414
rect 19984 14350 20036 14356
rect 19524 14340 19576 14346
rect 19524 14282 19576 14288
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19064 13728 19116 13734
rect 19064 13670 19116 13676
rect 18972 12776 19024 12782
rect 18972 12718 19024 12724
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18984 12170 19012 12718
rect 19076 12306 19104 13670
rect 19536 13530 19564 14282
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 19524 12640 19576 12646
rect 19524 12582 19576 12588
rect 19536 12374 19564 12582
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19996 12374 20024 14350
rect 20088 14006 20116 17734
rect 20180 14414 20208 20198
rect 20260 19916 20312 19922
rect 20260 19858 20312 19864
rect 20272 19174 20300 19858
rect 20352 19712 20404 19718
rect 20352 19654 20404 19660
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 20272 18873 20300 19110
rect 20258 18864 20314 18873
rect 20258 18799 20314 18808
rect 20260 18080 20312 18086
rect 20260 18022 20312 18028
rect 20272 17882 20300 18022
rect 20260 17876 20312 17882
rect 20260 17818 20312 17824
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 20272 17202 20300 17682
rect 20260 17196 20312 17202
rect 20260 17138 20312 17144
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 20076 14000 20128 14006
rect 20076 13942 20128 13948
rect 20272 13814 20300 17138
rect 20088 13786 20300 13814
rect 19524 12368 19576 12374
rect 19524 12310 19576 12316
rect 19984 12368 20036 12374
rect 19984 12310 20036 12316
rect 19064 12300 19116 12306
rect 19064 12242 19116 12248
rect 18972 12164 19024 12170
rect 18972 12106 19024 12112
rect 19536 11898 19564 12310
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 18972 11688 19024 11694
rect 18972 11630 19024 11636
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18800 11354 18828 11494
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18984 11286 19012 11630
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 18972 11280 19024 11286
rect 18972 11222 19024 11228
rect 19248 11212 19300 11218
rect 19248 11154 19300 11160
rect 19260 10606 19288 11154
rect 19248 10600 19300 10606
rect 18524 10526 18736 10554
rect 19248 10542 19300 10548
rect 18512 10464 18564 10470
rect 18512 10406 18564 10412
rect 18524 10198 18552 10406
rect 18512 10192 18564 10198
rect 18512 10134 18564 10140
rect 18604 10192 18656 10198
rect 18604 10134 18656 10140
rect 18524 9178 18552 10134
rect 18616 9382 18644 10134
rect 18604 9376 18656 9382
rect 18604 9318 18656 9324
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 18604 4480 18656 4486
rect 18602 4448 18604 4457
rect 18656 4448 18658 4457
rect 18602 4383 18658 4392
rect 18418 4176 18474 4185
rect 18616 4146 18644 4383
rect 18418 4111 18474 4120
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 18236 4004 18288 4010
rect 18236 3946 18288 3952
rect 18248 3670 18276 3946
rect 18708 3670 18736 10526
rect 18880 10056 18932 10062
rect 18880 9998 18932 10004
rect 18892 9654 18920 9998
rect 19260 9926 19288 10542
rect 19444 10538 19472 11290
rect 20088 11218 20116 13786
rect 20168 13320 20220 13326
rect 20168 13262 20220 13268
rect 20180 12986 20208 13262
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 20364 11830 20392 19654
rect 20456 14346 20484 20810
rect 20628 20800 20680 20806
rect 20628 20742 20680 20748
rect 20536 20324 20588 20330
rect 20536 20266 20588 20272
rect 20548 15026 20576 20266
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20548 14618 20576 14962
rect 20536 14612 20588 14618
rect 20536 14554 20588 14560
rect 20444 14340 20496 14346
rect 20444 14282 20496 14288
rect 20640 14226 20668 20742
rect 20812 20528 20864 20534
rect 20812 20470 20864 20476
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20732 19145 20760 20198
rect 20718 19136 20774 19145
rect 20718 19071 20774 19080
rect 20720 18692 20772 18698
rect 20720 18634 20772 18640
rect 20732 18222 20760 18634
rect 20720 18216 20772 18222
rect 20720 18158 20772 18164
rect 20732 17746 20760 18158
rect 20720 17740 20772 17746
rect 20720 17682 20772 17688
rect 20824 17678 20852 20470
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 20732 16794 20760 17138
rect 20812 16992 20864 16998
rect 20812 16934 20864 16940
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20824 15570 20852 16934
rect 20916 16114 20944 21422
rect 21548 21344 21600 21350
rect 21548 21286 21600 21292
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 20996 17876 21048 17882
rect 20996 17818 21048 17824
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20812 15564 20864 15570
rect 20812 15506 20864 15512
rect 20824 14890 20852 15506
rect 20812 14884 20864 14890
rect 20812 14826 20864 14832
rect 20640 14198 20852 14226
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20732 13190 20760 13874
rect 20536 13184 20588 13190
rect 20536 13126 20588 13132
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20548 12238 20576 13126
rect 20824 12850 20852 14198
rect 21008 13326 21036 17818
rect 21100 17202 21128 20198
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 21088 17196 21140 17202
rect 21088 17138 21140 17144
rect 21088 14544 21140 14550
rect 21088 14486 21140 14492
rect 21100 14074 21128 14486
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21088 13796 21140 13802
rect 21088 13738 21140 13744
rect 21100 13530 21128 13738
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 21100 12850 21128 13126
rect 20812 12844 20864 12850
rect 20812 12786 20864 12792
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20168 11824 20220 11830
rect 20168 11766 20220 11772
rect 20352 11824 20404 11830
rect 20352 11766 20404 11772
rect 20076 11212 20128 11218
rect 20076 11154 20128 11160
rect 19616 11144 19668 11150
rect 19616 11086 19668 11092
rect 19628 10606 19656 11086
rect 20180 11082 20208 11766
rect 20260 11552 20312 11558
rect 20260 11494 20312 11500
rect 20272 11150 20300 11494
rect 20364 11354 20392 11766
rect 20548 11762 20576 12174
rect 20536 11756 20588 11762
rect 20536 11698 20588 11704
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 20812 11212 20864 11218
rect 20812 11154 20864 11160
rect 20260 11144 20312 11150
rect 20260 11086 20312 11092
rect 20168 11076 20220 11082
rect 20168 11018 20220 11024
rect 20076 11008 20128 11014
rect 20076 10950 20128 10956
rect 19616 10600 19668 10606
rect 19536 10560 19616 10588
rect 19432 10532 19484 10538
rect 19432 10474 19484 10480
rect 19536 10266 19564 10560
rect 19616 10542 19668 10548
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19524 10260 19576 10266
rect 19524 10202 19576 10208
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 18880 9648 18932 9654
rect 18880 9590 18932 9596
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 18800 8022 18828 8978
rect 18892 8498 18920 9590
rect 18972 9444 19024 9450
rect 18972 9386 19024 9392
rect 18984 8566 19012 9386
rect 19156 9104 19208 9110
rect 19156 9046 19208 9052
rect 19168 8634 19196 9046
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 18972 8560 19024 8566
rect 18972 8502 19024 8508
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18788 8016 18840 8022
rect 18788 7958 18840 7964
rect 18984 7818 19012 8502
rect 19168 8294 19196 8570
rect 19156 8288 19208 8294
rect 19156 8230 19208 8236
rect 18788 7812 18840 7818
rect 18788 7754 18840 7760
rect 18972 7812 19024 7818
rect 18972 7754 19024 7760
rect 17868 3664 17920 3670
rect 17868 3606 17920 3612
rect 18236 3664 18288 3670
rect 18236 3606 18288 3612
rect 18696 3664 18748 3670
rect 18696 3606 18748 3612
rect 17880 3194 17908 3606
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18248 3194 18276 3470
rect 17868 3188 17920 3194
rect 17868 3130 17920 3136
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 17132 2508 17184 2514
rect 17132 2450 17184 2456
rect 16948 2100 17000 2106
rect 16948 2042 17000 2048
rect 15934 54 16252 82
rect 16960 82 16988 2042
rect 17038 82 17094 480
rect 16960 54 17094 82
rect 15934 0 15990 54
rect 17038 0 17094 54
rect 18050 82 18106 480
rect 18708 82 18736 3606
rect 18050 54 18736 82
rect 18800 82 18828 7754
rect 18984 7410 19012 7754
rect 18972 7404 19024 7410
rect 18972 7346 19024 7352
rect 19260 6322 19288 9862
rect 19536 9722 19564 10202
rect 19524 9716 19576 9722
rect 19524 9658 19576 9664
rect 20088 9586 20116 10950
rect 20824 10470 20852 11154
rect 21088 11144 21140 11150
rect 21088 11086 21140 11092
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 21100 10198 21128 11086
rect 21088 10192 21140 10198
rect 21088 10134 21140 10140
rect 20076 9580 20128 9586
rect 20076 9522 20128 9528
rect 20352 9580 20404 9586
rect 20352 9522 20404 9528
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19996 9042 20024 9318
rect 20088 9110 20116 9522
rect 20076 9104 20128 9110
rect 20076 9046 20128 9052
rect 19984 9036 20036 9042
rect 19984 8978 20036 8984
rect 19996 8634 20024 8978
rect 20364 8974 20392 9522
rect 21100 9178 21128 10134
rect 21192 10062 21220 19110
rect 21272 18624 21324 18630
rect 21272 18566 21324 18572
rect 21284 18154 21312 18566
rect 21560 18193 21588 21286
rect 21640 21004 21692 21010
rect 21640 20946 21692 20952
rect 21652 20602 21680 20946
rect 21640 20596 21692 20602
rect 21640 20538 21692 20544
rect 21732 19304 21784 19310
rect 21732 19246 21784 19252
rect 21640 18828 21692 18834
rect 21640 18770 21692 18776
rect 21652 18426 21680 18770
rect 21640 18420 21692 18426
rect 21640 18362 21692 18368
rect 21546 18184 21602 18193
rect 21272 18148 21324 18154
rect 21546 18119 21602 18128
rect 21272 18090 21324 18096
rect 21284 17338 21312 18090
rect 21364 18080 21416 18086
rect 21364 18022 21416 18028
rect 21376 17882 21404 18022
rect 21364 17876 21416 17882
rect 21364 17818 21416 17824
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 21560 17202 21588 18119
rect 21652 17746 21680 18362
rect 21640 17740 21692 17746
rect 21640 17682 21692 17688
rect 21652 17270 21680 17682
rect 21640 17264 21692 17270
rect 21640 17206 21692 17212
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 21548 17196 21600 17202
rect 21548 17138 21600 17144
rect 21284 11218 21312 17138
rect 21640 17060 21692 17066
rect 21640 17002 21692 17008
rect 21652 16726 21680 17002
rect 21364 16720 21416 16726
rect 21364 16662 21416 16668
rect 21640 16720 21692 16726
rect 21640 16662 21692 16668
rect 21376 15978 21404 16662
rect 21548 16108 21600 16114
rect 21548 16050 21600 16056
rect 21364 15972 21416 15978
rect 21364 15914 21416 15920
rect 21376 15706 21404 15914
rect 21560 15706 21588 16050
rect 21364 15700 21416 15706
rect 21364 15642 21416 15648
rect 21548 15700 21600 15706
rect 21548 15642 21600 15648
rect 21548 15496 21600 15502
rect 21548 15438 21600 15444
rect 21560 14822 21588 15438
rect 21548 14816 21600 14822
rect 21548 14758 21600 14764
rect 21456 13456 21508 13462
rect 21560 13444 21588 14758
rect 21652 14550 21680 16662
rect 21640 14544 21692 14550
rect 21640 14486 21692 14492
rect 21652 14006 21680 14486
rect 21640 14000 21692 14006
rect 21640 13942 21692 13948
rect 21744 13814 21772 19246
rect 21824 18760 21876 18766
rect 21824 18702 21876 18708
rect 21836 15570 21864 18702
rect 21916 15972 21968 15978
rect 21916 15914 21968 15920
rect 21824 15564 21876 15570
rect 21824 15506 21876 15512
rect 21836 14550 21864 15506
rect 21928 15026 21956 15914
rect 22020 15094 22048 21626
rect 22848 21418 22876 27520
rect 24320 25650 24348 27520
rect 25134 26752 25190 26761
rect 25134 26687 25190 26696
rect 24228 25622 24348 25650
rect 24032 24268 24084 24274
rect 24032 24210 24084 24216
rect 24044 23526 24072 24210
rect 24228 23633 24256 25622
rect 24766 25528 24822 25537
rect 24766 25463 24822 25472
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24780 23866 24808 25463
rect 25148 24954 25176 26687
rect 25136 24948 25188 24954
rect 25136 24890 25188 24896
rect 25148 24750 25176 24890
rect 25136 24744 25188 24750
rect 25136 24686 25188 24692
rect 25792 24410 25820 27520
rect 25780 24404 25832 24410
rect 25780 24346 25832 24352
rect 24768 23860 24820 23866
rect 24768 23802 24820 23808
rect 24214 23624 24270 23633
rect 24214 23559 24270 23568
rect 24032 23520 24084 23526
rect 24032 23462 24084 23468
rect 25320 23520 25372 23526
rect 25320 23462 25372 23468
rect 22836 21412 22888 21418
rect 22836 21354 22888 21360
rect 22652 21140 22704 21146
rect 22652 21082 22704 21088
rect 22284 20392 22336 20398
rect 22284 20334 22336 20340
rect 22296 19417 22324 20334
rect 22560 19848 22612 19854
rect 22560 19790 22612 19796
rect 22282 19408 22338 19417
rect 22282 19343 22338 19352
rect 22192 19168 22244 19174
rect 22192 19110 22244 19116
rect 22100 18896 22152 18902
rect 22100 18838 22152 18844
rect 22112 18086 22140 18838
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 22008 15088 22060 15094
rect 22008 15030 22060 15036
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 21824 14544 21876 14550
rect 21824 14486 21876 14492
rect 21916 14408 21968 14414
rect 21916 14350 21968 14356
rect 21928 14074 21956 14350
rect 22020 14346 22048 15030
rect 22008 14340 22060 14346
rect 22008 14282 22060 14288
rect 21916 14068 21968 14074
rect 21916 14010 21968 14016
rect 22020 13870 22048 14282
rect 21508 13416 21588 13444
rect 21652 13786 21772 13814
rect 22008 13864 22060 13870
rect 22008 13806 22060 13812
rect 21456 13398 21508 13404
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21376 12442 21404 13262
rect 21468 12986 21496 13398
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 21456 12980 21508 12986
rect 21456 12922 21508 12928
rect 21364 12436 21416 12442
rect 21364 12378 21416 12384
rect 21456 12300 21508 12306
rect 21456 12242 21508 12248
rect 21468 11558 21496 12242
rect 21456 11552 21508 11558
rect 21456 11494 21508 11500
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 21364 11008 21416 11014
rect 21364 10950 21416 10956
rect 21376 10674 21404 10950
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 21468 10606 21496 11494
rect 21456 10600 21508 10606
rect 21456 10542 21508 10548
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 21088 9172 21140 9178
rect 21088 9114 21140 9120
rect 21192 9110 21220 9998
rect 21364 9376 21416 9382
rect 21364 9318 21416 9324
rect 21180 9104 21232 9110
rect 21180 9046 21232 9052
rect 20352 8968 20404 8974
rect 20352 8910 20404 8916
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 19996 8362 20024 8570
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 19984 8356 20036 8362
rect 19984 8298 20036 8304
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19432 8016 19484 8022
rect 19432 7958 19484 7964
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19352 7188 19380 7822
rect 19444 7546 19472 7958
rect 20088 7750 20116 8434
rect 20364 8090 20392 8910
rect 21180 8900 21232 8906
rect 21180 8842 21232 8848
rect 20996 8288 21048 8294
rect 20996 8230 21048 8236
rect 20352 8084 20404 8090
rect 20352 8026 20404 8032
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20076 7744 20128 7750
rect 20076 7686 20128 7692
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19432 7200 19484 7206
rect 19352 7160 19432 7188
rect 19432 7142 19484 7148
rect 19444 6458 19472 7142
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 20088 7002 20116 7686
rect 20350 7440 20406 7449
rect 20260 7404 20312 7410
rect 20350 7375 20406 7384
rect 20260 7346 20312 7352
rect 20076 6996 20128 7002
rect 20076 6938 20128 6944
rect 20272 6934 20300 7346
rect 20260 6928 20312 6934
rect 20166 6896 20222 6905
rect 19524 6860 19576 6866
rect 19524 6802 19576 6808
rect 19616 6860 19668 6866
rect 20260 6870 20312 6876
rect 20166 6831 20222 6840
rect 19616 6802 19668 6808
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 19248 6316 19300 6322
rect 19248 6258 19300 6264
rect 18972 6248 19024 6254
rect 18972 6190 19024 6196
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18892 2446 18920 5646
rect 18984 3913 19012 6190
rect 19432 6180 19484 6186
rect 19432 6122 19484 6128
rect 19248 5908 19300 5914
rect 19248 5850 19300 5856
rect 19156 5160 19208 5166
rect 19156 5102 19208 5108
rect 18970 3904 19026 3913
rect 18970 3839 19026 3848
rect 19168 2496 19196 5102
rect 19260 4690 19288 5850
rect 19340 5160 19392 5166
rect 19340 5102 19392 5108
rect 19352 4826 19380 5102
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19248 4684 19300 4690
rect 19248 4626 19300 4632
rect 19260 4282 19288 4626
rect 19248 4276 19300 4282
rect 19248 4218 19300 4224
rect 19352 4214 19380 4762
rect 19444 4214 19472 6122
rect 19536 6118 19564 6802
rect 19628 6254 19656 6802
rect 19616 6248 19668 6254
rect 19616 6190 19668 6196
rect 19984 6248 20036 6254
rect 19984 6190 20036 6196
rect 19524 6112 19576 6118
rect 19524 6054 19576 6060
rect 19340 4208 19392 4214
rect 19340 4150 19392 4156
rect 19432 4208 19484 4214
rect 19432 4150 19484 4156
rect 19430 3904 19486 3913
rect 19430 3839 19486 3848
rect 19444 3058 19472 3839
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19536 2632 19564 6054
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19996 5778 20024 6190
rect 20076 6180 20128 6186
rect 20076 6122 20128 6128
rect 20088 5914 20116 6122
rect 20076 5908 20128 5914
rect 20076 5850 20128 5856
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 19996 5302 20024 5714
rect 19984 5296 20036 5302
rect 19984 5238 20036 5244
rect 20088 5234 20116 5850
rect 20076 5228 20128 5234
rect 20076 5170 20128 5176
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 20088 4010 20116 4082
rect 20076 4004 20128 4010
rect 20076 3946 20128 3952
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 20088 3738 20116 3946
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 19616 3596 19668 3602
rect 19616 3538 19668 3544
rect 19628 3126 19656 3538
rect 19616 3120 19668 3126
rect 19616 3062 19668 3068
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19536 2604 19656 2632
rect 19524 2508 19576 2514
rect 19168 2468 19524 2496
rect 19524 2450 19576 2456
rect 19628 2446 19656 2604
rect 18880 2440 18932 2446
rect 18880 2382 18932 2388
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 19628 2106 19656 2382
rect 19616 2100 19668 2106
rect 19616 2042 19668 2048
rect 19062 82 19118 480
rect 18800 54 19118 82
rect 18050 0 18106 54
rect 19062 0 19118 54
rect 20074 82 20130 480
rect 20180 82 20208 6831
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 20272 3738 20300 3878
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 20364 3602 20392 7375
rect 20628 7268 20680 7274
rect 20628 7210 20680 7216
rect 20640 7002 20668 7210
rect 20628 6996 20680 7002
rect 20628 6938 20680 6944
rect 20628 6656 20680 6662
rect 20732 6644 20760 7822
rect 21008 6934 21036 8230
rect 21088 8016 21140 8022
rect 21088 7958 21140 7964
rect 21100 7546 21128 7958
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 21192 7274 21220 8842
rect 21272 8832 21324 8838
rect 21272 8774 21324 8780
rect 21284 7478 21312 8774
rect 21376 8294 21404 9318
rect 21468 8537 21496 10542
rect 21560 9518 21588 13262
rect 21652 10169 21680 13786
rect 22112 13326 22140 18022
rect 22204 16130 22232 19110
rect 22284 18624 22336 18630
rect 22284 18566 22336 18572
rect 22296 16590 22324 18566
rect 22284 16584 22336 16590
rect 22284 16526 22336 16532
rect 22296 16250 22324 16526
rect 22284 16244 22336 16250
rect 22284 16186 22336 16192
rect 22204 16102 22324 16130
rect 22192 15360 22244 15366
rect 22192 15302 22244 15308
rect 22204 14890 22232 15302
rect 22192 14884 22244 14890
rect 22192 14826 22244 14832
rect 22204 14618 22232 14826
rect 22192 14612 22244 14618
rect 22192 14554 22244 14560
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 22192 12912 22244 12918
rect 22192 12854 22244 12860
rect 21824 12640 21876 12646
rect 21824 12582 21876 12588
rect 21732 11552 21784 11558
rect 21732 11494 21784 11500
rect 21744 10810 21772 11494
rect 21732 10804 21784 10810
rect 21732 10746 21784 10752
rect 21836 10577 21864 12582
rect 21916 12096 21968 12102
rect 21916 12038 21968 12044
rect 21928 11608 21956 12038
rect 22204 11801 22232 12854
rect 22190 11792 22246 11801
rect 22190 11727 22246 11736
rect 22008 11620 22060 11626
rect 21928 11580 22008 11608
rect 21822 10568 21878 10577
rect 21822 10503 21878 10512
rect 21732 10464 21784 10470
rect 21732 10406 21784 10412
rect 21638 10160 21694 10169
rect 21638 10095 21694 10104
rect 21548 9512 21600 9518
rect 21548 9454 21600 9460
rect 21640 9104 21692 9110
rect 21640 9046 21692 9052
rect 21652 8634 21680 9046
rect 21640 8628 21692 8634
rect 21640 8570 21692 8576
rect 21454 8528 21510 8537
rect 21454 8463 21510 8472
rect 21364 8288 21416 8294
rect 21364 8230 21416 8236
rect 21272 7472 21324 7478
rect 21272 7414 21324 7420
rect 21180 7268 21232 7274
rect 21180 7210 21232 7216
rect 20996 6928 21048 6934
rect 20996 6870 21048 6876
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20680 6616 20760 6644
rect 20628 6598 20680 6604
rect 20640 5370 20668 6598
rect 20824 6186 20852 6734
rect 21008 6458 21036 6870
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 20812 6180 20864 6186
rect 20812 6122 20864 6128
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 21008 5166 21036 6394
rect 21192 5302 21220 7210
rect 21376 5846 21404 8230
rect 21364 5840 21416 5846
rect 21364 5782 21416 5788
rect 21272 5772 21324 5778
rect 21272 5714 21324 5720
rect 21180 5296 21232 5302
rect 21180 5238 21232 5244
rect 20996 5160 21048 5166
rect 20996 5102 21048 5108
rect 20444 5024 20496 5030
rect 20444 4966 20496 4972
rect 20456 4146 20484 4966
rect 20904 4820 20956 4826
rect 20904 4762 20956 4768
rect 20916 4282 20944 4762
rect 20996 4616 21048 4622
rect 20996 4558 21048 4564
rect 20904 4276 20956 4282
rect 20904 4218 20956 4224
rect 21008 4154 21036 4558
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 20824 4126 21036 4154
rect 20352 3596 20404 3602
rect 20352 3538 20404 3544
rect 20824 3534 20852 4126
rect 21008 4010 21036 4126
rect 20996 4004 21048 4010
rect 20996 3946 21048 3952
rect 21192 3602 21220 5238
rect 21284 5030 21312 5714
rect 21272 5024 21324 5030
rect 21272 4966 21324 4972
rect 21284 4729 21312 4966
rect 21270 4720 21326 4729
rect 21270 4655 21326 4664
rect 21272 4616 21324 4622
rect 21272 4558 21324 4564
rect 21284 4146 21312 4558
rect 21272 4140 21324 4146
rect 21272 4082 21324 4088
rect 21180 3596 21232 3602
rect 21180 3538 21232 3544
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 20352 3392 20404 3398
rect 20352 3334 20404 3340
rect 20364 3194 20392 3334
rect 20352 3188 20404 3194
rect 20352 3130 20404 3136
rect 20996 2984 21048 2990
rect 20996 2926 21048 2932
rect 21008 2854 21036 2926
rect 20996 2848 21048 2854
rect 20996 2790 21048 2796
rect 21088 2848 21140 2854
rect 21088 2790 21140 2796
rect 21008 2009 21036 2790
rect 21100 2582 21128 2790
rect 21192 2650 21220 3538
rect 21180 2644 21232 2650
rect 21180 2586 21232 2592
rect 21088 2576 21140 2582
rect 21088 2518 21140 2524
rect 21272 2372 21324 2378
rect 21272 2314 21324 2320
rect 20994 2000 21050 2009
rect 20994 1935 21050 1944
rect 20074 54 20208 82
rect 21178 82 21234 480
rect 21284 82 21312 2314
rect 21744 134 21772 10406
rect 21928 10062 21956 11580
rect 22008 11562 22060 11568
rect 22192 11348 22244 11354
rect 22192 11290 22244 11296
rect 22204 10538 22232 11290
rect 22296 11234 22324 16102
rect 22376 13864 22428 13870
rect 22376 13806 22428 13812
rect 22388 13190 22416 13806
rect 22376 13184 22428 13190
rect 22376 13126 22428 13132
rect 22388 12918 22416 13126
rect 22376 12912 22428 12918
rect 22376 12854 22428 12860
rect 22468 12368 22520 12374
rect 22468 12310 22520 12316
rect 22376 12232 22428 12238
rect 22376 12174 22428 12180
rect 22388 11830 22416 12174
rect 22480 11898 22508 12310
rect 22468 11892 22520 11898
rect 22468 11834 22520 11840
rect 22376 11824 22428 11830
rect 22376 11766 22428 11772
rect 22296 11206 22416 11234
rect 22284 11144 22336 11150
rect 22284 11086 22336 11092
rect 22192 10532 22244 10538
rect 22192 10474 22244 10480
rect 22296 10470 22324 11086
rect 22284 10464 22336 10470
rect 22284 10406 22336 10412
rect 21916 10056 21968 10062
rect 21916 9998 21968 10004
rect 21916 9716 21968 9722
rect 21916 9658 21968 9664
rect 21824 7336 21876 7342
rect 21822 7304 21824 7313
rect 21876 7304 21878 7313
rect 21822 7239 21878 7248
rect 21836 7206 21864 7239
rect 21824 7200 21876 7206
rect 21824 7142 21876 7148
rect 21928 6254 21956 9658
rect 22296 9586 22324 10406
rect 22284 9580 22336 9586
rect 22284 9522 22336 9528
rect 22388 8430 22416 11206
rect 22468 8900 22520 8906
rect 22468 8842 22520 8848
rect 22376 8424 22428 8430
rect 22376 8366 22428 8372
rect 22008 7744 22060 7750
rect 22008 7686 22060 7692
rect 22020 7324 22048 7686
rect 22100 7336 22152 7342
rect 22020 7296 22100 7324
rect 22020 6254 22048 7296
rect 22100 7278 22152 7284
rect 21916 6248 21968 6254
rect 21916 6190 21968 6196
rect 22008 6248 22060 6254
rect 22008 6190 22060 6196
rect 21824 6112 21876 6118
rect 21824 6054 21876 6060
rect 21836 5234 21864 6054
rect 21928 5710 21956 6190
rect 22020 5778 22048 6190
rect 22008 5772 22060 5778
rect 22008 5714 22060 5720
rect 22284 5772 22336 5778
rect 22284 5714 22336 5720
rect 21916 5704 21968 5710
rect 21916 5646 21968 5652
rect 21824 5228 21876 5234
rect 21824 5170 21876 5176
rect 21836 4826 21864 5170
rect 22296 4826 22324 5714
rect 21824 4820 21876 4826
rect 21824 4762 21876 4768
rect 22284 4820 22336 4826
rect 22284 4762 22336 4768
rect 22006 4720 22062 4729
rect 22006 4655 22062 4664
rect 22020 4078 22048 4655
rect 21824 4072 21876 4078
rect 21824 4014 21876 4020
rect 22008 4072 22060 4078
rect 22008 4014 22060 4020
rect 21836 3670 21864 4014
rect 22100 4004 22152 4010
rect 22100 3946 22152 3952
rect 22008 3936 22060 3942
rect 22008 3878 22060 3884
rect 21824 3664 21876 3670
rect 22020 3641 22048 3878
rect 21824 3606 21876 3612
rect 22006 3632 22062 3641
rect 22112 3602 22140 3946
rect 22006 3567 22062 3576
rect 22100 3596 22152 3602
rect 22100 3538 22152 3544
rect 22112 3194 22140 3538
rect 22192 3460 22244 3466
rect 22192 3402 22244 3408
rect 22100 3188 22152 3194
rect 22100 3130 22152 3136
rect 21916 3120 21968 3126
rect 21916 3062 21968 3068
rect 21178 54 21312 82
rect 21732 128 21784 134
rect 21732 70 21784 76
rect 21928 82 21956 3062
rect 22008 2848 22060 2854
rect 22008 2790 22060 2796
rect 22020 1873 22048 2790
rect 22204 2310 22232 3402
rect 22480 3398 22508 8842
rect 22572 7002 22600 19790
rect 22664 15609 22692 21082
rect 23664 19848 23716 19854
rect 23664 19790 23716 19796
rect 22836 18828 22888 18834
rect 22836 18770 22888 18776
rect 22848 18086 22876 18770
rect 22836 18080 22888 18086
rect 22836 18022 22888 18028
rect 22744 17536 22796 17542
rect 22744 17478 22796 17484
rect 22756 17134 22784 17478
rect 22744 17128 22796 17134
rect 22744 17070 22796 17076
rect 22848 16794 22876 18022
rect 23020 17740 23072 17746
rect 23020 17682 23072 17688
rect 23032 17338 23060 17682
rect 23480 17672 23532 17678
rect 23480 17614 23532 17620
rect 23020 17332 23072 17338
rect 23020 17274 23072 17280
rect 22928 17128 22980 17134
rect 22928 17070 22980 17076
rect 22836 16788 22888 16794
rect 22836 16730 22888 16736
rect 22836 16652 22888 16658
rect 22940 16640 22968 17070
rect 22888 16612 22968 16640
rect 22836 16594 22888 16600
rect 22848 15910 22876 16594
rect 22836 15904 22888 15910
rect 22836 15846 22888 15852
rect 22650 15600 22706 15609
rect 22650 15535 22706 15544
rect 22664 13938 22692 15535
rect 22848 14278 22876 15846
rect 22928 14476 22980 14482
rect 23032 14464 23060 17274
rect 23112 16652 23164 16658
rect 23112 16594 23164 16600
rect 23124 16250 23152 16594
rect 23388 16584 23440 16590
rect 23388 16526 23440 16532
rect 23112 16244 23164 16250
rect 23112 16186 23164 16192
rect 23124 15162 23152 16186
rect 23296 16040 23348 16046
rect 23296 15982 23348 15988
rect 23204 15904 23256 15910
rect 23204 15846 23256 15852
rect 23216 15638 23244 15846
rect 23204 15632 23256 15638
rect 23204 15574 23256 15580
rect 23112 15156 23164 15162
rect 23112 15098 23164 15104
rect 23124 14482 23152 15098
rect 23216 15094 23244 15574
rect 23204 15088 23256 15094
rect 23204 15030 23256 15036
rect 23308 14550 23336 15982
rect 23400 15570 23428 16526
rect 23388 15564 23440 15570
rect 23388 15506 23440 15512
rect 23400 15162 23428 15506
rect 23388 15156 23440 15162
rect 23388 15098 23440 15104
rect 23492 14618 23520 17614
rect 23572 16992 23624 16998
rect 23572 16934 23624 16940
rect 23480 14612 23532 14618
rect 23480 14554 23532 14560
rect 23296 14544 23348 14550
rect 23296 14486 23348 14492
rect 22980 14436 23060 14464
rect 23112 14476 23164 14482
rect 22928 14418 22980 14424
rect 23112 14418 23164 14424
rect 22836 14272 22888 14278
rect 22836 14214 22888 14220
rect 22652 13932 22704 13938
rect 22652 13874 22704 13880
rect 22848 13814 22876 14214
rect 22940 14074 22968 14418
rect 22928 14068 22980 14074
rect 22928 14010 22980 14016
rect 23124 14006 23152 14418
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 23112 14000 23164 14006
rect 23112 13942 23164 13948
rect 23020 13932 23072 13938
rect 23020 13874 23072 13880
rect 22848 13786 22968 13814
rect 22940 12288 22968 13786
rect 22756 12260 22968 12288
rect 22652 12232 22704 12238
rect 22652 12174 22704 12180
rect 22664 12102 22692 12174
rect 22652 12096 22704 12102
rect 22652 12038 22704 12044
rect 22664 11762 22692 12038
rect 22652 11756 22704 11762
rect 22652 11698 22704 11704
rect 22756 10130 22784 12260
rect 22928 12164 22980 12170
rect 22928 12106 22980 12112
rect 22836 11892 22888 11898
rect 22836 11834 22888 11840
rect 22848 11354 22876 11834
rect 22836 11348 22888 11354
rect 22836 11290 22888 11296
rect 22834 10704 22890 10713
rect 22834 10639 22890 10648
rect 22848 10606 22876 10639
rect 22836 10600 22888 10606
rect 22836 10542 22888 10548
rect 22744 10124 22796 10130
rect 22744 10066 22796 10072
rect 22756 9722 22784 10066
rect 22744 9716 22796 9722
rect 22744 9658 22796 9664
rect 22940 9586 22968 12106
rect 22928 9580 22980 9586
rect 22928 9522 22980 9528
rect 22744 9512 22796 9518
rect 22744 9454 22796 9460
rect 22836 9512 22888 9518
rect 22836 9454 22888 9460
rect 22756 9178 22784 9454
rect 22744 9172 22796 9178
rect 22744 9114 22796 9120
rect 22756 8974 22784 9114
rect 22744 8968 22796 8974
rect 22744 8910 22796 8916
rect 22744 8356 22796 8362
rect 22744 8298 22796 8304
rect 22756 8022 22784 8298
rect 22744 8016 22796 8022
rect 22744 7958 22796 7964
rect 22756 7546 22784 7958
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 22652 7268 22704 7274
rect 22652 7210 22704 7216
rect 22560 6996 22612 7002
rect 22560 6938 22612 6944
rect 22664 6798 22692 7210
rect 22756 6934 22784 7482
rect 22744 6928 22796 6934
rect 22744 6870 22796 6876
rect 22652 6792 22704 6798
rect 22652 6734 22704 6740
rect 22664 6458 22692 6734
rect 22652 6452 22704 6458
rect 22652 6394 22704 6400
rect 22756 6390 22784 6870
rect 22848 6866 22876 9454
rect 22928 9036 22980 9042
rect 22928 8978 22980 8984
rect 22940 8294 22968 8978
rect 23032 8906 23060 13874
rect 23296 13728 23348 13734
rect 23296 13670 23348 13676
rect 23308 13462 23336 13670
rect 23296 13456 23348 13462
rect 23296 13398 23348 13404
rect 23112 12640 23164 12646
rect 23112 12582 23164 12588
rect 23124 9500 23152 12582
rect 23296 12164 23348 12170
rect 23296 12106 23348 12112
rect 23204 10124 23256 10130
rect 23204 10066 23256 10072
rect 23216 9654 23244 10066
rect 23204 9648 23256 9654
rect 23204 9590 23256 9596
rect 23124 9472 23244 9500
rect 23112 9172 23164 9178
rect 23112 9114 23164 9120
rect 23020 8900 23072 8906
rect 23020 8842 23072 8848
rect 23124 8634 23152 9114
rect 23216 8922 23244 9472
rect 23308 9110 23336 12106
rect 23400 10130 23428 14010
rect 23492 13938 23520 14554
rect 23480 13932 23532 13938
rect 23480 13874 23532 13880
rect 23584 13394 23612 16934
rect 23676 16726 23704 19790
rect 24044 19514 24072 23462
rect 24676 23180 24728 23186
rect 24676 23122 24728 23128
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24688 22778 24716 23122
rect 24676 22772 24728 22778
rect 24676 22714 24728 22720
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24688 20466 24716 22714
rect 25042 21720 25098 21729
rect 25042 21655 25098 21664
rect 24676 20460 24728 20466
rect 24676 20402 24728 20408
rect 25056 20398 25084 21655
rect 24216 20392 24268 20398
rect 24216 20334 24268 20340
rect 25044 20392 25096 20398
rect 25044 20334 25096 20340
rect 24124 19848 24176 19854
rect 24124 19790 24176 19796
rect 24032 19508 24084 19514
rect 24032 19450 24084 19456
rect 23754 19136 23810 19145
rect 23754 19071 23810 19080
rect 23664 16720 23716 16726
rect 23664 16662 23716 16668
rect 23664 16448 23716 16454
rect 23664 16390 23716 16396
rect 23572 13388 23624 13394
rect 23572 13330 23624 13336
rect 23584 12986 23612 13330
rect 23676 13258 23704 16390
rect 23768 13394 23796 19071
rect 23848 17740 23900 17746
rect 23848 17682 23900 17688
rect 23860 17066 23888 17682
rect 23848 17060 23900 17066
rect 23848 17002 23900 17008
rect 23860 16454 23888 17002
rect 23848 16448 23900 16454
rect 23848 16390 23900 16396
rect 24032 16448 24084 16454
rect 24032 16390 24084 16396
rect 24044 16114 24072 16390
rect 24032 16108 24084 16114
rect 24032 16050 24084 16056
rect 23940 16040 23992 16046
rect 23940 15982 23992 15988
rect 23848 13456 23900 13462
rect 23848 13398 23900 13404
rect 23756 13388 23808 13394
rect 23756 13330 23808 13336
rect 23664 13252 23716 13258
rect 23664 13194 23716 13200
rect 23860 12986 23888 13398
rect 23572 12980 23624 12986
rect 23572 12922 23624 12928
rect 23848 12980 23900 12986
rect 23848 12922 23900 12928
rect 23480 11280 23532 11286
rect 23480 11222 23532 11228
rect 23492 10810 23520 11222
rect 23664 11144 23716 11150
rect 23664 11086 23716 11092
rect 23480 10804 23532 10810
rect 23480 10746 23532 10752
rect 23492 10538 23520 10746
rect 23480 10532 23532 10538
rect 23480 10474 23532 10480
rect 23676 10198 23704 11086
rect 23756 10532 23808 10538
rect 23756 10474 23808 10480
rect 23768 10266 23796 10474
rect 23756 10260 23808 10266
rect 23756 10202 23808 10208
rect 23664 10192 23716 10198
rect 23664 10134 23716 10140
rect 23388 10124 23440 10130
rect 23388 10066 23440 10072
rect 23400 9466 23428 10066
rect 23572 10056 23624 10062
rect 23572 9998 23624 10004
rect 23400 9450 23520 9466
rect 23400 9444 23532 9450
rect 23400 9438 23480 9444
rect 23480 9386 23532 9392
rect 23296 9104 23348 9110
rect 23296 9046 23348 9052
rect 23480 9036 23532 9042
rect 23480 8978 23532 8984
rect 23216 8894 23336 8922
rect 23112 8628 23164 8634
rect 23112 8570 23164 8576
rect 23112 8424 23164 8430
rect 23112 8366 23164 8372
rect 22928 8288 22980 8294
rect 22928 8230 22980 8236
rect 22836 6860 22888 6866
rect 22836 6802 22888 6808
rect 22744 6384 22796 6390
rect 22744 6326 22796 6332
rect 22756 5846 22784 6326
rect 22744 5840 22796 5846
rect 22744 5782 22796 5788
rect 22756 5370 22784 5782
rect 22744 5364 22796 5370
rect 22744 5306 22796 5312
rect 22744 5024 22796 5030
rect 22744 4966 22796 4972
rect 22756 4758 22784 4966
rect 22744 4752 22796 4758
rect 22744 4694 22796 4700
rect 22756 4282 22784 4694
rect 22928 4616 22980 4622
rect 22928 4558 22980 4564
rect 22744 4276 22796 4282
rect 22744 4218 22796 4224
rect 22836 4140 22888 4146
rect 22940 4128 22968 4558
rect 22888 4100 22968 4128
rect 22836 4082 22888 4088
rect 22742 4040 22798 4049
rect 22742 3975 22798 3984
rect 22756 3942 22784 3975
rect 22744 3936 22796 3942
rect 22744 3878 22796 3884
rect 22940 3738 22968 4100
rect 22928 3732 22980 3738
rect 22928 3674 22980 3680
rect 22468 3392 22520 3398
rect 22468 3334 22520 3340
rect 22652 3392 22704 3398
rect 22652 3334 22704 3340
rect 22664 2990 22692 3334
rect 22652 2984 22704 2990
rect 22652 2926 22704 2932
rect 22664 2582 22692 2926
rect 22652 2576 22704 2582
rect 22652 2518 22704 2524
rect 23124 2417 23152 8366
rect 23204 5568 23256 5574
rect 23204 5510 23256 5516
rect 23216 5370 23244 5510
rect 23204 5364 23256 5370
rect 23204 5306 23256 5312
rect 23308 5137 23336 8894
rect 23386 8664 23442 8673
rect 23386 8599 23442 8608
rect 23400 8566 23428 8599
rect 23388 8560 23440 8566
rect 23388 8502 23440 8508
rect 23400 8294 23428 8502
rect 23492 8294 23520 8978
rect 23584 8974 23612 9998
rect 23664 9376 23716 9382
rect 23664 9318 23716 9324
rect 23572 8968 23624 8974
rect 23572 8910 23624 8916
rect 23388 8288 23440 8294
rect 23388 8230 23440 8236
rect 23480 8288 23532 8294
rect 23480 8230 23532 8236
rect 23400 7274 23428 8230
rect 23676 7834 23704 9318
rect 23952 9058 23980 15982
rect 24032 15972 24084 15978
rect 24032 15914 24084 15920
rect 24044 15706 24072 15914
rect 24032 15700 24084 15706
rect 24032 15642 24084 15648
rect 24032 15564 24084 15570
rect 24032 15506 24084 15512
rect 24044 11150 24072 15506
rect 24136 11898 24164 19790
rect 24228 15570 24256 20334
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24952 19236 25004 19242
rect 24952 19178 25004 19184
rect 24860 19168 24912 19174
rect 24766 19136 24822 19145
rect 24860 19110 24912 19116
rect 24766 19071 24822 19080
rect 24676 18624 24728 18630
rect 24676 18566 24728 18572
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24688 18222 24716 18566
rect 24780 18426 24808 19071
rect 24768 18420 24820 18426
rect 24768 18362 24820 18368
rect 24676 18216 24728 18222
rect 24676 18158 24728 18164
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24688 17270 24716 17682
rect 24676 17264 24728 17270
rect 24676 17206 24728 17212
rect 24768 16788 24820 16794
rect 24768 16730 24820 16736
rect 24676 16720 24728 16726
rect 24676 16662 24728 16668
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24688 16250 24716 16662
rect 24676 16244 24728 16250
rect 24676 16186 24728 16192
rect 24780 16182 24808 16730
rect 24768 16176 24820 16182
rect 24768 16118 24820 16124
rect 24216 15564 24268 15570
rect 24216 15506 24268 15512
rect 24676 15360 24728 15366
rect 24676 15302 24728 15308
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24688 15162 24716 15302
rect 24676 15156 24728 15162
rect 24872 15144 24900 19110
rect 24964 18290 24992 19178
rect 25044 18828 25096 18834
rect 25044 18770 25096 18776
rect 24952 18284 25004 18290
rect 24952 18226 25004 18232
rect 24964 16590 24992 18226
rect 25056 18086 25084 18770
rect 25136 18624 25188 18630
rect 25136 18566 25188 18572
rect 25044 18080 25096 18086
rect 25044 18022 25096 18028
rect 24952 16584 25004 16590
rect 24952 16526 25004 16532
rect 24952 15360 25004 15366
rect 24952 15302 25004 15308
rect 24676 15098 24728 15104
rect 24780 15116 24900 15144
rect 24688 14890 24716 15098
rect 24676 14884 24728 14890
rect 24676 14826 24728 14832
rect 24780 14618 24808 15116
rect 24964 15026 24992 15302
rect 24952 15020 25004 15026
rect 24952 14962 25004 14968
rect 24860 14816 24912 14822
rect 24860 14758 24912 14764
rect 24768 14612 24820 14618
rect 24768 14554 24820 14560
rect 24676 14544 24728 14550
rect 24676 14486 24728 14492
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24688 14074 24716 14486
rect 24780 14074 24808 14554
rect 24676 14068 24728 14074
rect 24676 14010 24728 14016
rect 24768 14068 24820 14074
rect 24768 14010 24820 14016
rect 24688 13530 24716 14010
rect 24676 13524 24728 13530
rect 24676 13466 24728 13472
rect 24216 13252 24268 13258
rect 24216 13194 24268 13200
rect 24124 11892 24176 11898
rect 24124 11834 24176 11840
rect 24032 11144 24084 11150
rect 24032 11086 24084 11092
rect 24124 9512 24176 9518
rect 24228 9500 24256 13194
rect 24676 13184 24728 13190
rect 24676 13126 24728 13132
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24688 12714 24716 13126
rect 24492 12708 24544 12714
rect 24492 12650 24544 12656
rect 24676 12708 24728 12714
rect 24676 12650 24728 12656
rect 24504 12442 24532 12650
rect 24492 12436 24544 12442
rect 24492 12378 24544 12384
rect 24768 12368 24820 12374
rect 24768 12310 24820 12316
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24584 11620 24636 11626
rect 24584 11562 24636 11568
rect 24596 11354 24624 11562
rect 24780 11558 24808 12310
rect 24768 11552 24820 11558
rect 24768 11494 24820 11500
rect 24584 11348 24636 11354
rect 24636 11308 24716 11336
rect 24584 11290 24636 11296
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24688 10810 24716 11308
rect 24780 11218 24808 11494
rect 24768 11212 24820 11218
rect 24768 11154 24820 11160
rect 24676 10804 24728 10810
rect 24676 10746 24728 10752
rect 24584 10600 24636 10606
rect 24584 10542 24636 10548
rect 24596 10266 24624 10542
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24176 9472 24256 9500
rect 24124 9454 24176 9460
rect 24136 9178 24164 9454
rect 24124 9172 24176 9178
rect 24124 9114 24176 9120
rect 23952 9030 24072 9058
rect 24872 9042 24900 14758
rect 24952 14408 25004 14414
rect 24952 14350 25004 14356
rect 24964 12918 24992 14350
rect 24952 12912 25004 12918
rect 24952 12854 25004 12860
rect 25056 12374 25084 18022
rect 25148 13530 25176 18566
rect 25226 18184 25282 18193
rect 25226 18119 25282 18128
rect 25240 17134 25268 18119
rect 25228 17128 25280 17134
rect 25228 17070 25280 17076
rect 25228 16584 25280 16590
rect 25228 16526 25280 16532
rect 25240 15026 25268 16526
rect 25228 15020 25280 15026
rect 25228 14962 25280 14968
rect 25226 14920 25282 14929
rect 25226 14855 25282 14864
rect 25240 13870 25268 14855
rect 25228 13864 25280 13870
rect 25228 13806 25280 13812
rect 25136 13524 25188 13530
rect 25136 13466 25188 13472
rect 25148 12850 25176 13466
rect 25226 13424 25282 13433
rect 25226 13359 25282 13368
rect 25136 12844 25188 12850
rect 25136 12786 25188 12792
rect 25044 12368 25096 12374
rect 25044 12310 25096 12316
rect 25056 12102 25084 12310
rect 25044 12096 25096 12102
rect 25044 12038 25096 12044
rect 25056 11830 25084 12038
rect 25044 11824 25096 11830
rect 25044 11766 25096 11772
rect 25240 11234 25268 13359
rect 25148 11206 25268 11234
rect 25044 10056 25096 10062
rect 25044 9998 25096 10004
rect 25056 9722 25084 9998
rect 25044 9716 25096 9722
rect 25044 9658 25096 9664
rect 25148 9518 25176 11206
rect 25228 11144 25280 11150
rect 25228 11086 25280 11092
rect 25240 10810 25268 11086
rect 25228 10804 25280 10810
rect 25228 10746 25280 10752
rect 25136 9512 25188 9518
rect 25136 9454 25188 9460
rect 23940 8832 23992 8838
rect 23940 8774 23992 8780
rect 23952 8498 23980 8774
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 23848 8356 23900 8362
rect 23848 8298 23900 8304
rect 23860 7954 23888 8298
rect 24044 8090 24072 9030
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24872 8294 24900 8978
rect 25228 8424 25280 8430
rect 25042 8392 25098 8401
rect 25228 8366 25280 8372
rect 25042 8327 25098 8336
rect 24124 8288 24176 8294
rect 24124 8230 24176 8236
rect 24860 8288 24912 8294
rect 24860 8230 24912 8236
rect 24032 8084 24084 8090
rect 24032 8026 24084 8032
rect 23848 7948 23900 7954
rect 23848 7890 23900 7896
rect 23584 7806 23704 7834
rect 23584 7410 23612 7806
rect 24136 7750 24164 8230
rect 24676 7948 24728 7954
rect 24676 7890 24728 7896
rect 23756 7744 23808 7750
rect 23662 7712 23718 7721
rect 23756 7686 23808 7692
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 23662 7647 23718 7656
rect 23572 7404 23624 7410
rect 23572 7346 23624 7352
rect 23388 7268 23440 7274
rect 23388 7210 23440 7216
rect 23294 5128 23350 5137
rect 23294 5063 23350 5072
rect 23676 3194 23704 7647
rect 23768 7206 23796 7686
rect 23848 7336 23900 7342
rect 23848 7278 23900 7284
rect 23756 7200 23808 7206
rect 23756 7142 23808 7148
rect 23860 6662 23888 7278
rect 24032 6792 24084 6798
rect 24032 6734 24084 6740
rect 23848 6656 23900 6662
rect 23848 6598 23900 6604
rect 23860 6254 23888 6598
rect 23938 6352 23994 6361
rect 23938 6287 23994 6296
rect 23848 6248 23900 6254
rect 23848 6190 23900 6196
rect 23756 5636 23808 5642
rect 23756 5578 23808 5584
rect 23768 5098 23796 5578
rect 23848 5364 23900 5370
rect 23848 5306 23900 5312
rect 23860 5098 23888 5306
rect 23756 5092 23808 5098
rect 23756 5034 23808 5040
rect 23848 5092 23900 5098
rect 23848 5034 23900 5040
rect 23768 4826 23796 5034
rect 23756 4820 23808 4826
rect 23756 4762 23808 4768
rect 23664 3188 23716 3194
rect 23664 3130 23716 3136
rect 23952 3058 23980 6287
rect 24044 4622 24072 6734
rect 24136 5234 24164 7686
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24688 7206 24716 7890
rect 25056 7342 25084 8327
rect 25044 7336 25096 7342
rect 25044 7278 25096 7284
rect 24676 7200 24728 7206
rect 24676 7142 24728 7148
rect 24216 6928 24268 6934
rect 24216 6870 24268 6876
rect 24228 6458 24256 6870
rect 24688 6798 24716 7142
rect 24952 6928 25004 6934
rect 24952 6870 25004 6876
rect 24676 6792 24728 6798
rect 24676 6734 24728 6740
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24964 6458 24992 6870
rect 25134 6760 25190 6769
rect 25134 6695 25190 6704
rect 24216 6452 24268 6458
rect 24216 6394 24268 6400
rect 24952 6452 25004 6458
rect 24952 6394 25004 6400
rect 25148 6254 25176 6695
rect 24308 6248 24360 6254
rect 25136 6248 25188 6254
rect 24308 6190 24360 6196
rect 24950 6216 25006 6225
rect 24320 5846 24348 6190
rect 25136 6190 25188 6196
rect 24950 6151 25006 6160
rect 24308 5840 24360 5846
rect 24308 5782 24360 5788
rect 24216 5772 24268 5778
rect 24216 5714 24268 5720
rect 24228 5370 24256 5714
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24216 5364 24268 5370
rect 24216 5306 24268 5312
rect 24124 5228 24176 5234
rect 24124 5170 24176 5176
rect 24582 5128 24638 5137
rect 24582 5063 24638 5072
rect 24766 5128 24822 5137
rect 24766 5063 24822 5072
rect 24596 4690 24624 5063
rect 24780 4826 24808 5063
rect 24768 4820 24820 4826
rect 24768 4762 24820 4768
rect 24584 4684 24636 4690
rect 24636 4644 24716 4672
rect 24584 4626 24636 4632
rect 24032 4616 24084 4622
rect 24032 4558 24084 4564
rect 24216 4548 24268 4554
rect 24216 4490 24268 4496
rect 24030 4448 24086 4457
rect 24030 4383 24086 4392
rect 24044 4282 24072 4383
rect 24032 4276 24084 4282
rect 24032 4218 24084 4224
rect 24228 4214 24256 4490
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24688 4214 24716 4644
rect 24216 4208 24268 4214
rect 24216 4150 24268 4156
rect 24676 4208 24728 4214
rect 24676 4150 24728 4156
rect 24964 3602 24992 6151
rect 25136 5772 25188 5778
rect 25136 5714 25188 5720
rect 25148 4486 25176 5714
rect 25136 4480 25188 4486
rect 25136 4422 25188 4428
rect 25148 3738 25176 4422
rect 25240 4282 25268 8366
rect 25332 6458 25360 23462
rect 27264 23322 27292 27520
rect 27252 23316 27304 23322
rect 27252 23258 27304 23264
rect 27618 20904 27674 20913
rect 27618 20839 27674 20848
rect 27632 20534 27660 20839
rect 27620 20528 27672 20534
rect 27620 20470 27672 20476
rect 25504 18828 25556 18834
rect 25504 18770 25556 18776
rect 25516 18086 25544 18770
rect 25504 18080 25556 18086
rect 25504 18022 25556 18028
rect 25410 17912 25466 17921
rect 25410 17847 25466 17856
rect 25424 17338 25452 17847
rect 25412 17332 25464 17338
rect 25412 17274 25464 17280
rect 25412 15564 25464 15570
rect 25412 15506 25464 15512
rect 25424 14822 25452 15506
rect 25412 14816 25464 14822
rect 25412 14758 25464 14764
rect 25410 14512 25466 14521
rect 25410 14447 25466 14456
rect 25424 14074 25452 14447
rect 25412 14068 25464 14074
rect 25412 14010 25464 14016
rect 25516 13433 25544 18022
rect 27620 17536 27672 17542
rect 27620 17478 27672 17484
rect 25594 16552 25650 16561
rect 25594 16487 25650 16496
rect 25608 16250 25636 16487
rect 25596 16244 25648 16250
rect 25596 16186 25648 16192
rect 25502 13424 25558 13433
rect 25412 13388 25464 13394
rect 25502 13359 25558 13368
rect 25412 13330 25464 13336
rect 25424 12986 25452 13330
rect 27632 13297 27660 17478
rect 27710 14648 27766 14657
rect 27710 14583 27766 14592
rect 27724 13394 27752 14583
rect 27712 13388 27764 13394
rect 27712 13330 27764 13336
rect 27618 13288 27674 13297
rect 27618 13223 27674 13232
rect 25504 13184 25556 13190
rect 25504 13126 25556 13132
rect 25412 12980 25464 12986
rect 25412 12922 25464 12928
rect 25412 12232 25464 12238
rect 25412 12174 25464 12180
rect 25424 11898 25452 12174
rect 25412 11892 25464 11898
rect 25412 11834 25464 11840
rect 25410 10160 25466 10169
rect 25410 10095 25466 10104
rect 25424 9722 25452 10095
rect 25412 9716 25464 9722
rect 25412 9658 25464 9664
rect 25410 8936 25466 8945
rect 25410 8871 25466 8880
rect 25424 8634 25452 8871
rect 25412 8628 25464 8634
rect 25412 8570 25464 8576
rect 25412 8288 25464 8294
rect 25412 8230 25464 8236
rect 25320 6452 25372 6458
rect 25320 6394 25372 6400
rect 25424 5001 25452 8230
rect 25410 4992 25466 5001
rect 25410 4927 25466 4936
rect 25228 4276 25280 4282
rect 25228 4218 25280 4224
rect 25136 3732 25188 3738
rect 25136 3674 25188 3680
rect 24216 3596 24268 3602
rect 24216 3538 24268 3544
rect 24952 3596 25004 3602
rect 24952 3538 25004 3544
rect 24228 3126 24256 3538
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24964 3194 24992 3538
rect 24952 3188 25004 3194
rect 24952 3130 25004 3136
rect 24216 3120 24268 3126
rect 24216 3062 24268 3068
rect 23940 3052 23992 3058
rect 23940 2994 23992 3000
rect 23110 2408 23166 2417
rect 23110 2343 23166 2352
rect 23940 2372 23992 2378
rect 23940 2314 23992 2320
rect 22192 2304 22244 2310
rect 22192 2246 22244 2252
rect 22006 1864 22062 1873
rect 22006 1799 22062 1808
rect 22190 82 22246 480
rect 21928 54 22246 82
rect 20074 0 20130 54
rect 21178 0 21234 54
rect 22190 0 22246 54
rect 23202 128 23258 480
rect 23202 76 23204 128
rect 23256 76 23258 128
rect 23202 0 23258 76
rect 23952 82 23980 2314
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24214 82 24270 480
rect 23952 54 24270 82
rect 24214 0 24270 54
rect 25318 82 25374 480
rect 25516 82 25544 13126
rect 25594 11520 25650 11529
rect 25594 11455 25650 11464
rect 25608 10810 25636 11455
rect 25596 10804 25648 10810
rect 25596 10746 25648 10752
rect 25596 10600 25648 10606
rect 25596 10542 25648 10548
rect 25608 4554 25636 10542
rect 25596 4548 25648 4554
rect 25596 4490 25648 4496
rect 27528 3120 27580 3126
rect 27618 3088 27674 3097
rect 27580 3068 27618 3074
rect 27528 3062 27618 3068
rect 27540 3046 27618 3062
rect 27618 3023 27674 3032
rect 26424 2372 26476 2378
rect 26424 2314 26476 2320
rect 25318 54 25544 82
rect 26330 82 26386 480
rect 26436 82 26464 2314
rect 27066 1728 27122 1737
rect 27066 1663 27122 1672
rect 26330 54 26464 82
rect 27080 82 27108 1663
rect 27342 82 27398 480
rect 27080 54 27398 82
rect 25318 0 25374 54
rect 26330 0 26386 54
rect 27342 0 27398 54
<< via2 >>
rect 1214 26832 1270 26888
rect 110 13912 166 13968
rect 110 11192 166 11248
rect 1582 24112 1638 24168
rect 1582 21256 1638 21312
rect 1582 20032 1638 20088
rect 1582 18672 1638 18728
rect 1306 15680 1362 15736
rect 1582 17448 1638 17504
rect 1582 16904 1638 16960
rect 1582 13776 1638 13832
rect 1858 25336 1914 25392
rect 1858 22616 1914 22672
rect 2042 20304 2098 20360
rect 2042 15988 2044 16008
rect 2044 15988 2096 16008
rect 2096 15988 2098 16008
rect 2042 15952 2098 15988
rect 2778 22344 2834 22400
rect 2318 15136 2374 15192
rect 1766 9832 1822 9888
rect 1582 7928 1638 7984
rect 2134 9968 2190 10024
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 3698 19896 3754 19952
rect 3238 18672 3294 18728
rect 3054 15136 3110 15192
rect 3330 14456 3386 14512
rect 3238 13912 3294 13968
rect 2870 12688 2926 12744
rect 2778 11328 2834 11384
rect 2870 9832 2926 9888
rect 1582 6704 1638 6760
rect 3054 9424 3110 9480
rect 3146 9288 3202 9344
rect 2594 8744 2650 8800
rect 1950 5344 2006 5400
rect 1858 2352 1914 2408
rect 2594 4256 2650 4312
rect 2778 4120 2834 4176
rect 2502 1672 2558 1728
rect 3330 12144 3386 12200
rect 3422 9696 3478 9752
rect 3882 12824 3938 12880
rect 3698 9560 3754 9616
rect 3606 9288 3662 9344
rect 4526 13776 4582 13832
rect 4158 11192 4214 11248
rect 4894 14728 4950 14784
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5814 19760 5870 19816
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 6274 19624 6330 19680
rect 6182 18536 6238 18592
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5354 13912 5410 13968
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5170 13640 5226 13696
rect 5078 12280 5134 12336
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 4802 11736 4858 11792
rect 4618 10104 4674 10160
rect 4158 9716 4214 9752
rect 4158 9696 4160 9716
rect 4160 9696 4212 9716
rect 4212 9696 4214 9716
rect 4342 9560 4398 9616
rect 3974 9016 4030 9072
rect 3330 7656 3386 7712
rect 4342 9288 4398 9344
rect 4342 8880 4398 8936
rect 4434 8744 4490 8800
rect 3698 7656 3754 7712
rect 3790 5344 3846 5400
rect 4618 5344 4674 5400
rect 3790 3168 3846 3224
rect 3974 2896 4030 2952
rect 5354 12144 5410 12200
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 6366 11328 6422 11384
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5354 9832 5410 9888
rect 5630 9968 5686 10024
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5354 7248 5410 7304
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 7470 17176 7526 17232
rect 7194 16632 7250 16688
rect 7010 13912 7066 13968
rect 6734 9424 6790 9480
rect 6458 9036 6514 9072
rect 6458 9016 6460 9036
rect 6460 9016 6512 9036
rect 6512 9016 6514 9036
rect 6642 7928 6698 7984
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5538 4664 5594 4720
rect 5446 3168 5502 3224
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 6182 2352 6238 2408
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6090 2080 6146 2136
rect 7470 14864 7526 14920
rect 7378 13776 7434 13832
rect 8758 22616 8814 22672
rect 8114 20304 8170 20360
rect 7746 13640 7802 13696
rect 8574 20168 8630 20224
rect 8574 19488 8630 19544
rect 9218 21664 9274 21720
rect 9126 17040 9182 17096
rect 7654 12144 7710 12200
rect 6366 1128 6422 1184
rect 9034 13368 9090 13424
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10782 21936 10838 21992
rect 9678 20848 9734 20904
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10138 18672 10194 18728
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10690 15952 10746 16008
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10690 13232 10746 13288
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 11058 13912 11114 13968
rect 9034 10512 9090 10568
rect 8022 5344 8078 5400
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 9034 2352 9090 2408
rect 9310 40 9366 96
rect 10046 10240 10102 10296
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 12070 19896 12126 19952
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 11702 14456 11758 14512
rect 11886 9832 11942 9888
rect 11610 7928 11666 7984
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 11058 5072 11114 5128
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 12070 12824 12126 12880
rect 12438 15952 12494 16008
rect 12070 4256 12126 4312
rect 11886 2896 11942 2952
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 12990 18536 13046 18592
rect 13358 22480 13414 22536
rect 13726 16632 13782 16688
rect 13266 14456 13322 14512
rect 12806 10512 12862 10568
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 13910 12144 13966 12200
rect 14554 21664 14610 21720
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14646 19624 14702 19680
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14738 18536 14794 18592
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14462 13776 14518 13832
rect 14094 6296 14150 6352
rect 14094 5344 14150 5400
rect 13634 5072 13690 5128
rect 12990 2896 13046 2952
rect 12070 1944 12126 2000
rect 12438 1808 12494 1864
rect 14462 9832 14518 9888
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 15198 13912 15254 13968
rect 14922 13776 14978 13832
rect 14738 13368 14794 13424
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 15106 12688 15162 12744
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 15290 6704 15346 6760
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15290 4936 15346 4992
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14738 4256 14794 4312
rect 14462 3576 14518 3632
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 16118 20304 16174 20360
rect 18234 23568 18290 23624
rect 18510 23432 18566 23488
rect 16394 19760 16450 19816
rect 16394 17176 16450 17232
rect 16670 15408 16726 15464
rect 15842 8608 15898 8664
rect 13818 2080 13874 2136
rect 14186 2080 14242 2136
rect 16578 6160 16634 6216
rect 16854 13912 16910 13968
rect 16854 3984 16910 4040
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 17498 21936 17554 21992
rect 17314 20848 17370 20904
rect 17222 15680 17278 15736
rect 17314 10648 17370 10704
rect 17682 14864 17738 14920
rect 17590 13776 17646 13832
rect 17866 11192 17922 11248
rect 17590 7656 17646 7712
rect 18602 21392 18658 21448
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 20902 24112 20958 24168
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 21270 22616 21326 22672
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 18510 17176 18566 17232
rect 18510 14864 18566 14920
rect 17314 4936 17370 4992
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19246 17040 19302 17096
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19982 15544 20038 15600
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 20258 18808 20314 18864
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 18602 4428 18604 4448
rect 18604 4428 18656 4448
rect 18656 4428 18658 4448
rect 18602 4392 18658 4428
rect 18418 4120 18474 4176
rect 20718 19080 20774 19136
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 21546 18128 21602 18184
rect 25134 26696 25190 26752
rect 24766 25472 24822 25528
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24214 23568 24270 23624
rect 22282 19352 22338 19408
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 20350 7384 20406 7440
rect 20166 6840 20222 6896
rect 18970 3848 19026 3904
rect 19430 3848 19486 3904
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 22190 11736 22246 11792
rect 21822 10512 21878 10568
rect 21638 10104 21694 10160
rect 21454 8472 21510 8528
rect 21270 4664 21326 4720
rect 20994 1944 21050 2000
rect 21822 7284 21824 7304
rect 21824 7284 21876 7304
rect 21876 7284 21878 7304
rect 21822 7248 21878 7284
rect 22006 4664 22062 4720
rect 22006 3576 22062 3632
rect 22650 15544 22706 15600
rect 22834 10648 22890 10704
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 25042 21664 25098 21720
rect 23754 19080 23810 19136
rect 22742 3984 22798 4040
rect 23386 8608 23442 8664
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24766 19080 24822 19136
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 25226 18128 25282 18184
rect 25226 14864 25282 14920
rect 25226 13368 25282 13424
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 25042 8336 25098 8392
rect 23662 7656 23718 7712
rect 23294 5072 23350 5128
rect 23938 6296 23994 6352
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 25134 6704 25190 6760
rect 24950 6160 25006 6216
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24582 5072 24638 5128
rect 24766 5072 24822 5128
rect 24030 4392 24086 4448
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 27618 20848 27674 20904
rect 25410 17856 25466 17912
rect 25410 14456 25466 14512
rect 25594 16496 25650 16552
rect 25502 13368 25558 13424
rect 27710 14592 27766 14648
rect 27618 13232 27674 13288
rect 25410 10104 25466 10160
rect 25410 8880 25466 8936
rect 25410 4936 25466 4992
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 23110 2352 23166 2408
rect 22006 1808 22062 1864
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 25594 11464 25650 11520
rect 27618 3032 27674 3088
rect 27066 1672 27122 1728
<< metal3 >>
rect 0 27208 480 27328
rect 27520 27208 28000 27328
rect 62 26890 122 27208
rect 1209 26890 1275 26893
rect 62 26888 1275 26890
rect 62 26832 1214 26888
rect 1270 26832 1275 26888
rect 62 26830 1275 26832
rect 1209 26827 1275 26830
rect 25129 26754 25195 26757
rect 27662 26754 27722 27208
rect 25129 26752 27722 26754
rect 25129 26696 25134 26752
rect 25190 26696 27722 26752
rect 25129 26694 27722 26696
rect 25129 26691 25195 26694
rect 27520 25984 28000 26104
rect 0 25848 480 25968
rect 62 25394 122 25848
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 24761 25530 24827 25533
rect 27662 25530 27722 25984
rect 24761 25528 27722 25530
rect 24761 25472 24766 25528
rect 24822 25472 27722 25528
rect 24761 25470 27722 25472
rect 24761 25467 24827 25470
rect 1853 25394 1919 25397
rect 62 25392 1919 25394
rect 62 25336 1858 25392
rect 1914 25336 1919 25392
rect 62 25334 1919 25336
rect 1853 25331 1919 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 27520 24624 28000 24744
rect 0 24488 480 24608
rect 10277 24512 10597 24513
rect 62 24170 122 24488
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 1577 24170 1643 24173
rect 62 24168 1643 24170
rect 62 24112 1582 24168
rect 1638 24112 1643 24168
rect 62 24110 1643 24112
rect 1577 24107 1643 24110
rect 20897 24170 20963 24173
rect 27662 24170 27722 24624
rect 20897 24168 27722 24170
rect 20897 24112 20902 24168
rect 20958 24112 27722 24168
rect 20897 24110 27722 24112
rect 20897 24107 20963 24110
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 18229 23626 18295 23629
rect 24209 23626 24275 23629
rect 18229 23624 24275 23626
rect 18229 23568 18234 23624
rect 18290 23568 24214 23624
rect 24270 23568 24275 23624
rect 18229 23566 24275 23568
rect 18229 23563 18295 23566
rect 24209 23563 24275 23566
rect 18505 23490 18571 23493
rect 18638 23490 18644 23492
rect 18505 23488 18644 23490
rect 18505 23432 18510 23488
rect 18566 23432 18644 23488
rect 18505 23430 18644 23432
rect 18505 23427 18571 23430
rect 18638 23428 18644 23430
rect 18708 23428 18714 23492
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 27520 23400 28000 23520
rect 19610 23359 19930 23360
rect 0 23128 480 23248
rect 62 22674 122 23128
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 1853 22674 1919 22677
rect 62 22672 1919 22674
rect 62 22616 1858 22672
rect 1914 22616 1919 22672
rect 62 22614 1919 22616
rect 1853 22611 1919 22614
rect 8753 22674 8819 22677
rect 21265 22674 21331 22677
rect 8753 22672 21331 22674
rect 8753 22616 8758 22672
rect 8814 22616 21270 22672
rect 21326 22616 21331 22672
rect 8753 22614 21331 22616
rect 8753 22611 8819 22614
rect 21265 22611 21331 22614
rect 13353 22538 13419 22541
rect 27662 22538 27722 23400
rect 13353 22536 27722 22538
rect 13353 22480 13358 22536
rect 13414 22480 27722 22536
rect 13353 22478 27722 22480
rect 13353 22475 13419 22478
rect 2773 22402 2839 22405
rect 2773 22400 4170 22402
rect 2773 22344 2778 22400
rect 2834 22344 4170 22400
rect 2773 22342 4170 22344
rect 2773 22339 2839 22342
rect 4110 22130 4170 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 27520 22176 28000 22296
rect 15510 22130 15516 22132
rect 4110 22070 15516 22130
rect 15510 22068 15516 22070
rect 15580 22068 15586 22132
rect 10777 21994 10843 21997
rect 17493 21994 17559 21997
rect 10777 21992 17559 21994
rect 10777 21936 10782 21992
rect 10838 21936 17498 21992
rect 17554 21936 17559 21992
rect 10777 21934 17559 21936
rect 10777 21931 10843 21934
rect 17493 21931 17559 21934
rect 0 21768 480 21888
rect 5610 21792 5930 21793
rect 62 21314 122 21768
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 9213 21722 9279 21725
rect 14549 21722 14615 21725
rect 9213 21720 14615 21722
rect 9213 21664 9218 21720
rect 9274 21664 14554 21720
rect 14610 21664 14615 21720
rect 9213 21662 14615 21664
rect 9213 21659 9279 21662
rect 14549 21659 14615 21662
rect 25037 21722 25103 21725
rect 27662 21722 27722 22176
rect 25037 21720 27722 21722
rect 25037 21664 25042 21720
rect 25098 21664 27722 21720
rect 25037 21662 27722 21664
rect 25037 21659 25103 21662
rect 18454 21388 18460 21452
rect 18524 21450 18530 21452
rect 18597 21450 18663 21453
rect 18524 21448 18663 21450
rect 18524 21392 18602 21448
rect 18658 21392 18663 21448
rect 18524 21390 18663 21392
rect 18524 21388 18530 21390
rect 18597 21387 18663 21390
rect 1577 21314 1643 21317
rect 62 21312 1643 21314
rect 62 21256 1582 21312
rect 1638 21256 1643 21312
rect 62 21254 1643 21256
rect 1577 21251 1643 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 9673 20906 9739 20909
rect 17309 20906 17375 20909
rect 9673 20904 17375 20906
rect 9673 20848 9678 20904
rect 9734 20848 17314 20904
rect 17370 20848 17375 20904
rect 9673 20846 17375 20848
rect 9673 20843 9739 20846
rect 17309 20843 17375 20846
rect 27520 20904 28000 20936
rect 27520 20848 27618 20904
rect 27674 20848 28000 20904
rect 27520 20816 28000 20848
rect 5610 20704 5930 20705
rect 0 20544 480 20664
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 62 20090 122 20544
rect 2037 20362 2103 20365
rect 8109 20362 8175 20365
rect 16113 20362 16179 20365
rect 2037 20360 4170 20362
rect 2037 20304 2042 20360
rect 2098 20304 4170 20360
rect 2037 20302 4170 20304
rect 2037 20299 2103 20302
rect 4110 20226 4170 20302
rect 8109 20360 16179 20362
rect 8109 20304 8114 20360
rect 8170 20304 16118 20360
rect 16174 20304 16179 20360
rect 8109 20302 16179 20304
rect 8109 20299 8175 20302
rect 16113 20299 16179 20302
rect 8569 20226 8635 20229
rect 4110 20224 8635 20226
rect 4110 20168 8574 20224
rect 8630 20168 8635 20224
rect 4110 20166 8635 20168
rect 8569 20163 8635 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 1577 20090 1643 20093
rect 62 20088 1643 20090
rect 62 20032 1582 20088
rect 1638 20032 1643 20088
rect 62 20030 1643 20032
rect 1577 20027 1643 20030
rect 3693 19954 3759 19957
rect 12065 19954 12131 19957
rect 3693 19952 12131 19954
rect 3693 19896 3698 19952
rect 3754 19896 12070 19952
rect 12126 19896 12131 19952
rect 3693 19894 12131 19896
rect 3693 19891 3759 19894
rect 12065 19891 12131 19894
rect 5809 19818 5875 19821
rect 16389 19818 16455 19821
rect 5809 19816 16455 19818
rect 5809 19760 5814 19816
rect 5870 19760 16394 19816
rect 16450 19760 16455 19816
rect 5809 19758 16455 19760
rect 5809 19755 5875 19758
rect 16389 19755 16455 19758
rect 6269 19682 6335 19685
rect 14641 19682 14707 19685
rect 6269 19680 14707 19682
rect 6269 19624 6274 19680
rect 6330 19624 14646 19680
rect 14702 19624 14707 19680
rect 6269 19622 14707 19624
rect 6269 19619 6335 19622
rect 14641 19619 14707 19622
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 27520 19592 28000 19712
rect 24277 19551 24597 19552
rect 8569 19546 8635 19549
rect 8569 19544 13830 19546
rect 8569 19488 8574 19544
rect 8630 19488 13830 19544
rect 8569 19486 13830 19488
rect 8569 19483 8635 19486
rect 13770 19410 13830 19486
rect 22277 19410 22343 19413
rect 13770 19408 22343 19410
rect 13770 19352 22282 19408
rect 22338 19352 22343 19408
rect 13770 19350 22343 19352
rect 22277 19347 22343 19350
rect 0 19184 480 19304
rect 62 18730 122 19184
rect 20713 19138 20779 19141
rect 23749 19138 23815 19141
rect 20713 19136 23815 19138
rect 20713 19080 20718 19136
rect 20774 19080 23754 19136
rect 23810 19080 23815 19136
rect 20713 19078 23815 19080
rect 20713 19075 20779 19078
rect 23749 19075 23815 19078
rect 24761 19138 24827 19141
rect 27662 19138 27722 19592
rect 24761 19136 27722 19138
rect 24761 19080 24766 19136
rect 24822 19080 27722 19136
rect 24761 19078 27722 19080
rect 24761 19075 24827 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 19374 18804 19380 18868
rect 19444 18866 19450 18868
rect 20253 18866 20319 18869
rect 19444 18864 20319 18866
rect 19444 18808 20258 18864
rect 20314 18808 20319 18864
rect 19444 18806 20319 18808
rect 19444 18804 19450 18806
rect 20253 18803 20319 18806
rect 1577 18730 1643 18733
rect 62 18728 1643 18730
rect 62 18672 1582 18728
rect 1638 18672 1643 18728
rect 62 18670 1643 18672
rect 1577 18667 1643 18670
rect 3233 18730 3299 18733
rect 10133 18730 10199 18733
rect 3233 18728 10199 18730
rect 3233 18672 3238 18728
rect 3294 18672 10138 18728
rect 10194 18672 10199 18728
rect 3233 18670 10199 18672
rect 3233 18667 3299 18670
rect 10133 18667 10199 18670
rect 6177 18594 6243 18597
rect 12985 18594 13051 18597
rect 14733 18594 14799 18597
rect 6177 18592 14799 18594
rect 6177 18536 6182 18592
rect 6238 18536 12990 18592
rect 13046 18536 14738 18592
rect 14794 18536 14799 18592
rect 6177 18534 14799 18536
rect 6177 18531 6243 18534
rect 12985 18531 13051 18534
rect 14733 18531 14799 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 27520 18368 28000 18488
rect 21541 18186 21607 18189
rect 25221 18186 25287 18189
rect 21541 18184 25287 18186
rect 21541 18128 21546 18184
rect 21602 18128 25226 18184
rect 25282 18128 25287 18184
rect 21541 18126 25287 18128
rect 21541 18123 21607 18126
rect 25221 18123 25287 18126
rect 10277 17984 10597 17985
rect 0 17824 480 17944
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 25405 17914 25471 17917
rect 27662 17914 27722 18368
rect 25405 17912 27722 17914
rect 25405 17856 25410 17912
rect 25466 17856 27722 17912
rect 25405 17854 27722 17856
rect 25405 17851 25471 17854
rect 62 17506 122 17824
rect 1577 17506 1643 17509
rect 62 17504 1643 17506
rect 62 17448 1582 17504
rect 1638 17448 1643 17504
rect 62 17446 1643 17448
rect 1577 17443 1643 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 7465 17234 7531 17237
rect 16389 17234 16455 17237
rect 7465 17232 16455 17234
rect 7465 17176 7470 17232
rect 7526 17176 16394 17232
rect 16450 17176 16455 17232
rect 7465 17174 16455 17176
rect 7465 17171 7531 17174
rect 16389 17171 16455 17174
rect 18505 17234 18571 17237
rect 18638 17234 18644 17236
rect 18505 17232 18644 17234
rect 18505 17176 18510 17232
rect 18566 17176 18644 17232
rect 18505 17174 18644 17176
rect 18505 17171 18571 17174
rect 18638 17172 18644 17174
rect 18708 17172 18714 17236
rect 9121 17098 9187 17101
rect 19241 17098 19307 17101
rect 9121 17096 19307 17098
rect 9121 17040 9126 17096
rect 9182 17040 19246 17096
rect 19302 17040 19307 17096
rect 9121 17038 19307 17040
rect 9121 17035 9187 17038
rect 19241 17035 19307 17038
rect 27520 17008 28000 17128
rect 54 16900 60 16964
rect 124 16962 130 16964
rect 1577 16962 1643 16965
rect 124 16960 1643 16962
rect 124 16904 1582 16960
rect 1638 16904 1643 16960
rect 124 16902 1643 16904
rect 124 16900 130 16902
rect 1577 16899 1643 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 7189 16690 7255 16693
rect 13721 16690 13787 16693
rect 7189 16688 13787 16690
rect 7189 16632 7194 16688
rect 7250 16632 13726 16688
rect 13782 16632 13787 16688
rect 7189 16630 13787 16632
rect 7189 16627 7255 16630
rect 13721 16627 13787 16630
rect 0 16556 480 16584
rect 0 16492 60 16556
rect 124 16492 480 16556
rect 0 16464 480 16492
rect 25589 16554 25655 16557
rect 27662 16554 27722 17008
rect 25589 16552 27722 16554
rect 25589 16496 25594 16552
rect 25650 16496 27722 16552
rect 25589 16494 27722 16496
rect 25589 16491 25655 16494
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 2037 16010 2103 16013
rect 10685 16010 10751 16013
rect 12433 16010 12499 16013
rect 2037 16008 12499 16010
rect 2037 15952 2042 16008
rect 2098 15952 10690 16008
rect 10746 15952 12438 16008
rect 12494 15952 12499 16008
rect 2037 15950 12499 15952
rect 2037 15947 2103 15950
rect 10685 15947 10751 15950
rect 12433 15947 12499 15950
rect 27520 15876 28000 15904
rect 27520 15812 27660 15876
rect 27724 15812 28000 15876
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 27520 15784 28000 15812
rect 19610 15743 19930 15744
rect 1301 15738 1367 15741
rect 62 15736 1367 15738
rect 62 15680 1306 15736
rect 1362 15680 1367 15736
rect 62 15678 1367 15680
rect 62 15224 122 15678
rect 1301 15675 1367 15678
rect 15510 15676 15516 15740
rect 15580 15738 15586 15740
rect 17217 15738 17283 15741
rect 15580 15736 17283 15738
rect 15580 15680 17222 15736
rect 17278 15680 17283 15736
rect 15580 15678 17283 15680
rect 15580 15676 15586 15678
rect 17217 15675 17283 15678
rect 19977 15602 20043 15605
rect 20294 15602 20300 15604
rect 19977 15600 20300 15602
rect 19977 15544 19982 15600
rect 20038 15544 20300 15600
rect 19977 15542 20300 15544
rect 19977 15539 20043 15542
rect 20294 15540 20300 15542
rect 20364 15540 20370 15604
rect 22645 15602 22711 15605
rect 27654 15602 27660 15604
rect 22645 15600 27660 15602
rect 22645 15544 22650 15600
rect 22706 15544 27660 15600
rect 22645 15542 27660 15544
rect 22645 15539 22711 15542
rect 27654 15540 27660 15542
rect 27724 15540 27730 15604
rect 16665 15466 16731 15469
rect 18454 15466 18460 15468
rect 16665 15464 18460 15466
rect 16665 15408 16670 15464
rect 16726 15408 18460 15464
rect 16665 15406 18460 15408
rect 16665 15403 16731 15406
rect 18454 15404 18460 15406
rect 18524 15404 18530 15468
rect 5610 15264 5930 15265
rect 0 15196 480 15224
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 0 15132 60 15196
rect 124 15132 480 15196
rect 0 15104 480 15132
rect 2313 15194 2379 15197
rect 3049 15194 3115 15197
rect 2313 15192 3115 15194
rect 2313 15136 2318 15192
rect 2374 15136 3054 15192
rect 3110 15136 3115 15192
rect 2313 15134 3115 15136
rect 2313 15131 2379 15134
rect 3049 15131 3115 15134
rect 7465 14922 7531 14925
rect 17677 14922 17743 14925
rect 7465 14920 17743 14922
rect 7465 14864 7470 14920
rect 7526 14864 17682 14920
rect 17738 14864 17743 14920
rect 7465 14862 17743 14864
rect 7465 14859 7531 14862
rect 17677 14859 17743 14862
rect 18505 14922 18571 14925
rect 25221 14922 25287 14925
rect 18505 14920 25287 14922
rect 18505 14864 18510 14920
rect 18566 14864 25226 14920
rect 25282 14864 25287 14920
rect 18505 14862 25287 14864
rect 18505 14859 18571 14862
rect 25221 14859 25287 14862
rect 4889 14786 4955 14789
rect 9254 14786 9260 14788
rect 4889 14784 9260 14786
rect 4889 14728 4894 14784
rect 4950 14728 9260 14784
rect 4889 14726 9260 14728
rect 4889 14723 4955 14726
rect 9254 14724 9260 14726
rect 9324 14724 9330 14788
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 27520 14648 28000 14680
rect 27520 14592 27710 14648
rect 27766 14592 28000 14648
rect 27520 14560 28000 14592
rect 3325 14514 3391 14517
rect 11697 14514 11763 14517
rect 3325 14512 11763 14514
rect 3325 14456 3330 14512
rect 3386 14456 11702 14512
rect 11758 14456 11763 14512
rect 3325 14454 11763 14456
rect 3325 14451 3391 14454
rect 11697 14451 11763 14454
rect 13261 14514 13327 14517
rect 25405 14514 25471 14517
rect 13261 14512 25471 14514
rect 13261 14456 13266 14512
rect 13322 14456 25410 14512
rect 25466 14456 25471 14512
rect 13261 14454 25471 14456
rect 13261 14451 13327 14454
rect 25405 14451 25471 14454
rect 19374 14378 19380 14380
rect 4110 14318 19380 14378
rect 0 13968 480 14000
rect 3233 13970 3299 13973
rect 0 13912 110 13968
rect 166 13912 480 13968
rect 0 13880 480 13912
rect 3190 13968 3299 13970
rect 3190 13912 3238 13968
rect 3294 13912 3299 13968
rect 3190 13907 3299 13912
rect 1577 13834 1643 13837
rect 3190 13834 3250 13907
rect 4110 13834 4170 14318
rect 19374 14316 19380 14318
rect 19444 14316 19450 14380
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 5349 13970 5415 13973
rect 7005 13970 7071 13973
rect 11053 13970 11119 13973
rect 15193 13970 15259 13973
rect 16849 13970 16915 13973
rect 5349 13968 7666 13970
rect 5349 13912 5354 13968
rect 5410 13912 7010 13968
rect 7066 13912 7666 13968
rect 5349 13910 7666 13912
rect 5349 13907 5415 13910
rect 7005 13907 7071 13910
rect 1577 13832 4170 13834
rect 1577 13776 1582 13832
rect 1638 13776 4170 13832
rect 1577 13774 4170 13776
rect 4521 13834 4587 13837
rect 7373 13834 7439 13837
rect 4521 13832 7439 13834
rect 4521 13776 4526 13832
rect 4582 13776 7378 13832
rect 7434 13776 7439 13832
rect 4521 13774 7439 13776
rect 7606 13834 7666 13910
rect 11053 13968 14980 13970
rect 11053 13912 11058 13968
rect 11114 13912 14980 13968
rect 11053 13910 14980 13912
rect 11053 13907 11119 13910
rect 14920 13837 14980 13910
rect 15193 13968 16915 13970
rect 15193 13912 15198 13968
rect 15254 13912 16854 13968
rect 16910 13912 16915 13968
rect 15193 13910 16915 13912
rect 15193 13907 15259 13910
rect 16849 13907 16915 13910
rect 14457 13834 14523 13837
rect 7606 13832 14523 13834
rect 7606 13776 14462 13832
rect 14518 13776 14523 13832
rect 7606 13774 14523 13776
rect 1577 13771 1643 13774
rect 4521 13771 4587 13774
rect 7373 13771 7439 13774
rect 14457 13771 14523 13774
rect 14917 13834 14983 13837
rect 17585 13834 17651 13837
rect 14917 13832 17651 13834
rect 14917 13776 14922 13832
rect 14978 13776 17590 13832
rect 17646 13776 17651 13832
rect 14917 13774 17651 13776
rect 14917 13771 14983 13774
rect 17585 13771 17651 13774
rect 5165 13698 5231 13701
rect 7741 13698 7807 13701
rect 5165 13696 7807 13698
rect 5165 13640 5170 13696
rect 5226 13640 7746 13696
rect 7802 13640 7807 13696
rect 5165 13638 7807 13640
rect 5165 13635 5231 13638
rect 7741 13635 7807 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 9029 13426 9095 13429
rect 14733 13426 14799 13429
rect 25221 13426 25287 13429
rect 25497 13426 25563 13429
rect 9029 13424 25563 13426
rect 9029 13368 9034 13424
rect 9090 13368 14738 13424
rect 14794 13368 25226 13424
rect 25282 13368 25502 13424
rect 25558 13368 25563 13424
rect 9029 13366 25563 13368
rect 9029 13363 9095 13366
rect 14733 13363 14799 13366
rect 25221 13363 25287 13366
rect 25497 13363 25563 13366
rect 54 13228 60 13292
rect 124 13290 130 13292
rect 10685 13290 10751 13293
rect 124 13288 10751 13290
rect 124 13232 10690 13288
rect 10746 13232 10751 13288
rect 124 13230 10751 13232
rect 124 13228 130 13230
rect 10685 13227 10751 13230
rect 27520 13288 28000 13320
rect 27520 13232 27618 13288
rect 27674 13232 28000 13288
rect 27520 13200 28000 13232
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 3877 12882 3943 12885
rect 12065 12882 12131 12885
rect 3877 12880 12131 12882
rect 3877 12824 3882 12880
rect 3938 12824 12070 12880
rect 12126 12824 12131 12880
rect 3877 12822 12131 12824
rect 3877 12819 3943 12822
rect 12065 12819 12131 12822
rect 2865 12746 2931 12749
rect 15101 12746 15167 12749
rect 2865 12744 15167 12746
rect 2865 12688 2870 12744
rect 2926 12688 15106 12744
rect 15162 12688 15167 12744
rect 2865 12686 15167 12688
rect 2865 12683 2931 12686
rect 15101 12683 15167 12686
rect 0 12612 480 12640
rect 0 12548 60 12612
rect 124 12548 480 12612
rect 0 12520 480 12548
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 54 12276 60 12340
rect 124 12338 130 12340
rect 5073 12338 5139 12341
rect 124 12336 5139 12338
rect 124 12280 5078 12336
rect 5134 12280 5139 12336
rect 124 12278 5139 12280
rect 124 12276 130 12278
rect 5073 12275 5139 12278
rect 3325 12202 3391 12205
rect 5349 12202 5415 12205
rect 3325 12200 5415 12202
rect 3325 12144 3330 12200
rect 3386 12144 5354 12200
rect 5410 12144 5415 12200
rect 3325 12142 5415 12144
rect 3325 12139 3391 12142
rect 5349 12139 5415 12142
rect 7649 12202 7715 12205
rect 13905 12202 13971 12205
rect 7649 12200 13971 12202
rect 7649 12144 7654 12200
rect 7710 12144 13910 12200
rect 13966 12144 13971 12200
rect 7649 12142 13971 12144
rect 7649 12139 7715 12142
rect 13905 12139 13971 12142
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 27520 11976 28000 12096
rect 24277 11935 24597 11936
rect 4797 11794 4863 11797
rect 22185 11794 22251 11797
rect 4797 11792 22251 11794
rect 4797 11736 4802 11792
rect 4858 11736 22190 11792
rect 22246 11736 22251 11792
rect 4797 11734 22251 11736
rect 4797 11731 4863 11734
rect 22185 11731 22251 11734
rect 25589 11522 25655 11525
rect 27662 11522 27722 11976
rect 25589 11520 27722 11522
rect 25589 11464 25594 11520
rect 25650 11464 27722 11520
rect 25589 11462 27722 11464
rect 25589 11459 25655 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 2773 11386 2839 11389
rect 6361 11386 6427 11389
rect 2773 11384 6427 11386
rect 2773 11328 2778 11384
rect 2834 11328 6366 11384
rect 6422 11328 6427 11384
rect 2773 11326 6427 11328
rect 2773 11323 2839 11326
rect 6361 11323 6427 11326
rect 0 11248 480 11280
rect 0 11192 110 11248
rect 166 11192 480 11248
rect 0 11160 480 11192
rect 4153 11250 4219 11253
rect 17861 11250 17927 11253
rect 4153 11248 17927 11250
rect 4153 11192 4158 11248
rect 4214 11192 17866 11248
rect 17922 11192 17927 11248
rect 4153 11190 17927 11192
rect 4153 11187 4219 11190
rect 17861 11187 17927 11190
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 17309 10706 17375 10709
rect 22829 10706 22895 10709
rect 17309 10704 22895 10706
rect 17309 10648 17314 10704
rect 17370 10648 22834 10704
rect 22890 10648 22895 10704
rect 17309 10646 22895 10648
rect 17309 10643 17375 10646
rect 22829 10643 22895 10646
rect 27520 10616 28000 10736
rect 54 10508 60 10572
rect 124 10570 130 10572
rect 9029 10570 9095 10573
rect 124 10568 9095 10570
rect 124 10512 9034 10568
rect 9090 10512 9095 10568
rect 124 10510 9095 10512
rect 124 10508 130 10510
rect 9029 10507 9095 10510
rect 12801 10570 12867 10573
rect 21817 10570 21883 10573
rect 12801 10568 21883 10570
rect 12801 10512 12806 10568
rect 12862 10512 21822 10568
rect 21878 10512 21883 10568
rect 12801 10510 21883 10512
rect 12801 10507 12867 10510
rect 21817 10507 21883 10510
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 9254 10236 9260 10300
rect 9324 10298 9330 10300
rect 10041 10298 10107 10301
rect 9324 10296 10107 10298
rect 9324 10240 10046 10296
rect 10102 10240 10107 10296
rect 9324 10238 10107 10240
rect 9324 10236 9330 10238
rect 10041 10235 10107 10238
rect 4613 10162 4679 10165
rect 21633 10162 21699 10165
rect 4613 10160 21699 10162
rect 4613 10104 4618 10160
rect 4674 10104 21638 10160
rect 21694 10104 21699 10160
rect 4613 10102 21699 10104
rect 4613 10099 4679 10102
rect 21633 10099 21699 10102
rect 25405 10162 25471 10165
rect 27662 10162 27722 10616
rect 25405 10160 27722 10162
rect 25405 10104 25410 10160
rect 25466 10104 27722 10160
rect 25405 10102 27722 10104
rect 25405 10099 25471 10102
rect 2129 10026 2195 10029
rect 5625 10026 5691 10029
rect 2129 10024 5691 10026
rect 2129 9968 2134 10024
rect 2190 9968 5630 10024
rect 5686 9968 5691 10024
rect 2129 9966 5691 9968
rect 2129 9963 2195 9966
rect 5625 9963 5691 9966
rect 0 9800 480 9920
rect 1761 9890 1827 9893
rect 2865 9890 2931 9893
rect 5349 9890 5415 9893
rect 1761 9888 5415 9890
rect 1761 9832 1766 9888
rect 1822 9832 2870 9888
rect 2926 9832 5354 9888
rect 5410 9832 5415 9888
rect 1761 9830 5415 9832
rect 1761 9827 1827 9830
rect 2865 9827 2931 9830
rect 5349 9827 5415 9830
rect 11881 9890 11947 9893
rect 14457 9890 14523 9893
rect 11881 9888 14523 9890
rect 11881 9832 11886 9888
rect 11942 9832 14462 9888
rect 14518 9832 14523 9888
rect 11881 9830 14523 9832
rect 11881 9827 11947 9830
rect 14457 9827 14523 9830
rect 5610 9824 5930 9825
rect 62 9346 122 9800
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 3417 9754 3483 9757
rect 3918 9754 3924 9756
rect 3417 9752 3924 9754
rect 3417 9696 3422 9752
rect 3478 9696 3924 9752
rect 3417 9694 3924 9696
rect 3417 9691 3483 9694
rect 3918 9692 3924 9694
rect 3988 9754 3994 9756
rect 4153 9754 4219 9757
rect 3988 9752 4219 9754
rect 3988 9696 4158 9752
rect 4214 9696 4219 9752
rect 3988 9694 4219 9696
rect 3988 9692 3994 9694
rect 4153 9691 4219 9694
rect 3693 9618 3759 9621
rect 4337 9618 4403 9621
rect 3693 9616 4403 9618
rect 3693 9560 3698 9616
rect 3754 9560 4342 9616
rect 4398 9560 4403 9616
rect 3693 9558 4403 9560
rect 3693 9555 3759 9558
rect 4337 9555 4403 9558
rect 3049 9482 3115 9485
rect 6729 9482 6795 9485
rect 3049 9480 6795 9482
rect 3049 9424 3054 9480
rect 3110 9424 6734 9480
rect 6790 9424 6795 9480
rect 3049 9422 6795 9424
rect 3049 9419 3115 9422
rect 6729 9419 6795 9422
rect 27520 9392 28000 9512
rect 3141 9346 3207 9349
rect 62 9344 3207 9346
rect 62 9288 3146 9344
rect 3202 9288 3207 9344
rect 62 9286 3207 9288
rect 3141 9283 3207 9286
rect 3601 9346 3667 9349
rect 4337 9346 4403 9349
rect 3601 9344 4403 9346
rect 3601 9288 3606 9344
rect 3662 9288 4342 9344
rect 4398 9288 4403 9344
rect 3601 9286 4403 9288
rect 3601 9283 3667 9286
rect 4337 9283 4403 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 3969 9074 4035 9077
rect 6453 9074 6519 9077
rect 3969 9072 6519 9074
rect 3969 9016 3974 9072
rect 4030 9016 6458 9072
rect 6514 9016 6519 9072
rect 3969 9014 6519 9016
rect 3969 9011 4035 9014
rect 6453 9011 6519 9014
rect 3918 8876 3924 8940
rect 3988 8938 3994 8940
rect 4337 8938 4403 8941
rect 3988 8936 4403 8938
rect 3988 8880 4342 8936
rect 4398 8880 4403 8936
rect 3988 8878 4403 8880
rect 3988 8876 3994 8878
rect 4337 8875 4403 8878
rect 25405 8938 25471 8941
rect 27662 8938 27722 9392
rect 25405 8936 27722 8938
rect 25405 8880 25410 8936
rect 25466 8880 27722 8936
rect 25405 8878 27722 8880
rect 25405 8875 25471 8878
rect 2589 8802 2655 8805
rect 4429 8802 4495 8805
rect 2589 8800 4495 8802
rect 2589 8744 2594 8800
rect 2650 8744 4434 8800
rect 4490 8744 4495 8800
rect 2589 8742 4495 8744
rect 2589 8739 2655 8742
rect 4429 8739 4495 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 15837 8666 15903 8669
rect 23381 8666 23447 8669
rect 15837 8664 23447 8666
rect 15837 8608 15842 8664
rect 15898 8608 23386 8664
rect 23442 8608 23447 8664
rect 15837 8606 23447 8608
rect 15837 8603 15903 8606
rect 23381 8603 23447 8606
rect 0 8440 480 8560
rect 21449 8530 21515 8533
rect 21449 8528 27722 8530
rect 21449 8472 21454 8528
rect 21510 8472 27722 8528
rect 21449 8470 27722 8472
rect 21449 8467 21515 8470
rect 62 7986 122 8440
rect 25037 8394 25103 8397
rect 13770 8392 25103 8394
rect 13770 8336 25042 8392
rect 25098 8336 25103 8392
rect 13770 8334 25103 8336
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 13770 8122 13830 8334
rect 25037 8331 25103 8334
rect 27662 8288 27722 8470
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 27520 8168 28000 8288
rect 19610 8127 19930 8128
rect 13540 8062 13830 8122
rect 1577 7986 1643 7989
rect 62 7984 1643 7986
rect 62 7928 1582 7984
rect 1638 7928 1643 7984
rect 62 7926 1643 7928
rect 1577 7923 1643 7926
rect 6637 7986 6703 7989
rect 11605 7986 11671 7989
rect 13540 7986 13600 8062
rect 6637 7984 13600 7986
rect 6637 7928 6642 7984
rect 6698 7928 11610 7984
rect 11666 7928 13600 7984
rect 6637 7926 13600 7928
rect 6637 7923 6703 7926
rect 11605 7923 11671 7926
rect 3325 7714 3391 7717
rect 3693 7714 3759 7717
rect 3325 7712 3759 7714
rect 3325 7656 3330 7712
rect 3386 7656 3698 7712
rect 3754 7656 3759 7712
rect 3325 7654 3759 7656
rect 3325 7651 3391 7654
rect 3693 7651 3759 7654
rect 17585 7714 17651 7717
rect 23657 7714 23723 7717
rect 17585 7712 23723 7714
rect 17585 7656 17590 7712
rect 17646 7656 23662 7712
rect 23718 7656 23723 7712
rect 17585 7654 23723 7656
rect 17585 7651 17651 7654
rect 23657 7651 23723 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 19374 7380 19380 7444
rect 19444 7442 19450 7444
rect 20345 7442 20411 7445
rect 19444 7440 27722 7442
rect 19444 7384 20350 7440
rect 20406 7384 27722 7440
rect 19444 7382 27722 7384
rect 19444 7380 19450 7382
rect 20345 7379 20411 7382
rect 0 7216 480 7336
rect 5349 7306 5415 7309
rect 21817 7306 21883 7309
rect 5349 7304 21883 7306
rect 5349 7248 5354 7304
rect 5410 7248 21822 7304
rect 21878 7248 21883 7304
rect 5349 7246 21883 7248
rect 5349 7243 5415 7246
rect 21817 7243 21883 7246
rect 62 6762 122 7216
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 27662 6928 27722 7382
rect 20161 6898 20227 6901
rect 20294 6898 20300 6900
rect 20161 6896 20300 6898
rect 20161 6840 20166 6896
rect 20222 6840 20300 6896
rect 20161 6838 20300 6840
rect 20161 6835 20227 6838
rect 20294 6836 20300 6838
rect 20364 6836 20370 6900
rect 27520 6808 28000 6928
rect 1577 6762 1643 6765
rect 62 6760 1643 6762
rect 62 6704 1582 6760
rect 1638 6704 1643 6760
rect 62 6702 1643 6704
rect 1577 6699 1643 6702
rect 15285 6762 15351 6765
rect 25129 6762 25195 6765
rect 15285 6760 25195 6762
rect 15285 6704 15290 6760
rect 15346 6704 25134 6760
rect 25190 6704 25195 6760
rect 15285 6702 25195 6704
rect 15285 6699 15351 6702
rect 25129 6699 25195 6702
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 14089 6354 14155 6357
rect 23933 6354 23999 6357
rect 14089 6352 23999 6354
rect 14089 6296 14094 6352
rect 14150 6296 23938 6352
rect 23994 6296 23999 6352
rect 14089 6294 23999 6296
rect 14089 6291 14155 6294
rect 23933 6291 23999 6294
rect 16573 6218 16639 6221
rect 24945 6218 25011 6221
rect 16573 6216 25011 6218
rect 16573 6160 16578 6216
rect 16634 6160 24950 6216
rect 25006 6160 25011 6216
rect 16573 6158 25011 6160
rect 16573 6155 16639 6158
rect 24945 6155 25011 6158
rect 10277 6016 10597 6017
rect 0 5948 480 5976
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 0 5884 60 5948
rect 124 5884 480 5948
rect 0 5856 480 5884
rect 62 5402 122 5856
rect 27520 5584 28000 5704
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 1945 5402 2011 5405
rect 62 5400 2011 5402
rect 62 5344 1950 5400
rect 2006 5344 2011 5400
rect 62 5342 2011 5344
rect 1945 5339 2011 5342
rect 3785 5402 3851 5405
rect 4613 5402 4679 5405
rect 3785 5400 4679 5402
rect 3785 5344 3790 5400
rect 3846 5344 4618 5400
rect 4674 5344 4679 5400
rect 3785 5342 4679 5344
rect 3785 5339 3851 5342
rect 4613 5339 4679 5342
rect 8017 5402 8083 5405
rect 14089 5402 14155 5405
rect 8017 5400 14155 5402
rect 8017 5344 8022 5400
rect 8078 5344 14094 5400
rect 14150 5344 14155 5400
rect 8017 5342 14155 5344
rect 8017 5339 8083 5342
rect 14089 5339 14155 5342
rect 11053 5130 11119 5133
rect 13629 5130 13695 5133
rect 23289 5130 23355 5133
rect 24577 5130 24643 5133
rect 11053 5128 24643 5130
rect 11053 5072 11058 5128
rect 11114 5072 13634 5128
rect 13690 5072 23294 5128
rect 23350 5072 24582 5128
rect 24638 5072 24643 5128
rect 11053 5070 24643 5072
rect 11053 5067 11119 5070
rect 13629 5067 13695 5070
rect 23289 5067 23355 5070
rect 24577 5067 24643 5070
rect 24761 5130 24827 5133
rect 27662 5130 27722 5584
rect 24761 5128 27722 5130
rect 24761 5072 24766 5128
rect 24822 5072 27722 5128
rect 24761 5070 27722 5072
rect 24761 5067 24827 5070
rect 15285 4994 15351 4997
rect 17309 4994 17375 4997
rect 15285 4992 17375 4994
rect 15285 4936 15290 4992
rect 15346 4936 17314 4992
rect 17370 4936 17375 4992
rect 15285 4934 17375 4936
rect 15285 4931 15351 4934
rect 17309 4931 17375 4934
rect 25405 4994 25471 4997
rect 25405 4992 27722 4994
rect 25405 4936 25410 4992
rect 25466 4936 27722 4992
rect 25405 4934 27722 4936
rect 25405 4931 25471 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 5533 4722 5599 4725
rect 21265 4722 21331 4725
rect 22001 4722 22067 4725
rect 5533 4720 22067 4722
rect 5533 4664 5538 4720
rect 5594 4664 21270 4720
rect 21326 4664 22006 4720
rect 22062 4664 22067 4720
rect 5533 4662 22067 4664
rect 5533 4659 5599 4662
rect 21265 4659 21331 4662
rect 22001 4659 22067 4662
rect 0 4496 480 4616
rect 62 4314 122 4496
rect 27662 4480 27722 4934
rect 18597 4450 18663 4453
rect 24025 4450 24091 4453
rect 18597 4448 24091 4450
rect 18597 4392 18602 4448
rect 18658 4392 24030 4448
rect 24086 4392 24091 4448
rect 18597 4390 24091 4392
rect 18597 4387 18663 4390
rect 24025 4387 24091 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 27520 4360 28000 4480
rect 24277 4319 24597 4320
rect 2589 4314 2655 4317
rect 62 4312 2655 4314
rect 62 4256 2594 4312
rect 2650 4256 2655 4312
rect 62 4254 2655 4256
rect 2589 4251 2655 4254
rect 12065 4314 12131 4317
rect 14733 4314 14799 4317
rect 12065 4312 14799 4314
rect 12065 4256 12070 4312
rect 12126 4256 14738 4312
rect 14794 4256 14799 4312
rect 12065 4254 14799 4256
rect 12065 4251 12131 4254
rect 14733 4251 14799 4254
rect 2773 4178 2839 4181
rect 18413 4178 18479 4181
rect 2773 4176 18479 4178
rect 2773 4120 2778 4176
rect 2834 4120 18418 4176
rect 18474 4120 18479 4176
rect 2773 4118 18479 4120
rect 2773 4115 2839 4118
rect 18413 4115 18479 4118
rect 16849 4042 16915 4045
rect 22737 4042 22803 4045
rect 4110 3982 13830 4042
rect 4110 3498 4170 3982
rect 13770 3906 13830 3982
rect 16849 4040 22803 4042
rect 16849 3984 16854 4040
rect 16910 3984 22742 4040
rect 22798 3984 22803 4040
rect 16849 3982 22803 3984
rect 16849 3979 16915 3982
rect 22737 3979 22803 3982
rect 18965 3906 19031 3909
rect 19425 3906 19491 3909
rect 13770 3904 19491 3906
rect 13770 3848 18970 3904
rect 19026 3848 19430 3904
rect 19486 3848 19491 3904
rect 13770 3846 19491 3848
rect 18965 3843 19031 3846
rect 19425 3843 19491 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 14457 3634 14523 3637
rect 22001 3634 22067 3637
rect 14457 3632 22067 3634
rect 14457 3576 14462 3632
rect 14518 3576 22006 3632
rect 22062 3576 22067 3632
rect 14457 3574 22067 3576
rect 14457 3571 14523 3574
rect 22001 3571 22067 3574
rect 62 3438 4170 3498
rect 62 3256 122 3438
rect 5610 3296 5930 3297
rect 0 3136 480 3256
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 3785 3226 3851 3229
rect 5441 3226 5507 3229
rect 3785 3224 5507 3226
rect 3785 3168 3790 3224
rect 3846 3168 5446 3224
rect 5502 3168 5507 3224
rect 3785 3166 5507 3168
rect 3785 3163 3851 3166
rect 5441 3163 5507 3166
rect 27520 3088 28000 3120
rect 27520 3032 27618 3088
rect 27674 3032 28000 3088
rect 27520 3000 28000 3032
rect 3969 2954 4035 2957
rect 11881 2954 11947 2957
rect 12985 2954 13051 2957
rect 3969 2952 13051 2954
rect 3969 2896 3974 2952
rect 4030 2896 11886 2952
rect 11942 2896 12990 2952
rect 13046 2896 13051 2952
rect 3969 2894 13051 2896
rect 3969 2891 4035 2894
rect 11881 2891 11947 2894
rect 12985 2891 13051 2894
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 1853 2410 1919 2413
rect 62 2408 1919 2410
rect 62 2352 1858 2408
rect 1914 2352 1919 2408
rect 62 2350 1919 2352
rect 62 1896 122 2350
rect 1853 2347 1919 2350
rect 6177 2410 6243 2413
rect 9029 2410 9095 2413
rect 6177 2408 9095 2410
rect 6177 2352 6182 2408
rect 6238 2352 9034 2408
rect 9090 2352 9095 2408
rect 6177 2350 9095 2352
rect 6177 2347 6243 2350
rect 9029 2347 9095 2350
rect 23105 2410 23171 2413
rect 23105 2408 27722 2410
rect 23105 2352 23110 2408
rect 23166 2352 27722 2408
rect 23105 2350 27722 2352
rect 23105 2347 23171 2350
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 6085 2138 6151 2141
rect 13813 2138 13879 2141
rect 14181 2138 14247 2141
rect 6085 2136 14247 2138
rect 6085 2080 6090 2136
rect 6146 2080 13818 2136
rect 13874 2080 14186 2136
rect 14242 2080 14247 2136
rect 6085 2078 14247 2080
rect 6085 2075 6151 2078
rect 13813 2075 13879 2078
rect 14181 2075 14247 2078
rect 12065 2002 12131 2005
rect 20989 2002 21055 2005
rect 12065 2000 21055 2002
rect 12065 1944 12070 2000
rect 12126 1944 20994 2000
rect 21050 1944 21055 2000
rect 12065 1942 21055 1944
rect 12065 1939 12131 1942
rect 20989 1939 21055 1942
rect 27662 1896 27722 2350
rect 0 1776 480 1896
rect 12433 1866 12499 1869
rect 22001 1866 22067 1869
rect 12433 1864 22067 1866
rect 12433 1808 12438 1864
rect 12494 1808 22006 1864
rect 22062 1808 22067 1864
rect 12433 1806 22067 1808
rect 12433 1803 12499 1806
rect 22001 1803 22067 1806
rect 27520 1776 28000 1896
rect 2497 1730 2563 1733
rect 27061 1730 27127 1733
rect 2497 1728 27127 1730
rect 2497 1672 2502 1728
rect 2558 1672 27066 1728
rect 27122 1672 27127 1728
rect 2497 1670 27127 1672
rect 2497 1667 2563 1670
rect 27061 1667 27127 1670
rect 6361 1186 6427 1189
rect 62 1184 6427 1186
rect 62 1128 6366 1184
rect 6422 1128 6427 1184
rect 62 1126 6427 1128
rect 62 672 122 1126
rect 6361 1123 6427 1126
rect 0 552 480 672
rect 27520 552 28000 672
rect 9305 98 9371 101
rect 27662 98 27722 552
rect 9305 96 27722 98
rect 9305 40 9310 96
rect 9366 40 27722 96
rect 9305 38 27722 40
rect 9305 35 9371 38
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 18644 23428 18708 23492
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 15516 22068 15580 22132
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 18460 21388 18524 21452
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 19380 18804 19444 18868
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 18644 17172 18708 17236
rect 60 16900 124 16964
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 60 16492 124 16556
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 27660 15812 27724 15876
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 15516 15676 15580 15740
rect 20300 15540 20364 15604
rect 27660 15540 27724 15604
rect 18460 15404 18524 15468
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 60 15132 124 15196
rect 9260 14724 9324 14788
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 19380 14316 19444 14380
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 60 13228 124 13292
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 60 12548 124 12612
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 60 12276 124 12340
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 60 10508 124 10572
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 9260 10236 9324 10300
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 3924 9692 3988 9756
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 3924 8876 3988 8940
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 19380 7380 19444 7444
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 20300 6836 20364 6900
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 60 5884 124 5948
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 59 16964 125 16965
rect 59 16900 60 16964
rect 124 16900 125 16964
rect 59 16899 125 16900
rect 62 16557 122 16899
rect 59 16556 125 16557
rect 59 16492 60 16556
rect 124 16492 125 16556
rect 59 16491 125 16492
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 59 15196 125 15197
rect 59 15132 60 15196
rect 124 15132 125 15196
rect 59 15131 125 15132
rect 62 13293 122 15131
rect 5610 14176 5931 15200
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 9259 14788 9325 14789
rect 9259 14724 9260 14788
rect 9324 14724 9325 14788
rect 9259 14723 9325 14724
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 59 13292 125 13293
rect 59 13228 60 13292
rect 124 13228 125 13292
rect 59 13227 125 13228
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 59 12612 125 12613
rect 59 12548 60 12612
rect 124 12548 125 12612
rect 59 12547 125 12548
rect 62 12341 122 12547
rect 59 12340 125 12341
rect 59 12276 60 12340
rect 124 12276 125 12340
rect 59 12275 125 12276
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 59 10572 125 10573
rect 59 10508 60 10572
rect 124 10508 125 10572
rect 59 10507 125 10508
rect 62 5949 122 10507
rect 5610 9824 5931 10848
rect 9262 10301 9322 14723
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 9259 10300 9325 10301
rect 9259 10236 9260 10300
rect 9324 10236 9325 10300
rect 9259 10235 9325 10236
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 3923 9756 3989 9757
rect 3923 9692 3924 9756
rect 3988 9692 3989 9756
rect 3923 9691 3989 9692
rect 3926 8941 3986 9691
rect 3923 8940 3989 8941
rect 3923 8876 3924 8940
rect 3988 8876 3989 8940
rect 3923 8875 3989 8876
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 59 5948 125 5949
rect 59 5884 60 5948
rect 124 5884 125 5948
rect 59 5883 125 5884
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 18643 23492 18709 23493
rect 18643 23428 18644 23492
rect 18708 23428 18709 23492
rect 18643 23427 18709 23428
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 15515 22132 15581 22133
rect 15515 22068 15516 22132
rect 15580 22068 15581 22132
rect 15515 22067 15581 22068
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 15518 15741 15578 22067
rect 18459 21452 18525 21453
rect 18459 21388 18460 21452
rect 18524 21388 18525 21452
rect 18459 21387 18525 21388
rect 15515 15740 15581 15741
rect 15515 15676 15516 15740
rect 15580 15676 15581 15740
rect 15515 15675 15581 15676
rect 18462 15469 18522 21387
rect 18646 17237 18706 23427
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19379 18868 19445 18869
rect 19379 18804 19380 18868
rect 19444 18804 19445 18868
rect 19379 18803 19445 18804
rect 18643 17236 18709 17237
rect 18643 17172 18644 17236
rect 18708 17172 18709 17236
rect 18643 17171 18709 17172
rect 18459 15468 18525 15469
rect 18459 15404 18460 15468
rect 18524 15404 18525 15468
rect 18459 15403 18525 15404
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 19382 14381 19442 18803
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 20299 15604 20365 15605
rect 20299 15540 20300 15604
rect 20364 15540 20365 15604
rect 20299 15539 20365 15540
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19379 14380 19445 14381
rect 19379 14316 19380 14380
rect 19444 14316 19445 14380
rect 19379 14315 19445 14316
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 19382 7445 19442 14315
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19379 7444 19445 7445
rect 19379 7380 19380 7444
rect 19444 7380 19445 7444
rect 19379 7379 19445 7380
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 20302 6901 20362 15539
rect 24277 15264 24597 16288
rect 27659 15876 27725 15877
rect 27659 15812 27660 15876
rect 27724 15812 27725 15876
rect 27659 15811 27725 15812
rect 27662 15605 27722 15811
rect 27659 15604 27725 15605
rect 27659 15540 27660 15604
rect 27724 15540 27725 15604
rect 27659 15539 27725 15540
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 20299 6900 20365 6901
rect 20299 6836 20300 6900
rect 20364 6836 20365 6900
rect 20299 6835 20365 6836
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_inv_1  mux_right_track_0.INVTX1_3_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__209__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_12 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_11
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_16 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2576 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_16
timestamp 1586364061
transform 1 0 2576 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 222 592
use scs8hd_conb_1  _249_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_22
timestamp 1586364061
transform 1 0 3128 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3312 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_31
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 4232 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4324 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_38
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_36
timestamp 1586364061
transform 1 0 4416 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_1  _110_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4784 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_43
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_47
timestamp 1586364061
transform 1 0 5428 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_6  FILLER_1_42
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _260_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use scs8hd_nor2_4  _114_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _258_
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__260__A
timestamp 1586364061
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_67
timestamp 1586364061
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_71
timestamp 1586364061
transform 1 0 7636 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_71
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_75
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _214_
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__258__A
timestamp 1586364061
transform 1 0 8556 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__214__A
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__214__B
timestamp 1586364061
transform 1 0 9016 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_79
timestamp 1586364061
transform 1 0 8372 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_83
timestamp 1586364061
transform 1 0 8740 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_0_88
timestamp 1586364061
transform 1 0 9200 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_79
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_83 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8740 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__213__B
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_99
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_95
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_97
timestamp 1586364061
transform 1 0 10028 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__213__A
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_101
timestamp 1586364061
transform 1 0 10396 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12880 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12696 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13248 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13892 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_130
timestamp 1586364061
transform 1 0 13064 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_137
timestamp 1586364061
transform 1 0 13708 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_141
timestamp 1586364061
transform 1 0 14076 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _268_
timestamp 1586364061
transform 1 0 14444 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__268__A
timestamp 1586364061
transform 1 0 14996 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_143
timestamp 1586364061
transform 1 0 14260 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_147 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_149
timestamp 1586364061
transform 1 0 14812 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_153
timestamp 1586364061
transform 1 0 15180 0 1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_162
timestamp 1586364061
transform 1 0 16008 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_158
timestamp 1586364061
transform 1 0 15640 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17204 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17572 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_173
timestamp 1586364061
transform 1 0 17020 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_177
timestamp 1586364061
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_169
timestamp 1586364061
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_173
timestamp 1586364061
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_177
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_181
timestamp 1586364061
transform 1 0 17756 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_188
timestamp 1586364061
transform 1 0 18400 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__265__A
timestamp 1586364061
transform 1 0 18768 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_buf_2  _265_
timestamp 1586364061
transform 1 0 18952 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _273_
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_198
timestamp 1586364061
transform 1 0 19320 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_202
timestamp 1586364061
transform 1 0 19688 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_210
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__273__A
timestamp 1586364061
transform 1 0 20424 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _270_
timestamp 1586364061
transform 1 0 20056 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_214
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_212
timestamp 1586364061
transform 1 0 20608 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__270__A
timestamp 1586364061
transform 1 0 20608 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20976 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 774 592
use scs8hd_buf_2  _286_
timestamp 1586364061
transform 1 0 22080 0 -1 2720
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21896 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_226
timestamp 1586364061
transform 1 0 21896 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_221
timestamp 1586364061
transform 1 0 21436 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_225
timestamp 1586364061
transform 1 0 21804 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_228
timestamp 1586364061
transform 1 0 22080 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22908 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__286__A
timestamp 1586364061
transform 1 0 22632 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_232
timestamp 1586364061
transform 1 0 22448 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_236 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 22816 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_239
timestamp 1586364061
transform 1 0 23092 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_243
timestamp 1586364061
transform 1 0 23460 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_248
timestamp 1586364061
transform 1 0 23920 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_252
timestamp 1586364061
transform 1 0 24288 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _280_
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_6  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__280__A
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 25116 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25484 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_259
timestamp 1586364061
transform 1 0 24932 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_263
timestamp 1586364061
transform 1 0 25300 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_259
timestamp 1586364061
transform 1 0 24932 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_263
timestamp 1586364061
transform 1 0 25300 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_267
timestamp 1586364061
transform 1 0 25668 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_275
timestamp 1586364061
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_275
timestamp 1586364061
transform 1 0 26404 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _209_
timestamp 1586364061
transform 1 0 1932 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_6  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_8  FILLER_2_12
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 774 592
use scs8hd_buf_1  _104_
timestamp 1586364061
transform 1 0 2944 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 774 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_41
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_45
timestamp 1586364061
transform 1 0 5244 0 -1 3808
box -38 -48 774 592
use scs8hd_nor2_4  _108_
timestamp 1586364061
transform 1 0 6164 0 -1 3808
box -38 -48 866 592
use scs8hd_fill_2  FILLER_2_53
timestamp 1586364061
transform 1 0 5980 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_64
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7544 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_72
timestamp 1586364061
transform 1 0 7728 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_83
timestamp 1586364061
transform 1 0 8740 0 -1 3808
box -38 -48 774 592
use scs8hd_nor2_4  _213_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_91
timestamp 1586364061
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_106
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_121
timestamp 1586364061
transform 1 0 12236 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_128
timestamp 1586364061
transform 1 0 12880 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_4  FILLER_2_138
timestamp 1586364061
transform 1 0 13800 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_142
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15456 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_167
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_171
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_2_179
timestamp 1586364061
transform 1 0 17572 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17756 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_8  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19320 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19872 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_201
timestamp 1586364061
transform 1 0 19596 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_206
timestamp 1586364061
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_210
timestamp 1586364061
transform 1 0 20424 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_218
timestamp 1586364061
transform 1 0 21160 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21896 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22356 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_229
timestamp 1586364061
transform 1 0 22172 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22908 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_2_233
timestamp 1586364061
transform 1 0 22540 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_240
timestamp 1586364061
transform 1 0 23184 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23920 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 774 592
use scs8hd_buf_1  _154_
timestamp 1586364061
transform 1 0 24932 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_262
timestamp 1586364061
transform 1 0 25208 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_274
timestamp 1586364061
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2116 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use scs8hd_buf_1  _107_
timestamp 1586364061
transform 1 0 3128 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_14
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_18
timestamp 1586364061
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_25
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4140 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_29
timestamp 1586364061
transform 1 0 3772 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5336 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_44
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_48
timestamp 1586364061
transform 1 0 5520 0 1 3808
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6992 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_54
timestamp 1586364061
transform 1 0 6072 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_75
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__212__A
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__212__B
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_92
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_97
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_101
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_139
timestamp 1586364061
transform 1 0 13892 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_152
timestamp 1586364061
transform 1 0 15088 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_169
timestamp 1586364061
transform 1 0 16652 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_174
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_178
timestamp 1586364061
transform 1 0 17480 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19872 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 19320 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19688 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_200
timestamp 1586364061
transform 1 0 19504 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_213
timestamp 1586364061
transform 1 0 20700 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_217
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21436 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21896 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22264 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_224
timestamp 1586364061
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_228
timestamp 1586364061
transform 1 0 22080 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22908 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23276 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_235
timestamp 1586364061
transform 1 0 22724 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_239
timestamp 1586364061
transform 1 0 23092 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_243
timestamp 1586364061
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__257__A
timestamp 1586364061
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_248
timestamp 1586364061
transform 1 0 23920 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_252
timestamp 1586364061
transform 1 0 24288 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_259
timestamp 1586364061
transform 1 0 24932 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_263
timestamp 1586364061
transform 1 0 25300 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_275
timestamp 1586364061
transform 1 0 26404 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1932 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__256__A
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_12
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_16
timestamp 1586364061
transform 1 0 2576 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_36
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_4  FILLER_4_48
timestamp 1586364061
transform 1 0 5520 0 -1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_54
timestamp 1586364061
transform 1 0 6072 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_62
timestamp 1586364061
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_75
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_79
timestamp 1586364061
transform 1 0 8372 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_6  FILLER_4_85
timestamp 1586364061
transform 1 0 8924 0 -1 4896
box -38 -48 590 592
use scs8hd_nor2_4  _212_
timestamp 1586364061
transform 1 0 9844 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_91
timestamp 1586364061
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11408 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_104
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_108
timestamp 1586364061
transform 1 0 11040 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_123
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_127
timestamp 1586364061
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_131
timestamp 1586364061
transform 1 0 13156 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_142
timestamp 1586364061
transform 1 0 14168 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_146
timestamp 1586364061
transform 1 0 14536 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_152
timestamp 1586364061
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15548 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 17296 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_168
timestamp 1586364061
transform 1 0 16560 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_172
timestamp 1586364061
transform 1 0 16928 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_187
timestamp 1586364061
transform 1 0 18308 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_191
timestamp 1586364061
transform 1 0 18676 0 -1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 4896
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22264 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_224
timestamp 1586364061
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_228
timestamp 1586364061
transform 1 0 22080 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22816 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_4  FILLER_4_232
timestamp 1586364061
transform 1 0 22448 0 -1 4896
box -38 -48 406 592
use scs8hd_buf_2  _257_
timestamp 1586364061
transform 1 0 24564 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 24012 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24380 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_245
timestamp 1586364061
transform 1 0 23644 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_259
timestamp 1586364061
transform 1 0 24932 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_271
timestamp 1586364061
transform 1 0 26036 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_buf_2  _259_
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__259__A
timestamp 1586364061
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_11
timestamp 1586364061
transform 1 0 2116 0 1 4896
box -38 -48 314 592
use scs8hd_nor2_4  _102_
timestamp 1586364061
transform 1 0 3128 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_16
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 4140 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_31
timestamp 1586364061
transform 1 0 3956 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_35
timestamp 1586364061
transform 1 0 4324 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 866 592
use scs8hd_decap_4  FILLER_5_48
timestamp 1586364061
transform 1 0 5520 0 1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5888 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_54
timestamp 1586364061
transform 1 0 6072 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_58
timestamp 1586364061
transform 1 0 6440 0 1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7728 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_66
timestamp 1586364061
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_70
timestamp 1586364061
transform 1 0 7544 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_83
timestamp 1586364061
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_87
timestamp 1586364061
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9476 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_100
timestamp 1586364061
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _132_
timestamp 1586364061
transform 1 0 11040 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 10856 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_104
timestamp 1586364061
transform 1 0 10672 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_111
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_115
timestamp 1586364061
transform 1 0 11684 0 1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_134
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_138
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_151
timestamp 1586364061
transform 1 0 14996 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_156
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_160
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_173
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18400 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 18216 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_191
timestamp 1586364061
transform 1 0 18676 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19504 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19320 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_195
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 20700 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_211
timestamp 1586364061
transform 1 0 20516 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_215
timestamp 1586364061
transform 1 0 20884 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21252 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_221
timestamp 1586364061
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_conb_1  _248_
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_5_265
timestamp 1586364061
transform 1 0 25484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_6
timestamp 1586364061
transform 1 0 1656 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_6_6
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_10
timestamp 1586364061
transform 1 0 2024 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_10
timestamp 1586364061
transform 1 0 2024 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2116 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _138_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_13
timestamp 1586364061
transform 1 0 2300 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_13
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_23
timestamp 1586364061
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_31
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4140 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4324 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5336 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5704 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_48
timestamp 1586364061
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_46
timestamp 1586364061
transform 1 0 5336 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_50
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_61
timestamp 1586364061
transform 1 0 6716 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6992 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_66
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_71
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_79
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _215_
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__210__A
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__210__B
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_92
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_96
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_99
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__215__A
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_108
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 11776 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_127
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_134
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_145
timestamp 1586364061
transform 1 0 14444 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_144
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_149
timestamp 1586364061
transform 1 0 14812 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_6_148
timestamp 1586364061
transform 1 0 14720 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_152
timestamp 1586364061
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 15456 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_166
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _171_
timestamp 1586364061
transform 1 0 17388 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_169
timestamp 1586364061
transform 1 0 16652 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_170
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_174
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_178
timestamp 1586364061
transform 1 0 17480 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_181
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_186
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18124 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_192
timestamp 1586364061
transform 1 0 18768 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_188
timestamp 1586364061
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18584 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 590 592
use scs8hd_nor2_4  _168_
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 19136 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 18952 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_205
timestamp 1586364061
transform 1 0 19964 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_205
timestamp 1586364061
transform 1 0 19964 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_209
timestamp 1586364061
transform 1 0 20332 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_209
timestamp 1586364061
transform 1 0 20332 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20148 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20148 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_213
timestamp 1586364061
transform 1 0 20700 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_213
timestamp 1586364061
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20516 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_217
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 314 592
use scs8hd_nor2_4  _167_
timestamp 1586364061
transform 1 0 21528 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_6_.latch
timestamp 1586364061
transform 1 0 22264 0 -1 5984
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21252 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_222
timestamp 1586364061
transform 1 0 21528 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_226
timestamp 1586364061
transform 1 0 21896 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_231
timestamp 1586364061
transform 1 0 22356 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 22632 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_241
timestamp 1586364061
transform 1 0 23276 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 24012 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 23644 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_247
timestamp 1586364061
transform 1 0 23828 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_254
timestamp 1586364061
transform 1 0 24472 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25024 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_258
timestamp 1586364061
transform 1 0 24840 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_258
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_265
timestamp 1586364061
transform 1 0 25484 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_270
timestamp 1586364061
transform 1 0 25944 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_274
timestamp 1586364061
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 2116 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 1564 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_7
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 3312 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_22
timestamp 1586364061
transform 1 0 3128 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 4232 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 4600 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 3680 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_26
timestamp 1586364061
transform 1 0 3496 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_30
timestamp 1586364061
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_36
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4968 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_2  FILLER_8_40
timestamp 1586364061
transform 1 0 4784 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_51
timestamp 1586364061
transform 1 0 5796 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 6532 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 6348 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__C
timestamp 1586364061
transform 1 0 5980 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_55
timestamp 1586364061
transform 1 0 6164 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_1  _128_
timestamp 1586364061
transform 1 0 8096 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 7912 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_72
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__C
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 8924 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_79
timestamp 1586364061
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_83
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_87
timestamp 1586364061
transform 1 0 9108 0 -1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _210_
timestamp 1586364061
transform 1 0 10028 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_91
timestamp 1586364061
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 11592 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__215__B
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__226__B
timestamp 1586364061
transform 1 0 11408 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_106
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_110
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_123
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_127
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_140
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 774 592
use scs8hd_nor2_4  _170_
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__173__B
timestamp 1586364061
transform 1 0 14904 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_148
timestamp 1586364061
transform 1 0 14720 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_152
timestamp 1586364061
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_163
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 17572 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_175
timestamp 1586364061
transform 1 0 17204 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18768 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19504 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 19136 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_194
timestamp 1586364061
transform 1 0 18952 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_198
timestamp 1586364061
transform 1 0 19320 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_203
timestamp 1586364061
transform 1 0 19780 0 -1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_207
timestamp 1586364061
transform 1 0 20148 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_210
timestamp 1586364061
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_226
timestamp 1586364061
transform 1 0 21896 0 -1 7072
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 22632 0 -1 7072
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24380 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 23828 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_245
timestamp 1586364061
transform 1 0 23644 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_249
timestamp 1586364061
transform 1 0 24012 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_262
timestamp 1586364061
transform 1 0 25208 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_274
timestamp 1586364061
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_2  _256_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_11
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 314 592
use scs8hd_nor2_4  _099_
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_25
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_29
timestamp 1586364061
transform 1 0 3772 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _098_
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_42
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_46
timestamp 1586364061
transform 1 0 5336 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 6440 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_60
timestamp 1586364061
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use scs8hd_buf_1  _126_
timestamp 1586364061
transform 1 0 7268 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 7084 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_70
timestamp 1586364061
transform 1 0 7544 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_77
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use scs8hd_or3_4  _109_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8280 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_87
timestamp 1586364061
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__211__A
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_91
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_95
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_101
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _211_
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12604 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__211__B
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_127
timestamp 1586364061
transform 1 0 12788 0 1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _173_
timestamp 1586364061
transform 1 0 14904 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 14720 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_142
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_146
timestamp 1586364061
transform 1 0 14536 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 15916 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 16284 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_163
timestamp 1586364061
transform 1 0 16100 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16652 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17480 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_167
timestamp 1586364061
transform 1 0 16468 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_172
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_176
timestamp 1586364061
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_180
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_197
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_201
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_205
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20424 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _166_
timestamp 1586364061
transform 1 0 21988 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_219
timestamp 1586364061
transform 1 0 21252 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_223
timestamp 1586364061
transform 1 0 21620 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_236
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_240
timestamp 1586364061
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _155_
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_254
timestamp 1586364061
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_265
timestamp 1586364061
transform 1 0 25484 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_buf_1  _091_
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_6
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_10
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__208__D
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__C
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_43
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_47
timestamp 1586364061
transform 1 0 5428 0 -1 8160
box -38 -48 314 592
use scs8hd_or3_4  _106_
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_52
timestamp 1586364061
transform 1 0 5888 0 -1 8160
box -38 -48 406 592
use scs8hd_or3_4  _115_
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__C
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_67
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_71
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__228__B
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 406 592
use scs8hd_buf_1  _113_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_90
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_96
timestamp 1586364061
transform 1 0 9936 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _226_
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_114
timestamp 1586364061
transform 1 0 11592 0 -1 8160
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 12328 0 -1 8160
box -38 -48 1050 592
use scs8hd_buf_1  _116_
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13524 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13892 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_133
timestamp 1586364061
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_137
timestamp 1586364061
transform 1 0 13708 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _172_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_144
timestamp 1586364061
transform 1 0 14352 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_150
timestamp 1586364061
transform 1 0 14904 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 17388 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_167
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18768 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_188
timestamp 1586364061
transform 1 0 18400 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 -1 8160
box -38 -48 866 592
use scs8hd_fill_2  FILLER_10_194
timestamp 1586364061
transform 1 0 18952 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_205
timestamp 1586364061
transform 1 0 19964 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_209
timestamp 1586364061
transform 1 0 20332 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_224
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_10_229
timestamp 1586364061
transform 1 0 22172 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_7_.latch
timestamp 1586364061
transform 1 0 22724 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22540 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24472 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23920 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24288 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_246
timestamp 1586364061
transform 1 0 23736 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_250
timestamp 1586364061
transform 1 0 24104 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_257
timestamp 1586364061
transform 1 0 24748 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_10_269
timestamp 1586364061
transform 1 0 25852 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_8  _090_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_12
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _255_
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__093__D
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_16
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_24
timestamp 1586364061
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__255__A
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__208__B
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_28
timestamp 1586364061
transform 1 0 3680 0 1 8160
box -38 -48 314 592
use scs8hd_buf_1  _130_
timestamp 1586364061
transform 1 0 5704 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__208__C
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_42
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_46
timestamp 1586364061
transform 1 0 5336 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _083_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__C
timestamp 1586364061
transform 1 0 6440 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_60
timestamp 1586364061
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_77
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _228_
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_81
timestamp 1586364061
transform 1 0 8556 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_85
timestamp 1586364061
transform 1 0 8924 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_97
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_101
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_134
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 866 592
use scs8hd_decap_4  FILLER_11_151
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_155
timestamp 1586364061
transform 1 0 15364 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_158
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_173
timestamp 1586364061
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_177
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_181
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19688 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_194
timestamp 1586364061
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_198
timestamp 1586364061
transform 1 0 19320 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_211
timestamp 1586364061
transform 1 0 20516 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_216
timestamp 1586364061
transform 1 0 20976 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_11_231
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22540 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_235
timestamp 1586364061
transform 1 0 22724 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_240
timestamp 1586364061
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_254
timestamp 1586364061
transform 1 0 24472 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _267_
timestamp 1586364061
transform 1 0 25208 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__267__A
timestamp 1586364061
transform 1 0 25760 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_258
timestamp 1586364061
transform 1 0 24840 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_266
timestamp 1586364061
transform 1 0 25576 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_11_270
timestamp 1586364061
transform 1 0 25944 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_276
timestamp 1586364061
transform 1 0 26496 0 1 8160
box -38 -48 130 592
use scs8hd_buf_1  _094_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 2116 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_10
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 130 592
use scs8hd_or3_4  _085_
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_12_13
timestamp 1586364061
transform 1 0 2300 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 406 592
use scs8hd_or4_4  _208_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 3680 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_30
timestamp 1586364061
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 5428 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__D
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_41
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_45
timestamp 1586364061
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_49
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use scs8hd_or3_4  _103_
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__207__B
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_53
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 314 592
use scs8hd_or3_4  _112_
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 7452 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_67
timestamp 1586364061
transform 1 0 7268 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_71
timestamp 1586364061
transform 1 0 7636 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use scs8hd_buf_1  _136_
timestamp 1586364061
transform 1 0 9844 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10304 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_98
timestamp 1586364061
transform 1 0 10120 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12696 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_121
timestamp 1586364061
transform 1 0 12236 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_137
timestamp 1586364061
transform 1 0 13708 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_144
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_148
timestamp 1586364061
transform 1 0 14720 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_152
timestamp 1586364061
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _160_
timestamp 1586364061
transform 1 0 15456 0 -1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_12_165
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17020 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_169
timestamp 1586364061
transform 1 0 16652 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18768 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_184
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_188
timestamp 1586364061
transform 1 0 18400 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_203
timestamp 1586364061
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21068 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_207
timestamp 1586364061
transform 1 0 20148 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_211
timestamp 1586364061
transform 1 0 20516 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21436 0 -1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_12_219
timestamp 1586364061
transform 1 0 21252 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_230
timestamp 1586364061
transform 1 0 22264 0 -1 9248
box -38 -48 406 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 23000 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__178__B
timestamp 1586364061
transform 1 0 22724 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_234
timestamp 1586364061
transform 1 0 22632 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_237
timestamp 1586364061
transform 1 0 22908 0 -1 9248
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 24012 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_247
timestamp 1586364061
transform 1 0 23828 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_258
timestamp 1586364061
transform 1 0 24840 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_270
timestamp 1586364061
transform 1 0 25944 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_274
timestamp 1586364061
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_buf_1  _119_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_10
timestamp 1586364061
transform 1 0 2024 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__C
timestamp 1586364061
transform 1 0 2116 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_or4_4  _093_
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 866 592
use scs8hd_inv_8  _084_
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__C
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_20
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_24
timestamp 1586364061
transform 1 0 3312 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_13
timestamp 1586364061
transform 1 0 2300 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_or4_4  _163_
timestamp 1586364061
transform 1 0 3680 0 1 9248
box -38 -48 866 592
use scs8hd_or4_4  _197_
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__224__B
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_37
timestamp 1586364061
transform 1 0 4508 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_41
timestamp 1586364061
transform 1 0 4876 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__C
timestamp 1586364061
transform 1 0 5060 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__B
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_48
timestamp 1586364061
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_45
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 222 592
use scs8hd_buf_2  _254_
timestamp 1586364061
transform 1 0 5244 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_49
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 5704 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__254__A
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _206_
timestamp 1586364061
transform 1 0 6348 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _207_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__224__D
timestamp 1586364061
transform 1 0 6072 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_52
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 130 592
use scs8hd_or3_4  _097_
timestamp 1586364061
transform 1 0 7912 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__097__C
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__B
timestamp 1586364061
transform 1 0 7728 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_76
timestamp 1586364061
transform 1 0 8096 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_66
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_70
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 222 592
use scs8hd_or3_4  _100_
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 8924 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__C
timestamp 1586364061
transform 1 0 9292 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_88
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_83
timestamp 1586364061
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_87
timestamp 1586364061
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_91
timestamp 1586364061
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_96
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_92
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__229__B
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 9384 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_97
timestamp 1586364061
transform 1 0 10028 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_100
timestamp 1586364061
transform 1 0 10304 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _229_
timestamp 1586364061
transform 1 0 10120 0 -1 10336
box -38 -48 866 592
use scs8hd_buf_1  _134_
timestamp 1586364061
transform 1 0 11684 0 -1 10336
box -38 -48 314 592
use scs8hd_nor2_4  _227_
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__227__B
timestamp 1586364061
transform 1 0 11132 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11500 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_107
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_111
timestamp 1586364061
transform 1 0 11316 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_118
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_127
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_123
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13892 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_134
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_138
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_137
timestamp 1586364061
transform 1 0 13708 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_151
timestamp 1586364061
transform 1 0 14996 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_159
timestamp 1586364061
transform 1 0 15732 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_158
timestamp 1586364061
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_155
timestamp 1586364061
transform 1 0 15364 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15456 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_165
timestamp 1586364061
transform 1 0 16284 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_162
timestamp 1586364061
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 16376 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16468 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_6  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 590 592
use scs8hd_decap_8  FILLER_14_176
timestamp 1586364061
transform 1 0 17296 0 -1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_184
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_197
timestamp 1586364061
transform 1 0 19228 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_195
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_201
timestamp 1586364061
transform 1 0 19596 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_199
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19780 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__B
timestamp 1586364061
transform 1 0 19780 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 19412 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_205
timestamp 1586364061
transform 1 0 19964 0 -1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19964 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__180__B
timestamp 1586364061
transform 1 0 20976 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_214
timestamp 1586364061
transform 1 0 20792 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_218
timestamp 1586364061
transform 1 0 21160 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_nor2_4  _180_
timestamp 1586364061
transform 1 0 21528 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_231
timestamp 1586364061
transform 1 0 22356 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 774 592
use scs8hd_nor2_4  _178_
timestamp 1586364061
transform 1 0 22724 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 22724 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_237
timestamp 1586364061
transform 1 0 22908 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_241
timestamp 1586364061
transform 1 0 23276 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_232
timestamp 1586364061
transform 1 0 22448 0 -1 10336
box -38 -48 314 592
use scs8hd_nor2_4  _146_
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _177_
timestamp 1586364061
transform 1 0 24288 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 23736 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24104 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_254
timestamp 1586364061
transform 1 0 24472 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_244
timestamp 1586364061
transform 1 0 23552 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_248
timestamp 1586364061
transform 1 0 23920 0 -1 10336
box -38 -48 222 592
use scs8hd_buf_2  _264_
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__264__A
timestamp 1586364061
transform 1 0 25760 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_258
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_266
timestamp 1586364061
transform 1 0 25576 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_261
timestamp 1586364061
transform 1 0 25116 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_13_270
timestamp 1586364061
transform 1 0 25944 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_276
timestamp 1586364061
transform 1 0 26496 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_273
timestamp 1586364061
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_8  _082_
timestamp 1586364061
transform 1 0 2208 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 2024 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_21
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_25
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use scs8hd_or4_4  _224_
timestamp 1586364061
transform 1 0 3772 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__224__A
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_38
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_or2_4  _092_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5336 0 1 10336
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_42
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7084 0 1 10336
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_15_76
timestamp 1586364061
transform 1 0 8096 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8832 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_81
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_93
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_99
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_139
timestamp 1586364061
transform 1 0 13892 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  FILLER_15_152
timestamp 1586364061
transform 1 0 15088 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 16100 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_157
timestamp 1586364061
transform 1 0 15548 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17296 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_174
timestamp 1586364061
transform 1 0 17112 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_178
timestamp 1586364061
transform 1 0 17480 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18124 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18584 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_188
timestamp 1586364061
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_192
timestamp 1586364061
transform 1 0 18768 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _179_
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 18952 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_205
timestamp 1586364061
transform 1 0 19964 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 20700 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20516 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 20148 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_209
timestamp 1586364061
transform 1 0 20332 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 21896 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22264 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_224
timestamp 1586364061
transform 1 0 21712 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_228
timestamp 1586364061
transform 1 0 22080 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22908 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_235
timestamp 1586364061
transform 1 0 22724 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_239
timestamp 1586364061
transform 1 0 23092 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_7_.latch
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_256
timestamp 1586364061
transform 1 0 24656 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _263_
timestamp 1586364061
transform 1 0 25392 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25208 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24840 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_260
timestamp 1586364061
transform 1 0 25024 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_268
timestamp 1586364061
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__263__A
timestamp 1586364061
transform 1 0 25944 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_272
timestamp 1586364061
transform 1 0 26128 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_276
timestamp 1586364061
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use scs8hd_buf_1  _089_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__C
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_10
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _231_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__186__C
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_or4_4  _174_
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__224__C
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_1  _088_
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__D
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_41
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_45
timestamp 1586364061
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6624 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__204__B
timestamp 1586364061
transform 1 0 6072 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__231__B
timestamp 1586364061
transform 1 0 6440 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_52
timestamp 1586364061
transform 1 0 5888 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_71
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_75
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_1  _101_
timestamp 1586364061
transform 1 0 8372 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_82
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_86
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_90
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__230__B
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_107
timestamp 1586364061
transform 1 0 10948 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_121
timestamp 1586364061
transform 1 0 12236 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_127
timestamp 1586364061
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_138
timestamp 1586364061
transform 1 0 13800 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__184__B
timestamp 1586364061
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_142
timestamp 1586364061
transform 1 0 14168 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_4  FILLER_16_148
timestamp 1586364061
transform 1 0 14720 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_152
timestamp 1586364061
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_158
timestamp 1586364061
transform 1 0 15640 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_162
timestamp 1586364061
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_165
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_175
timestamp 1586364061
transform 1 0 17204 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_179
timestamp 1586364061
transform 1 0 17572 0 -1 11424
box -38 -48 406 592
use scs8hd_buf_1  _140_
timestamp 1586364061
transform 1 0 17940 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__182__B
timestamp 1586364061
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_191
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20332 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_211
timestamp 1586364061
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_218
timestamp 1586364061
transform 1 0 21160 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 21896 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21344 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_222
timestamp 1586364061
transform 1 0 21528 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_237
timestamp 1586364061
transform 1 0 22908 0 -1 11424
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_6_.latch
timestamp 1586364061
transform 1 0 23644 0 -1 11424
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_16_256
timestamp 1586364061
transform 1 0 24656 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_260
timestamp 1586364061
transform 1 0 25024 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_267
timestamp 1586364061
transform 1 0 25668 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_or4_4  _120_
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 2024 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__D
timestamp 1586364061
transform 1 0 1656 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_8
timestamp 1586364061
transform 1 0 1840 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__216__B
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_21
timestamp 1586364061
transform 1 0 3036 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_25
timestamp 1586364061
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use scs8hd_or4_4  _216_
timestamp 1586364061
transform 1 0 3772 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__216__A
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_38
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use scs8hd_or2_4  _185_
timestamp 1586364061
transform 1 0 5336 0 1 11424
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__B
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_42
timestamp 1586364061
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_67
timestamp 1586364061
transform 1 0 7268 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9200 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_80
timestamp 1586364061
transform 1 0 8464 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_84
timestamp 1586364061
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_97
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_101
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _230_
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__195__B
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_134
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_138
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _184_
timestamp 1586364061
transform 1 0 14536 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_142
timestamp 1586364061
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_155
timestamp 1586364061
transform 1 0 15364 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_162
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__B
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_172
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_177
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _182_
timestamp 1586364061
transform 1 0 18492 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 18308 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_181
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19504 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_198
timestamp 1586364061
transform 1 0 19320 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_202
timestamp 1586364061
transform 1 0 19688 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20332 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20148 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_206
timestamp 1586364061
transform 1 0 20056 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_218
timestamp 1586364061
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21896 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_222
timestamp 1586364061
transform 1 0 21528 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22908 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23276 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_235
timestamp 1586364061
transform 1 0 22724 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_239
timestamp 1586364061
transform 1 0 23092 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_243
timestamp 1586364061
transform 1 0 23460 0 1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24380 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24196 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23828 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_249
timestamp 1586364061
transform 1 0 24012 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25392 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_262
timestamp 1586364061
transform 1 0 25208 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_266
timestamp 1586364061
transform 1 0 25576 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_274
timestamp 1586364061
transform 1 0 26312 0 1 11424
box -38 -48 314 592
use scs8hd_inv_8  _118_
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__232__C
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_8
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_21
timestamp 1586364061
transform 1 0 3036 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_25
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 406 592
use scs8hd_or4_4  _186_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__216__C
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__B
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__D
timestamp 1586364061
transform 1 0 5704 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_41
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_45
timestamp 1586364061
transform 1 0 5244 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_48
timestamp 1586364061
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _204_
timestamp 1586364061
transform 1 0 5980 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_52
timestamp 1586364061
transform 1 0 5888 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_62
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7636 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_66
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_82
timestamp 1586364061
transform 1 0 8648 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_86
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _195_
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_106
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_119
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__B
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_136
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_140
timestamp 1586364061
transform 1 0 13984 0 -1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_143
timestamp 1586364061
transform 1 0 14260 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_147
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 590 592
use scs8hd_decap_4  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15824 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15640 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _183_
timestamp 1586364061
transform 1 0 17572 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_171
timestamp 1586364061
transform 1 0 16836 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_175
timestamp 1586364061
transform 1 0 17204 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_188
timestamp 1586364061
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_192
timestamp 1586364061
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18952 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_196
timestamp 1586364061
transform 1 0 19136 0 -1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_218
timestamp 1586364061
transform 1 0 21160 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22264 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21344 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_222
timestamp 1586364061
transform 1 0 21528 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_228
timestamp 1586364061
transform 1 0 22080 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24472 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24288 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_nand2_4  _151_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 -1 13600
box -38 -48 866 592
use scs8hd_or4_4  _232_
timestamp 1586364061
transform 1 0 1656 0 1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__232__B
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_8
timestamp 1586364061
transform 1 0 1840 0 -1 13600
box -38 -48 130 592
use scs8hd_nor2_4  _201_
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 2944 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__D
timestamp 1586364061
transform 1 0 3312 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_19
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_18
timestamp 1586364061
transform 1 0 2760 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_22
timestamp 1586364061
transform 1 0 3128 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _200_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__216__D
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__201__B
timestamp 1586364061
transform 1 0 3680 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_32
timestamp 1586364061
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_36
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_26
timestamp 1586364061
transform 1 0 3496 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_30
timestamp 1586364061
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use scs8hd_nor2_4  _202_
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__203__B
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__B
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_41
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_46
timestamp 1586364061
transform 1 0 5336 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_51
timestamp 1586364061
transform 1 0 5796 0 -1 13600
box -38 -48 406 592
use scs8hd_buf_1  _124_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6348 0 -1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_69
timestamp 1586364061
transform 1 0 7452 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_65
timestamp 1586364061
transform 1 0 7084 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7544 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_72
timestamp 1586364061
transform 1 0 7728 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_72
timestamp 1586364061
transform 1 0 7728 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7912 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _086_
timestamp 1586364061
transform 1 0 8096 0 -1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 8096 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_87
timestamp 1586364061
transform 1 0 9108 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_79
timestamp 1586364061
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_83
timestamp 1586364061
transform 1 0 8740 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_91
timestamp 1586364061
transform 1 0 9476 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_104
timestamp 1586364061
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_108
timestamp 1586364061
transform 1 0 11040 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_112
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_115
timestamp 1586364061
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_119
timestamp 1586364061
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_116
timestamp 1586364061
transform 1 0 11776 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_128
timestamp 1586364061
transform 1 0 12880 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _181_
timestamp 1586364061
transform 1 0 14076 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 13892 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_137
timestamp 1586364061
transform 1 0 13708 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_132
timestamp 1586364061
transform 1 0 13248 0 -1 13600
box -38 -48 222 592
use scs8hd_buf_1  _121_
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_150
timestamp 1586364061
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_154
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15732 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_157
timestamp 1586364061
transform 1 0 15548 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_161
timestamp 1586364061
transform 1 0 15916 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_165
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16652 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_169
timestamp 1586364061
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_173
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_177
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_178
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 18768 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18216 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_188
timestamp 1586364061
transform 1 0 18400 0 1 12512
box -38 -48 406 592
use scs8hd_buf_1  _141_
timestamp 1586364061
transform 1 0 19780 0 -1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18952 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_205
timestamp 1586364061
transform 1 0 19964 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_195
timestamp 1586364061
transform 1 0 19044 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20700 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20516 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_209
timestamp 1586364061
transform 1 0 20332 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22264 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 21712 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_222
timestamp 1586364061
transform 1 0 21528 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_226
timestamp 1586364061
transform 1 0 21896 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_226
timestamp 1586364061
transform 1 0 21896 0 -1 13600
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 23460 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22724 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 22448 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_233
timestamp 1586364061
transform 1 0 22540 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_237
timestamp 1586364061
transform 1 0 22908 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_241
timestamp 1586364061
transform 1 0 23276 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_234
timestamp 1586364061
transform 1 0 22632 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_242
timestamp 1586364061
transform 1 0 23368 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24288 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 23828 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_249
timestamp 1586364061
transform 1 0 24012 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_254
timestamp 1586364061
transform 1 0 24472 0 -1 13600
box -38 -48 222 592
use scs8hd_buf_2  _285_
timestamp 1586364061
transform 1 0 25208 0 -1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__285__A
timestamp 1586364061
transform 1 0 25300 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_261
timestamp 1586364061
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_265
timestamp 1586364061
transform 1 0 25484 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_20_258
timestamp 1586364061
transform 1 0 24840 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_266
timestamp 1586364061
transform 1 0 25576 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_274
timestamp 1586364061
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_6_.latch
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 1050 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 1564 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_18
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_22
timestamp 1586364061
transform 1 0 3128 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_7_.latch
timestamp 1586364061
transform 1 0 3496 0 1 13600
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_21_37
timestamp 1586364061
transform 1 0 4508 0 1 13600
box -38 -48 222 592
use scs8hd_buf_1  _087_
timestamp 1586364061
transform 1 0 5244 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 5704 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__200__B
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_41
timestamp 1586364061
transform 1 0 4876 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_48
timestamp 1586364061
transform 1 0 5520 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 6072 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_52
timestamp 1586364061
transform 1 0 5888 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_56
timestamp 1586364061
transform 1 0 6256 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_73
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_77
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9936 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_90
timestamp 1586364061
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_94
timestamp 1586364061
transform 1 0 9752 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_107
timestamp 1586364061
transform 1 0 10948 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_111
timestamp 1586364061
transform 1 0 11316 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_134
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_138
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_151
timestamp 1586364061
transform 1 0 14996 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_156
timestamp 1586364061
transform 1 0 15456 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_160
timestamp 1586364061
transform 1 0 15824 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 17480 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_172
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_176
timestamp 1586364061
transform 1 0 17296 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18584 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_180
timestamp 1586364061
transform 1 0 17664 0 1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19780 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_201
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_205
timestamp 1586364061
transform 1 0 19964 0 1 13600
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20700 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20332 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_211
timestamp 1586364061
transform 1 0 20516 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 22264 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_224
timestamp 1586364061
transform 1 0 21712 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_228
timestamp 1586364061
transform 1 0 22080 0 1 13600
box -38 -48 222 592
use scs8hd_buf_1  _175_
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 22908 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_235
timestamp 1586364061
transform 1 0 22724 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_239
timestamp 1586364061
transform 1 0 23092 0 1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_256
timestamp 1586364061
transform 1 0 24656 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24840 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_260
timestamp 1586364061
transform 1 0 25024 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_267
timestamp 1586364061
transform 1 0 25668 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_6  FILLER_21_271
timestamp 1586364061
transform 1 0 26036 0 1 13600
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__225__A
timestamp 1586364061
transform 1 0 2944 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_17
timestamp 1586364061
transform 1 0 2668 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_22_22
timestamp 1586364061
transform 1 0 3128 0 -1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__205__B
timestamp 1586364061
transform 1 0 3496 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_28
timestamp 1586364061
transform 1 0 3680 0 -1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _203_
timestamp 1586364061
transform 1 0 5612 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__189__B
timestamp 1586364061
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5428 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_41
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_45
timestamp 1586364061
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_58
timestamp 1586364061
transform 1 0 6440 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_64
timestamp 1586364061
transform 1 0 6992 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_78
timestamp 1586364061
transform 1 0 8280 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_82
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_86
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_102
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11592 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__196__B
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_107
timestamp 1586364061
transform 1 0 10948 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_113
timestamp 1586364061
transform 1 0 11500 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_123
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 -1 14688
box -38 -48 866 592
use scs8hd_fill_2  FILLER_22_140
timestamp 1586364061
transform 1 0 13984 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_144
timestamp 1586364061
transform 1 0 14352 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_148
timestamp 1586364061
transform 1 0 14720 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_152
timestamp 1586364061
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _137_
timestamp 1586364061
transform 1 0 16836 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_180
timestamp 1586364061
transform 1 0 17664 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_188
timestamp 1586364061
transform 1 0 18400 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_192
timestamp 1586364061
transform 1 0 18768 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18952 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_196
timestamp 1586364061
transform 1 0 19136 0 -1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_206
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_212
timestamp 1586364061
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22356 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_224
timestamp 1586364061
transform 1 0 21712 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_229
timestamp 1586364061
transform 1 0 22172 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 22540 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  FILLER_22_242
timestamp 1586364061
transform 1 0 23368 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23644 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_247
timestamp 1586364061
transform 1 0 23828 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_259
timestamp 1586364061
transform 1 0 24932 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_271
timestamp 1586364061
transform 1 0 26036 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_or4_4  _139_
timestamp 1586364061
transform 1 0 1932 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_18
timestamp 1586364061
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_22
timestamp 1586364061
transform 1 0 3128 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _205_
timestamp 1586364061
transform 1 0 3496 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_35
timestamp 1586364061
transform 1 0 4324 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _189_
timestamp 1586364061
transform 1 0 5060 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 4876 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 6072 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_52
timestamp 1586364061
transform 1 0 5888 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_56
timestamp 1586364061
transform 1 0 6256 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_71
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_75
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_91
timestamp 1586364061
transform 1 0 9476 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_95
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_23_98
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_102
timestamp 1586364061
transform 1 0 10488 0 1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _196_
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_126
timestamp 1586364061
transform 1 0 12696 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_130
timestamp 1586364061
transform 1 0 13064 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 15088 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_145
timestamp 1586364061
transform 1 0 14444 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_150
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_154
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 15640 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 17296 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_167
timestamp 1586364061
transform 1 0 16468 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_23_178
timestamp 1586364061
transform 1 0 17480 0 1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 18584 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 18400 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19596 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_199
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_203
timestamp 1586364061
transform 1 0 19780 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20424 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_207
timestamp 1586364061
transform 1 0 20148 0 1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_219
timestamp 1586364061
transform 1 0 21252 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_223
timestamp 1586364061
transform 1 0 21620 0 1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_23_226
timestamp 1586364061
transform 1 0 21896 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_236
timestamp 1586364061
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_240
timestamp 1586364061
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24472 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 23828 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24288 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_249
timestamp 1586364061
transform 1 0 24012 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25484 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_263
timestamp 1586364061
transform 1 0 25300 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_267
timestamp 1586364061
transform 1 0 25668 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_275
timestamp 1586364061
transform 1 0 26404 0 1 14688
box -38 -48 222 592
use scs8hd_inv_8  _150_
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_12
timestamp 1586364061
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_1  _225_
timestamp 1586364061
transform 1 0 2944 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__139__D
timestamp 1586364061
transform 1 0 2392 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__C
timestamp 1586364061
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_16
timestamp 1586364061
transform 1 0 2576 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4324 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_29
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_38
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 5336 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__190__B
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__217__A
timestamp 1586364061
transform 1 0 4784 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_42
timestamp 1586364061
transform 1 0 4968 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__192__B
timestamp 1586364061
transform 1 0 6900 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_57
timestamp 1586364061
transform 1 0 6348 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_61
timestamp 1586364061
transform 1 0 6716 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 7084 0 -1 15776
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_24_76
timestamp 1586364061
transform 1 0 8096 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__B
timestamp 1586364061
transform 1 0 8280 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8648 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9936 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 11684 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11500 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_107
timestamp 1586364061
transform 1 0 10948 0 -1 15776
box -38 -48 590 592
use scs8hd_decap_6  FILLER_24_126
timestamp 1586364061
transform 1 0 12696 0 -1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_143
timestamp 1586364061
transform 1 0 14260 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_147
timestamp 1586364061
transform 1 0 14628 0 -1 15776
box -38 -48 590 592
use scs8hd_decap_4  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 15732 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_1  FILLER_24_158
timestamp 1586364061
transform 1 0 15640 0 -1 15776
box -38 -48 130 592
use scs8hd_buf_1  _122_
timestamp 1586364061
transform 1 0 17296 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16744 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_168
timestamp 1586364061
transform 1 0 16560 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_172
timestamp 1586364061
transform 1 0 16928 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_3  FILLER_24_179
timestamp 1586364061
transform 1 0 17572 0 -1 15776
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18492 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17848 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_184
timestamp 1586364061
transform 1 0 18032 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_188
timestamp 1586364061
transform 1 0 18400 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_200
timestamp 1586364061
transform 1 0 19504 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_204
timestamp 1586364061
transform 1 0 19872 0 -1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21160 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_212
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 21712 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21528 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_220
timestamp 1586364061
transform 1 0 21344 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_235
timestamp 1586364061
transform 1 0 22724 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_243
timestamp 1586364061
transform 1 0 23460 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_6_.latch
timestamp 1586364061
transform 1 0 23644 0 -1 15776
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_24_256
timestamp 1586364061
transform 1 0 24656 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24840 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_260
timestamp 1586364061
transform 1 0 25024 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_24_267
timestamp 1586364061
transform 1 0 25668 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_buf_2  _262_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__262__A
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_11
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__276__A
timestamp 1586364061
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_19
timestamp 1586364061
transform 1 0 2852 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_23
timestamp 1586364061
transform 1 0 3220 0 1 15776
box -38 -48 222 592
use scs8hd_or4_4  _152_
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__152__C
timestamp 1586364061
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_36
timestamp 1586364061
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _190_
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_40
timestamp 1586364061
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _192_
timestamp 1586364061
transform 1 0 6900 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_72
timestamp 1586364061
transform 1 0 7728 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_76
timestamp 1586364061
transform 1 0 8096 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 8464 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8280 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _222_
timestamp 1586364061
transform 1 0 10488 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__222__A
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__222__B
timestamp 1586364061
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_91
timestamp 1586364061
transform 1 0 9476 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_95
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_111
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_115
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_119
timestamp 1586364061
transform 1 0 12052 0 1 15776
box -38 -48 130 592
use scs8hd_nor2_4  _194_
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__194__B
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_132
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_136
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_149
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_153
timestamp 1586364061
transform 1 0 15180 0 1 15776
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_158
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_173
timestamp 1586364061
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_177
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 406 592
use scs8hd_buf_1  _176_
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 18492 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_187
timestamp 1586364061
transform 1 0 18308 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_191
timestamp 1586364061
transform 1 0 18676 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 19412 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_195
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_210
timestamp 1586364061
transform 1 0 20424 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_214
timestamp 1586364061
transform 1 0 20792 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_217
timestamp 1586364061
transform 1 0 21068 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22172 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_227
timestamp 1586364061
transform 1 0 21988 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_231
timestamp 1586364061
transform 1 0 22356 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 22632 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_236
timestamp 1586364061
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_240
timestamp 1586364061
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_7_.latch
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_256
timestamp 1586364061
transform 1 0 24656 0 1 15776
box -38 -48 222 592
use scs8hd_buf_2  _278_
timestamp 1586364061
transform 1 0 25392 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24840 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25208 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_260
timestamp 1586364061
transform 1 0 25024 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_268
timestamp 1586364061
transform 1 0 25760 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__278__A
timestamp 1586364061
transform 1 0 25944 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_272
timestamp 1586364061
transform 1 0 26128 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_276
timestamp 1586364061
transform 1 0 26496 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_2  _276_
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use scs8hd_buf_2  _272_
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_11
timestamp 1586364061
transform 1 0 2116 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_7
timestamp 1586364061
transform 1 0 1748 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1932 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__272__A
timestamp 1586364061
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_11
timestamp 1586364061
transform 1 0 2116 0 1 16864
box -38 -48 774 592
use scs8hd_buf_1  _188_
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__238__B
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2300 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_19
timestamp 1586364061
transform 1 0 2852 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_24
timestamp 1586364061
transform 1 0 3312 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_28
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_29
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_buf_1  _199_
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_35
timestamp 1586364061
transform 1 0 4324 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_36
timestamp 1586364061
transform 1 0 4416 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__152__D
timestamp 1586364061
transform 1 0 4232 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 4508 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  _217_
timestamp 1586364061
transform 1 0 4692 0 -1 16864
box -38 -48 314 592
use scs8hd_nor2_4  _235_
timestamp 1586364061
transform 1 0 5060 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5704 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 4876 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__235__B
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_42
timestamp 1586364061
transform 1 0 4968 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_46
timestamp 1586364061
transform 1 0 5336 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6072 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 6992 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6440 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_59
timestamp 1586364061
transform 1 0 6532 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_52
timestamp 1586364061
transform 1 0 5888 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_56
timestamp 1586364061
transform 1 0 6256 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_60
timestamp 1586364061
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _191_
timestamp 1586364061
transform 1 0 7176 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _193_
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__191__B
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7544 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_65
timestamp 1586364061
transform 1 0 7084 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_72
timestamp 1586364061
transform 1 0 7728 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_75
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_79
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__219__B
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__218__B
timestamp 1586364061
transform 1 0 9844 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_92
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_97
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_101
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _219_
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11500 0 -1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__218__A
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__219__A
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_107
timestamp 1586364061
transform 1 0 10948 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_124
timestamp 1586364061
transform 1 0 12512 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_126
timestamp 1586364061
transform 1 0 12696 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_128
timestamp 1586364061
transform 1 0 12880 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12696 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_130
timestamp 1586364061
transform 1 0 13064 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14536 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_143
timestamp 1586364061
transform 1 0 14260 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_151
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_144
timestamp 1586364061
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_148
timestamp 1586364061
transform 1 0 14720 0 1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_27_154
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16192 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_162
timestamp 1586364061
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_158
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_162
timestamp 1586364061
transform 1 0 16008 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_174
timestamp 1586364061
transform 1 0 17112 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_175
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17848 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_191
timestamp 1586364061
transform 1 0 18676 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_187
timestamp 1586364061
transform 1 0 18308 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_191
timestamp 1586364061
transform 1 0 18676 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 19044 0 1 16864
box -38 -48 1050 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 19044 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19872 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_197
timestamp 1586364061
transform 1 0 19228 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20792 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 20608 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_206
timestamp 1586364061
transform 1 0 20056 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_206
timestamp 1586364061
transform 1 0 20056 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_210
timestamp 1586364061
transform 1 0 20424 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 22356 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_224
timestamp 1586364061
transform 1 0 21712 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_223
timestamp 1586364061
transform 1 0 21620 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_227
timestamp 1586364061
transform 1 0 21988 0 1 16864
box -38 -48 406 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 22632 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_232
timestamp 1586364061
transform 1 0 22448 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_243
timestamp 1586364061
transform 1 0 23460 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_236
timestamp 1586364061
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_240
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 23644 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24012 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__261__A
timestamp 1586364061
transform 1 0 24656 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_247
timestamp 1586364061
transform 1 0 23828 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_254
timestamp 1586364061
transform 1 0 24472 0 1 16864
box -38 -48 222 592
use scs8hd_buf_2  _277_
timestamp 1586364061
transform 1 0 25208 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__277__A
timestamp 1586364061
transform 1 0 25760 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_260
timestamp 1586364061
transform 1 0 25024 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_258
timestamp 1586364061
transform 1 0 24840 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_266
timestamp 1586364061
transform 1 0 25576 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_26_272
timestamp 1586364061
transform 1 0 26128 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_27_270
timestamp 1586364061
transform 1 0 25944 0 1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_27_276
timestamp 1586364061
transform 1 0 26496 0 1 16864
box -38 -48 130 592
use scs8hd_conb_1  _245_
timestamp 1586364061
transform 1 0 1932 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__287__A
timestamp 1586364061
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_7
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_12
timestamp 1586364061
transform 1 0 2208 0 -1 17952
box -38 -48 774 592
use scs8hd_buf_1  _187_
timestamp 1586364061
transform 1 0 2944 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__239__B
timestamp 1586364061
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _238_
timestamp 1586364061
transform 1 0 4232 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 5796 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__234__B
timestamp 1586364061
transform 1 0 5244 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_43
timestamp 1586364061
transform 1 0 5060 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_47
timestamp 1586364061
transform 1 0 5428 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_6  FILLER_28_62
timestamp 1586364061
transform 1 0 6808 0 -1 17952
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7544 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_81
timestamp 1586364061
transform 1 0 8556 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_85
timestamp 1586364061
transform 1 0 8924 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_89
timestamp 1586364061
transform 1 0 9292 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_97
timestamp 1586364061
transform 1 0 10028 0 -1 17952
box -38 -48 590 592
use scs8hd_nor2_4  _218_
timestamp 1586364061
transform 1 0 10580 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_112
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12144 0 -1 17952
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13892 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13708 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_131
timestamp 1586364061
transform 1 0 13156 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_135
timestamp 1586364061
transform 1 0 13524 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_142
timestamp 1586364061
transform 1 0 14168 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_146
timestamp 1586364061
transform 1 0 14536 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_152
timestamp 1586364061
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15640 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_161
timestamp 1586364061
transform 1 0 15916 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_165
timestamp 1586364061
transform 1 0 16284 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16652 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_182
timestamp 1586364061
transform 1 0 17848 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18860 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_206
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_210
timestamp 1586364061
transform 1 0 20424 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_224
timestamp 1586364061
transform 1 0 21712 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_228
timestamp 1586364061
transform 1 0 22080 0 -1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 22724 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22540 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_232
timestamp 1586364061
transform 1 0 22448 0 -1 17952
box -38 -48 130 592
use scs8hd_buf_2  _261_
timestamp 1586364061
transform 1 0 24564 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_8  FILLER_28_244
timestamp 1586364061
transform 1 0 23552 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_28_252
timestamp 1586364061
transform 1 0 24288 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_259
timestamp 1586364061
transform 1 0 24932 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_271
timestamp 1586364061
transform 1 0 26036 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_buf_2  _271_
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__271__A
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_11
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _239_
timestamp 1586364061
transform 1 0 3220 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 2576 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_18
timestamp 1586364061
transform 1 0 2760 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_22
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_32
timestamp 1586364061
transform 1 0 4048 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_38
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _234_
timestamp 1586364061
transform 1 0 4784 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_49
timestamp 1586364061
transform 1 0 5612 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 406 592
use scs8hd_decap_4  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7360 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7176 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9108 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_79
timestamp 1586364061
transform 1 0 8372 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_83
timestamp 1586364061
transform 1 0 8740 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_96
timestamp 1586364061
transform 1 0 9936 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_100
timestamp 1586364061
transform 1 0 10304 0 1 17952
box -38 -48 314 592
use scs8hd_nor2_4  _220_
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__220__A
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_134
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_138
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 866 592
use scs8hd_decap_4  FILLER_29_151
timestamp 1586364061
transform 1 0 14996 0 1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 16008 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 15824 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_155
timestamp 1586364061
transform 1 0 15364 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_158
timestamp 1586364061
transform 1 0 15640 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17480 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_173
timestamp 1586364061
transform 1 0 17020 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_177
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_180
timestamp 1586364061
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_187
timestamp 1586364061
transform 1 0 18308 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_191
timestamp 1586364061
transform 1 0 18676 0 1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19504 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_197
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 20516 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_209
timestamp 1586364061
transform 1 0 20332 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_213
timestamp 1586364061
transform 1 0 20700 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 22080 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_226
timestamp 1586364061
transform 1 0 21896 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_230
timestamp 1586364061
transform 1 0 22264 0 1 17952
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_238
timestamp 1586364061
transform 1 0 23000 0 1 17952
box -38 -48 590 592
use scs8hd_buf_2  _274_
timestamp 1586364061
transform 1 0 24564 0 1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24380 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__274__A
timestamp 1586364061
transform 1 0 24012 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_251
timestamp 1586364061
transform 1 0 24196 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_259
timestamp 1586364061
transform 1 0 24932 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_263
timestamp 1586364061
transform 1 0 25300 0 1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_29_266
timestamp 1586364061
transform 1 0 25576 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_274
timestamp 1586364061
transform 1 0 26312 0 1 17952
box -38 -48 314 592
use scs8hd_buf_2  _287_
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_30_19
timestamp 1586364061
transform 1 0 2852 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4416 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 5428 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 4876 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5244 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_39
timestamp 1586364061
transform 1 0 4692 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_43
timestamp 1586364061
transform 1 0 5060 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_58
timestamp 1586364061
transform 1 0 6440 0 -1 19040
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_66
timestamp 1586364061
transform 1 0 7176 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_70
timestamp 1586364061
transform 1 0 7544 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_88
timestamp 1586364061
transform 1 0 9200 0 -1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11684 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__220__B
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_107
timestamp 1586364061
transform 1 0 10948 0 -1 19040
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12696 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_124
timestamp 1586364061
transform 1 0 12512 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_128
timestamp 1586364061
transform 1 0 12880 0 -1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 -1 19040
box -38 -48 866 592
use scs8hd_fill_2  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14260 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_149
timestamp 1586364061
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_3  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15732 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15548 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_170
timestamp 1586364061
transform 1 0 16744 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_174
timestamp 1586364061
transform 1 0 17112 0 -1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_187
timestamp 1586364061
transform 1 0 18308 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_192
timestamp 1586364061
transform 1 0 18768 0 -1 19040
box -38 -48 314 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 19044 0 -1 19040
box -38 -48 866 592
use scs8hd_fill_2  FILLER_30_204
timestamp 1586364061
transform 1 0 19872 0 -1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21068 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20056 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_208
timestamp 1586364061
transform 1 0 20240 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_2  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 21252 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_228
timestamp 1586364061
transform 1 0 22080 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22816 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24380 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_256
timestamp 1586364061
transform 1 0 24656 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_267
timestamp 1586364061
transform 1 0 25668 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_6
timestamp 1586364061
transform 1 0 1656 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_10
timestamp 1586364061
transform 1 0 2024 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3128 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_14
timestamp 1586364061
transform 1 0 2392 0 1 19040
box -38 -48 590 592
use scs8hd_fill_2  FILLER_31_25
timestamp 1586364061
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use scs8hd_conb_1  _243_
timestamp 1586364061
transform 1 0 4140 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_29
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_36
timestamp 1586364061
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_40
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8096 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8648 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8464 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_78
timestamp 1586364061
transform 1 0 8280 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _223_
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__223__A
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_91
timestamp 1586364061
transform 1 0 9476 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_95
timestamp 1586364061
transform 1 0 9844 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 11408 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_134
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_138
timestamp 1586364061
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_151
timestamp 1586364061
transform 1 0 14996 0 1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_156
timestamp 1586364061
transform 1 0 15456 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_162
timestamp 1586364061
transform 1 0 16008 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 19596 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_193
timestamp 1586364061
transform 1 0 18860 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_197
timestamp 1586364061
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_210
timestamp 1586364061
transform 1 0 20424 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_214
timestamp 1586364061
transform 1 0 20792 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_217
timestamp 1586364061
transform 1 0 21068 0 1 19040
box -38 -48 130 592
use scs8hd_buf_1  _164_
timestamp 1586364061
transform 1 0 22172 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_221
timestamp 1586364061
transform 1 0 21436 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_225
timestamp 1586364061
transform 1 0 21804 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 22632 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_236
timestamp 1586364061
transform 1 0 22816 0 1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23828 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24288 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_250
timestamp 1586364061
transform 1 0 24104 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_254
timestamp 1586364061
transform 1 0 24472 0 1 19040
box -38 -48 406 592
use scs8hd_conb_1  _246_
timestamp 1586364061
transform 1 0 24840 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_261
timestamp 1586364061
transform 1 0 25116 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_31_273
timestamp 1586364061
transform 1 0 26220 0 1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_6
timestamp 1586364061
transform 1 0 1656 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_18
timestamp 1586364061
transform 1 0 2760 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 774 592
use scs8hd_buf_1  _198_
timestamp 1586364061
transform 1 0 4600 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_6  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 5612 0 -1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__237__B
timestamp 1586364061
transform 1 0 5060 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_41
timestamp 1586364061
transform 1 0 4876 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_45
timestamp 1586364061
transform 1 0 5244 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_60
timestamp 1586364061
transform 1 0 6624 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_64
timestamp 1586364061
transform 1 0 6992 0 -1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_67
timestamp 1586364061
transform 1 0 7268 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_77
timestamp 1586364061
transform 1 0 8188 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_81
timestamp 1586364061
transform 1 0 8556 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_86
timestamp 1586364061
transform 1 0 9016 0 -1 20128
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__223__B
timestamp 1586364061
transform 1 0 10396 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_96
timestamp 1586364061
transform 1 0 9936 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_100
timestamp 1586364061
transform 1 0 10304 0 -1 20128
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 11408 0 -1 20128
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_32_103
timestamp 1586364061
transform 1 0 10580 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_111
timestamp 1586364061
transform 1 0 11316 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12604 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_123
timestamp 1586364061
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_127
timestamp 1586364061
transform 1 0 12788 0 -1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13156 0 -1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_142
timestamp 1586364061
transform 1 0 14168 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_146
timestamp 1586364061
transform 1 0 14536 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_149
timestamp 1586364061
transform 1 0 14812 0 -1 20128
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16192 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_157
timestamp 1586364061
transform 1 0 15548 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_163
timestamp 1586364061
transform 1 0 16100 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_175
timestamp 1586364061
transform 1 0 17204 0 -1 20128
box -38 -48 774 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 18400 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_183
timestamp 1586364061
transform 1 0 17940 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_186
timestamp 1586364061
transform 1 0 18216 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 19596 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_199
timestamp 1586364061
transform 1 0 19412 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_203
timestamp 1586364061
transform 1 0 19780 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_32_211
timestamp 1586364061
transform 1 0 20516 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_218
timestamp 1586364061
transform 1 0 21160 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_230
timestamp 1586364061
transform 1 0 22264 0 -1 20128
box -38 -48 406 592
use scs8hd_conb_1  _240_
timestamp 1586364061
transform 1 0 22632 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_237
timestamp 1586364061
transform 1 0 22908 0 -1 20128
box -38 -48 774 592
use scs8hd_conb_1  _242_
timestamp 1586364061
transform 1 0 24656 0 -1 20128
box -38 -48 314 592
use scs8hd_conb_1  _251_
timestamp 1586364061
transform 1 0 23644 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_248
timestamp 1586364061
transform 1 0 23920 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_32_259
timestamp 1586364061
transform 1 0 24932 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_271
timestamp 1586364061
transform 1 0 26036 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_buf_2  _282_
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1472 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__282__A
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_11
timestamp 1586364061
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_7
timestamp 1586364061
transform 1 0 1748 0 -1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2300 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_19
timestamp 1586364061
transform 1 0 2852 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_1  _233_
timestamp 1586364061
transform 1 0 3864 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 4324 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 3680 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_33
timestamp 1586364061
transform 1 0 4140 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_37
timestamp 1586364061
transform 1 0 4508 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 774 592
use scs8hd_nor2_4  _236_
timestamp 1586364061
transform 1 0 5796 0 -1 21216
box -38 -48 866 592
use scs8hd_nor2_4  _237_
timestamp 1586364061
transform 1 0 4876 0 1 20128
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4784 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__236__B
timestamp 1586364061
transform 1 0 5612 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_50
timestamp 1586364061
transform 1 0 5704 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_43
timestamp 1586364061
transform 1 0 5060 0 -1 21216
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 5888 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_54
timestamp 1586364061
transform 1 0 6072 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_58
timestamp 1586364061
transform 1 0 6440 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_60
timestamp 1586364061
transform 1 0 6624 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_64
timestamp 1586364061
transform 1 0 6992 0 -1 21216
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_73
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_77
timestamp 1586364061
transform 1 0 8188 0 1 20128
box -38 -48 406 592
use scs8hd_decap_3  FILLER_34_72
timestamp 1586364061
transform 1 0 7728 0 -1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8832 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_81
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_84
timestamp 1586364061
transform 1 0 8832 0 -1 21216
box -38 -48 774 592
use scs8hd_nor2_4  _221_
timestamp 1586364061
transform 1 0 10396 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__221__A
timestamp 1586364061
transform 1 0 10212 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__221__B
timestamp 1586364061
transform 1 0 9844 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_93
timestamp 1586364061
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_97
timestamp 1586364061
transform 1 0 10028 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_102
timestamp 1586364061
transform 1 0 10488 0 -1 21216
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_114
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_110
timestamp 1586364061
transform 1 0 11224 0 -1 21216
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_127
timestamp 1586364061
transform 1 0 12788 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_122
timestamp 1586364061
transform 1 0 12328 0 -1 21216
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_139
timestamp 1586364061
transform 1 0 13892 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_139
timestamp 1586364061
transform 1 0 13892 0 -1 21216
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_143
timestamp 1586364061
transform 1 0 14260 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_151
timestamp 1586364061
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 130 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 15364 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 15640 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 16008 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_156
timestamp 1586364061
transform 1 0 15456 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_160
timestamp 1586364061
transform 1 0 15824 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_164
timestamp 1586364061
transform 1 0 16192 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_164
timestamp 1586364061
transform 1 0 16192 0 -1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_174
timestamp 1586364061
transform 1 0 17112 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_178
timestamp 1586364061
transform 1 0 17480 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_168
timestamp 1586364061
transform 1 0 16560 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_175
timestamp 1586364061
transform 1 0 17204 0 -1 21216
box -38 -48 774 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17940 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_186
timestamp 1586364061
transform 1 0 18216 0 -1 21216
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18952 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_193
timestamp 1586364061
transform 1 0 18860 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_197
timestamp 1586364061
transform 1 0 19228 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_197
timestamp 1586364061
transform 1 0 19228 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_209
timestamp 1586364061
transform 1 0 20332 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_33_210
timestamp 1586364061
transform 1 0 20424 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_206
timestamp 1586364061
transform 1 0 20056 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_213
timestamp 1586364061
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_217
timestamp 1586364061
transform 1 0 21068 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20792 0 1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_218
timestamp 1586364061
transform 1 0 21160 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21804 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21252 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22264 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_221
timestamp 1586364061
transform 1 0 21436 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_228
timestamp 1586364061
transform 1 0 22080 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_230
timestamp 1586364061
transform 1 0 22264 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_242
timestamp 1586364061
transform 1 0 23368 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_254
timestamp 1586364061
transform 1 0 24472 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_34_266
timestamp 1586364061
transform 1 0 25576 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_274
timestamp 1586364061
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_conb_1  _244_
timestamp 1586364061
transform 1 0 5704 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_35_47
timestamp 1586364061
transform 1 0 5428 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6992 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7544 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_66
timestamp 1586364061
transform 1 0 7176 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_73
timestamp 1586364061
transform 1 0 7820 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_77
timestamp 1586364061
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_90
timestamp 1586364061
transform 1 0 9384 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_95
timestamp 1586364061
transform 1 0 9844 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_101
timestamp 1586364061
transform 1 0 10396 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11132 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10948 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10580 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_105
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_112
timestamp 1586364061
transform 1 0 11408 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12788 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_116
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_120
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13156 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_129
timestamp 1586364061
transform 1 0 12972 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14904 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_142
timestamp 1586364061
transform 1 0 14168 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_146
timestamp 1586364061
transform 1 0 14536 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_153
timestamp 1586364061
transform 1 0 15180 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15916 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15364 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16376 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_157
timestamp 1586364061
transform 1 0 15548 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_164
timestamp 1586364061
transform 1 0 16192 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16744 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_168
timestamp 1586364061
transform 1 0 16560 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_175
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_179
timestamp 1586364061
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use scs8hd_buf_1  _165_
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_187
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_191
timestamp 1586364061
transform 1 0 18676 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 18860 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_198
timestamp 1586364061
transform 1 0 19320 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_202
timestamp 1586364061
transform 1 0 19688 0 1 21216
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20424 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_213
timestamp 1586364061
transform 1 0 20700 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_217
timestamp 1586364061
transform 1 0 21068 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21252 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_221
timestamp 1586364061
transform 1 0 21436 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_233
timestamp 1586364061
transform 1 0 22540 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_35_241
timestamp 1586364061
transform 1 0 23276 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6716 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_60
timestamp 1586364061
transform 1 0 6624 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_64
timestamp 1586364061
transform 1 0 6992 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7912 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_72
timestamp 1586364061
transform 1 0 7728 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_77
timestamp 1586364061
transform 1 0 8188 0 -1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_83
timestamp 1586364061
transform 1 0 8740 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_87
timestamp 1586364061
transform 1 0 9108 0 -1 22304
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_91
timestamp 1586364061
transform 1 0 9476 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_96
timestamp 1586364061
transform 1 0 9936 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__269__A
timestamp 1586364061
transform 1 0 10672 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_106
timestamp 1586364061
transform 1 0 10856 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_110
timestamp 1586364061
transform 1 0 11224 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11960 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_121
timestamp 1586364061
transform 1 0 12236 0 -1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_138
timestamp 1586364061
transform 1 0 13800 0 -1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_142
timestamp 1586364061
transform 1 0 14168 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  FILLER_36_150
timestamp 1586364061
transform 1 0 14904 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 130 592
use scs8hd_buf_1  _153_
timestamp 1586364061
transform 1 0 15364 0 -1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_158
timestamp 1586364061
transform 1 0 15640 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17388 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_169
timestamp 1586364061
transform 1 0 16652 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18400 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_180
timestamp 1586364061
transform 1 0 17664 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_12  FILLER_36_191
timestamp 1586364061
transform 1 0 18676 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_36_203
timestamp 1586364061
transform 1 0 19780 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_36_211
timestamp 1586364061
transform 1 0 20516 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_218
timestamp 1586364061
transform 1 0 21160 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_230
timestamp 1586364061
transform 1 0 22264 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_242
timestamp 1586364061
transform 1 0 23368 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_254
timestamp 1586364061
transform 1 0 24472 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_36_266
timestamp 1586364061
transform 1 0 25576 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_274
timestamp 1586364061
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_19
timestamp 1586364061
transform 1 0 2852 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_31
timestamp 1586364061
transform 1 0 3956 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_43
timestamp 1586364061
transform 1 0 5060 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_37_55
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 590 592
use scs8hd_decap_6  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 590 592
use scs8hd_buf_2  _252_
timestamp 1586364061
transform 1 0 7452 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__252__A
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_68
timestamp 1586364061
transform 1 0 7360 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_73
timestamp 1586364061
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_77
timestamp 1586364061
transform 1 0 8188 0 1 22304
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8648 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9108 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_81
timestamp 1586364061
transform 1 0 8556 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_85
timestamp 1586364061
transform 1 0 8924 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_89
timestamp 1586364061
transform 1 0 9292 0 1 22304
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10488 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_96
timestamp 1586364061
transform 1 0 9936 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_100
timestamp 1586364061
transform 1 0 10304 0 1 22304
box -38 -48 222 592
use scs8hd_buf_2  _269_
timestamp 1586364061
transform 1 0 10672 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_108
timestamp 1586364061
transform 1 0 11040 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_112
timestamp 1586364061
transform 1 0 11408 0 1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_120
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13616 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_130
timestamp 1586364061
transform 1 0 13064 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_134
timestamp 1586364061
transform 1 0 13432 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_138
timestamp 1586364061
transform 1 0 13800 0 1 22304
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15180 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_145
timestamp 1586364061
transform 1 0 14444 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_149
timestamp 1586364061
transform 1 0 14812 0 1 22304
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16192 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15640 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16008 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_156
timestamp 1586364061
transform 1 0 15456 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_160
timestamp 1586364061
transform 1 0 15824 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16652 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_167
timestamp 1586364061
transform 1 0 16468 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_171
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_175
timestamp 1586364061
transform 1 0 17204 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__281__A
timestamp 1586364061
transform 1 0 24564 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_37_253
timestamp 1586364061
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_6
timestamp 1586364061
transform 1 0 1656 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_18
timestamp 1586364061
transform 1 0 2760 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_30
timestamp 1586364061
transform 1 0 3864 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_96
timestamp 1586364061
transform 1 0 9936 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11132 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_108
timestamp 1586364061
transform 1 0 11040 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_112
timestamp 1586364061
transform 1 0 11408 0 -1 23392
box -38 -48 774 592
use scs8hd_conb_1  _247_
timestamp 1586364061
transform 1 0 12144 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_123
timestamp 1586364061
transform 1 0 12420 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13156 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_134
timestamp 1586364061
transform 1 0 13432 0 -1 23392
box -38 -48 774 592
use scs8hd_conb_1  _250_
timestamp 1586364061
transform 1 0 14168 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16284 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_157
timestamp 1586364061
transform 1 0 15548 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_38_168
timestamp 1586364061
transform 1 0 16560 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_180
timestamp 1586364061
transform 1 0 17664 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_192
timestamp 1586364061
transform 1 0 18768 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_204
timestamp 1586364061
transform 1 0 19872 0 -1 23392
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_212
timestamp 1586364061
transform 1 0 20608 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_2  _281_
timestamp 1586364061
transform 1 0 24564 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_259
timestamp 1586364061
transform 1 0 24932 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_271
timestamp 1586364061
transform 1 0 26036 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_22
timestamp 1586364061
transform 1 0 3128 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_6  FILLER_39_34
timestamp 1586364061
transform 1 0 4232 0 1 23392
box -38 -48 590 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4876 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5336 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_40
timestamp 1586364061
transform 1 0 4784 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_44
timestamp 1586364061
transform 1 0 5152 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_48
timestamp 1586364061
transform 1 0 5520 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _253_
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_39_60
timestamp 1586364061
transform 1 0 6624 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__253__A
timestamp 1586364061
transform 1 0 7360 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_66
timestamp 1586364061
transform 1 0 7176 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_70
timestamp 1586364061
transform 1 0 7544 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_82
timestamp 1586364061
transform 1 0 8648 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_94
timestamp 1586364061
transform 1 0 9752 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_106
timestamp 1586364061
transform 1 0 10856 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _266_
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_118
timestamp 1586364061
transform 1 0 11960 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_127
timestamp 1586364061
transform 1 0 12788 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_8  FILLER_40_128
timestamp 1586364061
transform 1 0 12880 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13616 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__266__A
timestamp 1586364061
transform 1 0 12972 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13340 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_131
timestamp 1586364061
transform 1 0 13156 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_138
timestamp 1586364061
transform 1 0 13800 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_139
timestamp 1586364061
transform 1 0 13892 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14536 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14996 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14352 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_142
timestamp 1586364061
transform 1 0 14168 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_149
timestamp 1586364061
transform 1 0 14812 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_153
timestamp 1586364061
transform 1 0 15180 0 1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_40_151
timestamp 1586364061
transform 1 0 14996 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _275_
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__275__A
timestamp 1586364061
transform 1 0 16284 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_163
timestamp 1586364061
transform 1 0 16100 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_167
timestamp 1586364061
transform 1 0 16468 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_39_179
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _284_
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__284__A
timestamp 1586364061
transform 1 0 18584 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_188
timestamp 1586364061
transform 1 0 18400 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_192
timestamp 1586364061
transform 1 0 18768 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_204
timestamp 1586364061
transform 1 0 19872 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_216
timestamp 1586364061
transform 1 0 20976 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_228
timestamp 1586364061
transform 1 0 22080 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_39_240
timestamp 1586364061
transform 1 0 23184 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _279_
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _283_
timestamp 1586364061
transform 1 0 24564 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__283__A
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_decap_4  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__279__A
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_259
timestamp 1586364061
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_263
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_259
timestamp 1586364061
transform 1 0 24932 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_275
timestamp 1586364061
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_271
timestamp 1586364061
transform 1 0 26036 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_conb_1  _241_
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_126
timestamp 1586364061
transform 1 0 12696 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_138
timestamp 1586364061
transform 1 0 13800 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_150
timestamp 1586364061
transform 1 0 14904 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_162
timestamp 1586364061
transform 1 0 16008 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_174
timestamp 1586364061
transform 1 0 17112 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_41_182
timestamp 1586364061
transform 1 0 17848 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_41_253
timestamp 1586364061
transform 1 0 24380 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_258
timestamp 1586364061
transform 1 0 24840 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_262
timestamp 1586364061
transform 1 0 25208 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_41_274
timestamp 1586364061
transform 1 0 26312 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal3 s 27520 552 28000 672 6 address[0]
port 0 nsew default input
rlabel metal2 s 754 27520 810 28000 6 address[1]
port 1 nsew default input
rlabel metal3 s 0 552 480 672 6 address[2]
port 2 nsew default input
rlabel metal2 s 2226 27520 2282 28000 6 address[3]
port 3 nsew default input
rlabel metal2 s 2502 0 2558 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 3698 27520 3754 28000 6 address[5]
port 5 nsew default input
rlabel metal3 s 0 1776 480 1896 6 address[6]
port 6 nsew default input
rlabel metal2 s 5170 27520 5226 28000 6 bottom_left_grid_pin_13_
port 7 nsew default input
rlabel metal2 s 3514 0 3570 480 6 bottom_right_grid_pin_11_
port 8 nsew default input
rlabel metal2 s 4618 0 4674 480 6 chanx_left_in[0]
port 9 nsew default input
rlabel metal3 s 0 3136 480 3256 6 chanx_left_in[1]
port 10 nsew default input
rlabel metal3 s 27520 1776 28000 1896 6 chanx_left_in[2]
port 11 nsew default input
rlabel metal3 s 0 4496 480 4616 6 chanx_left_in[3]
port 12 nsew default input
rlabel metal3 s 0 5856 480 5976 6 chanx_left_in[4]
port 13 nsew default input
rlabel metal2 s 5630 0 5686 480 6 chanx_left_in[5]
port 14 nsew default input
rlabel metal2 s 6642 0 6698 480 6 chanx_left_in[6]
port 15 nsew default input
rlabel metal3 s 27520 3000 28000 3120 6 chanx_left_in[7]
port 16 nsew default input
rlabel metal3 s 27520 4360 28000 4480 6 chanx_left_in[8]
port 17 nsew default input
rlabel metal2 s 7654 0 7710 480 6 chanx_left_out[0]
port 18 nsew default tristate
rlabel metal3 s 0 7216 480 7336 6 chanx_left_out[1]
port 19 nsew default tristate
rlabel metal2 s 8758 0 8814 480 6 chanx_left_out[2]
port 20 nsew default tristate
rlabel metal3 s 27520 5584 28000 5704 6 chanx_left_out[3]
port 21 nsew default tristate
rlabel metal3 s 0 8440 480 8560 6 chanx_left_out[4]
port 22 nsew default tristate
rlabel metal3 s 0 9800 480 9920 6 chanx_left_out[5]
port 23 nsew default tristate
rlabel metal3 s 0 11160 480 11280 6 chanx_left_out[6]
port 24 nsew default tristate
rlabel metal2 s 6642 27520 6698 28000 6 chanx_left_out[7]
port 25 nsew default tristate
rlabel metal2 s 8114 27520 8170 28000 6 chanx_left_out[8]
port 26 nsew default tristate
rlabel metal3 s 27520 6808 28000 6928 6 chanx_right_in[0]
port 27 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chanx_right_in[1]
port 28 nsew default input
rlabel metal2 s 10782 0 10838 480 6 chanx_right_in[2]
port 29 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chanx_right_in[3]
port 30 nsew default input
rlabel metal2 s 12898 0 12954 480 6 chanx_right_in[4]
port 31 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_right_in[5]
port 32 nsew default input
rlabel metal2 s 9586 27520 9642 28000 6 chanx_right_in[6]
port 33 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chanx_right_in[7]
port 34 nsew default input
rlabel metal3 s 27520 8168 28000 8288 6 chanx_right_in[8]
port 35 nsew default input
rlabel metal2 s 11058 27520 11114 28000 6 chanx_right_out[0]
port 36 nsew default tristate
rlabel metal2 s 14922 0 14978 480 6 chanx_right_out[1]
port 37 nsew default tristate
rlabel metal3 s 27520 9392 28000 9512 6 chanx_right_out[2]
port 38 nsew default tristate
rlabel metal2 s 12530 27520 12586 28000 6 chanx_right_out[3]
port 39 nsew default tristate
rlabel metal2 s 15934 0 15990 480 6 chanx_right_out[4]
port 40 nsew default tristate
rlabel metal3 s 27520 10616 28000 10736 6 chanx_right_out[5]
port 41 nsew default tristate
rlabel metal3 s 27520 11976 28000 12096 6 chanx_right_out[6]
port 42 nsew default tristate
rlabel metal3 s 0 13880 480 14000 6 chanx_right_out[7]
port 43 nsew default tristate
rlabel metal3 s 27520 13200 28000 13320 6 chanx_right_out[8]
port 44 nsew default tristate
rlabel metal2 s 17038 0 17094 480 6 chany_bottom_in[0]
port 45 nsew default input
rlabel metal3 s 27520 14560 28000 14680 6 chany_bottom_in[1]
port 46 nsew default input
rlabel metal2 s 18050 0 18106 480 6 chany_bottom_in[2]
port 47 nsew default input
rlabel metal2 s 19062 0 19118 480 6 chany_bottom_in[3]
port 48 nsew default input
rlabel metal3 s 0 15104 480 15224 6 chany_bottom_in[4]
port 49 nsew default input
rlabel metal2 s 14002 27520 14058 28000 6 chany_bottom_in[5]
port 50 nsew default input
rlabel metal3 s 27520 15784 28000 15904 6 chany_bottom_in[6]
port 51 nsew default input
rlabel metal2 s 20074 0 20130 480 6 chany_bottom_in[7]
port 52 nsew default input
rlabel metal2 s 15474 27520 15530 28000 6 chany_bottom_in[8]
port 53 nsew default input
rlabel metal3 s 27520 17008 28000 17128 6 chany_bottom_out[0]
port 54 nsew default tristate
rlabel metal3 s 27520 18368 28000 18488 6 chany_bottom_out[1]
port 55 nsew default tristate
rlabel metal3 s 0 16464 480 16584 6 chany_bottom_out[2]
port 56 nsew default tristate
rlabel metal2 s 16946 27520 17002 28000 6 chany_bottom_out[3]
port 57 nsew default tristate
rlabel metal3 s 27520 19592 28000 19712 6 chany_bottom_out[4]
port 58 nsew default tristate
rlabel metal2 s 21178 0 21234 480 6 chany_bottom_out[5]
port 59 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chany_bottom_out[6]
port 60 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chany_bottom_out[7]
port 61 nsew default tristate
rlabel metal2 s 22190 0 22246 480 6 chany_bottom_out[8]
port 62 nsew default tristate
rlabel metal2 s 23202 0 23258 480 6 chany_top_in[0]
port 63 nsew default input
rlabel metal2 s 18418 27520 18474 28000 6 chany_top_in[1]
port 64 nsew default input
rlabel metal3 s 27520 20816 28000 20936 6 chany_top_in[2]
port 65 nsew default input
rlabel metal2 s 19890 27520 19946 28000 6 chany_top_in[3]
port 66 nsew default input
rlabel metal2 s 21362 27520 21418 28000 6 chany_top_in[4]
port 67 nsew default input
rlabel metal2 s 22834 27520 22890 28000 6 chany_top_in[5]
port 68 nsew default input
rlabel metal3 s 27520 22176 28000 22296 6 chany_top_in[6]
port 69 nsew default input
rlabel metal3 s 27520 23400 28000 23520 6 chany_top_in[7]
port 70 nsew default input
rlabel metal3 s 27520 24624 28000 24744 6 chany_top_in[8]
port 71 nsew default input
rlabel metal3 s 0 20544 480 20664 6 chany_top_out[0]
port 72 nsew default tristate
rlabel metal2 s 24214 0 24270 480 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 25318 0 25374 480 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 24306 27520 24362 28000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 25778 27520 25834 28000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal3 s 0 21768 480 21888 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 27250 27520 27306 28000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 26330 0 26386 480 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal3 s 27520 25984 28000 26104 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 1490 0 1546 480 6 data_in
port 81 nsew default input
rlabel metal2 s 478 0 534 480 6 enable
port 82 nsew default input
rlabel metal3 s 0 23128 480 23248 6 left_bottom_grid_pin_12_
port 83 nsew default input
rlabel metal3 s 0 24488 480 24608 6 left_top_grid_pin_10_
port 84 nsew default input
rlabel metal3 s 0 25848 480 25968 6 right_bottom_grid_pin_12_
port 85 nsew default input
rlabel metal2 s 27342 0 27398 480 6 right_top_grid_pin_10_
port 86 nsew default input
rlabel metal3 s 27520 27208 28000 27328 6 top_left_grid_pin_13_
port 87 nsew default input
rlabel metal3 s 0 27208 480 27328 6 top_right_grid_pin_11_
port 88 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 89 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 90 nsew default input
<< end >>
