magic
tech sky130A
magscale 1 2
timestamp 1605016838
<< locali >>
rect 67885 235451 67919 235553
rect 65125 235247 65159 235417
rect 77453 235383 77487 235553
rect 116185 235451 116219 235553
rect 87205 235315 87239 235417
rect 91989 235247 92023 235417
rect 110113 235043 110147 235417
rect 125753 235315 125787 235553
rect 128513 235179 128547 235281
rect 133389 235179 133423 235349
rect 142313 235179 142347 235349
rect 134769 224027 134803 234465
rect 80305 151471 80339 151573
rect 59421 134539 59455 144025
rect 59329 115159 59363 132941
rect 84353 58311 84387 58481
rect 84445 58311 84479 58481
rect 88493 58107 88527 58345
rect 96865 58107 96899 58481
rect 99533 58311 99567 58413
rect 128605 58311 128639 58413
rect 147867 58345 147925 58379
rect 109687 58277 109745 58311
rect 135505 58175 135539 58277
rect 145073 58175 145107 58345
rect 198065 47499 198099 57053
rect 75981 18055 76015 18225
<< viali >>
rect 67885 235553 67919 235587
rect 65125 235417 65159 235451
rect 67885 235417 67919 235451
rect 77453 235553 77487 235587
rect 116185 235553 116219 235587
rect 77453 235349 77487 235383
rect 87205 235417 87239 235451
rect 87205 235281 87239 235315
rect 91989 235417 92023 235451
rect 65125 235213 65159 235247
rect 91989 235213 92023 235247
rect 110113 235417 110147 235451
rect 116185 235417 116219 235451
rect 125753 235553 125787 235587
rect 133389 235349 133423 235383
rect 125753 235281 125787 235315
rect 128513 235281 128547 235315
rect 128513 235145 128547 235179
rect 133389 235145 133423 235179
rect 142313 235349 142347 235383
rect 142313 235145 142347 235179
rect 110113 235009 110147 235043
rect 134769 234465 134803 234499
rect 134769 223993 134803 224027
rect 80305 151573 80339 151607
rect 80305 151437 80339 151471
rect 59421 144025 59455 144059
rect 59421 134505 59455 134539
rect 59329 132941 59363 132975
rect 59329 115125 59363 115159
rect 84353 58481 84387 58515
rect 84353 58277 84387 58311
rect 84445 58481 84479 58515
rect 96865 58481 96899 58515
rect 84445 58277 84479 58311
rect 88493 58345 88527 58379
rect 88493 58073 88527 58107
rect 99533 58413 99567 58447
rect 128605 58413 128639 58447
rect 145073 58345 145107 58379
rect 147833 58345 147867 58379
rect 147925 58345 147959 58379
rect 99533 58277 99567 58311
rect 109653 58277 109687 58311
rect 109745 58277 109779 58311
rect 128605 58277 128639 58311
rect 135505 58277 135539 58311
rect 135505 58141 135539 58175
rect 145073 58141 145107 58175
rect 96865 58073 96899 58107
rect 198065 57053 198099 57087
rect 198065 47465 198099 47499
rect 75981 18225 76015 18259
rect 75981 18021 76015 18055
<< metal1 >>
rect 99610 244248 99616 244300
rect 99668 244288 99674 244300
rect 99794 244288 99800 244300
rect 99668 244260 99800 244288
rect 99668 244248 99674 244260
rect 99794 244248 99800 244260
rect 99852 244248 99858 244300
rect 89858 241324 89864 241376
rect 89916 241364 89922 241376
rect 171830 241364 171836 241376
rect 89916 241336 171836 241364
rect 89916 241324 89922 241336
rect 171830 241324 171836 241336
rect 171888 241324 171894 241376
rect 174038 241324 174044 241376
rect 174096 241364 174102 241376
rect 207802 241364 207808 241376
rect 174096 241336 207808 241364
rect 174096 241324 174102 241336
rect 207802 241324 207808 241336
rect 207860 241324 207866 241376
rect 27850 241120 27856 241172
rect 27908 241160 27914 241172
rect 29138 241160 29144 241172
rect 27908 241132 29144 241160
rect 27908 241120 27914 241132
rect 29138 241120 29144 241132
rect 29196 241120 29202 241172
rect 63822 241120 63828 241172
rect 63880 241160 63886 241172
rect 65018 241160 65024 241172
rect 63880 241132 65024 241160
rect 63880 241120 63886 241132
rect 65018 241120 65024 241132
rect 65076 241120 65082 241172
rect 22698 236632 22704 236684
rect 22756 236672 22762 236684
rect 49838 236672 49844 236684
rect 22756 236644 49844 236672
rect 22756 236632 22762 236644
rect 49838 236632 49844 236644
rect 49896 236632 49902 236684
rect 72838 236632 72844 236684
rect 72896 236672 72902 236684
rect 121414 236672 121420 236684
rect 72896 236644 121420 236672
rect 72896 236632 72902 236644
rect 121414 236632 121420 236644
rect 121472 236632 121478 236684
rect 39442 236564 39448 236616
rect 39500 236604 39506 236616
rect 96114 236604 96120 236616
rect 39500 236576 96120 236604
rect 39500 236564 39506 236576
rect 96114 236564 96120 236576
rect 96172 236564 96178 236616
rect 29138 235884 29144 235936
rect 29196 235924 29202 235936
rect 82222 235924 82228 235936
rect 29196 235896 82228 235924
rect 29196 235884 29202 235896
rect 82222 235884 82228 235896
rect 82280 235884 82286 235936
rect 86178 235884 86184 235936
rect 86236 235924 86242 235936
rect 99610 235924 99616 235936
rect 86236 235896 99616 235924
rect 86236 235884 86242 235896
rect 99610 235884 99616 235896
rect 99668 235884 99674 235936
rect 135858 235884 135864 235936
rect 135916 235924 135922 235936
rect 169530 235924 169536 235936
rect 135916 235896 169536 235924
rect 135916 235884 135922 235896
rect 169530 235884 169536 235896
rect 169588 235884 169594 235936
rect 65018 235816 65024 235868
rect 65076 235856 65082 235868
rect 166218 235856 166224 235868
rect 65076 235828 166224 235856
rect 65076 235816 65082 235828
rect 166218 235816 166224 235828
rect 166276 235816 166282 235868
rect 67873 235587 67931 235593
rect 67873 235553 67885 235587
rect 67919 235584 67931 235587
rect 77441 235587 77499 235593
rect 77441 235584 77453 235587
rect 67919 235556 77453 235584
rect 67919 235553 67931 235556
rect 67873 235547 67931 235553
rect 77441 235553 77453 235556
rect 77487 235553 77499 235587
rect 77441 235547 77499 235553
rect 116173 235587 116231 235593
rect 116173 235553 116185 235587
rect 116219 235584 116231 235587
rect 125741 235587 125799 235593
rect 125741 235584 125753 235587
rect 116219 235556 125753 235584
rect 116219 235553 116231 235556
rect 116173 235547 116231 235553
rect 125741 235553 125753 235556
rect 125787 235553 125799 235587
rect 125741 235547 125799 235553
rect 65113 235451 65171 235457
rect 65113 235417 65125 235451
rect 65159 235448 65171 235451
rect 67873 235451 67931 235457
rect 67873 235448 67885 235451
rect 65159 235420 67885 235448
rect 65159 235417 65171 235420
rect 65113 235411 65171 235417
rect 67873 235417 67885 235420
rect 67919 235417 67931 235451
rect 67873 235411 67931 235417
rect 87193 235451 87251 235457
rect 87193 235417 87205 235451
rect 87239 235448 87251 235451
rect 91977 235451 92035 235457
rect 91977 235448 91989 235451
rect 87239 235420 91989 235448
rect 87239 235417 87251 235420
rect 87193 235411 87251 235417
rect 91977 235417 91989 235420
rect 92023 235417 92035 235451
rect 91977 235411 92035 235417
rect 110101 235451 110159 235457
rect 110101 235417 110113 235451
rect 110147 235448 110159 235451
rect 116173 235451 116231 235457
rect 116173 235448 116185 235451
rect 110147 235420 116185 235448
rect 110147 235417 110159 235420
rect 110101 235411 110159 235417
rect 116173 235417 116185 235420
rect 116219 235417 116231 235451
rect 116173 235411 116231 235417
rect 77441 235383 77499 235389
rect 77441 235349 77453 235383
rect 77487 235380 77499 235383
rect 107430 235380 107436 235392
rect 77487 235352 80244 235380
rect 77487 235349 77499 235352
rect 77441 235343 77499 235349
rect 47262 235272 47268 235324
rect 47320 235312 47326 235324
rect 65570 235312 65576 235324
rect 47320 235284 65576 235312
rect 47320 235272 47326 235284
rect 65570 235272 65576 235284
rect 65628 235272 65634 235324
rect 80216 235312 80244 235352
rect 99536 235352 107436 235380
rect 87193 235315 87251 235321
rect 87193 235312 87205 235315
rect 80216 235284 87205 235312
rect 87193 235281 87205 235284
rect 87239 235281 87251 235315
rect 87193 235275 87251 235281
rect 49838 235204 49844 235256
rect 49896 235244 49902 235256
rect 62534 235244 62540 235256
rect 49896 235216 62540 235244
rect 49896 235204 49902 235216
rect 62534 235204 62540 235216
rect 62592 235244 62598 235256
rect 65113 235247 65171 235253
rect 65113 235244 65125 235247
rect 62592 235216 65125 235244
rect 62592 235204 62598 235216
rect 65113 235213 65125 235216
rect 65159 235213 65171 235247
rect 65113 235207 65171 235213
rect 91977 235247 92035 235253
rect 91977 235213 91989 235247
rect 92023 235244 92035 235247
rect 99536 235244 99564 235352
rect 107430 235340 107436 235352
rect 107488 235340 107494 235392
rect 133377 235383 133435 235389
rect 133377 235349 133389 235383
rect 133423 235380 133435 235383
rect 139446 235380 139452 235392
rect 133423 235352 139452 235380
rect 133423 235349 133435 235352
rect 133377 235343 133435 235349
rect 139446 235340 139452 235352
rect 139504 235380 139510 235392
rect 142301 235383 142359 235389
rect 142301 235380 142313 235383
rect 139504 235352 142313 235380
rect 139504 235340 139510 235352
rect 142301 235349 142313 235352
rect 142347 235349 142359 235383
rect 142301 235343 142359 235349
rect 125741 235315 125799 235321
rect 125741 235281 125753 235315
rect 125787 235312 125799 235315
rect 128501 235315 128559 235321
rect 128501 235312 128513 235315
rect 125787 235284 128513 235312
rect 125787 235281 125799 235284
rect 125741 235275 125799 235281
rect 128501 235281 128513 235284
rect 128547 235281 128559 235315
rect 128501 235275 128559 235281
rect 92023 235216 99564 235244
rect 92023 235213 92035 235216
rect 91977 235207 92035 235213
rect 114422 235204 114428 235256
rect 114480 235244 114486 235256
rect 159502 235244 159508 235256
rect 114480 235216 159508 235244
rect 114480 235204 114486 235216
rect 159502 235204 159508 235216
rect 159560 235204 159566 235256
rect 173486 235204 173492 235256
rect 173544 235244 173550 235256
rect 174038 235244 174044 235256
rect 173544 235216 174044 235244
rect 173544 235204 173550 235216
rect 174038 235204 174044 235216
rect 174096 235204 174102 235256
rect 28218 235136 28224 235188
rect 28276 235176 28282 235188
rect 75506 235176 75512 235188
rect 28276 235148 75512 235176
rect 28276 235136 28282 235148
rect 75506 235136 75512 235148
rect 75564 235136 75570 235188
rect 128501 235179 128559 235185
rect 128501 235145 128513 235179
rect 128547 235176 128559 235179
rect 133377 235179 133435 235185
rect 133377 235176 133389 235179
rect 128547 235148 133389 235176
rect 128547 235145 128559 235148
rect 128501 235139 128559 235145
rect 133377 235145 133389 235148
rect 133423 235145 133435 235179
rect 133377 235139 133435 235145
rect 142301 235179 142359 235185
rect 142301 235145 142313 235179
rect 142347 235176 142359 235179
rect 146530 235176 146536 235188
rect 142347 235148 146536 235176
rect 142347 235145 142359 235148
rect 142301 235139 142359 235145
rect 146530 235136 146536 235148
rect 146588 235136 146594 235188
rect 156834 235136 156840 235188
rect 156892 235176 156898 235188
rect 215622 235176 215628 235188
rect 156892 235148 215628 235176
rect 156892 235136 156898 235148
rect 215622 235136 215628 235148
rect 215680 235136 215686 235188
rect 107430 235000 107436 235052
rect 107488 235040 107494 235052
rect 110101 235043 110159 235049
rect 110101 235040 110113 235043
rect 107488 235012 110113 235040
rect 107488 235000 107494 235012
rect 110101 235009 110113 235012
rect 110147 235009 110159 235043
rect 110101 235003 110159 235009
rect 134754 234496 134760 234508
rect 134715 234468 134760 234496
rect 134754 234456 134760 234468
rect 134812 234456 134818 234508
rect 51218 233912 51224 233964
rect 51276 233952 51282 233964
rect 58118 233952 58124 233964
rect 51276 233924 58124 233952
rect 51276 233912 51282 233924
rect 58118 233912 58124 233924
rect 58176 233912 58182 233964
rect 90226 233844 90232 233896
rect 90284 233884 90290 233896
rect 101174 233884 101180 233896
rect 90284 233856 101180 233884
rect 90284 233844 90290 233856
rect 101174 233844 101180 233856
rect 101232 233844 101238 233896
rect 134754 233844 134760 233896
rect 134812 233884 134818 233896
rect 142298 233884 142304 233896
rect 134812 233856 142304 233884
rect 134812 233844 134818 233856
rect 142298 233844 142304 233856
rect 142356 233844 142362 233896
rect 180294 233844 180300 233896
rect 180352 233884 180358 233896
rect 185170 233884 185176 233896
rect 180352 233856 185176 233884
rect 180352 233844 180358 233856
rect 185170 233844 185176 233856
rect 185228 233844 185234 233896
rect 13314 233776 13320 233828
rect 13372 233816 13378 233828
rect 185262 233816 185268 233828
rect 13372 233788 185268 233816
rect 13372 233776 13378 233788
rect 185262 233776 185268 233788
rect 185320 233776 185326 233828
rect 92710 233028 92716 233080
rect 92768 233068 92774 233080
rect 101358 233068 101364 233080
rect 92768 233040 101364 233068
rect 92768 233028 92774 233040
rect 101358 233028 101364 233040
rect 101416 233028 101422 233080
rect 177718 233028 177724 233080
rect 177776 233068 177782 233080
rect 185170 233068 185176 233080
rect 177776 233040 185176 233068
rect 177776 233028 177782 233040
rect 185170 233028 185176 233040
rect 185228 233028 185234 233080
rect 134754 232688 134760 232740
rect 134812 232728 134818 232740
rect 142206 232728 142212 232740
rect 134812 232700 142212 232728
rect 134812 232688 134818 232700
rect 142206 232688 142212 232700
rect 142264 232688 142270 232740
rect 134846 232620 134852 232672
rect 134904 232660 134910 232672
rect 142298 232660 142304 232672
rect 134904 232632 142304 232660
rect 134904 232620 134910 232632
rect 142298 232620 142304 232632
rect 142356 232620 142362 232672
rect 51218 232552 51224 232604
rect 51276 232592 51282 232604
rect 58026 232592 58032 232604
rect 51276 232564 58032 232592
rect 51276 232552 51282 232564
rect 58026 232552 58032 232564
rect 58084 232552 58090 232604
rect 50022 232416 50028 232468
rect 50080 232456 50086 232468
rect 58118 232456 58124 232468
rect 50080 232428 58124 232456
rect 50080 232416 50086 232428
rect 58118 232416 58124 232428
rect 58176 232416 58182 232468
rect 101726 232456 101732 232468
rect 98156 232428 101732 232456
rect 93998 232348 94004 232400
rect 94056 232388 94062 232400
rect 98156 232388 98184 232428
rect 101726 232416 101732 232428
rect 101784 232416 101790 232468
rect 185170 232456 185176 232468
rect 182336 232428 185176 232456
rect 94056 232360 98184 232388
rect 94056 232348 94062 232360
rect 177718 232348 177724 232400
rect 177776 232388 177782 232400
rect 182336 232388 182364 232428
rect 185170 232416 185176 232428
rect 185228 232416 185234 232468
rect 177776 232360 182364 232388
rect 177776 232348 177782 232360
rect 92710 231668 92716 231720
rect 92768 231708 92774 231720
rect 101266 231708 101272 231720
rect 92768 231680 101272 231708
rect 92768 231668 92774 231680
rect 101266 231668 101272 231680
rect 101324 231668 101330 231720
rect 177718 231668 177724 231720
rect 177776 231708 177782 231720
rect 185170 231708 185176 231720
rect 177776 231680 185176 231708
rect 177776 231668 177782 231680
rect 185170 231668 185176 231680
rect 185228 231668 185234 231720
rect 134754 231464 134760 231516
rect 134812 231504 134818 231516
rect 139630 231504 139636 231516
rect 134812 231476 139636 231504
rect 134812 231464 134818 231476
rect 139630 231464 139636 231476
rect 139688 231464 139694 231516
rect 50114 231124 50120 231176
rect 50172 231164 50178 231176
rect 56462 231164 56468 231176
rect 50172 231136 56468 231164
rect 50172 231124 50178 231136
rect 56462 231124 56468 231136
rect 56520 231124 56526 231176
rect 50758 231056 50764 231108
rect 50816 231096 50822 231108
rect 50816 231068 56784 231096
rect 50816 231056 50822 231068
rect 51218 230988 51224 231040
rect 51276 231028 51282 231040
rect 52690 231028 52696 231040
rect 51276 231000 52696 231028
rect 51276 230988 51282 231000
rect 52690 230988 52696 231000
rect 52748 230988 52754 231040
rect 56756 230960 56784 231068
rect 98874 231056 98880 231108
rect 98932 231096 98938 231108
rect 101450 231096 101456 231108
rect 98932 231068 101456 231096
rect 98932 231056 98938 231068
rect 101450 231056 101456 231068
rect 101508 231056 101514 231108
rect 134754 231056 134760 231108
rect 134812 231096 134818 231108
rect 136870 231096 136876 231108
rect 134812 231068 136876 231096
rect 134812 231056 134818 231068
rect 136870 231056 136876 231068
rect 136928 231056 136934 231108
rect 185262 231096 185268 231108
rect 183624 231068 185268 231096
rect 101726 231028 101732 231040
rect 98892 231000 101732 231028
rect 58210 230960 58216 230972
rect 56756 230932 58216 230960
rect 58210 230920 58216 230932
rect 58268 230920 58274 230972
rect 92710 230920 92716 230972
rect 92768 230960 92774 230972
rect 98892 230960 98920 231000
rect 101726 230988 101732 231000
rect 101784 230988 101790 231040
rect 134846 230988 134852 231040
rect 134904 231028 134910 231040
rect 134904 231000 139676 231028
rect 134904 230988 134910 231000
rect 92768 230932 98920 230960
rect 92768 230920 92774 230932
rect 93722 230852 93728 230904
rect 93780 230892 93786 230904
rect 98874 230892 98880 230904
rect 93780 230864 98880 230892
rect 93780 230852 93786 230864
rect 98874 230852 98880 230864
rect 98932 230852 98938 230904
rect 139648 230892 139676 231000
rect 143678 230892 143684 230904
rect 139648 230864 143684 230892
rect 143678 230852 143684 230864
rect 143736 230852 143742 230904
rect 177718 230852 177724 230904
rect 177776 230892 177782 230904
rect 183624 230892 183652 231068
rect 185262 231056 185268 231068
rect 185320 231056 185326 231108
rect 217554 231056 217560 231108
rect 217612 231096 217618 231108
rect 222338 231096 222344 231108
rect 217612 231068 222344 231096
rect 217612 231056 217618 231068
rect 222338 231056 222344 231068
rect 222396 231056 222402 231108
rect 183698 230988 183704 231040
rect 183756 231028 183762 231040
rect 185170 231028 185176 231040
rect 183756 231000 185176 231028
rect 183756 230988 183762 231000
rect 185170 230988 185176 231000
rect 185228 230988 185234 231040
rect 177776 230864 183652 230892
rect 177776 230852 177782 230864
rect 56462 230580 56468 230632
rect 56520 230620 56526 230632
rect 58210 230620 58216 230632
rect 56520 230592 58216 230620
rect 56520 230580 56526 230592
rect 58210 230580 58216 230592
rect 58268 230580 58274 230632
rect 139630 230580 139636 230632
rect 139688 230620 139694 230632
rect 142942 230620 142948 230632
rect 139688 230592 142948 230620
rect 139688 230580 139694 230592
rect 142942 230580 142948 230592
rect 143000 230580 143006 230632
rect 177718 230580 177724 230632
rect 177776 230620 177782 230632
rect 183698 230620 183704 230632
rect 177776 230592 183704 230620
rect 177776 230580 177782 230592
rect 183698 230580 183704 230592
rect 183756 230580 183762 230632
rect 134294 229968 134300 230020
rect 134352 230008 134358 230020
rect 139630 230008 139636 230020
rect 134352 229980 139636 230008
rect 134352 229968 134358 229980
rect 139630 229968 139636 229980
rect 139688 229968 139694 230020
rect 51218 229832 51224 229884
rect 51276 229872 51282 229884
rect 56462 229872 56468 229884
rect 51276 229844 56468 229872
rect 51276 229832 51282 229844
rect 56462 229832 56468 229844
rect 56520 229832 56526 229884
rect 51126 229696 51132 229748
rect 51184 229736 51190 229748
rect 56186 229736 56192 229748
rect 51184 229708 56192 229736
rect 51184 229696 51190 229708
rect 56186 229696 56192 229708
rect 56244 229696 56250 229748
rect 134386 229628 134392 229680
rect 134444 229668 134450 229680
rect 134444 229640 139676 229668
rect 134444 229628 134450 229640
rect 52690 229560 52696 229612
rect 52748 229600 52754 229612
rect 58210 229600 58216 229612
rect 52748 229572 58216 229600
rect 52748 229560 52754 229572
rect 58210 229560 58216 229572
rect 58268 229560 58274 229612
rect 92710 229560 92716 229612
rect 92768 229600 92774 229612
rect 101726 229600 101732 229612
rect 92768 229572 101732 229600
rect 92768 229560 92774 229572
rect 101726 229560 101732 229572
rect 101784 229560 101790 229612
rect 139648 229600 139676 229640
rect 143586 229600 143592 229612
rect 139648 229572 143592 229600
rect 143586 229560 143592 229572
rect 143644 229560 143650 229612
rect 177626 229560 177632 229612
rect 177684 229600 177690 229612
rect 185170 229600 185176 229612
rect 177684 229572 185176 229600
rect 177684 229560 177690 229572
rect 185170 229560 185176 229572
rect 185228 229560 185234 229612
rect 92802 229492 92808 229544
rect 92860 229532 92866 229544
rect 101542 229532 101548 229544
rect 92860 229504 101548 229532
rect 92860 229492 92866 229504
rect 101542 229492 101548 229504
rect 101600 229492 101606 229544
rect 136870 229492 136876 229544
rect 136928 229532 136934 229544
rect 143678 229532 143684 229544
rect 136928 229504 143684 229532
rect 136928 229492 136934 229504
rect 143678 229492 143684 229504
rect 143736 229492 143742 229544
rect 177718 229492 177724 229544
rect 177776 229532 177782 229544
rect 185262 229532 185268 229544
rect 177776 229504 185268 229532
rect 177776 229492 177782 229504
rect 185262 229492 185268 229504
rect 185320 229492 185326 229544
rect 139630 229424 139636 229476
rect 139688 229464 139694 229476
rect 143494 229464 143500 229476
rect 139688 229436 143500 229464
rect 139688 229424 139694 229436
rect 143494 229424 143500 229436
rect 143552 229424 143558 229476
rect 56186 229288 56192 229340
rect 56244 229328 56250 229340
rect 58210 229328 58216 229340
rect 56244 229300 58216 229328
rect 56244 229288 56250 229300
rect 58210 229288 58216 229300
rect 58268 229288 58274 229340
rect 56462 229016 56468 229068
rect 56520 229056 56526 229068
rect 58302 229056 58308 229068
rect 56520 229028 58308 229056
rect 56520 229016 56526 229028
rect 58302 229016 58308 229028
rect 58360 229016 58366 229068
rect 92710 228880 92716 228932
rect 92768 228920 92774 228932
rect 101726 228920 101732 228932
rect 92768 228892 101732 228920
rect 92768 228880 92774 228892
rect 101726 228880 101732 228892
rect 101784 228880 101790 228932
rect 176982 228880 176988 228932
rect 177040 228920 177046 228932
rect 185170 228920 185176 228932
rect 177040 228892 185176 228920
rect 177040 228880 177046 228892
rect 185170 228880 185176 228892
rect 185228 228880 185234 228932
rect 51034 228404 51040 228456
rect 51092 228444 51098 228456
rect 52690 228444 52696 228456
rect 51092 228416 52696 228444
rect 51092 228404 51098 228416
rect 52690 228404 52696 228416
rect 52748 228404 52754 228456
rect 134386 228404 134392 228456
rect 134444 228444 134450 228456
rect 134444 228416 140228 228444
rect 134444 228404 134450 228416
rect 51218 228336 51224 228388
rect 51276 228376 51282 228388
rect 55450 228376 55456 228388
rect 51276 228348 55456 228376
rect 51276 228336 51282 228348
rect 55450 228336 55456 228348
rect 55508 228336 55514 228388
rect 101450 228376 101456 228388
rect 99444 228348 101456 228376
rect 51126 228268 51132 228320
rect 51184 228308 51190 228320
rect 51184 228280 55496 228308
rect 51184 228268 51190 228280
rect 55468 228240 55496 228280
rect 58210 228240 58216 228252
rect 55468 228212 58216 228240
rect 58210 228200 58216 228212
rect 58268 228200 58274 228252
rect 93170 228200 93176 228252
rect 93228 228240 93234 228252
rect 99444 228240 99472 228348
rect 101450 228336 101456 228348
rect 101508 228336 101514 228388
rect 134754 228336 134760 228388
rect 134812 228376 134818 228388
rect 134812 228348 140136 228376
rect 134812 228336 134818 228348
rect 101726 228308 101732 228320
rect 93228 228212 99472 228240
rect 99536 228280 101732 228308
rect 93228 228200 93234 228212
rect 92710 228132 92716 228184
rect 92768 228172 92774 228184
rect 99536 228172 99564 228280
rect 101726 228268 101732 228280
rect 101784 228268 101790 228320
rect 134846 228268 134852 228320
rect 134904 228308 134910 228320
rect 136870 228308 136876 228320
rect 134904 228280 136876 228308
rect 134904 228268 134910 228280
rect 136870 228268 136876 228280
rect 136928 228268 136934 228320
rect 92768 228144 99564 228172
rect 140108 228172 140136 228348
rect 140200 228240 140228 228416
rect 185262 228376 185268 228388
rect 182428 228348 185268 228376
rect 143678 228240 143684 228252
rect 140200 228212 143684 228240
rect 143678 228200 143684 228212
rect 143736 228200 143742 228252
rect 177718 228200 177724 228252
rect 177776 228240 177782 228252
rect 182428 228240 182456 228348
rect 185262 228336 185268 228348
rect 185320 228336 185326 228388
rect 185170 228308 185176 228320
rect 177776 228212 182456 228240
rect 182520 228280 185176 228308
rect 177776 228200 177782 228212
rect 143310 228172 143316 228184
rect 140108 228144 143316 228172
rect 92768 228132 92774 228144
rect 143310 228132 143316 228144
rect 143368 228132 143374 228184
rect 177626 228132 177632 228184
rect 177684 228172 177690 228184
rect 182520 228172 182548 228280
rect 185170 228268 185176 228280
rect 185228 228268 185234 228320
rect 177684 228144 182548 228172
rect 177684 228132 177690 228144
rect 55450 227860 55456 227912
rect 55508 227900 55514 227912
rect 58302 227900 58308 227912
rect 55508 227872 58308 227900
rect 55508 227860 55514 227872
rect 58302 227860 58308 227872
rect 58360 227860 58366 227912
rect 50758 226840 50764 226892
rect 50816 226880 50822 226892
rect 55910 226880 55916 226892
rect 50816 226852 55916 226880
rect 50816 226840 50822 226852
rect 55910 226840 55916 226852
rect 55968 226840 55974 226892
rect 134754 226840 134760 226892
rect 134812 226880 134818 226892
rect 134812 226852 139676 226880
rect 134812 226840 134818 226852
rect 52690 226772 52696 226824
rect 52748 226812 52754 226824
rect 58210 226812 58216 226824
rect 52748 226784 58216 226812
rect 52748 226772 52754 226784
rect 58210 226772 58216 226784
rect 58268 226772 58274 226824
rect 92710 226772 92716 226824
rect 92768 226812 92774 226824
rect 101358 226812 101364 226824
rect 92768 226784 101364 226812
rect 92768 226772 92774 226784
rect 101358 226772 101364 226784
rect 101416 226772 101422 226824
rect 139648 226812 139676 226852
rect 143310 226812 143316 226824
rect 139648 226784 143316 226812
rect 143310 226772 143316 226784
rect 143368 226772 143374 226824
rect 177166 226772 177172 226824
rect 177224 226812 177230 226824
rect 185170 226812 185176 226824
rect 177224 226784 185176 226812
rect 177224 226772 177230 226784
rect 185170 226772 185176 226784
rect 185228 226772 185234 226824
rect 92802 226704 92808 226756
rect 92860 226744 92866 226756
rect 101450 226744 101456 226756
rect 92860 226716 101456 226744
rect 92860 226704 92866 226716
rect 101450 226704 101456 226716
rect 101508 226704 101514 226756
rect 136870 226704 136876 226756
rect 136928 226744 136934 226756
rect 143678 226744 143684 226756
rect 136928 226716 143684 226744
rect 136928 226704 136934 226716
rect 143678 226704 143684 226716
rect 143736 226704 143742 226756
rect 177718 226704 177724 226756
rect 177776 226744 177782 226756
rect 185262 226744 185268 226756
rect 177776 226716 185268 226744
rect 177776 226704 177782 226716
rect 185262 226704 185268 226716
rect 185320 226704 185326 226756
rect 55910 226364 55916 226416
rect 55968 226404 55974 226416
rect 58210 226404 58216 226416
rect 55968 226376 58216 226404
rect 55968 226364 55974 226376
rect 58210 226364 58216 226376
rect 58268 226364 58274 226416
rect 51218 225548 51224 225600
rect 51276 225588 51282 225600
rect 58302 225588 58308 225600
rect 51276 225560 58308 225588
rect 51276 225548 51282 225560
rect 58302 225548 58308 225560
rect 58360 225548 58366 225600
rect 134386 225548 134392 225600
rect 134444 225588 134450 225600
rect 143310 225588 143316 225600
rect 134444 225560 143316 225588
rect 134444 225548 134450 225560
rect 143310 225548 143316 225560
rect 143368 225548 143374 225600
rect 50022 225480 50028 225532
rect 50080 225520 50086 225532
rect 58394 225520 58400 225532
rect 50080 225492 58400 225520
rect 50080 225480 50086 225492
rect 58394 225480 58400 225492
rect 58452 225480 58458 225532
rect 134754 225480 134760 225532
rect 134812 225520 134818 225532
rect 142574 225520 142580 225532
rect 134812 225492 142580 225520
rect 134812 225480 134818 225492
rect 142574 225480 142580 225492
rect 142632 225480 142638 225532
rect 51310 225412 51316 225464
rect 51368 225452 51374 225464
rect 58210 225452 58216 225464
rect 51368 225424 58216 225452
rect 51368 225412 51374 225424
rect 58210 225412 58216 225424
rect 58268 225412 58274 225464
rect 93722 225412 93728 225464
rect 93780 225452 93786 225464
rect 101542 225452 101548 225464
rect 93780 225424 101548 225452
rect 93780 225412 93786 225424
rect 101542 225412 101548 225424
rect 101600 225412 101606 225464
rect 135490 225412 135496 225464
rect 135548 225452 135554 225464
rect 143678 225452 143684 225464
rect 135548 225424 143684 225452
rect 135548 225412 135554 225424
rect 143678 225412 143684 225424
rect 143736 225412 143742 225464
rect 177718 225412 177724 225464
rect 177776 225452 177782 225464
rect 185354 225452 185360 225464
rect 177776 225424 185360 225452
rect 177776 225412 177782 225424
rect 185354 225412 185360 225424
rect 185412 225412 185418 225464
rect 92802 225344 92808 225396
rect 92860 225384 92866 225396
rect 101818 225384 101824 225396
rect 92860 225356 101824 225384
rect 92860 225344 92866 225356
rect 101818 225344 101824 225356
rect 101876 225344 101882 225396
rect 177166 225344 177172 225396
rect 177224 225384 177230 225396
rect 185170 225384 185176 225396
rect 177224 225356 185176 225384
rect 177224 225344 177230 225356
rect 185170 225344 185176 225356
rect 185228 225344 185234 225396
rect 92710 225276 92716 225328
rect 92768 225316 92774 225328
rect 101634 225316 101640 225328
rect 92768 225288 101640 225316
rect 92768 225276 92774 225288
rect 101634 225276 101640 225288
rect 101692 225276 101698 225328
rect 177718 225276 177724 225328
rect 177776 225316 177782 225328
rect 185262 225316 185268 225328
rect 177776 225288 185268 225316
rect 177776 225276 177782 225288
rect 185262 225276 185268 225288
rect 185320 225276 185326 225328
rect 51126 224392 51132 224444
rect 51184 224432 51190 224444
rect 56738 224432 56744 224444
rect 51184 224404 56744 224432
rect 51184 224392 51190 224404
rect 56738 224392 56744 224404
rect 56796 224392 56802 224444
rect 51126 224256 51132 224308
rect 51184 224296 51190 224308
rect 52690 224296 52696 224308
rect 51184 224268 52696 224296
rect 51184 224256 51190 224268
rect 52690 224256 52696 224268
rect 52748 224256 52754 224308
rect 134662 224256 134668 224308
rect 134720 224296 134726 224308
rect 134720 224268 137008 224296
rect 134720 224256 134726 224268
rect 135398 224188 135404 224240
rect 135456 224228 135462 224240
rect 136870 224228 136876 224240
rect 135456 224200 136876 224228
rect 135456 224188 135462 224200
rect 136870 224188 136876 224200
rect 136928 224188 136934 224240
rect 136980 224228 137008 224268
rect 136980 224200 139860 224228
rect 51218 224120 51224 224172
rect 51276 224160 51282 224172
rect 51276 224132 56784 224160
rect 51276 224120 51282 224132
rect 56756 224092 56784 224132
rect 134294 224120 134300 224172
rect 134352 224160 134358 224172
rect 134352 224132 139768 224160
rect 134352 224120 134358 224132
rect 58210 224092 58216 224104
rect 56756 224064 58216 224092
rect 58210 224052 58216 224064
rect 58268 224052 58274 224104
rect 93906 224052 93912 224104
rect 93964 224092 93970 224104
rect 100990 224092 100996 224104
rect 93964 224064 100996 224092
rect 93964 224052 93970 224064
rect 100990 224052 100996 224064
rect 101048 224052 101054 224104
rect 56738 223984 56744 224036
rect 56796 224024 56802 224036
rect 58302 224024 58308 224036
rect 56796 223996 58308 224024
rect 56796 223984 56802 223996
rect 58302 223984 58308 223996
rect 58360 223984 58366 224036
rect 93722 223984 93728 224036
rect 93780 224024 93786 224036
rect 101082 224024 101088 224036
rect 93780 223996 101088 224024
rect 93780 223984 93786 223996
rect 101082 223984 101088 223996
rect 101140 223984 101146 224036
rect 134754 224024 134760 224036
rect 134715 223996 134760 224024
rect 134754 223984 134760 223996
rect 134812 223984 134818 224036
rect 139740 224024 139768 224132
rect 139832 224092 139860 224200
rect 143678 224092 143684 224104
rect 139832 224064 143684 224092
rect 143678 224052 143684 224064
rect 143736 224052 143742 224104
rect 177718 224052 177724 224104
rect 177776 224092 177782 224104
rect 185262 224092 185268 224104
rect 177776 224064 185268 224092
rect 177776 224052 177782 224064
rect 185262 224052 185268 224064
rect 185320 224052 185326 224104
rect 143310 224024 143316 224036
rect 139740 223996 143316 224024
rect 143310 223984 143316 223996
rect 143368 223984 143374 224036
rect 177626 223984 177632 224036
rect 177684 224024 177690 224036
rect 185170 224024 185176 224036
rect 177684 223996 185176 224024
rect 177684 223984 177690 223996
rect 185170 223984 185176 223996
rect 185228 223984 185234 224036
rect 51126 223032 51132 223084
rect 51184 223072 51190 223084
rect 52782 223072 52788 223084
rect 51184 223044 52788 223072
rect 51184 223032 51190 223044
rect 52782 223032 52788 223044
rect 52840 223032 52846 223084
rect 134478 223032 134484 223084
rect 134536 223072 134542 223084
rect 136962 223072 136968 223084
rect 134536 223044 136968 223072
rect 134536 223032 134542 223044
rect 136962 223032 136968 223044
rect 137020 223032 137026 223084
rect 51218 222896 51224 222948
rect 51276 222936 51282 222948
rect 55818 222936 55824 222948
rect 51276 222908 55824 222936
rect 51276 222896 51282 222908
rect 55818 222896 55824 222908
rect 55876 222896 55882 222948
rect 135398 222760 135404 222812
rect 135456 222800 135462 222812
rect 135456 222772 139676 222800
rect 135456 222760 135462 222772
rect 52690 222692 52696 222744
rect 52748 222732 52754 222744
rect 58210 222732 58216 222744
rect 52748 222704 58216 222732
rect 52748 222692 52754 222704
rect 58210 222692 58216 222704
rect 58268 222692 58274 222744
rect 92710 222692 92716 222744
rect 92768 222732 92774 222744
rect 101450 222732 101456 222744
rect 92768 222704 101456 222732
rect 92768 222692 92774 222704
rect 101450 222692 101456 222704
rect 101508 222692 101514 222744
rect 139648 222732 139676 222772
rect 143310 222732 143316 222744
rect 139648 222704 143316 222732
rect 143310 222692 143316 222704
rect 143368 222692 143374 222744
rect 177626 222692 177632 222744
rect 177684 222732 177690 222744
rect 185170 222732 185176 222744
rect 177684 222704 185176 222732
rect 177684 222692 177690 222704
rect 185170 222692 185176 222704
rect 185228 222692 185234 222744
rect 92986 222624 92992 222676
rect 93044 222664 93050 222676
rect 101358 222664 101364 222676
rect 93044 222636 101364 222664
rect 93044 222624 93050 222636
rect 101358 222624 101364 222636
rect 101416 222624 101422 222676
rect 136870 222624 136876 222676
rect 136928 222664 136934 222676
rect 143678 222664 143684 222676
rect 136928 222636 143684 222664
rect 136928 222624 136934 222636
rect 143678 222624 143684 222636
rect 143736 222624 143742 222676
rect 177718 222624 177724 222676
rect 177776 222664 177782 222676
rect 185262 222664 185268 222676
rect 177776 222636 185268 222664
rect 177776 222624 177782 222636
rect 185262 222624 185268 222636
rect 185320 222624 185326 222676
rect 55818 222284 55824 222336
rect 55876 222324 55882 222336
rect 58302 222324 58308 222336
rect 55876 222296 58308 222324
rect 55876 222284 55882 222296
rect 58302 222284 58308 222296
rect 58360 222284 58366 222336
rect 51218 221672 51224 221724
rect 51276 221712 51282 221724
rect 56002 221712 56008 221724
rect 51276 221684 56008 221712
rect 51276 221672 51282 221684
rect 56002 221672 56008 221684
rect 56060 221672 56066 221724
rect 134846 221672 134852 221724
rect 134904 221712 134910 221724
rect 139630 221712 139636 221724
rect 134904 221684 139636 221712
rect 134904 221672 134910 221684
rect 139630 221672 139636 221684
rect 139688 221672 139694 221724
rect 51126 221400 51132 221452
rect 51184 221440 51190 221452
rect 56462 221440 56468 221452
rect 51184 221412 56468 221440
rect 51184 221400 51190 221412
rect 56462 221400 56468 221412
rect 56520 221400 56526 221452
rect 134662 221400 134668 221452
rect 134720 221440 134726 221452
rect 139722 221440 139728 221452
rect 134720 221412 139728 221440
rect 134720 221400 134726 221412
rect 139722 221400 139728 221412
rect 139780 221400 139786 221452
rect 51218 221332 51224 221384
rect 51276 221372 51282 221384
rect 52690 221372 52696 221384
rect 51276 221344 52696 221372
rect 51276 221332 51282 221344
rect 52690 221332 52696 221344
rect 52748 221332 52754 221384
rect 135398 221332 135404 221384
rect 135456 221372 135462 221384
rect 136870 221372 136876 221384
rect 135456 221344 136876 221372
rect 135456 221332 135462 221344
rect 136870 221332 136876 221344
rect 136928 221332 136934 221384
rect 52782 221264 52788 221316
rect 52840 221304 52846 221316
rect 58210 221304 58216 221316
rect 52840 221276 58216 221304
rect 52840 221264 52846 221276
rect 58210 221264 58216 221276
rect 58268 221264 58274 221316
rect 92802 221264 92808 221316
rect 92860 221304 92866 221316
rect 101542 221304 101548 221316
rect 92860 221276 101548 221304
rect 92860 221264 92866 221276
rect 101542 221264 101548 221276
rect 101600 221264 101606 221316
rect 136962 221264 136968 221316
rect 137020 221304 137026 221316
rect 143678 221304 143684 221316
rect 137020 221276 143684 221304
rect 137020 221264 137026 221276
rect 143678 221264 143684 221276
rect 143736 221264 143742 221316
rect 177166 221264 177172 221316
rect 177224 221304 177230 221316
rect 185170 221304 185176 221316
rect 177224 221276 185176 221304
rect 177224 221264 177230 221276
rect 185170 221264 185176 221276
rect 185228 221264 185234 221316
rect 93722 221196 93728 221248
rect 93780 221236 93786 221248
rect 101634 221236 101640 221248
rect 93780 221208 101640 221236
rect 93780 221196 93786 221208
rect 101634 221196 101640 221208
rect 101692 221196 101698 221248
rect 177626 221196 177632 221248
rect 177684 221236 177690 221248
rect 185262 221236 185268 221248
rect 177684 221208 185268 221236
rect 177684 221196 177690 221208
rect 185262 221196 185268 221208
rect 185320 221196 185326 221248
rect 92710 221128 92716 221180
rect 92768 221168 92774 221180
rect 100898 221168 100904 221180
rect 92768 221140 100904 221168
rect 92768 221128 92774 221140
rect 100898 221128 100904 221140
rect 100956 221128 100962 221180
rect 177718 221128 177724 221180
rect 177776 221168 177782 221180
rect 185078 221168 185084 221180
rect 177776 221140 185084 221168
rect 177776 221128 177782 221140
rect 185078 221128 185084 221140
rect 185136 221128 185142 221180
rect 56002 221060 56008 221112
rect 56060 221100 56066 221112
rect 58210 221100 58216 221112
rect 56060 221072 58216 221100
rect 56060 221060 56066 221072
rect 58210 221060 58216 221072
rect 58268 221060 58274 221112
rect 139630 220924 139636 220976
rect 139688 220964 139694 220976
rect 143310 220964 143316 220976
rect 139688 220936 143316 220964
rect 139688 220924 139694 220936
rect 143310 220924 143316 220936
rect 143368 220924 143374 220976
rect 56462 220652 56468 220704
rect 56520 220692 56526 220704
rect 58302 220692 58308 220704
rect 56520 220664 58308 220692
rect 56520 220652 56526 220664
rect 58302 220652 58308 220664
rect 58360 220652 58366 220704
rect 139722 220584 139728 220636
rect 139780 220624 139786 220636
rect 143678 220624 143684 220636
rect 139780 220596 143684 220624
rect 139780 220584 139786 220596
rect 143678 220584 143684 220596
rect 143736 220584 143742 220636
rect 135306 220108 135312 220160
rect 135364 220148 135370 220160
rect 138158 220148 138164 220160
rect 135364 220120 138164 220148
rect 135364 220108 135370 220120
rect 138158 220108 138164 220120
rect 138216 220108 138222 220160
rect 51126 220040 51132 220092
rect 51184 220080 51190 220092
rect 52782 220080 52788 220092
rect 51184 220052 52788 220080
rect 51184 220040 51190 220052
rect 52782 220040 52788 220052
rect 52840 220040 52846 220092
rect 51218 219972 51224 220024
rect 51276 220012 51282 220024
rect 55818 220012 55824 220024
rect 51276 219984 55824 220012
rect 51276 219972 51282 219984
rect 55818 219972 55824 219984
rect 55876 219972 55882 220024
rect 135398 219972 135404 220024
rect 135456 220012 135462 220024
rect 135456 219984 139676 220012
rect 135456 219972 135462 219984
rect 52690 219904 52696 219956
rect 52748 219944 52754 219956
rect 58210 219944 58216 219956
rect 52748 219916 58216 219944
rect 52748 219904 52754 219916
rect 58210 219904 58216 219916
rect 58268 219904 58274 219956
rect 93722 219904 93728 219956
rect 93780 219944 93786 219956
rect 101818 219944 101824 219956
rect 93780 219916 101824 219944
rect 93780 219904 93786 219916
rect 101818 219904 101824 219916
rect 101876 219904 101882 219956
rect 139648 219944 139676 219984
rect 143126 219944 143132 219956
rect 139648 219916 143132 219944
rect 143126 219904 143132 219916
rect 143184 219904 143190 219956
rect 177166 219904 177172 219956
rect 177224 219944 177230 219956
rect 185170 219944 185176 219956
rect 177224 219916 185176 219944
rect 177224 219904 177230 219916
rect 185170 219904 185176 219916
rect 185228 219904 185234 219956
rect 93906 219836 93912 219888
rect 93964 219876 93970 219888
rect 101266 219876 101272 219888
rect 93964 219848 101272 219876
rect 93964 219836 93970 219848
rect 101266 219836 101272 219848
rect 101324 219836 101330 219888
rect 136870 219836 136876 219888
rect 136928 219876 136934 219888
rect 143678 219876 143684 219888
rect 136928 219848 143684 219876
rect 136928 219836 136934 219848
rect 143678 219836 143684 219848
rect 143736 219836 143742 219888
rect 177718 219836 177724 219888
rect 177776 219876 177782 219888
rect 185354 219876 185360 219888
rect 177776 219848 185360 219876
rect 177776 219836 177782 219848
rect 185354 219836 185360 219848
rect 185412 219836 185418 219888
rect 55818 219292 55824 219344
rect 55876 219332 55882 219344
rect 58302 219332 58308 219344
rect 55876 219304 58308 219332
rect 55876 219292 55882 219304
rect 58302 219292 58308 219304
rect 58360 219292 58366 219344
rect 51218 218816 51224 218868
rect 51276 218856 51282 218868
rect 53334 218856 53340 218868
rect 51276 218828 53340 218856
rect 51276 218816 51282 218828
rect 53334 218816 53340 218828
rect 53392 218816 53398 218868
rect 135030 218816 135036 218868
rect 135088 218856 135094 218868
rect 137514 218856 137520 218868
rect 135088 218828 137520 218856
rect 135088 218816 135094 218828
rect 137514 218816 137520 218828
rect 137572 218816 137578 218868
rect 51218 218680 51224 218732
rect 51276 218720 51282 218732
rect 52782 218720 52788 218732
rect 51276 218692 52788 218720
rect 51276 218680 51282 218692
rect 52782 218680 52788 218692
rect 52840 218680 52846 218732
rect 135398 218680 135404 218732
rect 135456 218720 135462 218732
rect 135456 218692 140228 218720
rect 135456 218680 135462 218692
rect 50850 218612 50856 218664
rect 50908 218652 50914 218664
rect 55450 218652 55456 218664
rect 50908 218624 55456 218652
rect 50908 218612 50914 218624
rect 55450 218612 55456 218624
rect 55508 218612 55514 218664
rect 93538 218612 93544 218664
rect 93596 218652 93602 218664
rect 101726 218652 101732 218664
rect 93596 218624 101732 218652
rect 93596 218612 93602 218624
rect 101726 218612 101732 218624
rect 101784 218612 101790 218664
rect 135306 218612 135312 218664
rect 135364 218652 135370 218664
rect 137974 218652 137980 218664
rect 135364 218624 137980 218652
rect 135364 218612 135370 218624
rect 137974 218612 137980 218624
rect 138032 218612 138038 218664
rect 52690 218544 52696 218596
rect 52748 218584 52754 218596
rect 58210 218584 58216 218596
rect 52748 218556 58216 218584
rect 52748 218544 52754 218556
rect 58210 218544 58216 218556
rect 58268 218544 58274 218596
rect 93722 218544 93728 218596
rect 93780 218584 93786 218596
rect 101358 218584 101364 218596
rect 93780 218556 101364 218584
rect 93780 218544 93786 218556
rect 101358 218544 101364 218556
rect 101416 218544 101422 218596
rect 140200 218584 140228 218692
rect 177994 218612 178000 218664
rect 178052 218652 178058 218664
rect 185170 218652 185176 218664
rect 178052 218624 185176 218652
rect 178052 218612 178058 218624
rect 185170 218612 185176 218624
rect 185228 218612 185234 218664
rect 143494 218584 143500 218596
rect 140200 218556 143500 218584
rect 143494 218544 143500 218556
rect 143552 218544 143558 218596
rect 177166 218544 177172 218596
rect 177224 218584 177230 218596
rect 185814 218584 185820 218596
rect 177224 218556 185820 218584
rect 177224 218544 177230 218556
rect 185814 218544 185820 218556
rect 185872 218544 185878 218596
rect 93170 218476 93176 218528
rect 93228 218516 93234 218528
rect 100898 218516 100904 218528
rect 93228 218488 100904 218516
rect 93228 218476 93234 218488
rect 100898 218476 100904 218488
rect 100956 218476 100962 218528
rect 138158 218476 138164 218528
rect 138216 218516 138222 218528
rect 143678 218516 143684 218528
rect 138216 218488 143684 218516
rect 138216 218476 138222 218488
rect 143678 218476 143684 218488
rect 143736 218476 143742 218528
rect 177718 218476 177724 218528
rect 177776 218516 177782 218528
rect 185078 218516 185084 218528
rect 177776 218488 185084 218516
rect 177776 218476 177782 218488
rect 185078 218476 185084 218488
rect 185136 218476 185142 218528
rect 55450 218000 55456 218052
rect 55508 218040 55514 218052
rect 58210 218040 58216 218052
rect 55508 218012 58216 218040
rect 55508 218000 55514 218012
rect 58210 218000 58216 218012
rect 58268 218000 58274 218052
rect 51218 217320 51224 217372
rect 51276 217360 51282 217372
rect 52874 217360 52880 217372
rect 51276 217332 52880 217360
rect 51276 217320 51282 217332
rect 52874 217320 52880 217332
rect 52932 217320 52938 217372
rect 134478 217320 134484 217372
rect 134536 217360 134542 217372
rect 137606 217360 137612 217372
rect 134536 217332 137612 217360
rect 134536 217320 134542 217332
rect 137606 217320 137612 217332
rect 137664 217320 137670 217372
rect 135398 217252 135404 217304
rect 135456 217292 135462 217304
rect 137698 217292 137704 217304
rect 135456 217264 137704 217292
rect 135456 217252 135462 217264
rect 137698 217252 137704 217264
rect 137756 217252 137762 217304
rect 50758 217184 50764 217236
rect 50816 217224 50822 217236
rect 52690 217224 52696 217236
rect 50816 217196 52696 217224
rect 50816 217184 50822 217196
rect 52690 217184 52696 217196
rect 52748 217184 52754 217236
rect 101174 217224 101180 217236
rect 98892 217196 101180 217224
rect 53334 217116 53340 217168
rect 53392 217156 53398 217168
rect 58210 217156 58216 217168
rect 53392 217128 58216 217156
rect 53392 217116 53398 217128
rect 58210 217116 58216 217128
rect 58268 217116 58274 217168
rect 92710 217116 92716 217168
rect 92768 217156 92774 217168
rect 98892 217156 98920 217196
rect 101174 217184 101180 217196
rect 101232 217184 101238 217236
rect 185170 217224 185176 217236
rect 183440 217196 185176 217224
rect 92768 217128 98920 217156
rect 92768 217116 92774 217128
rect 137514 217116 137520 217168
rect 137572 217156 137578 217168
rect 143678 217156 143684 217168
rect 137572 217128 143684 217156
rect 137572 217116 137578 217128
rect 143678 217116 143684 217128
rect 143736 217116 143742 217168
rect 177718 217116 177724 217168
rect 177776 217156 177782 217168
rect 183440 217156 183468 217196
rect 185170 217184 185176 217196
rect 185228 217184 185234 217236
rect 177776 217128 183468 217156
rect 177776 217116 177782 217128
rect 52782 217048 52788 217100
rect 52840 217088 52846 217100
rect 58302 217088 58308 217100
rect 52840 217060 58308 217088
rect 52840 217048 52846 217060
rect 58302 217048 58308 217060
rect 58360 217048 58366 217100
rect 137974 217048 137980 217100
rect 138032 217088 138038 217100
rect 143126 217088 143132 217100
rect 138032 217060 143132 217088
rect 138032 217048 138038 217060
rect 143126 217048 143132 217060
rect 143184 217048 143190 217100
rect 51126 215824 51132 215876
rect 51184 215864 51190 215876
rect 56462 215864 56468 215876
rect 51184 215836 56468 215864
rect 51184 215824 51190 215836
rect 56462 215824 56468 215836
rect 56520 215824 56526 215876
rect 135398 215824 135404 215876
rect 135456 215864 135462 215876
rect 135456 215836 139676 215864
rect 135456 215824 135462 215836
rect 52690 215756 52696 215808
rect 52748 215796 52754 215808
rect 58210 215796 58216 215808
rect 52748 215768 58216 215796
rect 52748 215756 52754 215768
rect 58210 215756 58216 215768
rect 58268 215756 58274 215808
rect 93538 215756 93544 215808
rect 93596 215796 93602 215808
rect 101358 215796 101364 215808
rect 93596 215768 101364 215796
rect 93596 215756 93602 215768
rect 101358 215756 101364 215768
rect 101416 215756 101422 215808
rect 139648 215796 139676 215836
rect 143494 215796 143500 215808
rect 139648 215768 143500 215796
rect 143494 215756 143500 215768
rect 143552 215756 143558 215808
rect 177166 215756 177172 215808
rect 177224 215796 177230 215808
rect 185170 215796 185176 215808
rect 177224 215768 185176 215796
rect 177224 215756 177230 215768
rect 185170 215756 185176 215768
rect 185228 215756 185234 215808
rect 52874 215688 52880 215740
rect 52932 215728 52938 215740
rect 58302 215728 58308 215740
rect 52932 215700 58308 215728
rect 52932 215688 52938 215700
rect 58302 215688 58308 215700
rect 58360 215688 58366 215740
rect 92710 215688 92716 215740
rect 92768 215728 92774 215740
rect 100806 215728 100812 215740
rect 92768 215700 100812 215728
rect 92768 215688 92774 215700
rect 100806 215688 100812 215700
rect 100864 215688 100870 215740
rect 137698 215688 137704 215740
rect 137756 215728 137762 215740
rect 143126 215728 143132 215740
rect 137756 215700 143132 215728
rect 137756 215688 137762 215700
rect 143126 215688 143132 215700
rect 143184 215688 143190 215740
rect 177718 215688 177724 215740
rect 177776 215728 177782 215740
rect 184986 215728 184992 215740
rect 177776 215700 184992 215728
rect 177776 215688 177782 215700
rect 184986 215688 184992 215700
rect 185044 215688 185050 215740
rect 92802 215620 92808 215672
rect 92860 215660 92866 215672
rect 100898 215660 100904 215672
rect 92860 215632 100904 215660
rect 92860 215620 92866 215632
rect 100898 215620 100904 215632
rect 100956 215620 100962 215672
rect 137606 215620 137612 215672
rect 137664 215660 137670 215672
rect 142942 215660 142948 215672
rect 137664 215632 142948 215660
rect 137664 215620 137670 215632
rect 142942 215620 142948 215632
rect 143000 215620 143006 215672
rect 177626 215620 177632 215672
rect 177684 215660 177690 215672
rect 185078 215660 185084 215672
rect 177684 215632 185084 215660
rect 177684 215620 177690 215632
rect 185078 215620 185084 215632
rect 185136 215620 185142 215672
rect 56462 215144 56468 215196
rect 56520 215184 56526 215196
rect 58210 215184 58216 215196
rect 56520 215156 58216 215184
rect 56520 215144 56526 215156
rect 58210 215144 58216 215156
rect 58268 215144 58274 215196
rect 50390 214872 50396 214924
rect 50448 214912 50454 214924
rect 52782 214912 52788 214924
rect 50448 214884 52788 214912
rect 50448 214872 50454 214884
rect 52782 214872 52788 214884
rect 52840 214872 52846 214924
rect 134846 214872 134852 214924
rect 134904 214912 134910 214924
rect 137606 214912 137612 214924
rect 134904 214884 137612 214912
rect 134904 214872 134910 214884
rect 137606 214872 137612 214884
rect 137664 214872 137670 214924
rect 51126 214532 51132 214584
rect 51184 214572 51190 214584
rect 52690 214572 52696 214584
rect 51184 214544 52696 214572
rect 51184 214532 51190 214544
rect 52690 214532 52696 214544
rect 52748 214532 52754 214584
rect 135306 214532 135312 214584
rect 135364 214572 135370 214584
rect 136870 214572 136876 214584
rect 135364 214544 136876 214572
rect 135364 214532 135370 214544
rect 136870 214532 136876 214544
rect 136928 214532 136934 214584
rect 51218 214464 51224 214516
rect 51276 214504 51282 214516
rect 58302 214504 58308 214516
rect 51276 214476 58308 214504
rect 51276 214464 51282 214476
rect 58302 214464 58308 214476
rect 58360 214464 58366 214516
rect 135398 214464 135404 214516
rect 135456 214504 135462 214516
rect 143678 214504 143684 214516
rect 135456 214476 143684 214504
rect 135456 214464 135462 214476
rect 143678 214464 143684 214476
rect 143736 214464 143742 214516
rect 51310 214396 51316 214448
rect 51368 214436 51374 214448
rect 58210 214436 58216 214448
rect 51368 214408 58216 214436
rect 51368 214396 51374 214408
rect 58210 214396 58216 214408
rect 58268 214396 58274 214448
rect 93354 214396 93360 214448
rect 93412 214436 93418 214448
rect 100990 214436 100996 214448
rect 93412 214408 100996 214436
rect 93412 214396 93418 214408
rect 100990 214396 100996 214408
rect 101048 214396 101054 214448
rect 134754 214396 134760 214448
rect 134812 214436 134818 214448
rect 135306 214436 135312 214448
rect 134812 214408 135312 214436
rect 134812 214396 134818 214408
rect 135306 214396 135312 214408
rect 135364 214396 135370 214448
rect 135490 214396 135496 214448
rect 135548 214436 135554 214448
rect 142942 214436 142948 214448
rect 135548 214408 142948 214436
rect 135548 214396 135554 214408
rect 142942 214396 142948 214408
rect 143000 214396 143006 214448
rect 177626 214396 177632 214448
rect 177684 214436 177690 214448
rect 185170 214436 185176 214448
rect 177684 214408 185176 214436
rect 177684 214396 177690 214408
rect 185170 214396 185176 214408
rect 185228 214396 185234 214448
rect 92710 214328 92716 214380
rect 92768 214368 92774 214380
rect 100714 214368 100720 214380
rect 92768 214340 100720 214368
rect 92768 214328 92774 214340
rect 100714 214328 100720 214340
rect 100772 214328 100778 214380
rect 177718 214328 177724 214380
rect 177776 214368 177782 214380
rect 184802 214368 184808 214380
rect 177776 214340 184808 214368
rect 177776 214328 177782 214340
rect 184802 214328 184808 214340
rect 184860 214328 184866 214380
rect 134478 213512 134484 213564
rect 134536 213552 134542 213564
rect 137054 213552 137060 213564
rect 134536 213524 137060 213552
rect 134536 213512 134542 213524
rect 137054 213512 137060 213524
rect 137112 213512 137118 213564
rect 51218 213376 51224 213428
rect 51276 213416 51282 213428
rect 52874 213416 52880 213428
rect 51276 213388 52880 213416
rect 51276 213376 51282 213388
rect 52874 213376 52880 213388
rect 52932 213376 52938 213428
rect 50390 213104 50396 213156
rect 50448 213144 50454 213156
rect 52966 213144 52972 213156
rect 50448 213116 52972 213144
rect 50448 213104 50454 213116
rect 52966 213104 52972 213116
rect 53024 213104 53030 213156
rect 134478 213104 134484 213156
rect 134536 213144 134542 213156
rect 136962 213144 136968 213156
rect 134536 213116 136968 213144
rect 134536 213104 134542 213116
rect 136962 213104 136968 213116
rect 137020 213104 137026 213156
rect 52782 213036 52788 213088
rect 52840 213076 52846 213088
rect 58210 213076 58216 213088
rect 52840 213048 58216 213076
rect 52840 213036 52846 213048
rect 58210 213036 58216 213048
rect 58268 213036 58274 213088
rect 93354 213036 93360 213088
rect 93412 213076 93418 213088
rect 100990 213076 100996 213088
rect 93412 213048 100996 213076
rect 93412 213036 93418 213048
rect 100990 213036 100996 213048
rect 101048 213036 101054 213088
rect 137606 213036 137612 213088
rect 137664 213076 137670 213088
rect 143678 213076 143684 213088
rect 137664 213048 143684 213076
rect 137664 213036 137670 213048
rect 143678 213036 143684 213048
rect 143736 213036 143742 213088
rect 177166 213036 177172 213088
rect 177224 213076 177230 213088
rect 185262 213076 185268 213088
rect 177224 213048 185268 213076
rect 177224 213036 177230 213048
rect 185262 213036 185268 213048
rect 185320 213036 185326 213088
rect 52690 212968 52696 213020
rect 52748 213008 52754 213020
rect 58302 213008 58308 213020
rect 52748 212980 58308 213008
rect 52748 212968 52754 212980
rect 58302 212968 58308 212980
rect 58360 212968 58366 213020
rect 92710 212968 92716 213020
rect 92768 213008 92774 213020
rect 100806 213008 100812 213020
rect 92768 212980 100812 213008
rect 92768 212968 92774 212980
rect 100806 212968 100812 212980
rect 100864 212968 100870 213020
rect 136870 212968 136876 213020
rect 136928 213008 136934 213020
rect 143494 213008 143500 213020
rect 136928 212980 143500 213008
rect 136928 212968 136934 212980
rect 143494 212968 143500 212980
rect 143552 212968 143558 213020
rect 177718 212968 177724 213020
rect 177776 213008 177782 213020
rect 184894 213008 184900 213020
rect 177776 212980 184900 213008
rect 177776 212968 177782 212980
rect 184894 212968 184900 212980
rect 184952 212968 184958 213020
rect 51126 212016 51132 212068
rect 51184 212056 51190 212068
rect 52690 212056 52696 212068
rect 51184 212028 52696 212056
rect 51184 212016 51190 212028
rect 52690 212016 52696 212028
rect 52748 212016 52754 212068
rect 97494 211948 97500 212000
rect 97552 211988 97558 212000
rect 100990 211988 100996 212000
rect 97552 211960 100996 211988
rect 97552 211948 97558 211960
rect 100990 211948 100996 211960
rect 101048 211948 101054 212000
rect 134478 211880 134484 211932
rect 134536 211920 134542 211932
rect 139630 211920 139636 211932
rect 134536 211892 139636 211920
rect 134536 211880 134542 211892
rect 139630 211880 139636 211892
rect 139688 211880 139694 211932
rect 51218 211744 51224 211796
rect 51276 211784 51282 211796
rect 56278 211784 56284 211796
rect 51276 211756 56284 211784
rect 51276 211744 51282 211756
rect 56278 211744 56284 211756
rect 56336 211744 56342 211796
rect 134662 211744 134668 211796
rect 134720 211784 134726 211796
rect 136870 211784 136876 211796
rect 134720 211756 136876 211784
rect 134720 211744 134726 211756
rect 136870 211744 136876 211756
rect 136928 211744 136934 211796
rect 181766 211676 181772 211728
rect 181824 211716 181830 211728
rect 185170 211716 185176 211728
rect 181824 211688 185176 211716
rect 181824 211676 181830 211688
rect 185170 211676 185176 211688
rect 185228 211676 185234 211728
rect 52966 211608 52972 211660
rect 53024 211648 53030 211660
rect 58210 211648 58216 211660
rect 53024 211620 58216 211648
rect 53024 211608 53030 211620
rect 58210 211608 58216 211620
rect 58268 211608 58274 211660
rect 92802 211608 92808 211660
rect 92860 211648 92866 211660
rect 100898 211648 100904 211660
rect 92860 211620 100904 211648
rect 92860 211608 92866 211620
rect 100898 211608 100904 211620
rect 100956 211608 100962 211660
rect 137054 211608 137060 211660
rect 137112 211648 137118 211660
rect 143678 211648 143684 211660
rect 137112 211620 143684 211648
rect 137112 211608 137118 211620
rect 143678 211608 143684 211620
rect 143736 211608 143742 211660
rect 177718 211608 177724 211660
rect 177776 211648 177782 211660
rect 184986 211648 184992 211660
rect 177776 211620 184992 211648
rect 177776 211608 177782 211620
rect 184986 211608 184992 211620
rect 185044 211608 185050 211660
rect 52874 211540 52880 211592
rect 52932 211580 52938 211592
rect 58302 211580 58308 211592
rect 52932 211552 58308 211580
rect 52932 211540 52938 211552
rect 58302 211540 58308 211552
rect 58360 211540 58366 211592
rect 92710 211540 92716 211592
rect 92768 211580 92774 211592
rect 100714 211580 100720 211592
rect 92768 211552 100720 211580
rect 92768 211540 92774 211552
rect 100714 211540 100720 211552
rect 100772 211540 100778 211592
rect 177166 211540 177172 211592
rect 177224 211580 177230 211592
rect 185078 211580 185084 211592
rect 177224 211552 185084 211580
rect 177224 211540 177230 211552
rect 185078 211540 185084 211552
rect 185136 211540 185142 211592
rect 92894 211472 92900 211524
rect 92952 211512 92958 211524
rect 97494 211512 97500 211524
rect 92952 211484 97500 211512
rect 92952 211472 92958 211484
rect 97494 211472 97500 211484
rect 97552 211472 97558 211524
rect 136962 211336 136968 211388
rect 137020 211376 137026 211388
rect 143678 211376 143684 211388
rect 137020 211348 143684 211376
rect 137020 211336 137026 211348
rect 143678 211336 143684 211348
rect 143736 211336 143742 211388
rect 56278 210996 56284 211048
rect 56336 211036 56342 211048
rect 58394 211036 58400 211048
rect 56336 211008 58400 211036
rect 56336 210996 56342 211008
rect 58394 210996 58400 211008
rect 58452 210996 58458 211048
rect 139630 210928 139636 210980
rect 139688 210968 139694 210980
rect 143586 210968 143592 210980
rect 139688 210940 143592 210968
rect 139688 210928 139694 210940
rect 143586 210928 143592 210940
rect 143644 210928 143650 210980
rect 177718 210792 177724 210844
rect 177776 210832 177782 210844
rect 181766 210832 181772 210844
rect 177776 210804 181772 210832
rect 177776 210792 177782 210804
rect 181766 210792 181772 210804
rect 181824 210792 181830 210844
rect 51218 210520 51224 210572
rect 51276 210560 51282 210572
rect 56094 210560 56100 210572
rect 51276 210532 56100 210560
rect 51276 210520 51282 210532
rect 56094 210520 56100 210532
rect 56152 210520 56158 210572
rect 93998 210384 94004 210436
rect 94056 210424 94062 210436
rect 101082 210424 101088 210436
rect 94056 210396 101088 210424
rect 94056 210384 94062 210396
rect 101082 210384 101088 210396
rect 101140 210384 101146 210436
rect 178178 210384 178184 210436
rect 178236 210424 178242 210436
rect 185262 210424 185268 210436
rect 178236 210396 185268 210424
rect 178236 210384 178242 210396
rect 185262 210384 185268 210396
rect 185320 210384 185326 210436
rect 92618 210316 92624 210368
rect 92676 210356 92682 210368
rect 100990 210356 100996 210368
rect 92676 210328 100996 210356
rect 92676 210316 92682 210328
rect 100990 210316 100996 210328
rect 101048 210316 101054 210368
rect 134570 210316 134576 210368
rect 134628 210356 134634 210368
rect 134628 210328 139676 210356
rect 134628 210316 134634 210328
rect 52690 210248 52696 210300
rect 52748 210288 52754 210300
rect 58210 210288 58216 210300
rect 52748 210260 58216 210288
rect 52748 210248 52754 210260
rect 58210 210248 58216 210260
rect 58268 210248 58274 210300
rect 93170 210248 93176 210300
rect 93228 210288 93234 210300
rect 101266 210288 101272 210300
rect 93228 210260 101272 210288
rect 93228 210248 93234 210260
rect 101266 210248 101272 210260
rect 101324 210248 101330 210300
rect 139648 210288 139676 210328
rect 176798 210316 176804 210368
rect 176856 210356 176862 210368
rect 185170 210356 185176 210368
rect 176856 210328 185176 210356
rect 176856 210316 176862 210328
rect 185170 210316 185176 210328
rect 185228 210316 185234 210368
rect 143678 210288 143684 210300
rect 139648 210260 143684 210288
rect 143678 210248 143684 210260
rect 143736 210248 143742 210300
rect 177166 210248 177172 210300
rect 177224 210288 177230 210300
rect 185446 210288 185452 210300
rect 177224 210260 185452 210288
rect 177224 210248 177230 210260
rect 185446 210248 185452 210260
rect 185504 210248 185510 210300
rect 92710 210180 92716 210232
rect 92768 210220 92774 210232
rect 101174 210220 101180 210232
rect 92768 210192 101180 210220
rect 92768 210180 92774 210192
rect 101174 210180 101180 210192
rect 101232 210180 101238 210232
rect 136870 210180 136876 210232
rect 136928 210220 136934 210232
rect 142942 210220 142948 210232
rect 136928 210192 142948 210220
rect 136928 210180 136934 210192
rect 142942 210180 142948 210192
rect 143000 210180 143006 210232
rect 177718 210180 177724 210232
rect 177776 210220 177782 210232
rect 185354 210220 185360 210232
rect 177776 210192 185360 210220
rect 177776 210180 177782 210192
rect 185354 210180 185360 210192
rect 185412 210180 185418 210232
rect 56094 209840 56100 209892
rect 56152 209880 56158 209892
rect 58302 209880 58308 209892
rect 56152 209852 58308 209880
rect 56152 209840 56158 209852
rect 58302 209840 58308 209852
rect 58360 209840 58366 209892
rect 83050 208956 83056 209008
rect 83108 208996 83114 209008
rect 84246 208996 84252 209008
rect 83108 208968 84252 208996
rect 83108 208956 83114 208968
rect 84246 208956 84252 208968
rect 84304 208956 84310 209008
rect 91238 208956 91244 209008
rect 91296 208996 91302 209008
rect 100990 208996 100996 209008
rect 91296 208968 100996 208996
rect 91296 208956 91302 208968
rect 100990 208956 100996 208968
rect 101048 208956 101054 209008
rect 175418 208956 175424 209008
rect 175476 208996 175482 209008
rect 185170 208996 185176 209008
rect 175476 208968 185176 208996
rect 175476 208956 175482 208968
rect 185170 208956 185176 208968
rect 185228 208956 185234 209008
rect 134202 207664 134208 207716
rect 134260 207704 134266 207716
rect 140274 207704 140280 207716
rect 134260 207676 140280 207704
rect 134260 207664 134266 207676
rect 140274 207664 140280 207676
rect 140332 207664 140338 207716
rect 50574 207460 50580 207512
rect 50632 207500 50638 207512
rect 61246 207500 61252 207512
rect 50632 207472 61252 207500
rect 50632 207460 50638 207472
rect 61246 207460 61252 207472
rect 61304 207460 61310 207512
rect 135306 207460 135312 207512
rect 135364 207500 135370 207512
rect 145334 207500 145340 207512
rect 135364 207472 145340 207500
rect 135364 207460 135370 207472
rect 145334 207460 145340 207472
rect 145392 207460 145398 207512
rect 174038 207460 174044 207512
rect 174096 207500 174102 207512
rect 180294 207500 180300 207512
rect 174096 207472 180300 207500
rect 174096 207460 174102 207472
rect 180294 207460 180300 207472
rect 180352 207460 180358 207512
rect 76794 206304 76800 206356
rect 76852 206344 76858 206356
rect 78358 206344 78364 206356
rect 76852 206316 78364 206344
rect 76852 206304 76858 206316
rect 78358 206304 78364 206316
rect 78416 206304 78422 206356
rect 73206 206236 73212 206288
rect 73264 206276 73270 206288
rect 75506 206276 75512 206288
rect 73264 206248 75512 206276
rect 73264 206236 73270 206248
rect 75506 206236 75512 206248
rect 75564 206236 75570 206288
rect 78174 206236 78180 206288
rect 78232 206276 78238 206288
rect 79738 206276 79744 206288
rect 78232 206248 79744 206276
rect 78232 206236 78238 206248
rect 79738 206236 79744 206248
rect 79796 206236 79802 206288
rect 157478 206236 157484 206288
rect 157536 206276 157542 206288
rect 159502 206276 159508 206288
rect 157536 206248 159508 206276
rect 157536 206236 157542 206248
rect 159502 206236 159508 206248
rect 159560 206236 159566 206288
rect 160974 206236 160980 206288
rect 161032 206276 161038 206288
rect 162446 206276 162452 206288
rect 161032 206248 162452 206276
rect 161032 206236 161038 206248
rect 162446 206236 162452 206248
rect 162504 206236 162510 206288
rect 73298 206168 73304 206220
rect 73356 206208 73362 206220
rect 74034 206208 74040 206220
rect 73356 206180 74040 206208
rect 73356 206168 73362 206180
rect 74034 206168 74040 206180
rect 74092 206168 74098 206220
rect 74678 206168 74684 206220
rect 74736 206208 74742 206220
rect 76886 206208 76892 206220
rect 74736 206180 76892 206208
rect 74736 206168 74742 206180
rect 76886 206168 76892 206180
rect 76944 206168 76950 206220
rect 79554 206168 79560 206220
rect 79612 206208 79618 206220
rect 81210 206208 81216 206220
rect 79612 206180 81216 206208
rect 79612 206168 79618 206180
rect 81210 206168 81216 206180
rect 81268 206168 81274 206220
rect 85718 206168 85724 206220
rect 85776 206208 85782 206220
rect 100990 206208 100996 206220
rect 85776 206180 100996 206208
rect 85776 206168 85782 206180
rect 100990 206168 100996 206180
rect 101048 206168 101054 206220
rect 147266 206168 147272 206220
rect 147324 206208 147330 206220
rect 147818 206208 147824 206220
rect 147324 206180 147824 206208
rect 147324 206168 147330 206180
rect 147818 206168 147824 206180
rect 147876 206168 147882 206220
rect 156834 206168 156840 206220
rect 156892 206208 156898 206220
rect 158030 206208 158036 206220
rect 156892 206180 158036 206208
rect 156892 206168 156898 206180
rect 158030 206168 158036 206180
rect 158088 206168 158094 206220
rect 158858 206168 158864 206220
rect 158916 206208 158922 206220
rect 160882 206208 160888 206220
rect 158916 206180 160888 206208
rect 158916 206168 158922 206180
rect 160882 206168 160888 206180
rect 160940 206168 160946 206220
rect 162354 206168 162360 206220
rect 162412 206208 162418 206220
rect 163734 206208 163740 206220
rect 162412 206180 163740 206208
rect 162412 206168 162418 206180
rect 163734 206168 163740 206180
rect 163792 206168 163798 206220
rect 169898 206168 169904 206220
rect 169956 206208 169962 206220
rect 185170 206208 185176 206220
rect 169956 206180 185176 206208
rect 169956 206168 169962 206180
rect 185170 206168 185176 206180
rect 185228 206168 185234 206220
rect 216174 204808 216180 204860
rect 216232 204848 216238 204860
rect 222338 204848 222344 204860
rect 216232 204820 222344 204848
rect 216232 204808 216238 204820
rect 222338 204808 222344 204820
rect 222396 204808 222402 204860
rect 148738 204740 148744 204792
rect 148796 204780 148802 204792
rect 215530 204780 215536 204792
rect 148796 204752 215536 204780
rect 148796 204740 148802 204752
rect 215530 204740 215536 204752
rect 215588 204740 215594 204792
rect 24078 204672 24084 204724
rect 24136 204712 24142 204724
rect 28126 204712 28132 204724
rect 24136 204684 28132 204712
rect 24136 204672 24142 204684
rect 28126 204672 28132 204684
rect 28184 204672 28190 204724
rect 21502 204604 21508 204656
rect 21560 204644 21566 204656
rect 26930 204644 26936 204656
rect 21560 204616 26936 204644
rect 21560 204604 21566 204616
rect 26930 204604 26936 204616
rect 26988 204604 26994 204656
rect 22790 204536 22796 204588
rect 22848 204576 22854 204588
rect 26838 204576 26844 204588
rect 22848 204548 26844 204576
rect 22848 204536 22854 204548
rect 26838 204536 26844 204548
rect 26896 204536 26902 204588
rect 121414 204536 121420 204588
rect 121472 204576 121478 204588
rect 123162 204576 123168 204588
rect 121472 204548 123168 204576
rect 121472 204536 121478 204548
rect 123162 204536 123168 204548
rect 123220 204536 123226 204588
rect 208538 204536 208544 204588
rect 208596 204576 208602 204588
rect 211114 204576 211120 204588
rect 208596 204548 211120 204576
rect 208596 204536 208602 204548
rect 211114 204536 211120 204548
rect 211172 204536 211178 204588
rect 23434 204468 23440 204520
rect 23492 204508 23498 204520
rect 26746 204508 26752 204520
rect 23492 204480 26752 204508
rect 23492 204468 23498 204480
rect 26746 204468 26752 204480
rect 26804 204468 26810 204520
rect 45054 204400 45060 204452
rect 45112 204440 45118 204452
rect 45882 204440 45888 204452
rect 45112 204412 45888 204440
rect 45112 204400 45118 204412
rect 45882 204400 45888 204412
rect 45940 204400 45946 204452
rect 98966 204400 98972 204452
rect 99024 204440 99030 204452
rect 104762 204440 104768 204452
rect 99024 204412 104768 204440
rect 99024 204400 99030 204412
rect 104762 204400 104768 204412
rect 104820 204400 104826 204452
rect 121598 204400 121604 204452
rect 121656 204440 121662 204452
rect 123714 204440 123720 204452
rect 121656 204412 123720 204440
rect 121656 204400 121662 204412
rect 123714 204400 123720 204412
rect 123772 204400 123778 204452
rect 207894 204400 207900 204452
rect 207952 204440 207958 204452
rect 210562 204440 210568 204452
rect 207952 204412 210568 204440
rect 207952 204400 207958 204412
rect 210562 204400 210568 204412
rect 210620 204400 210626 204452
rect 24722 204332 24728 204384
rect 24780 204372 24786 204384
rect 28034 204372 28040 204384
rect 24780 204344 28040 204372
rect 24780 204332 24786 204344
rect 28034 204332 28040 204344
rect 28092 204332 28098 204384
rect 120126 204332 120132 204384
rect 120184 204372 120190 204384
rect 121506 204372 121512 204384
rect 120184 204344 121512 204372
rect 120184 204332 120190 204344
rect 121506 204332 121512 204344
rect 121564 204332 121570 204384
rect 200258 204332 200264 204384
rect 200316 204372 200322 204384
rect 200994 204372 201000 204384
rect 200316 204344 201000 204372
rect 200316 204332 200322 204344
rect 200994 204332 201000 204344
rect 201052 204332 201058 204384
rect 22146 204264 22152 204316
rect 22204 204304 22210 204316
rect 26654 204304 26660 204316
rect 22204 204276 26660 204304
rect 22204 204264 22210 204276
rect 26654 204264 26660 204276
rect 26712 204264 26718 204316
rect 99426 204264 99432 204316
rect 99484 204304 99490 204316
rect 107522 204304 107528 204316
rect 99484 204276 107528 204304
rect 99484 204264 99490 204276
rect 107522 204264 107528 204276
rect 107580 204264 107586 204316
rect 208078 204264 208084 204316
rect 208136 204304 208142 204316
rect 210010 204304 210016 204316
rect 208136 204276 210016 204304
rect 208136 204264 208142 204276
rect 210010 204264 210016 204276
rect 210068 204264 210074 204316
rect 121506 204196 121512 204248
rect 121564 204236 121570 204248
rect 124266 204236 124272 204248
rect 121564 204208 124272 204236
rect 121564 204196 121570 204208
rect 124266 204196 124272 204208
rect 124324 204196 124330 204248
rect 183606 204196 183612 204248
rect 183664 204236 183670 204248
rect 191518 204236 191524 204248
rect 183664 204208 191524 204236
rect 183664 204196 183670 204208
rect 191518 204196 191524 204208
rect 191576 204196 191582 204248
rect 208446 204196 208452 204248
rect 208504 204236 208510 204248
rect 211666 204236 211672 204248
rect 208504 204208 211672 204236
rect 208504 204196 208510 204208
rect 211666 204196 211672 204208
rect 211724 204196 211730 204248
rect 99242 204128 99248 204180
rect 99300 204168 99306 204180
rect 106970 204168 106976 204180
rect 99300 204140 106976 204168
rect 99300 204128 99306 204140
rect 106970 204128 106976 204140
rect 107028 204128 107034 204180
rect 183698 204128 183704 204180
rect 183756 204168 183762 204180
rect 192070 204168 192076 204180
rect 183756 204140 192076 204168
rect 183756 204128 183762 204140
rect 192070 204128 192076 204140
rect 192128 204128 192134 204180
rect 208354 204128 208360 204180
rect 208412 204168 208418 204180
rect 212218 204168 212224 204180
rect 208412 204140 212224 204168
rect 208412 204128 208418 204140
rect 212218 204128 212224 204140
rect 212276 204128 212282 204180
rect 20214 204060 20220 204112
rect 20272 204100 20278 204112
rect 41742 204100 41748 204112
rect 20272 204072 41748 204100
rect 20272 204060 20278 204072
rect 41742 204060 41748 204072
rect 41800 204060 41806 204112
rect 99518 204060 99524 204112
rect 99576 204100 99582 204112
rect 108074 204100 108080 204112
rect 99576 204072 108080 204100
rect 99576 204060 99582 204072
rect 108074 204060 108080 204072
rect 108132 204060 108138 204112
rect 183422 204060 183428 204112
rect 183480 204100 183486 204112
rect 190966 204100 190972 204112
rect 183480 204072 190972 204100
rect 183480 204060 183486 204072
rect 190966 204060 190972 204072
rect 191024 204060 191030 204112
rect 191978 204060 191984 204112
rect 192036 204100 192042 204112
rect 214978 204100 214984 204112
rect 192036 204072 214984 204100
rect 192036 204060 192042 204072
rect 214978 204060 214984 204072
rect 215036 204060 215042 204112
rect 99150 203788 99156 203840
rect 99208 203828 99214 203840
rect 106418 203828 106424 203840
rect 99208 203800 106424 203828
rect 99208 203788 99214 203800
rect 106418 203788 106424 203800
rect 106476 203788 106482 203840
rect 117458 203788 117464 203840
rect 117516 203828 117522 203840
rect 118746 203828 118752 203840
rect 117516 203800 118752 203828
rect 117516 203788 117522 203800
rect 118746 203788 118752 203800
rect 118804 203788 118810 203840
rect 124266 203788 124272 203840
rect 124324 203828 124330 203840
rect 128222 203828 128228 203840
rect 124324 203800 128228 203828
rect 124324 203788 124330 203800
rect 128222 203788 128228 203800
rect 128280 203788 128286 203840
rect 123714 203720 123720 203772
rect 123772 203760 123778 203772
rect 125462 203760 125468 203772
rect 123772 203732 125468 203760
rect 123772 203720 123778 203732
rect 125462 203720 125468 203732
rect 125520 203720 125526 203772
rect 205686 203720 205692 203772
rect 205744 203760 205750 203772
rect 208814 203760 208820 203772
rect 205744 203732 208820 203760
rect 205744 203720 205750 203732
rect 208814 203720 208820 203732
rect 208872 203720 208878 203772
rect 110282 203652 110288 203704
rect 110340 203692 110346 203704
rect 111018 203692 111024 203704
rect 110340 203664 111024 203692
rect 110340 203652 110346 203664
rect 111018 203652 111024 203664
rect 111076 203652 111082 203704
rect 118746 203652 118752 203704
rect 118804 203692 118810 203704
rect 120954 203692 120960 203704
rect 118804 203664 120960 203692
rect 118804 203652 118810 203664
rect 120954 203652 120960 203664
rect 121012 203652 121018 203704
rect 123898 203652 123904 203704
rect 123956 203692 123962 203704
rect 126566 203692 126572 203704
rect 123956 203664 126572 203692
rect 123956 203652 123962 203664
rect 126566 203652 126572 203664
rect 126624 203652 126630 203704
rect 183330 203652 183336 203704
rect 183388 203692 183394 203704
rect 189862 203692 189868 203704
rect 183388 203664 189868 203692
rect 183388 203652 183394 203664
rect 189862 203652 189868 203664
rect 189920 203652 189926 203704
rect 204306 203652 204312 203704
rect 204364 203692 204370 203704
rect 206606 203692 206612 203704
rect 204364 203664 206612 203692
rect 204364 203652 204370 203664
rect 206606 203652 206612 203664
rect 206664 203652 206670 203704
rect 99334 203584 99340 203636
rect 99392 203624 99398 203636
rect 105866 203624 105872 203636
rect 99392 203596 105872 203624
rect 99392 203584 99398 203596
rect 105866 203584 105872 203596
rect 105924 203584 105930 203636
rect 124174 203584 124180 203636
rect 124232 203624 124238 203636
rect 127118 203624 127124 203636
rect 124232 203596 127124 203624
rect 124232 203584 124238 203596
rect 127118 203584 127124 203596
rect 127176 203584 127182 203636
rect 127946 203584 127952 203636
rect 128004 203624 128010 203636
rect 130430 203624 130436 203636
rect 128004 203596 130436 203624
rect 128004 203584 128010 203596
rect 130430 203584 130436 203596
rect 130488 203584 130494 203636
rect 183238 203584 183244 203636
rect 183296 203624 183302 203636
rect 189310 203624 189316 203636
rect 183296 203596 189316 203624
rect 183296 203584 183302 203596
rect 189310 203584 189316 203596
rect 189368 203584 189374 203636
rect 201454 203584 201460 203636
rect 201512 203624 201518 203636
rect 203294 203624 203300 203636
rect 201512 203596 203300 203624
rect 201512 203584 201518 203596
rect 203294 203584 203300 203596
rect 203352 203584 203358 203636
rect 204214 203584 204220 203636
rect 204272 203624 204278 203636
rect 206054 203624 206060 203636
rect 204272 203596 206060 203624
rect 204272 203584 204278 203596
rect 206054 203584 206060 203596
rect 206112 203584 206118 203636
rect 40914 203516 40920 203568
rect 40972 203556 40978 203568
rect 43030 203556 43036 203568
rect 40972 203528 43036 203556
rect 40972 203516 40978 203528
rect 43030 203516 43036 203528
rect 43088 203516 43094 203568
rect 99058 203516 99064 203568
rect 99116 203556 99122 203568
rect 105314 203556 105320 203568
rect 99116 203528 105320 203556
rect 99116 203516 99122 203528
rect 105314 203516 105320 203528
rect 105372 203516 105378 203568
rect 109270 203516 109276 203568
rect 109328 203556 109334 203568
rect 110282 203556 110288 203568
rect 109328 203528 110288 203556
rect 109328 203516 109334 203528
rect 110282 203516 110288 203528
rect 110340 203516 110346 203568
rect 116354 203516 116360 203568
rect 116412 203556 116418 203568
rect 117550 203556 117556 203568
rect 116412 203528 117556 203556
rect 116412 203516 116418 203528
rect 117550 203516 117556 203528
rect 117608 203516 117614 203568
rect 118838 203516 118844 203568
rect 118896 203556 118902 203568
rect 120402 203556 120408 203568
rect 118896 203528 120408 203556
rect 118896 203516 118902 203528
rect 120402 203516 120408 203528
rect 120460 203516 120466 203568
rect 123990 203516 123996 203568
rect 124048 203556 124054 203568
rect 126014 203556 126020 203568
rect 124048 203528 126020 203556
rect 124048 203516 124054 203528
rect 126014 203516 126020 203528
rect 126072 203516 126078 203568
rect 127854 203516 127860 203568
rect 127912 203556 127918 203568
rect 128774 203556 128780 203568
rect 127912 203528 128780 203556
rect 127912 203516 127918 203528
rect 128774 203516 128780 203528
rect 128832 203516 128838 203568
rect 183146 203516 183152 203568
rect 183204 203556 183210 203568
rect 188758 203556 188764 203568
rect 183204 203528 188764 203556
rect 183204 203516 183210 203528
rect 188758 203516 188764 203528
rect 188816 203516 188822 203568
rect 202926 203516 202932 203568
rect 202984 203556 202990 203568
rect 204398 203556 204404 203568
rect 202984 203528 204404 203556
rect 202984 203516 202990 203528
rect 204398 203516 204404 203528
rect 204456 203516 204462 203568
rect 205778 203516 205784 203568
rect 205836 203556 205842 203568
rect 208262 203556 208268 203568
rect 205836 203528 208268 203556
rect 205836 203516 205842 203528
rect 208262 203516 208268 203528
rect 208320 203516 208326 203568
rect 20858 203448 20864 203500
rect 20916 203488 20922 203500
rect 25458 203488 25464 203500
rect 20916 203460 25464 203488
rect 20916 203448 20922 203460
rect 25458 203448 25464 203460
rect 25516 203448 25522 203500
rect 41098 203448 41104 203500
rect 41156 203488 41162 203500
rect 42294 203488 42300 203500
rect 41156 203460 42300 203488
rect 41156 203448 41162 203460
rect 42294 203448 42300 203460
rect 42352 203448 42358 203500
rect 43766 203448 43772 203500
rect 43824 203488 43830 203500
rect 44870 203488 44876 203500
rect 43824 203460 44876 203488
rect 43824 203448 43830 203460
rect 44870 203448 44876 203460
rect 44928 203448 44934 203500
rect 98874 203448 98880 203500
rect 98932 203488 98938 203500
rect 104210 203488 104216 203500
rect 98932 203460 104216 203488
rect 98932 203448 98938 203460
rect 104210 203448 104216 203460
rect 104268 203448 104274 203500
rect 116078 203448 116084 203500
rect 116136 203488 116142 203500
rect 116998 203488 117004 203500
rect 116136 203460 117004 203488
rect 116136 203448 116142 203460
rect 116998 203448 117004 203460
rect 117056 203448 117062 203500
rect 117642 203448 117648 203500
rect 117700 203488 117706 203500
rect 117700 203460 118332 203488
rect 117700 203448 117706 203460
rect 25366 203380 25372 203432
rect 25424 203420 25430 203432
rect 26102 203420 26108 203432
rect 25424 203392 26108 203420
rect 25424 203380 25430 203392
rect 26102 203380 26108 203392
rect 26160 203380 26166 203432
rect 27206 203380 27212 203432
rect 27264 203420 27270 203432
rect 27666 203420 27672 203432
rect 27264 203392 27672 203420
rect 27264 203380 27270 203392
rect 27666 203380 27672 203392
rect 27724 203380 27730 203432
rect 28586 203380 28592 203432
rect 28644 203420 28650 203432
rect 29138 203420 29144 203432
rect 28644 203392 29144 203420
rect 28644 203380 28650 203392
rect 29138 203380 29144 203392
rect 29196 203380 29202 203432
rect 29966 203380 29972 203432
rect 30024 203420 30030 203432
rect 30518 203420 30524 203432
rect 30024 203392 30524 203420
rect 30024 203380 30030 203392
rect 30518 203380 30524 203392
rect 30576 203380 30582 203432
rect 31254 203380 31260 203432
rect 31312 203420 31318 203432
rect 31806 203420 31812 203432
rect 31312 203392 31812 203420
rect 31312 203380 31318 203392
rect 31806 203380 31812 203392
rect 31864 203380 31870 203432
rect 37418 203380 37424 203432
rect 37476 203420 37482 203432
rect 38430 203420 38436 203432
rect 37476 203392 38436 203420
rect 37476 203380 37482 203392
rect 38430 203380 38436 203392
rect 38488 203380 38494 203432
rect 39534 203380 39540 203432
rect 39592 203420 39598 203432
rect 40362 203420 40368 203432
rect 39592 203392 40368 203420
rect 39592 203380 39598 203392
rect 40362 203380 40368 203392
rect 40420 203380 40426 203432
rect 41006 203380 41012 203432
rect 41064 203420 41070 203432
rect 41650 203420 41656 203432
rect 41064 203392 41656 203420
rect 41064 203380 41070 203392
rect 41650 203380 41656 203392
rect 41708 203380 41714 203432
rect 43674 203380 43680 203432
rect 43732 203420 43738 203432
rect 44410 203420 44416 203432
rect 43732 203392 44416 203420
rect 43732 203380 43738 203392
rect 44410 203380 44416 203392
rect 44468 203380 44474 203432
rect 108626 203380 108632 203432
rect 108684 203420 108690 203432
rect 109270 203420 109276 203432
rect 108684 203392 109276 203420
rect 108684 203380 108690 203392
rect 109270 203380 109276 203392
rect 109328 203380 109334 203432
rect 109730 203380 109736 203432
rect 109788 203420 109794 203432
rect 110742 203420 110748 203432
rect 109788 203392 110748 203420
rect 109788 203380 109794 203392
rect 110742 203380 110748 203392
rect 110800 203380 110806 203432
rect 111478 203380 111484 203432
rect 111536 203420 111542 203432
rect 112306 203420 112312 203432
rect 111536 203392 112312 203420
rect 111536 203380 111542 203392
rect 112306 203380 112312 203392
rect 112364 203380 112370 203432
rect 114606 203380 114612 203432
rect 114664 203420 114670 203432
rect 114790 203420 114796 203432
rect 114664 203392 114796 203420
rect 114664 203380 114670 203392
rect 114790 203380 114796 203392
rect 114848 203380 114854 203432
rect 115986 203380 115992 203432
rect 116044 203420 116050 203432
rect 116446 203420 116452 203432
rect 116044 203392 116452 203420
rect 116044 203380 116050 203392
rect 116446 203380 116452 203392
rect 116504 203380 116510 203432
rect 117366 203380 117372 203432
rect 117424 203420 117430 203432
rect 118194 203420 118200 203432
rect 117424 203392 118200 203420
rect 117424 203380 117430 203392
rect 118194 203380 118200 203392
rect 118252 203380 118258 203432
rect 118304 203420 118332 203460
rect 118654 203448 118660 203500
rect 118712 203488 118718 203500
rect 119850 203488 119856 203500
rect 118712 203460 119856 203488
rect 118712 203448 118718 203460
rect 119850 203448 119856 203460
rect 119908 203448 119914 203500
rect 120034 203448 120040 203500
rect 120092 203488 120098 203500
rect 122058 203488 122064 203500
rect 120092 203460 122064 203488
rect 120092 203448 120098 203460
rect 122058 203448 122064 203460
rect 122116 203448 122122 203500
rect 123806 203448 123812 203500
rect 123864 203488 123870 203500
rect 124818 203488 124824 203500
rect 123864 203460 124824 203488
rect 123864 203448 123870 203460
rect 124818 203448 124824 203460
rect 124876 203448 124882 203500
rect 128130 203448 128136 203500
rect 128188 203488 128194 203500
rect 129878 203488 129884 203500
rect 128188 203460 129884 203488
rect 128188 203448 128194 203460
rect 129878 203448 129884 203460
rect 129936 203448 129942 203500
rect 183054 203448 183060 203500
rect 183112 203488 183118 203500
rect 188206 203488 188212 203500
rect 183112 203460 188212 203488
rect 183112 203448 183118 203460
rect 188206 203448 188212 203460
rect 188264 203448 188270 203500
rect 203018 203448 203024 203500
rect 203076 203488 203082 203500
rect 204950 203488 204956 203500
rect 203076 203460 204956 203488
rect 203076 203448 203082 203460
rect 204950 203448 204956 203460
rect 205008 203448 205014 203500
rect 205410 203448 205416 203500
rect 205468 203488 205474 203500
rect 207158 203488 207164 203500
rect 205468 203460 207164 203488
rect 205468 203448 205474 203460
rect 207158 203448 207164 203460
rect 207216 203448 207222 203500
rect 119298 203420 119304 203432
rect 118304 203392 119304 203420
rect 119298 203380 119304 203392
rect 119356 203380 119362 203432
rect 120218 203380 120224 203432
rect 120276 203420 120282 203432
rect 122610 203420 122616 203432
rect 120276 203392 122616 203420
rect 120276 203380 120282 203392
rect 122610 203380 122616 203392
rect 122668 203380 122674 203432
rect 124358 203380 124364 203432
rect 124416 203420 124422 203432
rect 127670 203420 127676 203432
rect 124416 203392 127676 203420
rect 124416 203380 124422 203392
rect 127670 203380 127676 203392
rect 127728 203380 127734 203432
rect 128038 203380 128044 203432
rect 128096 203420 128102 203432
rect 129326 203420 129332 203432
rect 128096 203392 129332 203420
rect 128096 203380 128102 203392
rect 129326 203380 129332 203392
rect 129384 203380 129390 203432
rect 183514 203380 183520 203432
rect 183572 203420 183578 203432
rect 190414 203420 190420 203432
rect 183572 203392 190420 203420
rect 183572 203380 183578 203392
rect 190414 203380 190420 203392
rect 190472 203380 190478 203432
rect 192622 203380 192628 203432
rect 192680 203420 192686 203432
rect 193358 203420 193364 203432
rect 192680 203392 193364 203420
rect 192680 203380 192686 203392
rect 193358 203380 193364 203392
rect 193416 203380 193422 203432
rect 193726 203380 193732 203432
rect 193784 203420 193790 203432
rect 194738 203420 194744 203432
rect 193784 203392 194744 203420
rect 193784 203380 193790 203392
rect 194738 203380 194744 203392
rect 194796 203380 194802 203432
rect 201546 203380 201552 203432
rect 201604 203420 201610 203432
rect 202742 203420 202748 203432
rect 201604 203392 202748 203420
rect 201604 203380 201610 203392
rect 202742 203380 202748 203392
rect 202800 203380 202806 203432
rect 202834 203380 202840 203432
rect 202892 203420 202898 203432
rect 203846 203420 203852 203432
rect 202892 203392 203852 203420
rect 202892 203380 202898 203392
rect 203846 203380 203852 203392
rect 203904 203380 203910 203432
rect 204398 203380 204404 203432
rect 204456 203420 204462 203432
rect 205502 203420 205508 203432
rect 204456 203392 205508 203420
rect 204456 203380 204462 203392
rect 205502 203380 205508 203392
rect 205560 203380 205566 203432
rect 205594 203380 205600 203432
rect 205652 203420 205658 203432
rect 207710 203420 207716 203432
rect 205652 203392 207716 203420
rect 205652 203380 205658 203392
rect 207710 203380 207716 203392
rect 207768 203380 207774 203432
rect 207986 203380 207992 203432
rect 208044 203420 208050 203432
rect 209458 203420 209464 203432
rect 208044 203392 209464 203420
rect 208044 203380 208050 203392
rect 209458 203380 209464 203392
rect 209516 203380 209522 203432
rect 213414 203380 213420 203432
rect 213472 203420 213478 203432
rect 214426 203420 214432 203432
rect 213472 203392 214432 203420
rect 213472 203380 213478 203392
rect 214426 203380 214432 203392
rect 214484 203380 214490 203432
rect 33370 203040 33376 203092
rect 33428 203080 33434 203092
rect 33830 203080 33836 203092
rect 33428 203052 33836 203080
rect 33428 203040 33434 203052
rect 33830 203040 33836 203052
rect 33888 203040 33894 203092
rect 212862 203040 212868 203092
rect 212920 203080 212926 203092
rect 213046 203080 213052 203092
rect 212920 203052 213052 203080
rect 212920 203040 212926 203052
rect 213046 203040 213052 203052
rect 213104 203040 213110 203092
rect 197498 202836 197504 202888
rect 197556 202876 197562 202888
rect 197774 202876 197780 202888
rect 197556 202848 197780 202876
rect 197556 202836 197562 202848
rect 197774 202836 197780 202848
rect 197832 202836 197838 202888
rect 196210 201408 196216 201460
rect 196268 201448 196274 201460
rect 196854 201448 196860 201460
rect 196268 201420 196860 201448
rect 196268 201408 196274 201420
rect 196854 201408 196860 201420
rect 196912 201408 196918 201460
rect 50482 196444 50488 196496
rect 50540 196484 50546 196496
rect 57566 196484 57572 196496
rect 50540 196456 57572 196484
rect 50540 196444 50546 196456
rect 57566 196444 57572 196456
rect 57624 196444 57630 196496
rect 110834 196444 110840 196496
rect 110892 196484 110898 196496
rect 111662 196484 111668 196496
rect 110892 196456 111668 196484
rect 110892 196444 110898 196456
rect 111662 196444 111668 196456
rect 111720 196444 111726 196496
rect 112030 196444 112036 196496
rect 112088 196484 112094 196496
rect 112490 196484 112496 196496
rect 112088 196456 112496 196484
rect 112088 196444 112094 196456
rect 112490 196444 112496 196456
rect 112548 196444 112554 196496
rect 114882 196444 114888 196496
rect 114940 196484 114946 196496
rect 115342 196484 115348 196496
rect 114940 196456 115348 196484
rect 114940 196444 114946 196456
rect 115342 196444 115348 196456
rect 115400 196444 115406 196496
rect 123622 196444 123628 196496
rect 123680 196484 123686 196496
rect 124358 196484 124364 196496
rect 123680 196456 124364 196484
rect 123680 196444 123686 196456
rect 124358 196444 124364 196456
rect 124416 196444 124422 196496
rect 26746 196376 26752 196428
rect 26804 196416 26810 196428
rect 27390 196416 27396 196428
rect 26804 196388 27396 196416
rect 26804 196376 26810 196388
rect 27390 196376 27396 196388
rect 27448 196376 27454 196428
rect 27758 196376 27764 196428
rect 27816 196416 27822 196428
rect 30150 196416 30156 196428
rect 27816 196388 30156 196416
rect 27816 196376 27822 196388
rect 30150 196376 30156 196388
rect 30208 196376 30214 196428
rect 72010 196376 72016 196428
rect 72068 196416 72074 196428
rect 73298 196416 73304 196428
rect 72068 196388 73304 196416
rect 72068 196376 72074 196388
rect 73298 196376 73304 196388
rect 73356 196376 73362 196428
rect 115250 196376 115256 196428
rect 115308 196416 115314 196428
rect 115894 196416 115900 196428
rect 115308 196388 115900 196416
rect 115308 196376 115314 196388
rect 115894 196376 115900 196388
rect 115952 196376 115958 196428
rect 120862 196376 120868 196428
rect 120920 196416 120926 196428
rect 121598 196416 121604 196428
rect 120920 196388 121604 196416
rect 120920 196376 120926 196388
rect 121598 196376 121604 196388
rect 121656 196376 121662 196428
rect 121690 196376 121696 196428
rect 121748 196416 121754 196428
rect 123806 196416 123812 196428
rect 121748 196388 123812 196416
rect 121748 196376 121754 196388
rect 123806 196376 123812 196388
rect 123864 196376 123870 196428
rect 135306 196376 135312 196428
rect 135364 196416 135370 196428
rect 140458 196416 140464 196428
rect 135364 196388 140464 196416
rect 135364 196376 135370 196388
rect 140458 196376 140464 196388
rect 140516 196376 140522 196428
rect 196302 196376 196308 196428
rect 196360 196416 196366 196428
rect 196854 196416 196860 196428
rect 196360 196388 196860 196416
rect 196360 196376 196366 196388
rect 196854 196376 196860 196388
rect 196912 196376 196918 196428
rect 200810 196376 200816 196428
rect 200868 196416 200874 196428
rect 201638 196416 201644 196428
rect 200868 196388 201644 196416
rect 200868 196376 200874 196388
rect 201638 196376 201644 196388
rect 201696 196376 201702 196428
rect 203662 196376 203668 196428
rect 203720 196416 203726 196428
rect 204214 196416 204220 196428
rect 203720 196388 204220 196416
rect 203720 196376 203726 196388
rect 204214 196376 204220 196388
rect 204272 196376 204278 196428
rect 204490 196376 204496 196428
rect 204548 196416 204554 196428
rect 205502 196416 205508 196428
rect 204548 196388 205508 196416
rect 204548 196376 204554 196388
rect 205502 196376 205508 196388
rect 205560 196376 205566 196428
rect 26562 196308 26568 196360
rect 26620 196348 26626 196360
rect 26930 196348 26936 196360
rect 26620 196320 26936 196348
rect 26620 196308 26626 196320
rect 26930 196308 26936 196320
rect 26988 196308 26994 196360
rect 28034 196308 28040 196360
rect 28092 196348 28098 196360
rect 28218 196348 28224 196360
rect 28092 196320 28224 196348
rect 28092 196308 28098 196320
rect 28218 196308 28224 196320
rect 28276 196308 28282 196360
rect 38430 196308 38436 196360
rect 38488 196348 38494 196360
rect 39534 196348 39540 196360
rect 38488 196320 39540 196348
rect 38488 196308 38494 196320
rect 39534 196308 39540 196320
rect 39592 196308 39598 196360
rect 40086 196308 40092 196360
rect 40144 196348 40150 196360
rect 40914 196348 40920 196360
rect 40144 196320 40920 196348
rect 40144 196308 40150 196320
rect 40914 196308 40920 196320
rect 40972 196308 40978 196360
rect 41650 196308 41656 196360
rect 41708 196348 41714 196360
rect 45054 196348 45060 196360
rect 41708 196320 45060 196348
rect 41708 196308 41714 196320
rect 45054 196308 45060 196320
rect 45112 196308 45118 196360
rect 69802 196308 69808 196360
rect 69860 196348 69866 196360
rect 70630 196348 70636 196360
rect 69860 196320 70636 196348
rect 69860 196308 69866 196320
rect 70630 196308 70636 196320
rect 70688 196308 70694 196360
rect 70906 196308 70912 196360
rect 70964 196348 70970 196360
rect 72194 196348 72200 196360
rect 70964 196320 72200 196348
rect 70964 196308 70970 196320
rect 72194 196308 72200 196320
rect 72252 196308 72258 196360
rect 75322 196308 75328 196360
rect 75380 196348 75386 196360
rect 76794 196348 76800 196360
rect 75380 196320 76800 196348
rect 75380 196308 75386 196320
rect 76794 196308 76800 196320
rect 76852 196308 76858 196360
rect 78634 196308 78640 196360
rect 78692 196348 78698 196360
rect 81670 196348 81676 196360
rect 78692 196320 81676 196348
rect 78692 196308 78698 196320
rect 81670 196308 81676 196320
rect 81728 196308 81734 196360
rect 93078 196308 93084 196360
rect 93136 196348 93142 196360
rect 93998 196348 94004 196360
rect 93136 196320 94004 196348
rect 93136 196308 93142 196320
rect 93998 196308 94004 196320
rect 94056 196308 94062 196360
rect 119666 196308 119672 196360
rect 119724 196348 119730 196360
rect 120034 196348 120040 196360
rect 119724 196320 120040 196348
rect 119724 196308 119730 196320
rect 120034 196308 120040 196320
rect 120092 196308 120098 196360
rect 120494 196308 120500 196360
rect 120552 196348 120558 196360
rect 121414 196348 121420 196360
rect 120552 196320 121420 196348
rect 120552 196308 120558 196320
rect 121414 196308 121420 196320
rect 121472 196308 121478 196360
rect 123254 196308 123260 196360
rect 123312 196348 123318 196360
rect 124174 196348 124180 196360
rect 123312 196320 124180 196348
rect 123312 196308 123318 196320
rect 124174 196308 124180 196320
rect 124232 196308 124238 196360
rect 140274 196308 140280 196360
rect 140332 196348 140338 196360
rect 141562 196348 141568 196360
rect 140332 196320 141568 196348
rect 140332 196308 140338 196320
rect 141562 196308 141568 196320
rect 141620 196308 141626 196360
rect 152602 196308 152608 196360
rect 152660 196348 152666 196360
rect 153430 196348 153436 196360
rect 152660 196320 153436 196348
rect 152660 196308 152666 196320
rect 153430 196308 153436 196320
rect 153488 196308 153494 196360
rect 153798 196308 153804 196360
rect 153856 196348 153862 196360
rect 154810 196348 154816 196360
rect 153856 196320 154816 196348
rect 153856 196308 153862 196320
rect 154810 196308 154816 196320
rect 154868 196308 154874 196360
rect 156006 196308 156012 196360
rect 156064 196348 156070 196360
rect 156834 196348 156840 196360
rect 156064 196320 156840 196348
rect 156064 196308 156070 196320
rect 156834 196308 156840 196320
rect 156892 196308 156898 196360
rect 162630 196308 162636 196360
rect 162688 196348 162694 196360
rect 165850 196348 165856 196360
rect 162688 196320 165856 196348
rect 162688 196308 162694 196320
rect 165850 196308 165856 196320
rect 165908 196308 165914 196360
rect 165942 196308 165948 196360
rect 166000 196348 166006 196360
rect 169990 196348 169996 196360
rect 166000 196320 169996 196348
rect 166000 196308 166006 196320
rect 169990 196308 169996 196320
rect 170048 196308 170054 196360
rect 175970 196308 175976 196360
rect 176028 196348 176034 196360
rect 176798 196348 176804 196360
rect 176028 196320 176804 196348
rect 176028 196308 176034 196320
rect 176798 196308 176804 196320
rect 176856 196308 176862 196360
rect 177074 196308 177080 196360
rect 177132 196348 177138 196360
rect 178178 196348 178184 196360
rect 177132 196320 178184 196348
rect 177132 196308 177138 196320
rect 178178 196308 178184 196320
rect 178236 196308 178242 196360
rect 195106 196308 195112 196360
rect 195164 196348 195170 196360
rect 196026 196348 196032 196360
rect 195164 196320 196032 196348
rect 195164 196308 195170 196320
rect 196026 196308 196032 196320
rect 196084 196308 196090 196360
rect 196210 196308 196216 196360
rect 196268 196348 196274 196360
rect 197222 196348 197228 196360
rect 196268 196320 197228 196348
rect 196268 196308 196274 196320
rect 197222 196308 197228 196320
rect 197280 196308 197286 196360
rect 203294 196308 203300 196360
rect 203352 196348 203358 196360
rect 204398 196348 204404 196360
rect 203352 196320 204404 196348
rect 203352 196308 203358 196320
rect 204398 196308 204404 196320
rect 204456 196308 204462 196360
rect 204858 196308 204864 196360
rect 204916 196348 204922 196360
rect 205594 196348 205600 196360
rect 204916 196320 205600 196348
rect 204916 196308 204922 196320
rect 205594 196308 205600 196320
rect 205652 196308 205658 196360
rect 207618 196308 207624 196360
rect 207676 196348 207682 196360
rect 208446 196348 208452 196360
rect 207676 196320 208452 196348
rect 207676 196308 207682 196320
rect 208446 196308 208452 196320
rect 208504 196308 208510 196360
rect 27666 196240 27672 196292
rect 27724 196280 27730 196292
rect 30058 196280 30064 196292
rect 27724 196252 30064 196280
rect 27724 196240 27730 196252
rect 30058 196240 30064 196252
rect 30116 196240 30122 196292
rect 80842 196240 80848 196292
rect 80900 196280 80906 196292
rect 84522 196280 84528 196292
rect 80900 196252 84528 196280
rect 80900 196240 80906 196252
rect 84522 196240 84528 196252
rect 84580 196240 84586 196292
rect 122426 196240 122432 196292
rect 122484 196280 122490 196292
rect 123990 196280 123996 196292
rect 122484 196252 123996 196280
rect 122484 196240 122490 196252
rect 123990 196240 123996 196252
rect 124048 196240 124054 196292
rect 201454 196240 201460 196292
rect 201512 196280 201518 196292
rect 201638 196280 201644 196292
rect 201512 196252 201644 196280
rect 201512 196240 201518 196252
rect 201638 196240 201644 196252
rect 201696 196240 201702 196292
rect 205226 196240 205232 196292
rect 205284 196280 205290 196292
rect 205778 196280 205784 196292
rect 205284 196252 205784 196280
rect 205284 196240 205290 196252
rect 205778 196240 205784 196252
rect 205836 196240 205842 196292
rect 39626 196172 39632 196224
rect 39684 196212 39690 196224
rect 41098 196212 41104 196224
rect 39684 196184 41104 196212
rect 39684 196172 39690 196184
rect 41098 196172 41104 196184
rect 41156 196172 41162 196224
rect 30518 196104 30524 196156
rect 30576 196144 30582 196156
rect 31622 196144 31628 196156
rect 30576 196116 31628 196144
rect 30576 196104 30582 196116
rect 31622 196104 31628 196116
rect 31680 196104 31686 196156
rect 51034 196104 51040 196156
rect 51092 196144 51098 196156
rect 59774 196144 59780 196156
rect 51092 196116 59780 196144
rect 51092 196104 51098 196116
rect 59774 196104 59780 196116
rect 59832 196104 59838 196156
rect 135398 196104 135404 196156
rect 135456 196144 135462 196156
rect 143770 196144 143776 196156
rect 135456 196116 143776 196144
rect 135456 196104 135462 196116
rect 143770 196104 143776 196116
rect 143828 196104 143834 196156
rect 154902 196104 154908 196156
rect 154960 196144 154966 196156
rect 156190 196144 156196 196156
rect 154960 196116 156196 196144
rect 154960 196104 154966 196116
rect 156190 196104 156196 196116
rect 156248 196104 156254 196156
rect 160422 196104 160428 196156
rect 160480 196144 160486 196156
rect 162354 196144 162360 196156
rect 160480 196116 162360 196144
rect 160480 196104 160486 196116
rect 162354 196104 162360 196116
rect 162412 196104 162418 196156
rect 206422 196104 206428 196156
rect 206480 196144 206486 196156
rect 208078 196144 208084 196156
rect 206480 196116 208084 196144
rect 206480 196104 206486 196116
rect 208078 196104 208084 196116
rect 208136 196104 208142 196156
rect 51218 196036 51224 196088
rect 51276 196076 51282 196088
rect 58670 196076 58676 196088
rect 51276 196048 58676 196076
rect 51276 196036 51282 196048
rect 58670 196036 58676 196048
rect 58728 196036 58734 196088
rect 89766 196036 89772 196088
rect 89824 196076 89830 196088
rect 101634 196076 101640 196088
rect 89824 196048 101640 196076
rect 89824 196036 89830 196048
rect 101634 196036 101640 196048
rect 101692 196036 101698 196088
rect 135214 196036 135220 196088
rect 135272 196076 135278 196088
rect 142666 196076 142672 196088
rect 135272 196048 142672 196076
rect 135272 196036 135278 196048
rect 142666 196036 142672 196048
rect 142724 196036 142730 196088
rect 173762 196036 173768 196088
rect 173820 196076 173826 196088
rect 185814 196076 185820 196088
rect 173820 196048 185820 196076
rect 173820 196036 173826 196048
rect 185814 196036 185820 196048
rect 185872 196036 185878 196088
rect 39258 195968 39264 196020
rect 39316 196008 39322 196020
rect 41006 196008 41012 196020
rect 39316 195980 41012 196008
rect 39316 195968 39322 195980
rect 41006 195968 41012 195980
rect 41064 195968 41070 196020
rect 50942 195968 50948 196020
rect 51000 196008 51006 196020
rect 60878 196008 60884 196020
rect 51000 195980 60884 196008
rect 51000 195968 51006 195980
rect 60878 195968 60884 195980
rect 60936 195968 60942 196020
rect 88662 195968 88668 196020
rect 88720 196008 88726 196020
rect 101726 196008 101732 196020
rect 88720 195980 101732 196008
rect 88720 195968 88726 195980
rect 101726 195968 101732 195980
rect 101784 195968 101790 196020
rect 124450 195968 124456 196020
rect 124508 196008 124514 196020
rect 127854 196008 127860 196020
rect 124508 195980 127860 196008
rect 124508 195968 124514 195980
rect 127854 195968 127860 195980
rect 127912 195968 127918 196020
rect 134938 195968 134944 196020
rect 134996 196008 135002 196020
rect 144874 196008 144880 196020
rect 134996 195980 144880 196008
rect 134996 195968 135002 195980
rect 144874 195968 144880 195980
rect 144932 195968 144938 196020
rect 161526 195968 161532 196020
rect 161584 196008 161590 196020
rect 164470 196008 164476 196020
rect 161584 195980 164476 196008
rect 161584 195968 161590 195980
rect 164470 195968 164476 195980
rect 164528 195968 164534 196020
rect 164838 195968 164844 196020
rect 164896 196008 164902 196020
rect 168610 196008 168616 196020
rect 164896 195980 168616 196008
rect 164896 195968 164902 195980
rect 168610 195968 168616 195980
rect 168668 195968 168674 196020
rect 172658 195968 172664 196020
rect 172716 196008 172722 196020
rect 185906 196008 185912 196020
rect 172716 195980 185912 196008
rect 172716 195968 172722 195980
rect 185906 195968 185912 195980
rect 185964 195968 185970 196020
rect 193266 195968 193272 196020
rect 193324 196008 193330 196020
rect 194462 196008 194468 196020
rect 193324 195980 194468 196008
rect 193324 195968 193330 195980
rect 194462 195968 194468 195980
rect 194520 195968 194526 196020
rect 202098 195968 202104 196020
rect 202156 196008 202162 196020
rect 202834 196008 202840 196020
rect 202156 195980 202840 196008
rect 202156 195968 202162 195980
rect 202834 195968 202840 195980
rect 202892 195968 202898 196020
rect 209274 195968 209280 196020
rect 209332 196008 209338 196020
rect 213046 196008 213052 196020
rect 209332 195980 213052 196008
rect 209332 195968 209338 195980
rect 213046 195968 213052 195980
rect 213104 195968 213110 196020
rect 50758 195900 50764 195952
rect 50816 195940 50822 195952
rect 61982 195940 61988 195952
rect 50816 195912 61988 195940
rect 50816 195900 50822 195912
rect 61982 195900 61988 195912
rect 62040 195900 62046 195952
rect 81946 195900 81952 195952
rect 82004 195940 82010 195952
rect 87190 195940 87196 195952
rect 82004 195912 87196 195940
rect 82004 195900 82010 195912
rect 87190 195900 87196 195912
rect 87248 195900 87254 195952
rect 87558 195900 87564 195952
rect 87616 195940 87622 195952
rect 102094 195940 102100 195952
rect 87616 195912 102100 195940
rect 87616 195900 87622 195912
rect 102094 195900 102100 195912
rect 102152 195900 102158 195952
rect 135122 195900 135128 195952
rect 135180 195940 135186 195952
rect 145978 195940 145984 195952
rect 135180 195912 145984 195940
rect 135180 195900 135186 195912
rect 145978 195900 145984 195912
rect 146036 195900 146042 195952
rect 171554 195900 171560 195952
rect 171612 195940 171618 195952
rect 186274 195940 186280 195952
rect 171612 195912 186280 195940
rect 171612 195900 171618 195912
rect 186274 195900 186280 195912
rect 186332 195900 186338 195952
rect 208814 195900 208820 195952
rect 208872 195940 208878 195952
rect 212862 195940 212868 195952
rect 208872 195912 212868 195940
rect 208872 195900 208878 195912
rect 212862 195900 212868 195912
rect 212920 195900 212926 195952
rect 26378 195832 26384 195884
rect 26436 195872 26442 195884
rect 29690 195872 29696 195884
rect 26436 195844 29696 195872
rect 26436 195832 26442 195844
rect 29690 195832 29696 195844
rect 29748 195832 29754 195884
rect 31898 195832 31904 195884
rect 31956 195872 31962 195884
rect 32818 195872 32824 195884
rect 31956 195844 32824 195872
rect 31956 195832 31962 195844
rect 32818 195832 32824 195844
rect 32876 195832 32882 195884
rect 36866 195832 36872 195884
rect 36924 195872 36930 195884
rect 37326 195872 37332 195884
rect 36924 195844 37332 195872
rect 36924 195832 36930 195844
rect 37326 195832 37332 195844
rect 37384 195832 37390 195884
rect 41282 195832 41288 195884
rect 41340 195872 41346 195884
rect 43766 195872 43772 195884
rect 41340 195844 43772 195872
rect 41340 195832 41346 195844
rect 43766 195832 43772 195844
rect 43824 195832 43830 195884
rect 50666 195832 50672 195884
rect 50724 195872 50730 195884
rect 63086 195872 63092 195884
rect 50724 195844 63092 195872
rect 50724 195832 50730 195844
rect 63086 195832 63092 195844
rect 63144 195832 63150 195884
rect 86454 195832 86460 195884
rect 86512 195872 86518 195884
rect 101910 195872 101916 195884
rect 86512 195844 101916 195872
rect 86512 195832 86518 195844
rect 101910 195832 101916 195844
rect 101968 195832 101974 195884
rect 122058 195832 122064 195884
rect 122116 195872 122122 195884
rect 123714 195872 123720 195884
rect 122116 195844 123720 195872
rect 122116 195832 122122 195844
rect 123714 195832 123720 195844
rect 123772 195832 123778 195884
rect 135030 195832 135036 195884
rect 135088 195872 135094 195884
rect 148186 195872 148192 195884
rect 135088 195844 148192 195872
rect 135088 195832 135094 195844
rect 148186 195832 148192 195844
rect 148244 195832 148250 195884
rect 163734 195832 163740 195884
rect 163792 195872 163798 195884
rect 167230 195872 167236 195884
rect 163792 195844 167236 195872
rect 163792 195832 163798 195844
rect 167230 195832 167236 195844
rect 167288 195832 167294 195884
rect 170450 195832 170456 195884
rect 170508 195872 170514 195884
rect 186090 195872 186096 195884
rect 170508 195844 186096 195872
rect 170508 195832 170514 195844
rect 186090 195832 186096 195844
rect 186148 195832 186154 195884
rect 209642 195832 209648 195884
rect 209700 195872 209706 195884
rect 213414 195872 213420 195884
rect 209700 195844 213420 195872
rect 209700 195832 209706 195844
rect 213414 195832 213420 195844
rect 213472 195832 213478 195884
rect 26286 195764 26292 195816
rect 26344 195804 26350 195816
rect 29230 195804 29236 195816
rect 26344 195776 29236 195804
rect 26344 195764 26350 195776
rect 29230 195764 29236 195776
rect 29288 195764 29294 195816
rect 50850 195764 50856 195816
rect 50908 195804 50914 195816
rect 64190 195804 64196 195816
rect 50908 195776 64196 195804
rect 50908 195764 50914 195776
rect 64190 195764 64196 195776
rect 64248 195764 64254 195816
rect 65018 195764 65024 195816
rect 65076 195804 65082 195816
rect 94182 195804 94188 195816
rect 65076 195776 94188 195804
rect 65076 195764 65082 195776
rect 94182 195764 94188 195776
rect 94240 195764 94246 195816
rect 125646 195764 125652 195816
rect 125704 195804 125710 195816
rect 127946 195804 127952 195816
rect 125704 195776 127952 195804
rect 125704 195764 125710 195776
rect 127946 195764 127952 195776
rect 128004 195764 128010 195816
rect 134846 195764 134852 195816
rect 134904 195804 134910 195816
rect 147082 195804 147088 195816
rect 134904 195776 147088 195804
rect 134904 195764 134910 195776
rect 147082 195764 147088 195776
rect 147140 195764 147146 195816
rect 147818 195764 147824 195816
rect 147876 195804 147882 195816
rect 179282 195804 179288 195816
rect 147876 195776 179288 195804
rect 147876 195764 147882 195776
rect 179282 195764 179288 195776
rect 179340 195764 179346 195816
rect 208446 195764 208452 195816
rect 208504 195804 208510 195816
rect 212954 195804 212960 195816
rect 208504 195776 212960 195804
rect 208504 195764 208510 195776
rect 212954 195764 212960 195776
rect 213012 195764 213018 195816
rect 26194 195696 26200 195748
rect 26252 195736 26258 195748
rect 28862 195736 28868 195748
rect 26252 195708 28868 195736
rect 26252 195696 26258 195708
rect 28862 195696 28868 195708
rect 28920 195696 28926 195748
rect 31990 195696 31996 195748
rect 32048 195736 32054 195748
rect 32910 195736 32916 195748
rect 32048 195708 32916 195736
rect 32048 195696 32054 195708
rect 32910 195696 32916 195708
rect 32968 195696 32974 195748
rect 33370 195696 33376 195748
rect 33428 195736 33434 195748
rect 34474 195736 34480 195748
rect 33428 195708 34480 195736
rect 33428 195696 33434 195708
rect 34474 195696 34480 195708
rect 34532 195696 34538 195748
rect 79738 195696 79744 195748
rect 79796 195736 79802 195748
rect 83050 195736 83056 195748
rect 79796 195708 83056 195736
rect 79796 195696 79802 195708
rect 83050 195696 83056 195708
rect 83108 195696 83114 195748
rect 91974 195696 91980 195748
rect 92032 195736 92038 195748
rect 92618 195736 92624 195748
rect 92032 195708 92624 195736
rect 92032 195696 92038 195708
rect 92618 195696 92624 195708
rect 92676 195696 92682 195748
rect 122886 195696 122892 195748
rect 122944 195736 122950 195748
rect 123898 195736 123904 195748
rect 122944 195708 123904 195736
rect 122944 195696 122950 195708
rect 123898 195696 123904 195708
rect 123956 195696 123962 195748
rect 194922 195696 194928 195748
rect 194980 195736 194986 195748
rect 195658 195736 195664 195748
rect 194980 195708 195664 195736
rect 194980 195696 194986 195708
rect 195658 195696 195664 195708
rect 195716 195696 195722 195748
rect 206054 195696 206060 195748
rect 206112 195736 206118 195748
rect 207986 195736 207992 195748
rect 206112 195708 207992 195736
rect 206112 195696 206118 195708
rect 207986 195696 207992 195708
rect 208044 195696 208050 195748
rect 38062 195628 38068 195680
rect 38120 195668 38126 195680
rect 38982 195668 38988 195680
rect 38120 195640 38988 195668
rect 38120 195628 38126 195640
rect 38982 195628 38988 195640
rect 39040 195628 39046 195680
rect 40454 195628 40460 195680
rect 40512 195668 40518 195680
rect 43122 195668 43128 195680
rect 40512 195640 43128 195668
rect 40512 195628 40518 195640
rect 43122 195628 43128 195640
rect 43180 195628 43186 195680
rect 125278 195628 125284 195680
rect 125336 195668 125342 195680
rect 128130 195668 128136 195680
rect 125336 195640 128136 195668
rect 125336 195628 125342 195640
rect 128130 195628 128136 195640
rect 128188 195628 128194 195680
rect 207250 195628 207256 195680
rect 207308 195668 207314 195680
rect 208538 195668 208544 195680
rect 207308 195640 208544 195668
rect 207308 195628 207314 195640
rect 208538 195628 208544 195640
rect 208596 195628 208602 195680
rect 124818 195560 124824 195612
rect 124876 195600 124882 195612
rect 128038 195600 128044 195612
rect 124876 195572 128044 195600
rect 124876 195560 124882 195572
rect 128038 195560 128044 195572
rect 128096 195560 128102 195612
rect 206882 195560 206888 195612
rect 206940 195600 206946 195612
rect 207894 195600 207900 195612
rect 206940 195572 207900 195600
rect 206940 195560 206946 195572
rect 207894 195560 207900 195572
rect 207952 195560 207958 195612
rect 33462 195492 33468 195544
rect 33520 195532 33526 195544
rect 34106 195532 34112 195544
rect 33520 195504 34112 195532
rect 33520 195492 33526 195504
rect 34106 195492 34112 195504
rect 34164 195492 34170 195544
rect 77530 195492 77536 195544
rect 77588 195532 77594 195544
rect 79554 195532 79560 195544
rect 77588 195504 79560 195532
rect 77588 195492 77594 195504
rect 79554 195492 79560 195504
rect 79612 195492 79618 195544
rect 29138 195424 29144 195476
rect 29196 195464 29202 195476
rect 30886 195464 30892 195476
rect 29196 195436 30892 195464
rect 29196 195424 29202 195436
rect 30886 195424 30892 195436
rect 30944 195424 30950 195476
rect 37694 195424 37700 195476
rect 37752 195464 37758 195476
rect 38890 195464 38896 195476
rect 37752 195436 38896 195464
rect 37752 195424 37758 195436
rect 38890 195424 38896 195436
rect 38948 195424 38954 195476
rect 51126 195424 51132 195476
rect 51184 195464 51190 195476
rect 56462 195464 56468 195476
rect 51184 195436 56468 195464
rect 51184 195424 51190 195436
rect 56462 195424 56468 195436
rect 56520 195424 56526 195476
rect 76426 195424 76432 195476
rect 76484 195464 76490 195476
rect 78174 195464 78180 195476
rect 76484 195436 78180 195464
rect 76484 195424 76490 195436
rect 78174 195424 78180 195436
rect 78232 195424 78238 195476
rect 119298 195424 119304 195476
rect 119356 195464 119362 195476
rect 120126 195464 120132 195476
rect 119356 195436 120132 195464
rect 119356 195424 119362 195436
rect 120126 195424 120132 195436
rect 120184 195424 120190 195476
rect 197590 195356 197596 195408
rect 197648 195396 197654 195408
rect 198050 195396 198056 195408
rect 197648 195368 198056 195396
rect 197648 195356 197654 195368
rect 198050 195356 198056 195368
rect 198108 195356 198114 195408
rect 38890 195288 38896 195340
rect 38948 195328 38954 195340
rect 40822 195328 40828 195340
rect 38948 195300 40828 195328
rect 38948 195288 38954 195300
rect 40822 195288 40828 195300
rect 40880 195288 40886 195340
rect 159318 195288 159324 195340
rect 159376 195328 159382 195340
rect 160974 195328 160980 195340
rect 159376 195300 160980 195328
rect 159376 195288 159382 195300
rect 160974 195288 160980 195300
rect 161032 195288 161038 195340
rect 29046 195220 29052 195272
rect 29104 195260 29110 195272
rect 31254 195260 31260 195272
rect 29104 195232 31260 195260
rect 29104 195220 29110 195232
rect 31254 195220 31260 195232
rect 31312 195220 31318 195272
rect 194646 195220 194652 195272
rect 194704 195260 194710 195272
rect 195290 195260 195296 195272
rect 194704 195232 195296 195260
rect 194704 195220 194710 195232
rect 195290 195220 195296 195232
rect 195348 195220 195354 195272
rect 30426 195152 30432 195204
rect 30484 195192 30490 195204
rect 30484 195164 32128 195192
rect 30484 195152 30490 195164
rect 32100 195136 32128 195164
rect 40822 195152 40828 195204
rect 40880 195192 40886 195204
rect 43674 195192 43680 195204
rect 40880 195164 43680 195192
rect 40880 195152 40886 195164
rect 43674 195152 43680 195164
rect 43732 195152 43738 195204
rect 32082 195084 32088 195136
rect 32140 195084 32146 195136
rect 118654 194132 118660 194184
rect 118712 194172 118718 194184
rect 118838 194172 118844 194184
rect 118712 194144 118844 194172
rect 118712 194132 118718 194144
rect 118838 194132 118844 194144
rect 118896 194132 118902 194184
rect 211942 190596 211948 190648
rect 212000 190636 212006 190648
rect 217554 190636 217560 190648
rect 212000 190608 217560 190636
rect 212000 190596 212006 190608
rect 217554 190596 217560 190608
rect 217612 190596 217618 190648
rect 187930 188216 187936 188268
rect 187988 188256 187994 188268
rect 191978 188256 191984 188268
rect 187988 188228 191984 188256
rect 187988 188216 187994 188228
rect 191978 188216 191984 188228
rect 192036 188216 192042 188268
rect 99426 186856 99432 186908
rect 99484 186896 99490 186908
rect 106786 186896 106792 186908
rect 99484 186868 106792 186896
rect 99484 186856 99490 186868
rect 106786 186856 106792 186868
rect 106844 186856 106850 186908
rect 13314 186788 13320 186840
rect 13372 186828 13378 186840
rect 22790 186828 22796 186840
rect 13372 186800 22796 186828
rect 13372 186788 13378 186800
rect 22790 186788 22796 186800
rect 22848 186788 22854 186840
rect 104394 184068 104400 184120
rect 104452 184108 104458 184120
rect 106786 184108 106792 184120
rect 104452 184080 106792 184108
rect 104452 184068 104458 184080
rect 106786 184068 106792 184080
rect 106844 184068 106850 184120
rect 99518 184000 99524 184052
rect 99576 184040 99582 184052
rect 105774 184040 105780 184052
rect 99576 184012 105780 184040
rect 99576 184000 99582 184012
rect 105774 184000 105780 184012
rect 105832 184000 105838 184052
rect 182870 184000 182876 184052
rect 182928 184040 182934 184052
rect 187930 184040 187936 184052
rect 182928 184012 187936 184040
rect 182928 184000 182934 184012
rect 187930 184000 187936 184012
rect 187988 184000 187994 184052
rect 13406 182708 13412 182760
rect 13464 182748 13470 182760
rect 22330 182748 22336 182760
rect 13464 182720 22336 182748
rect 13464 182708 13470 182720
rect 22330 182708 22336 182720
rect 22388 182708 22394 182760
rect 104486 182708 104492 182760
rect 104544 182748 104550 182760
rect 107154 182748 107160 182760
rect 104544 182720 107160 182748
rect 104544 182708 104550 182720
rect 107154 182708 107160 182720
rect 107212 182708 107218 182760
rect 128498 182708 128504 182760
rect 128556 182748 128562 182760
rect 137514 182748 137520 182760
rect 128556 182720 137520 182748
rect 128556 182708 128562 182720
rect 137514 182708 137520 182720
rect 137572 182708 137578 182760
rect 212494 182708 212500 182760
rect 212552 182748 212558 182760
rect 220406 182748 220412 182760
rect 212552 182720 220412 182748
rect 212552 182708 212558 182720
rect 220406 182708 220412 182720
rect 220464 182708 220470 182760
rect 98598 182640 98604 182692
rect 98656 182680 98662 182692
rect 106970 182680 106976 182692
rect 98656 182652 106976 182680
rect 98656 182640 98662 182652
rect 106970 182640 106976 182652
rect 107028 182640 107034 182692
rect 183146 182640 183152 182692
rect 183204 182680 183210 182692
rect 191150 182680 191156 182692
rect 183204 182652 191156 182680
rect 183204 182640 183210 182652
rect 191150 182640 191156 182652
rect 191208 182640 191214 182692
rect 183698 181280 183704 181332
rect 183756 181320 183762 181332
rect 191978 181320 191984 181332
rect 183756 181292 191984 181320
rect 183756 181280 183762 181292
rect 191978 181280 191984 181292
rect 192036 181280 192042 181332
rect 105130 180328 105136 180380
rect 105188 180368 105194 180380
rect 106970 180368 106976 180380
rect 105188 180340 106976 180368
rect 105188 180328 105194 180340
rect 106970 180328 106976 180340
rect 107028 180328 107034 180380
rect 98414 179852 98420 179904
rect 98472 179892 98478 179904
rect 104486 179892 104492 179904
rect 98472 179864 104492 179892
rect 98472 179852 98478 179864
rect 104486 179852 104492 179864
rect 104544 179852 104550 179904
rect 182502 179852 182508 179904
rect 182560 179892 182566 179904
rect 190690 179892 190696 179904
rect 182560 179864 190696 179892
rect 182560 179852 182566 179864
rect 190690 179852 190696 179864
rect 190748 179852 190754 179904
rect 183698 179784 183704 179836
rect 183756 179824 183762 179836
rect 190598 179824 190604 179836
rect 183756 179796 190604 179824
rect 183756 179784 183762 179796
rect 190598 179784 190604 179796
rect 190656 179784 190662 179836
rect 99518 179512 99524 179564
rect 99576 179552 99582 179564
rect 104394 179552 104400 179564
rect 99576 179524 104400 179552
rect 99576 179512 99582 179524
rect 104394 179512 104400 179524
rect 104452 179512 104458 179564
rect 182502 178492 182508 178544
rect 182560 178532 182566 178544
rect 191978 178532 191984 178544
rect 182560 178504 191984 178532
rect 182560 178492 182566 178504
rect 191978 178492 191984 178504
rect 192036 178492 192042 178544
rect 99518 177336 99524 177388
rect 99576 177376 99582 177388
rect 105130 177376 105136 177388
rect 99576 177348 105136 177376
rect 99576 177336 99582 177348
rect 105130 177336 105136 177348
rect 105188 177336 105194 177388
rect 98598 177132 98604 177184
rect 98656 177172 98662 177184
rect 106786 177172 106792 177184
rect 98656 177144 106792 177172
rect 98656 177132 98662 177144
rect 106786 177132 106792 177144
rect 106844 177132 106850 177184
rect 183238 176452 183244 176504
rect 183296 176492 183302 176504
rect 191978 176492 191984 176504
rect 183296 176464 191984 176492
rect 183296 176452 183302 176464
rect 191978 176452 191984 176464
rect 192036 176452 192042 176504
rect 211758 176316 211764 176368
rect 211816 176356 211822 176368
rect 216266 176356 216272 176368
rect 211816 176328 216272 176356
rect 211816 176316 211822 176328
rect 216266 176316 216272 176328
rect 216324 176316 216330 176368
rect 13314 175840 13320 175892
rect 13372 175880 13378 175892
rect 22330 175880 22336 175892
rect 13372 175852 22336 175880
rect 13372 175840 13378 175852
rect 22330 175840 22336 175852
rect 22388 175840 22394 175892
rect 98230 175772 98236 175824
rect 98288 175812 98294 175824
rect 106602 175812 106608 175824
rect 98288 175784 106608 175812
rect 98288 175772 98294 175784
rect 106602 175772 106608 175784
rect 106660 175772 106666 175824
rect 183698 175092 183704 175144
rect 183756 175132 183762 175144
rect 191518 175132 191524 175144
rect 183756 175104 191524 175132
rect 183756 175092 183762 175104
rect 191518 175092 191524 175104
rect 191576 175092 191582 175144
rect 99518 173664 99524 173716
rect 99576 173704 99582 173716
rect 106786 173704 106792 173716
rect 99576 173676 106792 173704
rect 99576 173664 99582 173676
rect 106786 173664 106792 173676
rect 106844 173664 106850 173716
rect 183330 173052 183336 173104
rect 183388 173092 183394 173104
rect 191978 173092 191984 173104
rect 183388 173064 191984 173092
rect 183388 173052 183394 173064
rect 191978 173052 191984 173064
rect 192036 173052 192042 173104
rect 99518 171692 99524 171744
rect 99576 171732 99582 171744
rect 106786 171732 106792 171744
rect 99576 171704 106792 171732
rect 99576 171692 99582 171704
rect 106786 171692 106792 171704
rect 106844 171692 106850 171744
rect 183514 171692 183520 171744
rect 183572 171732 183578 171744
rect 191150 171732 191156 171744
rect 183572 171704 191156 171732
rect 183572 171692 183578 171704
rect 191150 171692 191156 171704
rect 191208 171692 191214 171744
rect 182686 171216 182692 171268
rect 182744 171256 182750 171268
rect 185078 171256 185084 171268
rect 182744 171228 185084 171256
rect 182744 171216 182750 171228
rect 185078 171216 185084 171228
rect 185136 171216 185142 171268
rect 99426 170264 99432 170316
rect 99484 170304 99490 170316
rect 99484 170276 99656 170304
rect 99484 170264 99490 170276
rect 99628 170236 99656 170276
rect 106786 170236 106792 170248
rect 99628 170208 106792 170236
rect 106786 170196 106792 170208
rect 106844 170196 106850 170248
rect 99518 168904 99524 168956
rect 99576 168944 99582 168956
rect 106694 168944 106700 168956
rect 99576 168916 106700 168944
rect 99576 168904 99582 168916
rect 106694 168904 106700 168916
rect 106752 168904 106758 168956
rect 182502 168904 182508 168956
rect 182560 168944 182566 168956
rect 191886 168944 191892 168956
rect 182560 168916 191892 168944
rect 182560 168904 182566 168916
rect 191886 168904 191892 168916
rect 191944 168904 191950 168956
rect 44410 168836 44416 168888
rect 44468 168876 44474 168888
rect 49838 168876 49844 168888
rect 44468 168848 49844 168876
rect 44468 168836 44474 168848
rect 49838 168836 49844 168848
rect 49896 168836 49902 168888
rect 185078 168836 185084 168888
rect 185136 168876 185142 168888
rect 191978 168876 191984 168888
rect 185136 168848 191984 168876
rect 185136 168836 185142 168848
rect 191978 168836 191984 168848
rect 192036 168836 192042 168888
rect 99518 167612 99524 167664
rect 99576 167652 99582 167664
rect 106878 167652 106884 167664
rect 99576 167624 106884 167652
rect 99576 167612 99582 167624
rect 106878 167612 106884 167624
rect 106936 167612 106942 167664
rect 49838 167544 49844 167596
rect 49896 167584 49902 167596
rect 53426 167584 53432 167596
rect 49896 167556 53432 167584
rect 49896 167544 49902 167556
rect 53426 167544 53432 167556
rect 53484 167544 53490 167596
rect 99426 167544 99432 167596
rect 99484 167584 99490 167596
rect 106786 167584 106792 167596
rect 99484 167556 106792 167584
rect 99484 167544 99490 167556
rect 106786 167544 106792 167556
rect 106844 167544 106850 167596
rect 183698 167544 183704 167596
rect 183756 167584 183762 167596
rect 191334 167584 191340 167596
rect 183756 167556 191340 167584
rect 183756 167544 183762 167556
rect 191334 167544 191340 167556
rect 191392 167544 191398 167596
rect 182870 166456 182876 166508
rect 182928 166496 182934 166508
rect 187930 166496 187936 166508
rect 182928 166468 187936 166496
rect 182928 166456 182934 166468
rect 187930 166456 187936 166468
rect 187988 166456 187994 166508
rect 99518 166184 99524 166236
rect 99576 166224 99582 166236
rect 107246 166224 107252 166236
rect 99576 166196 107252 166224
rect 99576 166184 99582 166196
rect 107246 166184 107252 166196
rect 107304 166184 107310 166236
rect 212678 165232 212684 165284
rect 212736 165272 212742 165284
rect 218290 165272 218296 165284
rect 212736 165244 218296 165272
rect 212736 165232 212742 165244
rect 218290 165232 218296 165244
rect 218348 165232 218354 165284
rect 183698 164960 183704 165012
rect 183756 165000 183762 165012
rect 190046 165000 190052 165012
rect 183756 164972 190052 165000
rect 183756 164960 183762 164972
rect 190046 164960 190052 164972
rect 190104 164960 190110 165012
rect 99518 164756 99524 164808
rect 99576 164796 99582 164808
rect 107154 164796 107160 164808
rect 99576 164768 107160 164796
rect 99576 164756 99582 164768
rect 107154 164756 107160 164768
rect 107212 164756 107218 164808
rect 211758 163600 211764 163652
rect 211816 163640 211822 163652
rect 218290 163640 218296 163652
rect 211816 163612 218296 163640
rect 211816 163600 211822 163612
rect 218290 163600 218296 163612
rect 218348 163600 218354 163652
rect 99518 163396 99524 163448
rect 99576 163436 99582 163448
rect 104394 163436 104400 163448
rect 99576 163408 104400 163436
rect 99576 163396 99582 163408
rect 104394 163396 104400 163408
rect 104452 163396 104458 163448
rect 128498 163396 128504 163448
rect 128556 163436 128562 163448
rect 138158 163436 138164 163448
rect 128556 163408 138164 163436
rect 128556 163396 128562 163408
rect 138158 163396 138164 163408
rect 138216 163396 138222 163448
rect 183054 163396 183060 163448
rect 183112 163436 183118 163448
rect 189954 163436 189960 163448
rect 183112 163408 189960 163436
rect 183112 163396 183118 163408
rect 189954 163396 189960 163408
rect 190012 163396 190018 163448
rect 183790 162988 183796 163040
rect 183848 163028 183854 163040
rect 191978 163028 191984 163040
rect 183848 163000 191984 163028
rect 183848 162988 183854 163000
rect 191978 162988 191984 163000
rect 192036 162988 192042 163040
rect 187930 161968 187936 162020
rect 187988 162008 187994 162020
rect 191334 162008 191340 162020
rect 187988 161980 191340 162008
rect 187988 161968 187994 161980
rect 191334 161968 191340 161980
rect 191392 161968 191398 162020
rect 211942 156460 211948 156512
rect 212000 156500 212006 156512
rect 212678 156500 212684 156512
rect 212000 156472 212684 156500
rect 212000 156460 212006 156472
rect 212678 156460 212684 156472
rect 212736 156500 212742 156512
rect 216910 156500 216916 156512
rect 212736 156472 216916 156500
rect 212736 156460 212742 156472
rect 216910 156460 216916 156472
rect 216968 156460 216974 156512
rect 182686 155440 182692 155492
rect 182744 155480 182750 155492
rect 188022 155480 188028 155492
rect 182744 155452 188028 155480
rect 182744 155440 182750 155452
rect 188022 155440 188028 155452
rect 188080 155440 188086 155492
rect 104394 155032 104400 155084
rect 104452 155072 104458 155084
rect 106510 155072 106516 155084
rect 104452 155044 106516 155072
rect 104452 155032 104458 155044
rect 106510 155032 106516 155044
rect 106568 155032 106574 155084
rect 27758 152312 27764 152364
rect 27816 152352 27822 152364
rect 29690 152352 29696 152364
rect 27816 152324 29696 152352
rect 27816 152312 27822 152324
rect 29690 152312 29696 152324
rect 29748 152312 29754 152364
rect 30518 152312 30524 152364
rect 30576 152352 30582 152364
rect 31254 152352 31260 152364
rect 30576 152324 31260 152352
rect 30576 152312 30582 152324
rect 31254 152312 31260 152324
rect 31312 152312 31318 152364
rect 32082 152312 32088 152364
rect 32140 152352 32146 152364
rect 32818 152352 32824 152364
rect 32140 152324 32824 152352
rect 32140 152312 32146 152324
rect 32818 152312 32824 152324
rect 32876 152312 32882 152364
rect 37234 152312 37240 152364
rect 37292 152352 37298 152364
rect 38982 152352 38988 152364
rect 37292 152324 38988 152352
rect 37292 152312 37298 152324
rect 38982 152312 38988 152324
rect 39040 152312 39046 152364
rect 39258 152312 39264 152364
rect 39316 152352 39322 152364
rect 40178 152352 40184 152364
rect 39316 152324 40184 152352
rect 39316 152312 39322 152324
rect 40178 152312 40184 152324
rect 40236 152312 40242 152364
rect 41650 152312 41656 152364
rect 41708 152352 41714 152364
rect 43674 152352 43680 152364
rect 41708 152324 43680 152352
rect 41708 152312 41714 152324
rect 43674 152312 43680 152324
rect 43732 152312 43738 152364
rect 109178 152312 109184 152364
rect 109236 152352 109242 152364
rect 110098 152352 110104 152364
rect 109236 152324 110104 152352
rect 109236 152312 109242 152324
rect 110098 152312 110104 152324
rect 110156 152312 110162 152364
rect 119666 152312 119672 152364
rect 119724 152352 119730 152364
rect 121966 152352 121972 152364
rect 119724 152324 121972 152352
rect 119724 152312 119730 152324
rect 121966 152312 121972 152324
rect 122024 152312 122030 152364
rect 124818 152312 124824 152364
rect 124876 152352 124882 152364
rect 129234 152352 129240 152364
rect 124876 152324 129240 152352
rect 124876 152312 124882 152324
rect 129234 152312 129240 152324
rect 129292 152312 129298 152364
rect 193266 152312 193272 152364
rect 193324 152352 193330 152364
rect 194462 152352 194468 152364
rect 193324 152324 194468 152352
rect 193324 152312 193330 152324
rect 194462 152312 194468 152324
rect 194520 152312 194526 152364
rect 194922 152312 194928 152364
rect 194980 152352 194986 152364
rect 195658 152352 195664 152364
rect 194980 152324 195664 152352
rect 194980 152312 194986 152324
rect 195658 152312 195664 152324
rect 195716 152312 195722 152364
rect 196578 152312 196584 152364
rect 196636 152352 196642 152364
rect 197222 152352 197228 152364
rect 196636 152324 197228 152352
rect 196636 152312 196642 152324
rect 197222 152312 197228 152324
rect 197280 152312 197286 152364
rect 197590 152312 197596 152364
rect 197648 152352 197654 152364
rect 198050 152352 198056 152364
rect 197648 152324 198056 152352
rect 197648 152312 197654 152324
rect 198050 152312 198056 152324
rect 198108 152312 198114 152364
rect 202098 152312 202104 152364
rect 202156 152352 202162 152364
rect 202926 152352 202932 152364
rect 202156 152324 202932 152352
rect 202156 152312 202162 152324
rect 202926 152312 202932 152324
rect 202984 152312 202990 152364
rect 203662 152312 203668 152364
rect 203720 152352 203726 152364
rect 205962 152352 205968 152364
rect 203720 152324 205968 152352
rect 203720 152312 203726 152324
rect 205962 152312 205968 152324
rect 206020 152312 206026 152364
rect 30426 152244 30432 152296
rect 30484 152284 30490 152296
rect 31622 152284 31628 152296
rect 30484 152256 31628 152284
rect 30484 152244 30490 152256
rect 31622 152244 31628 152256
rect 31680 152244 31686 152296
rect 38890 152244 38896 152296
rect 38948 152284 38954 152296
rect 39902 152284 39908 152296
rect 38948 152256 39908 152284
rect 38948 152244 38954 152256
rect 39902 152244 39908 152256
rect 39960 152244 39966 152296
rect 118470 152244 118476 152296
rect 118528 152284 118534 152296
rect 120586 152284 120592 152296
rect 118528 152256 120592 152284
rect 118528 152244 118534 152256
rect 120586 152244 120592 152256
rect 120644 152244 120650 152296
rect 124450 152244 124456 152296
rect 124508 152284 124514 152296
rect 128774 152284 128780 152296
rect 124508 152256 128780 152284
rect 124508 152244 124514 152256
rect 128774 152244 128780 152256
rect 128832 152244 128838 152296
rect 193358 152244 193364 152296
rect 193416 152284 193422 152296
rect 194094 152284 194100 152296
rect 193416 152256 194100 152284
rect 193416 152244 193422 152256
rect 194094 152244 194100 152256
rect 194152 152244 194158 152296
rect 203294 152244 203300 152296
rect 203352 152284 203358 152296
rect 206054 152284 206060 152296
rect 203352 152256 206060 152284
rect 203352 152244 203358 152256
rect 206054 152244 206060 152256
rect 206112 152244 206118 152296
rect 29138 152176 29144 152228
rect 29196 152216 29202 152228
rect 30886 152216 30892 152228
rect 29196 152188 30892 152216
rect 29196 152176 29202 152188
rect 30886 152176 30892 152188
rect 30944 152176 30950 152228
rect 38430 152176 38436 152228
rect 38488 152216 38494 152228
rect 41834 152216 41840 152228
rect 38488 152188 41840 152216
rect 38488 152176 38494 152188
rect 41834 152176 41840 152188
rect 41892 152176 41898 152228
rect 120494 152176 120500 152228
rect 120552 152216 120558 152228
rect 123162 152216 123168 152228
rect 120552 152188 123168 152216
rect 120552 152176 120558 152188
rect 123162 152176 123168 152188
rect 123220 152176 123226 152228
rect 123622 152176 123628 152228
rect 123680 152216 123686 152228
rect 127946 152216 127952 152228
rect 123680 152188 127952 152216
rect 123680 152176 123686 152188
rect 127946 152176 127952 152188
rect 128004 152176 128010 152228
rect 204858 152176 204864 152228
rect 204916 152216 204922 152228
rect 207342 152216 207348 152228
rect 204916 152188 207348 152216
rect 204916 152176 204922 152188
rect 207342 152176 207348 152188
rect 207400 152176 207406 152228
rect 36866 152108 36872 152160
rect 36924 152148 36930 152160
rect 38890 152148 38896 152160
rect 36924 152120 38896 152148
rect 36924 152108 36930 152120
rect 38890 152108 38896 152120
rect 38948 152108 38954 152160
rect 120034 152108 120040 152160
rect 120092 152148 120098 152160
rect 123070 152148 123076 152160
rect 120092 152120 123076 152148
rect 120092 152108 120098 152120
rect 123070 152108 123076 152120
rect 123128 152108 123134 152160
rect 204490 152108 204496 152160
rect 204548 152148 204554 152160
rect 207250 152148 207256 152160
rect 204548 152120 207256 152148
rect 204548 152108 204554 152120
rect 207250 152108 207256 152120
rect 207308 152108 207314 152160
rect 118838 152040 118844 152092
rect 118896 152080 118902 152092
rect 120954 152080 120960 152092
rect 118896 152052 120960 152080
rect 118896 152040 118902 152052
rect 120954 152040 120960 152052
rect 121012 152040 121018 152092
rect 205226 152040 205232 152092
rect 205284 152080 205290 152092
rect 207986 152080 207992 152092
rect 205284 152052 207992 152080
rect 205284 152040 205290 152052
rect 207986 152040 207992 152052
rect 208044 152040 208050 152092
rect 208814 152040 208820 152092
rect 208872 152080 208878 152092
rect 212862 152080 212868 152092
rect 208872 152052 212868 152080
rect 208872 152040 208878 152052
rect 212862 152040 212868 152052
rect 212920 152040 212926 152092
rect 119298 151972 119304 152024
rect 119356 152012 119362 152024
rect 121782 152012 121788 152024
rect 119356 151984 121788 152012
rect 119356 151972 119362 151984
rect 121782 151972 121788 151984
rect 121840 151972 121846 152024
rect 127302 151944 127308 151956
rect 123088 151916 127308 151944
rect 31806 151836 31812 151888
rect 31864 151876 31870 151888
rect 32450 151876 32456 151888
rect 31864 151848 32456 151876
rect 31864 151836 31870 151848
rect 32450 151836 32456 151848
rect 32508 151836 32514 151888
rect 40454 151836 40460 151888
rect 40512 151876 40518 151888
rect 44962 151876 44968 151888
rect 40512 151848 44968 151876
rect 40512 151836 40518 151848
rect 44962 151836 44968 151848
rect 45020 151836 45026 151888
rect 122886 151836 122892 151888
rect 122944 151876 122950 151888
rect 123088 151876 123116 151916
rect 127302 151904 127308 151916
rect 127360 151904 127366 151956
rect 206422 151904 206428 151956
rect 206480 151944 206486 151956
rect 210010 151944 210016 151956
rect 206480 151916 210016 151944
rect 206480 151904 206486 151916
rect 210010 151904 210016 151916
rect 210068 151904 210074 151956
rect 122944 151848 123116 151876
rect 122944 151836 122950 151848
rect 123254 151836 123260 151888
rect 123312 151876 123318 151888
rect 127210 151876 127216 151888
rect 123312 151848 127216 151876
rect 123312 151836 123318 151848
rect 127210 151836 127216 151848
rect 127268 151836 127274 151888
rect 206330 151836 206336 151888
rect 206388 151876 206394 151888
rect 208814 151876 208820 151888
rect 206388 151848 208820 151876
rect 206388 151836 206394 151848
rect 208814 151836 208820 151848
rect 208872 151836 208878 151888
rect 79186 151768 79192 151820
rect 79244 151808 79250 151820
rect 98230 151808 98236 151820
rect 79244 151780 98236 151808
rect 79244 151768 79250 151780
rect 98230 151768 98236 151780
rect 98288 151768 98294 151820
rect 207618 151768 207624 151820
rect 207676 151808 207682 151820
rect 210930 151808 210936 151820
rect 207676 151780 210936 151808
rect 207676 151768 207682 151780
rect 210930 151768 210936 151780
rect 210988 151768 210994 151820
rect 26286 151700 26292 151752
rect 26344 151740 26350 151752
rect 29230 151740 29236 151752
rect 26344 151712 29236 151740
rect 26344 151700 26350 151712
rect 29230 151700 29236 151712
rect 29288 151700 29294 151752
rect 38062 151700 38068 151752
rect 38120 151740 38126 151752
rect 40914 151740 40920 151752
rect 38120 151712 40920 151740
rect 38120 151700 38126 151712
rect 40914 151700 40920 151712
rect 40972 151700 40978 151752
rect 69158 151700 69164 151752
rect 69216 151740 69222 151752
rect 92526 151740 92532 151752
rect 69216 151712 92532 151740
rect 69216 151700 69222 151712
rect 92526 151700 92532 151712
rect 92584 151700 92590 151752
rect 95378 151740 95384 151752
rect 95120 151712 95384 151740
rect 41282 151632 41288 151684
rect 41340 151672 41346 151684
rect 45146 151672 45152 151684
rect 41340 151644 45152 151672
rect 41340 151632 41346 151644
rect 45146 151632 45152 151644
rect 45204 151632 45210 151684
rect 37694 151564 37700 151616
rect 37752 151604 37758 151616
rect 40270 151604 40276 151616
rect 37752 151576 40276 151604
rect 37752 151564 37758 151576
rect 40270 151564 40276 151576
rect 40328 151564 40334 151616
rect 72562 151564 72568 151616
rect 72620 151604 72626 151616
rect 80293 151607 80351 151613
rect 80293 151604 80305 151607
rect 72620 151576 80305 151604
rect 72620 151564 72626 151576
rect 80293 151573 80305 151576
rect 80339 151573 80351 151607
rect 80293 151567 80351 151573
rect 36038 151428 36044 151480
rect 36096 151468 36102 151480
rect 37602 151468 37608 151480
rect 36096 151440 37608 151468
rect 36096 151428 36102 151440
rect 37602 151428 37608 151440
rect 37660 151428 37666 151480
rect 80293 151471 80351 151477
rect 80293 151437 80305 151471
rect 80339 151468 80351 151471
rect 95120 151468 95148 151712
rect 95378 151700 95384 151712
rect 95436 151740 95442 151752
rect 156558 151740 156564 151752
rect 95436 151712 156564 151740
rect 95436 151700 95442 151712
rect 156558 151700 156564 151712
rect 156616 151700 156622 151752
rect 209642 151700 209648 151752
rect 209700 151740 209706 151752
rect 214242 151740 214248 151752
rect 209700 151712 214248 151740
rect 209700 151700 209706 151712
rect 214242 151700 214248 151712
rect 214300 151700 214306 151752
rect 98230 151632 98236 151684
rect 98288 151672 98294 151684
rect 98874 151672 98880 151684
rect 98288 151644 98880 151672
rect 98288 151632 98294 151644
rect 98874 151632 98880 151644
rect 98932 151672 98938 151684
rect 163182 151672 163188 151684
rect 98932 151644 163188 151672
rect 98932 151632 98938 151644
rect 163182 151632 163188 151644
rect 163240 151632 163246 151684
rect 200442 151632 200448 151684
rect 200500 151672 200506 151684
rect 201178 151672 201184 151684
rect 200500 151644 201184 151672
rect 200500 151632 200506 151644
rect 201178 151632 201184 151644
rect 201236 151632 201242 151684
rect 205686 151632 205692 151684
rect 205744 151672 205750 151684
rect 207894 151672 207900 151684
rect 205744 151644 207900 151672
rect 205744 151632 205750 151644
rect 207894 151632 207900 151644
rect 207952 151632 207958 151684
rect 209274 151632 209280 151684
rect 209332 151672 209338 151684
rect 214150 151672 214156 151684
rect 209332 151644 214156 151672
rect 209332 151632 209338 151644
rect 214150 151632 214156 151644
rect 214208 151632 214214 151684
rect 124082 151496 124088 151548
rect 124140 151536 124146 151548
rect 127854 151536 127860 151548
rect 124140 151508 127860 151536
rect 124140 151496 124146 151508
rect 127854 151496 127860 151508
rect 127912 151496 127918 151548
rect 195106 151496 195112 151548
rect 195164 151536 195170 151548
rect 196026 151536 196032 151548
rect 195164 151508 196032 151536
rect 195164 151496 195170 151508
rect 196026 151496 196032 151508
rect 196084 151496 196090 151548
rect 80339 151440 95148 151468
rect 80339 151437 80351 151440
rect 80293 151431 80351 151437
rect 122426 151428 122432 151480
rect 122484 151468 122490 151480
rect 125094 151468 125100 151480
rect 122484 151440 125100 151468
rect 122484 151428 122490 151440
rect 125094 151428 125100 151440
rect 125152 151428 125158 151480
rect 24998 151360 25004 151412
rect 25056 151400 25062 151412
rect 28494 151400 28500 151412
rect 25056 151372 28500 151400
rect 25056 151360 25062 151372
rect 28494 151360 28500 151372
rect 28552 151360 28558 151412
rect 29046 151360 29052 151412
rect 29104 151400 29110 151412
rect 30150 151400 30156 151412
rect 29104 151372 30156 151400
rect 29104 151360 29110 151372
rect 30150 151360 30156 151372
rect 30208 151360 30214 151412
rect 24906 151292 24912 151344
rect 24964 151332 24970 151344
rect 28034 151332 28040 151344
rect 24964 151304 28040 151332
rect 24964 151292 24970 151304
rect 28034 151292 28040 151304
rect 28092 151292 28098 151344
rect 121690 151292 121696 151344
rect 121748 151332 121754 151344
rect 124634 151332 124640 151344
rect 121748 151304 124640 151332
rect 121748 151292 121754 151304
rect 124634 151292 124640 151304
rect 124692 151292 124698 151344
rect 125646 151292 125652 151344
rect 125704 151332 125710 151344
rect 131350 151332 131356 151344
rect 125704 151304 131356 151332
rect 125704 151292 125710 151304
rect 131350 151292 131356 151304
rect 131408 151292 131414 151344
rect 208078 151292 208084 151344
rect 208136 151332 208142 151344
rect 210746 151332 210752 151344
rect 208136 151304 210752 151332
rect 208136 151292 208142 151304
rect 210746 151292 210752 151304
rect 210804 151292 210810 151344
rect 26378 151224 26384 151276
rect 26436 151264 26442 151276
rect 28862 151264 28868 151276
rect 26436 151236 28868 151264
rect 26436 151224 26442 151236
rect 28862 151224 28868 151236
rect 28920 151224 28926 151276
rect 31990 151224 31996 151276
rect 32048 151264 32054 151276
rect 33278 151264 33284 151276
rect 32048 151236 33284 151264
rect 32048 151224 32054 151236
rect 33278 151224 33284 151236
rect 33336 151224 33342 151276
rect 118102 151224 118108 151276
rect 118160 151264 118166 151276
rect 120310 151264 120316 151276
rect 118160 151236 120316 151264
rect 118160 151224 118166 151236
rect 120310 151224 120316 151236
rect 120368 151224 120374 151276
rect 121230 151224 121236 151276
rect 121288 151264 121294 151276
rect 123714 151264 123720 151276
rect 121288 151236 123720 151264
rect 121288 151224 121294 151236
rect 123714 151224 123720 151236
rect 123772 151224 123778 151276
rect 194646 151224 194652 151276
rect 194704 151264 194710 151276
rect 195290 151264 195296 151276
rect 194704 151236 195296 151264
rect 194704 151224 194710 151236
rect 195290 151224 195296 151236
rect 195348 151224 195354 151276
rect 25734 151156 25740 151208
rect 25792 151196 25798 151208
rect 27666 151196 27672 151208
rect 25792 151168 27672 151196
rect 25792 151156 25798 151168
rect 27666 151156 27672 151168
rect 27724 151156 27730 151208
rect 36498 151156 36504 151208
rect 36556 151196 36562 151208
rect 37418 151196 37424 151208
rect 36556 151168 37424 151196
rect 36556 151156 36562 151168
rect 37418 151156 37424 151168
rect 37476 151156 37482 151208
rect 206882 151156 206888 151208
rect 206940 151196 206946 151208
rect 210102 151196 210108 151208
rect 206940 151168 210108 151196
rect 206940 151156 206946 151168
rect 210102 151156 210108 151168
rect 210160 151156 210166 151208
rect 26010 151088 26016 151140
rect 26068 151128 26074 151140
rect 27298 151128 27304 151140
rect 26068 151100 27304 151128
rect 26068 151088 26074 151100
rect 27298 151088 27304 151100
rect 27356 151088 27362 151140
rect 35302 151088 35308 151140
rect 35360 151128 35366 151140
rect 36038 151128 36044 151140
rect 35360 151100 36044 151128
rect 35360 151088 35366 151100
rect 36038 151088 36044 151100
rect 36096 151088 36102 151140
rect 199614 151088 199620 151140
rect 199672 151128 199678 151140
rect 200166 151128 200172 151140
rect 199672 151100 200172 151128
rect 199672 151088 199678 151100
rect 200166 151088 200172 151100
rect 200224 151088 200230 151140
rect 25918 151020 25924 151072
rect 25976 151060 25982 151072
rect 26838 151060 26844 151072
rect 25976 151032 26844 151060
rect 25976 151020 25982 151032
rect 26838 151020 26844 151032
rect 26896 151020 26902 151072
rect 27666 151020 27672 151072
rect 27724 151060 27730 151072
rect 30058 151060 30064 151072
rect 27724 151032 30064 151060
rect 27724 151020 27730 151032
rect 30058 151020 30064 151032
rect 30116 151020 30122 151072
rect 40822 151020 40828 151072
rect 40880 151060 40886 151072
rect 45054 151060 45060 151072
rect 40880 151032 45060 151060
rect 40880 151020 40886 151032
rect 45054 151020 45060 151032
rect 45112 151020 45118 151072
rect 111294 151060 111300 151072
rect 110576 151032 111300 151060
rect 25826 150952 25832 151004
rect 25884 150992 25890 151004
rect 26470 150992 26476 151004
rect 25884 150964 26476 150992
rect 25884 150952 25890 150964
rect 26470 150952 26476 150964
rect 26528 150952 26534 151004
rect 33462 150952 33468 151004
rect 33520 150992 33526 151004
rect 34106 150992 34112 151004
rect 33520 150964 34112 150992
rect 33520 150952 33526 150964
rect 34106 150952 34112 150964
rect 34164 150952 34170 151004
rect 109546 150952 109552 151004
rect 109604 150992 109610 151004
rect 110466 150992 110472 151004
rect 109604 150964 110472 150992
rect 109604 150952 109610 150964
rect 110466 150952 110472 150964
rect 110524 150952 110530 151004
rect 110466 150816 110472 150868
rect 110524 150856 110530 150868
rect 110576 150856 110604 151032
rect 111294 151020 111300 151032
rect 111352 151020 111358 151072
rect 112490 151060 112496 151072
rect 112048 151032 112496 151060
rect 111662 150992 111668 151004
rect 110668 150964 111668 150992
rect 110668 150936 110696 150964
rect 111662 150952 111668 150964
rect 111720 150952 111726 151004
rect 112048 150936 112076 151032
rect 112490 151020 112496 151032
rect 112548 151020 112554 151072
rect 120862 151020 120868 151072
rect 120920 151060 120926 151072
rect 123806 151060 123812 151072
rect 120920 151032 123812 151060
rect 120920 151020 120926 151032
rect 123806 151020 123812 151032
rect 123864 151020 123870 151072
rect 125278 151020 125284 151072
rect 125336 151060 125342 151072
rect 129326 151060 129332 151072
rect 125336 151032 129332 151060
rect 125336 151020 125342 151032
rect 129326 151020 129332 151032
rect 129384 151020 129390 151072
rect 196854 151060 196860 151072
rect 196228 151032 196860 151060
rect 112122 150952 112128 151004
rect 112180 150992 112186 151004
rect 112858 150992 112864 151004
rect 112180 150964 112864 150992
rect 112180 150952 112186 150964
rect 112858 150952 112864 150964
rect 112916 150952 112922 151004
rect 115618 150952 115624 151004
rect 115676 150992 115682 151004
rect 115986 150992 115992 151004
rect 115676 150964 115992 150992
rect 115676 150952 115682 150964
rect 115986 150952 115992 150964
rect 116044 150952 116050 151004
rect 116446 150952 116452 151004
rect 116504 150992 116510 151004
rect 117458 150992 117464 151004
rect 116504 150964 117464 150992
rect 116504 150952 116510 150964
rect 117458 150952 117464 150964
rect 117516 150952 117522 151004
rect 117642 150952 117648 151004
rect 117700 150992 117706 151004
rect 118838 150992 118844 151004
rect 117700 150964 118844 150992
rect 117700 150952 117706 150964
rect 118838 150952 118844 150964
rect 118896 150952 118902 151004
rect 122058 150952 122064 151004
rect 122116 150992 122122 151004
rect 125186 150992 125192 151004
rect 122116 150964 125192 150992
rect 122116 150952 122122 150964
rect 125186 150952 125192 150964
rect 125244 150952 125250 151004
rect 194738 150952 194744 151004
rect 194796 150992 194802 151004
rect 195014 150992 195020 151004
rect 194796 150964 195020 150992
rect 194796 150952 194802 150964
rect 195014 150952 195020 150964
rect 195072 150952 195078 151004
rect 196228 150936 196256 151032
rect 196854 151020 196860 151032
rect 196912 151020 196918 151072
rect 208446 151020 208452 151072
rect 208504 151060 208510 151072
rect 210654 151060 210660 151072
rect 208504 151032 210660 151060
rect 208504 151020 208510 151032
rect 210654 151020 210660 151032
rect 210712 151020 210718 151072
rect 204030 150952 204036 151004
rect 204088 150992 204094 151004
rect 206238 150992 206244 151004
rect 204088 150964 206244 150992
rect 204088 150952 204094 150964
rect 206238 150952 206244 150964
rect 206296 150952 206302 151004
rect 207526 150952 207532 151004
rect 207584 150992 207590 151004
rect 210838 150992 210844 151004
rect 207584 150964 210844 150992
rect 207584 150952 207590 150964
rect 210838 150952 210844 150964
rect 210896 150952 210902 151004
rect 110650 150884 110656 150936
rect 110708 150884 110714 150936
rect 112030 150884 112036 150936
rect 112088 150884 112094 150936
rect 196210 150884 196216 150936
rect 196268 150884 196274 150936
rect 110524 150828 110604 150856
rect 110524 150816 110530 150828
rect 59222 146804 59228 146856
rect 59280 146804 59286 146856
rect 59240 146776 59268 146804
rect 59406 146776 59412 146788
rect 59240 146748 59412 146776
rect 59406 146736 59412 146748
rect 59464 146736 59470 146788
rect 127210 146124 127216 146176
rect 127268 146164 127274 146176
rect 127670 146164 127676 146176
rect 127268 146136 127676 146164
rect 127268 146124 127274 146136
rect 127670 146124 127676 146136
rect 127728 146124 127734 146176
rect 197590 146124 197596 146176
rect 197648 146164 197654 146176
rect 198142 146164 198148 146176
rect 197648 146136 198148 146164
rect 197648 146124 197654 146136
rect 198142 146124 198148 146136
rect 198200 146124 198206 146176
rect 40178 144016 40184 144068
rect 40236 144056 40242 144068
rect 43030 144056 43036 144068
rect 40236 144028 43036 144056
rect 40236 144016 40242 144028
rect 43030 144016 43036 144028
rect 43088 144016 43094 144068
rect 59406 144056 59412 144068
rect 59367 144028 59412 144056
rect 59406 144016 59412 144028
rect 59464 144016 59470 144068
rect 118838 144016 118844 144068
rect 118896 144056 118902 144068
rect 119574 144056 119580 144068
rect 118896 144028 119580 144056
rect 118896 144016 118902 144028
rect 119574 144016 119580 144028
rect 119632 144016 119638 144068
rect 120954 144016 120960 144068
rect 121012 144056 121018 144068
rect 121690 144056 121696 144068
rect 121012 144028 121696 144056
rect 121012 144016 121018 144028
rect 121690 144016 121696 144028
rect 121748 144016 121754 144068
rect 123806 144016 123812 144068
rect 123864 144056 123870 144068
rect 124450 144056 124456 144068
rect 123864 144028 124456 144056
rect 123864 144016 123870 144028
rect 124450 144016 124456 144028
rect 124508 144016 124514 144068
rect 125186 144016 125192 144068
rect 125244 144056 125250 144068
rect 126014 144056 126020 144068
rect 125244 144028 126020 144056
rect 125244 144016 125250 144028
rect 126014 144016 126020 144028
rect 126072 144016 126078 144068
rect 127946 144016 127952 144068
rect 128004 144056 128010 144068
rect 128590 144056 128596 144068
rect 128004 144028 128596 144056
rect 128004 144016 128010 144028
rect 128590 144016 128596 144028
rect 128648 144016 128654 144068
rect 129234 144016 129240 144068
rect 129292 144056 129298 144068
rect 130062 144056 130068 144068
rect 129292 144028 130068 144056
rect 129292 144016 129298 144028
rect 130062 144016 130068 144028
rect 130120 144016 130126 144068
rect 183606 144016 183612 144068
rect 183664 144056 183670 144068
rect 187930 144056 187936 144068
rect 183664 144028 187936 144056
rect 183664 144016 183670 144028
rect 187930 144016 187936 144028
rect 187988 144016 187994 144068
rect 193082 144016 193088 144068
rect 193140 144056 193146 144068
rect 193358 144056 193364 144068
rect 193140 144028 193364 144056
rect 193140 144016 193146 144028
rect 193358 144016 193364 144028
rect 193416 144016 193422 144068
rect 198418 144016 198424 144068
rect 198476 144056 198482 144068
rect 199062 144056 199068 144068
rect 198476 144028 199068 144056
rect 198476 144016 198482 144028
rect 199062 144016 199068 144028
rect 199120 144016 199126 144068
rect 201178 144016 201184 144068
rect 201236 144056 201242 144068
rect 201730 144056 201736 144068
rect 201236 144028 201736 144056
rect 201236 144016 201242 144028
rect 201730 144016 201736 144028
rect 201788 144016 201794 144068
rect 202926 144016 202932 144068
rect 202984 144056 202990 144068
rect 203846 144056 203852 144068
rect 202984 144028 203852 144056
rect 202984 144016 202990 144028
rect 203846 144016 203852 144028
rect 203904 144016 203910 144068
rect 39902 143948 39908 144000
rect 39960 143988 39966 144000
rect 42294 143988 42300 144000
rect 39960 143960 42300 143988
rect 39960 143948 39966 143960
rect 42294 143948 42300 143960
rect 42352 143948 42358 144000
rect 123714 143948 123720 144000
rect 123772 143988 123778 144000
rect 124542 143988 124548 144000
rect 123772 143960 124548 143988
rect 123772 143948 123778 143960
rect 124542 143948 124548 143960
rect 124600 143948 124606 144000
rect 125094 143948 125100 144000
rect 125152 143988 125158 144000
rect 126566 143988 126572 144000
rect 125152 143960 126572 143988
rect 125152 143948 125158 143960
rect 126566 143948 126572 143960
rect 126624 143948 126630 144000
rect 127854 143948 127860 144000
rect 127912 143988 127918 144000
rect 128682 143988 128688 144000
rect 127912 143960 128688 143988
rect 127912 143948 127918 143960
rect 128682 143948 128688 143960
rect 128740 143948 128746 144000
rect 129326 143948 129332 144000
rect 129384 143988 129390 144000
rect 130614 143988 130620 144000
rect 129384 143960 130620 143988
rect 129384 143948 129390 143960
rect 130614 143948 130620 143960
rect 130672 143948 130678 144000
rect 183422 143948 183428 144000
rect 183480 143988 183486 144000
rect 189402 143988 189408 144000
rect 183480 143960 189408 143988
rect 183480 143948 183486 143960
rect 189402 143948 189408 143960
rect 189460 143948 189466 144000
rect 198878 143948 198884 144000
rect 198936 143988 198942 144000
rect 199246 143988 199252 144000
rect 198936 143960 199252 143988
rect 198936 143948 198942 143960
rect 199246 143948 199252 143960
rect 199304 143948 199310 144000
rect 201270 143948 201276 144000
rect 201328 143988 201334 144000
rect 202742 143988 202748 144000
rect 201328 143960 202748 143988
rect 201328 143948 201334 143960
rect 202742 143948 202748 143960
rect 202800 143948 202806 144000
rect 203018 143948 203024 144000
rect 203076 143988 203082 144000
rect 204950 143988 204956 144000
rect 203076 143960 204956 143988
rect 203076 143948 203082 143960
rect 204950 143948 204956 143960
rect 205008 143948 205014 144000
rect 40086 143880 40092 143932
rect 40144 143920 40150 143932
rect 44410 143920 44416 143932
rect 40144 143892 44416 143920
rect 40144 143880 40150 143892
rect 44410 143880 44416 143892
rect 44468 143880 44474 143932
rect 117274 143880 117280 143932
rect 117332 143920 117338 143932
rect 119022 143920 119028 143932
rect 117332 143892 119028 143920
rect 117332 143880 117338 143892
rect 119022 143880 119028 143892
rect 119080 143880 119086 143932
rect 183514 143880 183520 143932
rect 183572 143920 183578 143932
rect 189494 143920 189500 143932
rect 183572 143892 189500 143920
rect 183572 143880 183578 143892
rect 189494 143880 189500 143892
rect 189552 143880 189558 143932
rect 200810 143880 200816 143932
rect 200868 143920 200874 143932
rect 202282 143920 202288 143932
rect 200868 143892 202288 143920
rect 200868 143880 200874 143892
rect 202282 143880 202288 143892
rect 202340 143880 202346 143932
rect 202466 143880 202472 143932
rect 202524 143920 202530 143932
rect 204490 143920 204496 143932
rect 202524 143892 204496 143920
rect 202524 143880 202530 143892
rect 204490 143880 204496 143892
rect 204548 143880 204554 143932
rect 23250 143812 23256 143864
rect 23308 143852 23314 143864
rect 26010 143852 26016 143864
rect 23308 143824 26016 143852
rect 23308 143812 23314 143824
rect 26010 143812 26016 143824
rect 26068 143812 26074 143864
rect 39626 143812 39632 143864
rect 39684 143852 39690 143864
rect 43766 143852 43772 143864
rect 39684 143824 43772 143852
rect 39684 143812 39690 143824
rect 43766 143812 43772 143824
rect 43824 143812 43830 143864
rect 183330 143812 183336 143864
rect 183388 143852 183394 143864
rect 190046 143852 190052 143864
rect 183388 143824 190052 143852
rect 183388 143812 183394 143824
rect 190046 143812 190052 143824
rect 190104 143812 190110 143864
rect 201638 143812 201644 143864
rect 201696 143852 201702 143864
rect 203294 143852 203300 143864
rect 201696 143824 203300 143852
rect 201696 143812 201702 143824
rect 203294 143812 203300 143824
rect 203352 143812 203358 143864
rect 22146 143744 22152 143796
rect 22204 143784 22210 143796
rect 25918 143784 25924 143796
rect 22204 143756 25924 143784
rect 22204 143744 22210 143756
rect 25918 143744 25924 143756
rect 25976 143744 25982 143796
rect 24446 143676 24452 143728
rect 24504 143716 24510 143728
rect 24906 143716 24912 143728
rect 24504 143688 24912 143716
rect 24504 143676 24510 143688
rect 24906 143676 24912 143688
rect 24964 143676 24970 143728
rect 20766 143608 20772 143660
rect 20824 143648 20830 143660
rect 25090 143648 25096 143660
rect 20824 143620 25096 143648
rect 20824 143608 20830 143620
rect 25090 143608 25096 143620
rect 25148 143608 25154 143660
rect 26010 143608 26016 143660
rect 26068 143648 26074 143660
rect 26378 143648 26384 143660
rect 26068 143620 26384 143648
rect 26068 143608 26074 143620
rect 26378 143608 26384 143620
rect 26436 143608 26442 143660
rect 27298 143608 27304 143660
rect 27356 143648 27362 143660
rect 27758 143648 27764 143660
rect 27356 143620 27764 143648
rect 27356 143608 27362 143620
rect 27758 143608 27764 143620
rect 27816 143608 27822 143660
rect 28586 143608 28592 143660
rect 28644 143648 28650 143660
rect 29046 143648 29052 143660
rect 28644 143620 29052 143648
rect 28644 143608 28650 143620
rect 29046 143608 29052 143620
rect 29104 143608 29110 143660
rect 30058 143608 30064 143660
rect 30116 143648 30122 143660
rect 30518 143648 30524 143660
rect 30116 143620 30524 143648
rect 30116 143608 30122 143620
rect 30518 143608 30524 143620
rect 30576 143608 30582 143660
rect 31990 143608 31996 143660
rect 32048 143648 32054 143660
rect 32726 143648 32732 143660
rect 32048 143620 32732 143648
rect 32048 143608 32054 143620
rect 32726 143608 32732 143620
rect 32784 143608 32790 143660
rect 34474 143608 34480 143660
rect 34532 143648 34538 143660
rect 34934 143648 34940 143660
rect 34532 143620 34940 143648
rect 34532 143608 34538 143620
rect 34934 143608 34940 143620
rect 34992 143608 34998 143660
rect 43674 143608 43680 143660
rect 43732 143648 43738 143660
rect 47170 143648 47176 143660
rect 43732 143620 47176 143648
rect 43732 143608 43738 143620
rect 47170 143608 47176 143620
rect 47228 143608 47234 143660
rect 114422 143608 114428 143660
rect 114480 143648 114486 143660
rect 114974 143648 114980 143660
rect 114480 143620 114980 143648
rect 114480 143608 114486 143620
rect 114974 143608 114980 143620
rect 115032 143608 115038 143660
rect 115986 143608 115992 143660
rect 116044 143648 116050 143660
rect 116630 143648 116636 143660
rect 116044 143620 116636 143648
rect 116044 143608 116050 143620
rect 116630 143608 116636 143620
rect 116688 143608 116694 143660
rect 117458 143608 117464 143660
rect 117516 143648 117522 143660
rect 117918 143648 117924 143660
rect 117516 143620 117924 143648
rect 117516 143608 117522 143620
rect 117918 143608 117924 143620
rect 117976 143608 117982 143660
rect 205962 143608 205968 143660
rect 206020 143648 206026 143660
rect 206146 143648 206152 143660
rect 206020 143620 206152 143648
rect 206020 143608 206026 143620
rect 206146 143608 206152 143620
rect 206204 143608 206210 143660
rect 207986 143608 207992 143660
rect 208044 143648 208050 143660
rect 208630 143648 208636 143660
rect 208044 143620 208636 143648
rect 208044 143608 208050 143620
rect 208630 143608 208636 143620
rect 208688 143608 208694 143660
rect 208814 143608 208820 143660
rect 208872 143648 208878 143660
rect 209550 143648 209556 143660
rect 208872 143620 209556 143648
rect 208872 143608 208878 143620
rect 209550 143608 209556 143620
rect 209608 143608 209614 143660
rect 210838 143608 210844 143660
rect 210896 143648 210902 143660
rect 211390 143648 211396 143660
rect 210896 143620 211396 143648
rect 210896 143608 210902 143620
rect 211390 143608 211396 143620
rect 211448 143608 211454 143660
rect 214242 143608 214248 143660
rect 214300 143648 214306 143660
rect 214702 143648 214708 143660
rect 214300 143620 214708 143648
rect 214300 143608 214306 143620
rect 214702 143608 214708 143620
rect 214760 143608 214766 143660
rect 23526 143540 23532 143592
rect 23584 143580 23590 143592
rect 25734 143580 25740 143592
rect 23584 143552 25740 143580
rect 23584 143540 23590 143552
rect 25734 143540 25740 143552
rect 25792 143540 25798 143592
rect 34842 143540 34848 143592
rect 34900 143580 34906 143592
rect 35486 143580 35492 143592
rect 34900 143552 35492 143580
rect 34900 143540 34906 143552
rect 35486 143540 35492 143552
rect 35544 143540 35550 143592
rect 99242 143540 99248 143592
rect 99300 143580 99306 143592
rect 106602 143580 106608 143592
rect 99300 143552 106608 143580
rect 99300 143540 99306 143552
rect 106602 143540 106608 143552
rect 106660 143540 106666 143592
rect 114882 143540 114888 143592
rect 114940 143580 114946 143592
rect 115526 143580 115532 143592
rect 114940 143552 115532 143580
rect 114940 143540 114946 143552
rect 115526 143540 115532 143552
rect 115584 143540 115590 143592
rect 115894 143540 115900 143592
rect 115952 143580 115958 143592
rect 117642 143580 117648 143592
rect 115952 143552 117648 143580
rect 115952 143540 115958 143552
rect 117642 143540 117648 143552
rect 117700 143540 117706 143592
rect 207894 143540 207900 143592
rect 207952 143580 207958 143592
rect 208998 143580 209004 143592
rect 207952 143552 209004 143580
rect 207952 143540 207958 143552
rect 208998 143540 209004 143552
rect 209056 143540 209062 143592
rect 35670 143472 35676 143524
rect 35728 143512 35734 143524
rect 36958 143512 36964 143524
rect 35728 143484 36964 143512
rect 35728 143472 35734 143484
rect 36958 143472 36964 143484
rect 37016 143472 37022 143524
rect 99150 143472 99156 143524
rect 99208 143512 99214 143524
rect 106786 143512 106792 143524
rect 99208 143484 106792 143512
rect 99208 143472 99214 143484
rect 106786 143472 106792 143484
rect 106844 143472 106850 143524
rect 183238 143472 183244 143524
rect 183296 143512 183302 143524
rect 190782 143512 190788 143524
rect 183296 143484 190788 143512
rect 183296 143472 183302 143484
rect 190782 143472 190788 143484
rect 190840 143472 190846 143524
rect 99058 143404 99064 143456
rect 99116 143444 99122 143456
rect 107430 143444 107436 143456
rect 99116 143416 107436 143444
rect 99116 143404 99122 143416
rect 107430 143404 107436 143416
rect 107488 143404 107494 143456
rect 183054 143404 183060 143456
rect 183112 143444 183118 143456
rect 192070 143444 192076 143456
rect 183112 143416 192076 143444
rect 183112 143404 183118 143416
rect 192070 143404 192076 143416
rect 192128 143404 192134 143456
rect 194186 143404 194192 143456
rect 194244 143444 194250 143456
rect 194738 143444 194744 143456
rect 194244 143416 194744 143444
rect 194244 143404 194250 143416
rect 194738 143404 194744 143416
rect 194796 143404 194802 143456
rect 20490 143336 20496 143388
rect 20548 143376 20554 143388
rect 44502 143376 44508 143388
rect 20548 143348 44508 143376
rect 20548 143336 20554 143348
rect 44502 143336 44508 143348
rect 44560 143336 44566 143388
rect 98966 143336 98972 143388
rect 99024 143376 99030 143388
rect 107982 143376 107988 143388
rect 99024 143348 107988 143376
rect 99024 143336 99030 143348
rect 107982 143336 107988 143348
rect 108040 143336 108046 143388
rect 183146 143336 183152 143388
rect 183204 143376 183210 143388
rect 191334 143376 191340 143388
rect 183204 143348 191340 143376
rect 183204 143336 183210 143348
rect 191334 143336 191340 143348
rect 191392 143336 191398 143388
rect 191978 143336 191984 143388
rect 192036 143376 192042 143388
rect 215622 143376 215628 143388
rect 192036 143348 215628 143376
rect 192036 143336 192042 143348
rect 215622 143336 215628 143348
rect 215680 143336 215686 143388
rect 45146 143200 45152 143252
rect 45204 143240 45210 143252
rect 46526 143240 46532 143252
rect 45204 143212 46532 143240
rect 45204 143200 45210 143212
rect 46526 143200 46532 143212
rect 46584 143200 46590 143252
rect 110282 143200 110288 143252
rect 110340 143240 110346 143252
rect 110558 143240 110564 143252
rect 110340 143212 110564 143240
rect 110340 143200 110346 143212
rect 110558 143200 110564 143212
rect 110616 143200 110622 143252
rect 116814 143064 116820 143116
rect 116872 143104 116878 143116
rect 118470 143104 118476 143116
rect 116872 143076 118476 143104
rect 116872 143064 116878 143076
rect 118470 143064 118476 143076
rect 118528 143064 118534 143116
rect 210930 143064 210936 143116
rect 210988 143104 210994 143116
rect 211758 143104 211764 143116
rect 210988 143076 211764 143104
rect 210988 143064 210994 143076
rect 211758 143064 211764 143076
rect 211816 143064 211822 143116
rect 45054 142928 45060 142980
rect 45112 142968 45118 142980
rect 45790 142968 45796 142980
rect 45112 142940 45796 142968
rect 45112 142928 45118 142940
rect 45790 142928 45796 142940
rect 45848 142928 45854 142980
rect 98782 142928 98788 142980
rect 98840 142968 98846 142980
rect 103934 142968 103940 142980
rect 98840 142940 103940 142968
rect 98840 142928 98846 142940
rect 103934 142928 103940 142940
rect 103992 142928 103998 142980
rect 210654 142928 210660 142980
rect 210712 142968 210718 142980
rect 212862 142968 212868 142980
rect 210712 142940 212868 142968
rect 210712 142928 210718 142940
rect 212862 142928 212868 142940
rect 212920 142928 212926 142980
rect 99426 142860 99432 142912
rect 99484 142900 99490 142912
rect 105590 142900 105596 142912
rect 99484 142872 105596 142900
rect 99484 142860 99490 142872
rect 105590 142860 105596 142872
rect 105648 142860 105654 142912
rect 200258 142860 200264 142912
rect 200316 142900 200322 142912
rect 200902 142900 200908 142912
rect 200316 142872 200908 142900
rect 200316 142860 200322 142872
rect 200902 142860 200908 142872
rect 200960 142860 200966 142912
rect 21778 142792 21784 142844
rect 21836 142832 21842 142844
rect 25826 142832 25832 142844
rect 21836 142804 25832 142832
rect 21836 142792 21842 142804
rect 25826 142792 25832 142804
rect 25884 142792 25890 142844
rect 31346 142792 31352 142844
rect 31404 142832 31410 142844
rect 31898 142832 31904 142844
rect 31404 142804 31904 142832
rect 31404 142792 31410 142804
rect 31898 142792 31904 142804
rect 31956 142792 31962 142844
rect 37418 142792 37424 142844
rect 37476 142832 37482 142844
rect 38246 142832 38252 142844
rect 37476 142804 38252 142832
rect 37476 142792 37482 142804
rect 38246 142792 38252 142804
rect 38304 142792 38310 142844
rect 99334 142792 99340 142844
rect 99392 142832 99398 142844
rect 105130 142832 105136 142844
rect 99392 142804 105136 142832
rect 99392 142792 99398 142804
rect 105130 142792 105136 142804
rect 105188 142792 105194 142844
rect 210746 142792 210752 142844
rect 210804 142832 210810 142844
rect 212310 142832 212316 142844
rect 210804 142804 212316 142832
rect 210804 142792 210810 142804
rect 212310 142792 212316 142804
rect 212368 142792 212374 142844
rect 99518 142724 99524 142776
rect 99576 142764 99582 142776
rect 104578 142764 104584 142776
rect 99576 142736 104584 142764
rect 99576 142724 99582 142736
rect 104578 142724 104584 142736
rect 104636 142724 104642 142776
rect 68698 142656 68704 142708
rect 68756 142696 68762 142708
rect 69158 142696 69164 142708
rect 68756 142668 69164 142696
rect 68756 142656 68762 142668
rect 69158 142656 69164 142668
rect 69216 142656 69222 142708
rect 167690 142452 167696 142504
rect 167748 142492 167754 142504
rect 169898 142492 169904 142504
rect 167748 142464 169904 142492
rect 167748 142452 167754 142464
rect 169898 142452 169904 142464
rect 169956 142452 169962 142504
rect 134846 140004 134852 140056
rect 134904 140044 134910 140056
rect 143586 140044 143592 140056
rect 134904 140016 143592 140044
rect 134904 140004 134910 140016
rect 143586 140004 143592 140016
rect 143644 140004 143650 140056
rect 49930 139936 49936 139988
rect 49988 139976 49994 139988
rect 56186 139976 56192 139988
rect 49988 139948 56192 139976
rect 49988 139936 49994 139948
rect 56186 139936 56192 139948
rect 56244 139936 56250 139988
rect 135398 139936 135404 139988
rect 135456 139976 135462 139988
rect 143310 139976 143316 139988
rect 135456 139948 143316 139976
rect 135456 139936 135462 139948
rect 143310 139936 143316 139948
rect 143368 139936 143374 139988
rect 135398 138712 135404 138764
rect 135456 138752 135462 138764
rect 139814 138752 139820 138764
rect 135456 138724 139820 138752
rect 135456 138712 135462 138724
rect 139814 138712 139820 138724
rect 139872 138712 139878 138764
rect 49930 138644 49936 138696
rect 49988 138684 49994 138696
rect 58486 138684 58492 138696
rect 49988 138656 58492 138684
rect 49988 138644 49994 138656
rect 58486 138644 58492 138656
rect 58544 138644 58550 138696
rect 50022 138576 50028 138628
rect 50080 138616 50086 138628
rect 58394 138616 58400 138628
rect 50080 138588 58400 138616
rect 50080 138576 50086 138588
rect 58394 138576 58400 138588
rect 58452 138576 58458 138628
rect 134662 138576 134668 138628
rect 134720 138616 134726 138628
rect 139630 138616 139636 138628
rect 134720 138588 139636 138616
rect 134720 138576 134726 138588
rect 139630 138576 139636 138588
rect 139688 138576 139694 138628
rect 51402 138508 51408 138560
rect 51460 138548 51466 138560
rect 59222 138548 59228 138560
rect 51460 138520 59228 138548
rect 51460 138508 51466 138520
rect 59222 138508 59228 138520
rect 59280 138508 59286 138560
rect 92710 138508 92716 138560
rect 92768 138548 92774 138560
rect 100806 138548 100812 138560
rect 92768 138520 100812 138548
rect 92768 138508 92774 138520
rect 100806 138508 100812 138520
rect 100864 138508 100870 138560
rect 177626 138508 177632 138560
rect 177684 138548 177690 138560
rect 185078 138548 185084 138560
rect 177684 138520 185084 138548
rect 177684 138508 177690 138520
rect 185078 138508 185084 138520
rect 185136 138508 185142 138560
rect 56186 138440 56192 138492
rect 56244 138480 56250 138492
rect 58670 138480 58676 138492
rect 56244 138452 58676 138480
rect 56244 138440 56250 138452
rect 58670 138440 58676 138452
rect 58728 138440 58734 138492
rect 92802 138440 92808 138492
rect 92860 138480 92866 138492
rect 100898 138480 100904 138492
rect 92860 138452 100904 138480
rect 92860 138440 92866 138452
rect 100898 138440 100904 138452
rect 100956 138440 100962 138492
rect 177718 138440 177724 138492
rect 177776 138480 177782 138492
rect 184986 138480 184992 138492
rect 177776 138452 184992 138480
rect 177776 138440 177782 138452
rect 184986 138440 184992 138452
rect 185044 138440 185050 138492
rect 134662 137352 134668 137404
rect 134720 137392 134726 137404
rect 139722 137392 139728 137404
rect 134720 137364 139728 137392
rect 134720 137352 134726 137364
rect 139722 137352 139728 137364
rect 139780 137352 139786 137404
rect 97862 137284 97868 137336
rect 97920 137324 97926 137336
rect 100990 137324 100996 137336
rect 97920 137296 100996 137324
rect 97920 137284 97926 137296
rect 100990 137284 100996 137296
rect 101048 137284 101054 137336
rect 49930 137216 49936 137268
rect 49988 137256 49994 137268
rect 58302 137256 58308 137268
rect 49988 137228 58308 137256
rect 49988 137216 49994 137228
rect 58302 137216 58308 137228
rect 58360 137216 58366 137268
rect 97954 137216 97960 137268
rect 98012 137256 98018 137268
rect 101266 137256 101272 137268
rect 98012 137228 101272 137256
rect 98012 137216 98018 137228
rect 101266 137216 101272 137228
rect 101324 137216 101330 137268
rect 181582 137216 181588 137268
rect 181640 137256 181646 137268
rect 185170 137256 185176 137268
rect 181640 137228 185176 137256
rect 181640 137216 181646 137228
rect 185170 137216 185176 137228
rect 185228 137216 185234 137268
rect 50022 137148 50028 137200
rect 50080 137188 50086 137200
rect 50080 137160 56784 137188
rect 50080 137148 50086 137160
rect 56756 137120 56784 137160
rect 135398 137148 135404 137200
rect 135456 137188 135462 137200
rect 143402 137188 143408 137200
rect 135456 137160 143408 137188
rect 135456 137148 135462 137160
rect 143402 137148 143408 137160
rect 143460 137148 143466 137200
rect 182226 137148 182232 137200
rect 182284 137188 182290 137200
rect 185446 137188 185452 137200
rect 182284 137160 185452 137188
rect 182284 137148 182290 137160
rect 185446 137148 185452 137160
rect 185504 137148 185510 137200
rect 58210 137120 58216 137132
rect 56756 137092 58216 137120
rect 58210 137080 58216 137092
rect 58268 137080 58274 137132
rect 92710 137080 92716 137132
rect 92768 137120 92774 137132
rect 101174 137120 101180 137132
rect 92768 137092 101180 137120
rect 92768 137080 92774 137092
rect 101174 137080 101180 137092
rect 101232 137080 101238 137132
rect 177626 137080 177632 137132
rect 177684 137120 177690 137132
rect 185262 137120 185268 137132
rect 177684 137092 185268 137120
rect 177684 137080 177690 137092
rect 185262 137080 185268 137092
rect 185320 137080 185326 137132
rect 92802 137012 92808 137064
rect 92860 137052 92866 137064
rect 101082 137052 101088 137064
rect 92860 137024 101088 137052
rect 92860 137012 92866 137024
rect 101082 137012 101088 137024
rect 101140 137012 101146 137064
rect 139630 137012 139636 137064
rect 139688 137052 139694 137064
rect 143586 137052 143592 137064
rect 139688 137024 143592 137052
rect 139688 137012 139694 137024
rect 143586 137012 143592 137024
rect 143644 137012 143650 137064
rect 177718 137012 177724 137064
rect 177776 137052 177782 137064
rect 185354 137052 185360 137064
rect 177776 137024 185360 137052
rect 177776 137012 177782 137024
rect 185354 137012 185360 137024
rect 185412 137012 185418 137064
rect 92710 136944 92716 136996
rect 92768 136984 92774 136996
rect 97862 136984 97868 136996
rect 92768 136956 97868 136984
rect 92768 136944 92774 136956
rect 97862 136944 97868 136956
rect 97920 136944 97926 136996
rect 139814 136944 139820 136996
rect 139872 136984 139878 136996
rect 143126 136984 143132 136996
rect 139872 136956 143132 136984
rect 139872 136944 139878 136956
rect 143126 136944 143132 136956
rect 143184 136944 143190 136996
rect 139722 136604 139728 136656
rect 139780 136644 139786 136656
rect 143494 136644 143500 136656
rect 139780 136616 143500 136644
rect 139780 136604 139786 136616
rect 143494 136604 143500 136616
rect 143552 136604 143558 136656
rect 177718 136604 177724 136656
rect 177776 136644 177782 136656
rect 181582 136644 181588 136656
rect 177776 136616 181588 136644
rect 177776 136604 177782 136616
rect 181582 136604 181588 136616
rect 181640 136604 181646 136656
rect 51218 136128 51224 136180
rect 51276 136168 51282 136180
rect 52782 136168 52788 136180
rect 51276 136140 52788 136168
rect 51276 136128 51282 136140
rect 52782 136128 52788 136140
rect 52840 136128 52846 136180
rect 51218 135992 51224 136044
rect 51276 136032 51282 136044
rect 52690 136032 52696 136044
rect 51276 136004 52696 136032
rect 51276 135992 51282 136004
rect 52690 135992 52696 136004
rect 52748 135992 52754 136044
rect 135030 135924 135036 135976
rect 135088 135964 135094 135976
rect 143310 135964 143316 135976
rect 135088 135936 143316 135964
rect 135088 135924 135094 135936
rect 143310 135924 143316 135936
rect 143368 135924 143374 135976
rect 98046 135856 98052 135908
rect 98104 135896 98110 135908
rect 101450 135896 101456 135908
rect 98104 135868 101456 135896
rect 98104 135856 98110 135868
rect 101450 135856 101456 135868
rect 101508 135856 101514 135908
rect 135306 135856 135312 135908
rect 135364 135896 135370 135908
rect 143586 135896 143592 135908
rect 135364 135868 143592 135896
rect 135364 135856 135370 135868
rect 143586 135856 143592 135868
rect 143644 135856 143650 135908
rect 182318 135856 182324 135908
rect 182376 135896 182382 135908
rect 185354 135896 185360 135908
rect 182376 135868 185360 135896
rect 182376 135856 182382 135868
rect 185354 135856 185360 135868
rect 185412 135856 185418 135908
rect 50390 135788 50396 135840
rect 50448 135828 50454 135840
rect 50448 135800 56784 135828
rect 50448 135788 50454 135800
rect 56756 135760 56784 135800
rect 98138 135788 98144 135840
rect 98196 135828 98202 135840
rect 101726 135828 101732 135840
rect 98196 135800 101732 135828
rect 98196 135788 98202 135800
rect 101726 135788 101732 135800
rect 101784 135788 101790 135840
rect 135398 135788 135404 135840
rect 135456 135828 135462 135840
rect 143218 135828 143224 135840
rect 135456 135800 143224 135828
rect 135456 135788 135462 135800
rect 143218 135788 143224 135800
rect 143276 135788 143282 135840
rect 181950 135788 181956 135840
rect 182008 135828 182014 135840
rect 185262 135828 185268 135840
rect 182008 135800 185268 135828
rect 182008 135788 182014 135800
rect 185262 135788 185268 135800
rect 185320 135788 185326 135840
rect 58210 135760 58216 135772
rect 56756 135732 58216 135760
rect 58210 135720 58216 135732
rect 58268 135720 58274 135772
rect 92802 135720 92808 135772
rect 92860 135760 92866 135772
rect 101818 135760 101824 135772
rect 92860 135732 101824 135760
rect 92860 135720 92866 135732
rect 101818 135720 101824 135732
rect 101876 135720 101882 135772
rect 177626 135720 177632 135772
rect 177684 135760 177690 135772
rect 185170 135760 185176 135772
rect 177684 135732 185176 135760
rect 177684 135720 177690 135732
rect 185170 135720 185176 135732
rect 185228 135720 185234 135772
rect 92710 135652 92716 135704
rect 92768 135692 92774 135704
rect 97954 135692 97960 135704
rect 92768 135664 97960 135692
rect 92768 135652 92774 135664
rect 97954 135652 97960 135664
rect 98012 135652 98018 135704
rect 177718 135652 177724 135704
rect 177776 135692 177782 135704
rect 182226 135692 182232 135704
rect 177776 135664 182232 135692
rect 177776 135652 177782 135664
rect 182226 135652 182232 135664
rect 182284 135652 182290 135704
rect 51218 134564 51224 134616
rect 51276 134604 51282 134616
rect 56738 134604 56744 134616
rect 51276 134576 56744 134604
rect 51276 134564 51282 134576
rect 56738 134564 56744 134576
rect 56796 134564 56802 134616
rect 134662 134564 134668 134616
rect 134720 134604 134726 134616
rect 136870 134604 136876 134616
rect 134720 134576 136876 134604
rect 134720 134564 134726 134576
rect 136870 134564 136876 134576
rect 136928 134564 136934 134616
rect 51126 134496 51132 134548
rect 51184 134536 51190 134548
rect 52874 134536 52880 134548
rect 51184 134508 52880 134536
rect 51184 134496 51190 134508
rect 52874 134496 52880 134508
rect 52932 134496 52938 134548
rect 59406 134536 59412 134548
rect 59367 134508 59412 134536
rect 59406 134496 59412 134508
rect 59464 134496 59470 134548
rect 134846 134496 134852 134548
rect 134904 134536 134910 134548
rect 139630 134536 139636 134548
rect 134904 134508 139636 134536
rect 134904 134496 134910 134508
rect 139630 134496 139636 134508
rect 139688 134496 139694 134548
rect 52782 134360 52788 134412
rect 52840 134400 52846 134412
rect 58210 134400 58216 134412
rect 52840 134372 58216 134400
rect 52840 134360 52846 134372
rect 58210 134360 58216 134372
rect 58268 134360 58274 134412
rect 92894 134360 92900 134412
rect 92952 134400 92958 134412
rect 101450 134400 101456 134412
rect 92952 134372 101456 134400
rect 92952 134360 92958 134372
rect 101450 134360 101456 134372
rect 101508 134360 101514 134412
rect 177626 134360 177632 134412
rect 177684 134400 177690 134412
rect 185170 134400 185176 134412
rect 177684 134372 185176 134400
rect 177684 134360 177690 134372
rect 185170 134360 185176 134372
rect 185228 134360 185234 134412
rect 52690 134292 52696 134344
rect 52748 134332 52754 134344
rect 58302 134332 58308 134344
rect 52748 134304 58308 134332
rect 52748 134292 52754 134304
rect 58302 134292 58308 134304
rect 58360 134292 58366 134344
rect 92710 134292 92716 134344
rect 92768 134332 92774 134344
rect 98046 134332 98052 134344
rect 92768 134304 98052 134332
rect 92768 134292 92774 134304
rect 98046 134292 98052 134304
rect 98104 134292 98110 134344
rect 177718 134292 177724 134344
rect 177776 134332 177782 134344
rect 181950 134332 181956 134344
rect 177776 134304 181956 134332
rect 177776 134292 177782 134304
rect 181950 134292 181956 134304
rect 182008 134292 182014 134344
rect 92802 134224 92808 134276
rect 92860 134264 92866 134276
rect 98138 134264 98144 134276
rect 92860 134236 98144 134264
rect 92860 134224 92866 134236
rect 98138 134224 98144 134236
rect 98196 134224 98202 134276
rect 177718 134020 177724 134072
rect 177776 134060 177782 134072
rect 182318 134060 182324 134072
rect 177776 134032 182324 134060
rect 177776 134020 177782 134032
rect 182318 134020 182324 134032
rect 182376 134020 182382 134072
rect 56738 133816 56744 133868
rect 56796 133856 56802 133868
rect 58210 133856 58216 133868
rect 56796 133828 58216 133856
rect 56796 133816 56802 133828
rect 58210 133816 58216 133828
rect 58268 133816 58274 133868
rect 139630 133748 139636 133800
rect 139688 133788 139694 133800
rect 142942 133788 142948 133800
rect 139688 133760 142948 133788
rect 139688 133748 139694 133760
rect 142942 133748 142948 133760
rect 143000 133748 143006 133800
rect 50942 133068 50948 133120
rect 51000 133108 51006 133120
rect 52690 133108 52696 133120
rect 51000 133080 52696 133108
rect 51000 133068 51006 133080
rect 52690 133068 52696 133080
rect 52748 133068 52754 133120
rect 134110 133068 134116 133120
rect 134168 133108 134174 133120
rect 138158 133108 138164 133120
rect 134168 133080 138164 133108
rect 134168 133068 134174 133080
rect 138158 133068 138164 133080
rect 138216 133068 138222 133120
rect 50206 133000 50212 133052
rect 50264 133040 50270 133052
rect 56094 133040 56100 133052
rect 50264 133012 56100 133040
rect 50264 133000 50270 133012
rect 56094 133000 56100 133012
rect 56152 133000 56158 133052
rect 135398 133000 135404 133052
rect 135456 133040 135462 133052
rect 135456 133012 139676 133040
rect 135456 133000 135462 133012
rect 52874 132932 52880 132984
rect 52932 132972 52938 132984
rect 58210 132972 58216 132984
rect 52932 132944 58216 132972
rect 52932 132932 52938 132944
rect 58210 132932 58216 132944
rect 58268 132932 58274 132984
rect 59317 132975 59375 132981
rect 59317 132941 59329 132975
rect 59363 132972 59375 132975
rect 59406 132972 59412 132984
rect 59363 132944 59412 132972
rect 59363 132941 59375 132944
rect 59317 132935 59375 132941
rect 59406 132932 59412 132944
rect 59464 132932 59470 132984
rect 92802 132932 92808 132984
rect 92860 132972 92866 132984
rect 101818 132972 101824 132984
rect 92860 132944 101824 132972
rect 92860 132932 92866 132944
rect 101818 132932 101824 132944
rect 101876 132932 101882 132984
rect 139648 132972 139676 133012
rect 143218 132972 143224 132984
rect 139648 132944 143224 132972
rect 143218 132932 143224 132944
rect 143276 132932 143282 132984
rect 177626 132932 177632 132984
rect 177684 132972 177690 132984
rect 185170 132972 185176 132984
rect 177684 132944 185176 132972
rect 177684 132932 177690 132944
rect 185170 132932 185176 132944
rect 185228 132932 185234 132984
rect 92710 132864 92716 132916
rect 92768 132904 92774 132916
rect 100898 132904 100904 132916
rect 92768 132876 100904 132904
rect 92768 132864 92774 132876
rect 100898 132864 100904 132876
rect 100956 132864 100962 132916
rect 177718 132864 177724 132916
rect 177776 132904 177782 132916
rect 185078 132904 185084 132916
rect 177776 132876 185084 132904
rect 177776 132864 177782 132876
rect 185078 132864 185084 132876
rect 185136 132864 185142 132916
rect 136870 132796 136876 132848
rect 136928 132836 136934 132848
rect 143586 132836 143592 132848
rect 136928 132808 143592 132836
rect 136928 132796 136934 132808
rect 143586 132796 143592 132808
rect 143644 132796 143650 132848
rect 56094 132388 56100 132440
rect 56152 132428 56158 132440
rect 58302 132428 58308 132440
rect 56152 132400 58308 132428
rect 56152 132388 56158 132400
rect 58302 132388 58308 132400
rect 58360 132388 58366 132440
rect 50390 131980 50396 132032
rect 50448 132020 50454 132032
rect 53426 132020 53432 132032
rect 50448 131992 53432 132020
rect 50448 131980 50454 131992
rect 53426 131980 53432 131992
rect 53484 131980 53490 132032
rect 51218 131912 51224 131964
rect 51276 131952 51282 131964
rect 55450 131952 55456 131964
rect 51276 131924 55456 131952
rect 51276 131912 51282 131924
rect 55450 131912 55456 131924
rect 55508 131912 55514 131964
rect 134478 131912 134484 131964
rect 134536 131952 134542 131964
rect 137146 131952 137152 131964
rect 134536 131924 137152 131952
rect 134536 131912 134542 131924
rect 137146 131912 137152 131924
rect 137204 131912 137210 131964
rect 135306 131708 135312 131760
rect 135364 131748 135370 131760
rect 137974 131748 137980 131760
rect 135364 131720 137980 131748
rect 135364 131708 135370 131720
rect 137974 131708 137980 131720
rect 138032 131708 138038 131760
rect 51218 131640 51224 131692
rect 51276 131680 51282 131692
rect 52782 131680 52788 131692
rect 51276 131652 52788 131680
rect 51276 131640 51282 131652
rect 52782 131640 52788 131652
rect 52840 131640 52846 131692
rect 135122 131640 135128 131692
rect 135180 131680 135186 131692
rect 135180 131652 140228 131680
rect 135180 131640 135186 131652
rect 52690 131572 52696 131624
rect 52748 131612 52754 131624
rect 58210 131612 58216 131624
rect 52748 131584 58216 131612
rect 52748 131572 52754 131584
rect 58210 131572 58216 131584
rect 58268 131572 58274 131624
rect 92710 131572 92716 131624
rect 92768 131612 92774 131624
rect 101726 131612 101732 131624
rect 92768 131584 101732 131612
rect 92768 131572 92774 131584
rect 101726 131572 101732 131584
rect 101784 131572 101790 131624
rect 140200 131612 140228 131652
rect 142482 131612 142488 131624
rect 140200 131584 142488 131612
rect 142482 131572 142488 131584
rect 142540 131572 142546 131624
rect 177626 131572 177632 131624
rect 177684 131612 177690 131624
rect 185906 131612 185912 131624
rect 177684 131584 185912 131612
rect 177684 131572 177690 131584
rect 185906 131572 185912 131584
rect 185964 131572 185970 131624
rect 92802 131504 92808 131556
rect 92860 131544 92866 131556
rect 101818 131544 101824 131556
rect 92860 131516 101824 131544
rect 92860 131504 92866 131516
rect 101818 131504 101824 131516
rect 101876 131504 101882 131556
rect 138158 131504 138164 131556
rect 138216 131544 138222 131556
rect 143586 131544 143592 131556
rect 138216 131516 143592 131544
rect 138216 131504 138222 131516
rect 143586 131504 143592 131516
rect 143644 131504 143650 131556
rect 177718 131504 177724 131556
rect 177776 131544 177782 131556
rect 185814 131544 185820 131556
rect 177776 131516 185820 131544
rect 177776 131504 177782 131516
rect 185814 131504 185820 131516
rect 185872 131504 185878 131556
rect 55450 131300 55456 131352
rect 55508 131340 55514 131352
rect 58302 131340 58308 131352
rect 55508 131312 58308 131340
rect 55508 131300 55514 131312
rect 58302 131300 58308 131312
rect 58360 131300 58366 131352
rect 51218 130688 51224 130740
rect 51276 130728 51282 130740
rect 52966 130728 52972 130740
rect 51276 130700 52972 130728
rect 51276 130688 51282 130700
rect 52966 130688 52972 130700
rect 53024 130688 53030 130740
rect 134662 130552 134668 130604
rect 134720 130592 134726 130604
rect 137606 130592 137612 130604
rect 134720 130564 137612 130592
rect 134720 130552 134726 130564
rect 137606 130552 137612 130564
rect 137664 130552 137670 130604
rect 51218 130280 51224 130332
rect 51276 130320 51282 130332
rect 52690 130320 52696 130332
rect 51276 130292 52696 130320
rect 51276 130280 51282 130292
rect 52690 130280 52696 130292
rect 52748 130280 52754 130332
rect 134846 130280 134852 130332
rect 134904 130320 134910 130332
rect 137422 130320 137428 130332
rect 134904 130292 137428 130320
rect 134904 130280 134910 130292
rect 137422 130280 137428 130292
rect 137480 130280 137486 130332
rect 53426 130212 53432 130264
rect 53484 130252 53490 130264
rect 58210 130252 58216 130264
rect 53484 130224 58216 130252
rect 53484 130212 53490 130224
rect 58210 130212 58216 130224
rect 58268 130212 58274 130264
rect 92710 130212 92716 130264
rect 92768 130252 92774 130264
rect 101174 130252 101180 130264
rect 92768 130224 101180 130252
rect 92768 130212 92774 130224
rect 101174 130212 101180 130224
rect 101232 130212 101238 130264
rect 137146 130212 137152 130264
rect 137204 130252 137210 130264
rect 143586 130252 143592 130264
rect 137204 130224 143592 130252
rect 137204 130212 137210 130224
rect 143586 130212 143592 130224
rect 143644 130212 143650 130264
rect 177626 130212 177632 130264
rect 177684 130252 177690 130264
rect 185538 130252 185544 130264
rect 177684 130224 185544 130252
rect 177684 130212 177690 130224
rect 185538 130212 185544 130224
rect 185596 130212 185602 130264
rect 52782 130144 52788 130196
rect 52840 130184 52846 130196
rect 58302 130184 58308 130196
rect 52840 130156 58308 130184
rect 52840 130144 52846 130156
rect 58302 130144 58308 130156
rect 58360 130144 58366 130196
rect 92802 130144 92808 130196
rect 92860 130184 92866 130196
rect 101542 130184 101548 130196
rect 92860 130156 101548 130184
rect 92860 130144 92866 130156
rect 101542 130144 101548 130156
rect 101600 130144 101606 130196
rect 137974 130144 137980 130196
rect 138032 130184 138038 130196
rect 143034 130184 143040 130196
rect 138032 130156 143040 130184
rect 138032 130144 138038 130156
rect 143034 130144 143040 130156
rect 143092 130144 143098 130196
rect 177718 130144 177724 130196
rect 177776 130184 177782 130196
rect 185722 130184 185728 130196
rect 177776 130156 185728 130184
rect 177776 130144 177782 130156
rect 185722 130144 185728 130156
rect 185780 130144 185786 130196
rect 134662 129328 134668 129380
rect 134720 129368 134726 129380
rect 137514 129368 137520 129380
rect 134720 129340 137520 129368
rect 134720 129328 134726 129340
rect 137514 129328 137520 129340
rect 137572 129328 137578 129380
rect 50390 129056 50396 129108
rect 50448 129096 50454 129108
rect 56462 129096 56468 129108
rect 50448 129068 56468 129096
rect 50448 129056 50454 129068
rect 56462 129056 56468 129068
rect 56520 129056 56526 129108
rect 51218 128920 51224 128972
rect 51276 128960 51282 128972
rect 52874 128960 52880 128972
rect 51276 128932 52880 128960
rect 51276 128920 51282 128932
rect 52874 128920 52880 128932
rect 52932 128920 52938 128972
rect 135398 128920 135404 128972
rect 135456 128960 135462 128972
rect 135456 128932 139676 128960
rect 135456 128920 135462 128932
rect 52690 128852 52696 128904
rect 52748 128892 52754 128904
rect 58302 128892 58308 128904
rect 52748 128864 58308 128892
rect 52748 128852 52754 128864
rect 58302 128852 58308 128864
rect 58360 128852 58366 128904
rect 92710 128852 92716 128904
rect 92768 128892 92774 128904
rect 101818 128892 101824 128904
rect 92768 128864 101824 128892
rect 92768 128852 92774 128864
rect 101818 128852 101824 128864
rect 101876 128852 101882 128904
rect 139648 128892 139676 128932
rect 143126 128892 143132 128904
rect 139648 128864 143132 128892
rect 143126 128852 143132 128864
rect 143184 128852 143190 128904
rect 177350 128852 177356 128904
rect 177408 128892 177414 128904
rect 185170 128892 185176 128904
rect 177408 128864 185176 128892
rect 177408 128852 177414 128864
rect 185170 128852 185176 128864
rect 185228 128852 185234 128904
rect 52966 128784 52972 128836
rect 53024 128824 53030 128836
rect 58210 128824 58216 128836
rect 53024 128796 58216 128824
rect 53024 128784 53030 128796
rect 58210 128784 58216 128796
rect 58268 128784 58274 128836
rect 92802 128784 92808 128836
rect 92860 128824 92866 128836
rect 101358 128824 101364 128836
rect 92860 128796 101364 128824
rect 92860 128784 92866 128796
rect 101358 128784 101364 128796
rect 101416 128784 101422 128836
rect 137422 128784 137428 128836
rect 137480 128824 137486 128836
rect 142758 128824 142764 128836
rect 137480 128796 142764 128824
rect 137480 128784 137486 128796
rect 142758 128784 142764 128796
rect 142816 128784 142822 128836
rect 177626 128784 177632 128836
rect 177684 128824 177690 128836
rect 185262 128824 185268 128836
rect 177684 128796 185268 128824
rect 177684 128784 177690 128796
rect 185262 128784 185268 128796
rect 185320 128784 185326 128836
rect 92710 128716 92716 128768
rect 92768 128756 92774 128768
rect 101726 128756 101732 128768
rect 92768 128728 101732 128756
rect 92768 128716 92774 128728
rect 101726 128716 101732 128728
rect 101784 128716 101790 128768
rect 137606 128716 137612 128768
rect 137664 128756 137670 128768
rect 143586 128756 143592 128768
rect 137664 128728 143592 128756
rect 137664 128716 137670 128728
rect 143586 128716 143592 128728
rect 143644 128716 143650 128768
rect 177718 128716 177724 128768
rect 177776 128756 177782 128768
rect 185354 128756 185360 128768
rect 177776 128728 185360 128756
rect 177776 128716 177782 128728
rect 185354 128716 185360 128728
rect 185412 128716 185418 128768
rect 56462 128308 56468 128360
rect 56520 128348 56526 128360
rect 58210 128348 58216 128360
rect 56520 128320 58216 128348
rect 56520 128308 56526 128320
rect 58210 128308 58216 128320
rect 58268 128308 58274 128360
rect 50942 127832 50948 127884
rect 51000 127872 51006 127884
rect 56738 127872 56744 127884
rect 51000 127844 56744 127872
rect 51000 127832 51006 127844
rect 56738 127832 56744 127844
rect 56796 127832 56802 127884
rect 134662 127832 134668 127884
rect 134720 127872 134726 127884
rect 137606 127872 137612 127884
rect 134720 127844 137612 127872
rect 134720 127832 134726 127844
rect 137606 127832 137612 127844
rect 137664 127832 137670 127884
rect 51218 127764 51224 127816
rect 51276 127804 51282 127816
rect 52782 127804 52788 127816
rect 51276 127776 52788 127804
rect 51276 127764 51282 127776
rect 52782 127764 52788 127776
rect 52840 127764 52846 127816
rect 134662 127696 134668 127748
rect 134720 127736 134726 127748
rect 136870 127736 136876 127748
rect 134720 127708 136876 127736
rect 134720 127696 134726 127708
rect 136870 127696 136876 127708
rect 136928 127696 136934 127748
rect 51218 127560 51224 127612
rect 51276 127600 51282 127612
rect 52690 127600 52696 127612
rect 51276 127572 52696 127600
rect 51276 127560 51282 127572
rect 52690 127560 52696 127572
rect 52748 127560 52754 127612
rect 135398 127492 135404 127544
rect 135456 127532 135462 127544
rect 135456 127504 139676 127532
rect 135456 127492 135462 127504
rect 52874 127424 52880 127476
rect 52932 127464 52938 127476
rect 58210 127464 58216 127476
rect 52932 127436 58216 127464
rect 52932 127424 52938 127436
rect 58210 127424 58216 127436
rect 58268 127424 58274 127476
rect 92802 127424 92808 127476
rect 92860 127464 92866 127476
rect 100990 127464 100996 127476
rect 92860 127436 100996 127464
rect 92860 127424 92866 127436
rect 100990 127424 100996 127436
rect 101048 127424 101054 127476
rect 139648 127464 139676 127504
rect 143310 127464 143316 127476
rect 139648 127436 143316 127464
rect 143310 127424 143316 127436
rect 143368 127424 143374 127476
rect 177718 127424 177724 127476
rect 177776 127464 177782 127476
rect 185170 127464 185176 127476
rect 177776 127436 185176 127464
rect 177776 127424 177782 127436
rect 185170 127424 185176 127436
rect 185228 127424 185234 127476
rect 216266 127424 216272 127476
rect 216324 127464 216330 127476
rect 222338 127464 222344 127476
rect 216324 127436 222344 127464
rect 216324 127424 216330 127436
rect 222338 127424 222344 127436
rect 222396 127424 222402 127476
rect 92710 127356 92716 127408
rect 92768 127396 92774 127408
rect 101266 127396 101272 127408
rect 92768 127368 101272 127396
rect 92768 127356 92774 127368
rect 101266 127356 101272 127368
rect 101324 127356 101330 127408
rect 137514 127356 137520 127408
rect 137572 127396 137578 127408
rect 142482 127396 142488 127408
rect 137572 127368 142488 127396
rect 137572 127356 137578 127368
rect 142482 127356 142488 127368
rect 142540 127356 142546 127408
rect 177166 127356 177172 127408
rect 177224 127396 177230 127408
rect 185446 127396 185452 127408
rect 177224 127368 185452 127396
rect 177224 127356 177230 127368
rect 185446 127356 185452 127368
rect 185504 127356 185510 127408
rect 56738 127152 56744 127204
rect 56796 127192 56802 127204
rect 58302 127192 58308 127204
rect 56796 127164 58308 127192
rect 56796 127152 56802 127164
rect 58302 127152 58308 127164
rect 58360 127152 58366 127204
rect 98046 126200 98052 126252
rect 98104 126240 98110 126252
rect 101818 126240 101824 126252
rect 98104 126212 101824 126240
rect 98104 126200 98110 126212
rect 101818 126200 101824 126212
rect 101876 126200 101882 126252
rect 182226 126200 182232 126252
rect 182284 126240 182290 126252
rect 185446 126240 185452 126252
rect 182284 126212 185452 126240
rect 182284 126200 182290 126212
rect 185446 126200 185452 126212
rect 185504 126200 185510 126252
rect 98138 126132 98144 126184
rect 98196 126172 98202 126184
rect 101726 126172 101732 126184
rect 98196 126144 101732 126172
rect 98196 126132 98202 126144
rect 101726 126132 101732 126144
rect 101784 126132 101790 126184
rect 182318 126132 182324 126184
rect 182376 126172 182382 126184
rect 185170 126172 185176 126184
rect 182376 126144 185176 126172
rect 182376 126132 182382 126144
rect 185170 126132 185176 126144
rect 185228 126132 185234 126184
rect 52690 126064 52696 126116
rect 52748 126104 52754 126116
rect 58302 126104 58308 126116
rect 52748 126076 58308 126104
rect 52748 126064 52754 126076
rect 58302 126064 58308 126076
rect 58360 126064 58366 126116
rect 92802 126064 92808 126116
rect 92860 126104 92866 126116
rect 101082 126104 101088 126116
rect 92860 126076 101088 126104
rect 92860 126064 92866 126076
rect 101082 126064 101088 126076
rect 101140 126064 101146 126116
rect 137606 126064 137612 126116
rect 137664 126104 137670 126116
rect 143586 126104 143592 126116
rect 137664 126076 143592 126104
rect 137664 126064 137670 126076
rect 143586 126064 143592 126076
rect 143644 126064 143650 126116
rect 177626 126064 177632 126116
rect 177684 126104 177690 126116
rect 185262 126104 185268 126116
rect 177684 126076 185268 126104
rect 177684 126064 177690 126076
rect 185262 126064 185268 126076
rect 185320 126064 185326 126116
rect 52782 125996 52788 126048
rect 52840 126036 52846 126048
rect 58210 126036 58216 126048
rect 52840 126008 58216 126036
rect 52840 125996 52846 126008
rect 58210 125996 58216 126008
rect 58268 125996 58274 126048
rect 92710 125996 92716 126048
rect 92768 126036 92774 126048
rect 101174 126036 101180 126048
rect 92768 126008 101180 126036
rect 92768 125996 92774 126008
rect 101174 125996 101180 126008
rect 101232 125996 101238 126048
rect 136870 125996 136876 126048
rect 136928 126036 136934 126048
rect 143034 126036 143040 126048
rect 136928 126008 143040 126036
rect 136928 125996 136934 126008
rect 143034 125996 143040 126008
rect 143092 125996 143098 126048
rect 177718 125996 177724 126048
rect 177776 126036 177782 126048
rect 185354 126036 185360 126048
rect 177776 126008 185360 126036
rect 177776 125996 177782 126008
rect 185354 125996 185360 126008
rect 185412 125996 185418 126048
rect 135030 125248 135036 125300
rect 135088 125288 135094 125300
rect 137606 125288 137612 125300
rect 135088 125260 137612 125288
rect 135088 125248 135094 125260
rect 137606 125248 137612 125260
rect 137664 125248 137670 125300
rect 51218 124976 51224 125028
rect 51276 125016 51282 125028
rect 52966 125016 52972 125028
rect 51276 124988 52972 125016
rect 51276 124976 51282 124988
rect 52966 124976 52972 124988
rect 53024 124976 53030 125028
rect 51218 124840 51224 124892
rect 51276 124880 51282 124892
rect 52874 124880 52880 124892
rect 51276 124852 52880 124880
rect 51276 124840 51282 124852
rect 52874 124840 52880 124852
rect 52932 124840 52938 124892
rect 135398 124840 135404 124892
rect 135456 124880 135462 124892
rect 136870 124880 136876 124892
rect 135456 124852 136876 124880
rect 135456 124840 135462 124852
rect 136870 124840 136876 124852
rect 136928 124840 136934 124892
rect 50206 124772 50212 124824
rect 50264 124812 50270 124824
rect 58394 124812 58400 124824
rect 50264 124784 58400 124812
rect 50264 124772 50270 124784
rect 58394 124772 58400 124784
rect 58452 124772 58458 124824
rect 135214 124772 135220 124824
rect 135272 124812 135278 124824
rect 142758 124812 142764 124824
rect 135272 124784 142764 124812
rect 135272 124772 135278 124784
rect 142758 124772 142764 124784
rect 142816 124772 142822 124824
rect 51310 124704 51316 124756
rect 51368 124744 51374 124756
rect 58302 124744 58308 124756
rect 51368 124716 58308 124744
rect 51368 124704 51374 124716
rect 58302 124704 58308 124716
rect 58360 124704 58366 124756
rect 92894 124704 92900 124756
rect 92952 124744 92958 124756
rect 101450 124744 101456 124756
rect 92952 124716 101456 124744
rect 92952 124704 92958 124716
rect 101450 124704 101456 124716
rect 101508 124704 101514 124756
rect 135582 124704 135588 124756
rect 135640 124744 135646 124756
rect 143586 124744 143592 124756
rect 135640 124716 143592 124744
rect 135640 124704 135646 124716
rect 143586 124704 143592 124716
rect 143644 124704 143650 124756
rect 177626 124704 177632 124756
rect 177684 124744 177690 124756
rect 185170 124744 185176 124756
rect 177684 124716 185176 124744
rect 177684 124704 177690 124716
rect 185170 124704 185176 124716
rect 185228 124704 185234 124756
rect 51402 124636 51408 124688
rect 51460 124676 51466 124688
rect 58210 124676 58216 124688
rect 51460 124648 58216 124676
rect 51460 124636 51466 124648
rect 58210 124636 58216 124648
rect 58268 124636 58274 124688
rect 92710 124636 92716 124688
rect 92768 124676 92774 124688
rect 98046 124676 98052 124688
rect 92768 124648 98052 124676
rect 92768 124636 92774 124648
rect 98046 124636 98052 124648
rect 98104 124636 98110 124688
rect 177718 124636 177724 124688
rect 177776 124676 177782 124688
rect 182226 124676 182232 124688
rect 177776 124648 182232 124676
rect 177776 124636 177782 124648
rect 182226 124636 182232 124648
rect 182284 124636 182290 124688
rect 92802 124568 92808 124620
rect 92860 124608 92866 124620
rect 98138 124608 98144 124620
rect 92860 124580 98144 124608
rect 92860 124568 92866 124580
rect 98138 124568 98144 124580
rect 98196 124568 98202 124620
rect 135490 124364 135496 124416
rect 135548 124404 135554 124416
rect 142482 124404 142488 124416
rect 135548 124376 142488 124404
rect 135548 124364 135554 124376
rect 142482 124364 142488 124376
rect 142540 124364 142546 124416
rect 177166 124364 177172 124416
rect 177224 124404 177230 124416
rect 182318 124404 182324 124416
rect 177224 124376 182324 124404
rect 177224 124364 177230 124376
rect 182318 124364 182324 124376
rect 182376 124364 182382 124416
rect 134478 123480 134484 123532
rect 134536 123520 134542 123532
rect 137698 123520 137704 123532
rect 134536 123492 137704 123520
rect 134536 123480 134542 123492
rect 137698 123480 137704 123492
rect 137756 123480 137762 123532
rect 50574 123412 50580 123464
rect 50632 123452 50638 123464
rect 52690 123452 52696 123464
rect 50632 123424 52696 123452
rect 50632 123412 50638 123424
rect 52690 123412 52696 123424
rect 52748 123412 52754 123464
rect 51126 123344 51132 123396
rect 51184 123384 51190 123396
rect 52782 123384 52788 123396
rect 51184 123356 52788 123384
rect 51184 123344 51190 123356
rect 52782 123344 52788 123356
rect 52840 123344 52846 123396
rect 134110 123344 134116 123396
rect 134168 123384 134174 123396
rect 138158 123384 138164 123396
rect 134168 123356 138164 123384
rect 134168 123344 134174 123356
rect 138158 123344 138164 123356
rect 138216 123344 138222 123396
rect 52966 123276 52972 123328
rect 53024 123316 53030 123328
rect 58210 123316 58216 123328
rect 53024 123288 58216 123316
rect 53024 123276 53030 123288
rect 58210 123276 58216 123288
rect 58268 123276 58274 123328
rect 92710 123276 92716 123328
rect 92768 123316 92774 123328
rect 101634 123316 101640 123328
rect 92768 123288 101640 123316
rect 92768 123276 92774 123288
rect 101634 123276 101640 123288
rect 101692 123276 101698 123328
rect 137606 123276 137612 123328
rect 137664 123316 137670 123328
rect 143586 123316 143592 123328
rect 137664 123288 143592 123316
rect 137664 123276 137670 123288
rect 143586 123276 143592 123288
rect 143644 123276 143650 123328
rect 177626 123276 177632 123328
rect 177684 123316 177690 123328
rect 185262 123316 185268 123328
rect 177684 123288 185268 123316
rect 177684 123276 177690 123288
rect 185262 123276 185268 123288
rect 185320 123276 185326 123328
rect 52874 123208 52880 123260
rect 52932 123248 52938 123260
rect 58302 123248 58308 123260
rect 52932 123220 58308 123248
rect 52932 123208 52938 123220
rect 58302 123208 58308 123220
rect 58360 123208 58366 123260
rect 92802 123208 92808 123260
rect 92860 123248 92866 123260
rect 101726 123248 101732 123260
rect 92860 123220 101732 123248
rect 92860 123208 92866 123220
rect 101726 123208 101732 123220
rect 101784 123208 101790 123260
rect 177718 123208 177724 123260
rect 177776 123248 177782 123260
rect 185354 123248 185360 123260
rect 177776 123220 185360 123248
rect 177776 123208 177782 123220
rect 185354 123208 185360 123220
rect 185412 123208 185418 123260
rect 136870 122868 136876 122920
rect 136928 122908 136934 122920
rect 142850 122908 142856 122920
rect 136928 122880 142856 122908
rect 136928 122868 136934 122880
rect 142850 122868 142856 122880
rect 142908 122868 142914 122920
rect 134478 122392 134484 122444
rect 134536 122432 134542 122444
rect 138066 122432 138072 122444
rect 134536 122404 138072 122432
rect 134536 122392 134542 122404
rect 138066 122392 138072 122404
rect 138124 122392 138130 122444
rect 50850 122324 50856 122376
rect 50908 122364 50914 122376
rect 52966 122364 52972 122376
rect 50908 122336 52972 122364
rect 50908 122324 50914 122336
rect 52966 122324 52972 122336
rect 53024 122324 53030 122376
rect 134938 122256 134944 122308
rect 134996 122296 135002 122308
rect 137238 122296 137244 122308
rect 134996 122268 137244 122296
rect 134996 122256 135002 122268
rect 137238 122256 137244 122268
rect 137296 122256 137302 122308
rect 50206 122188 50212 122240
rect 50264 122228 50270 122240
rect 52874 122228 52880 122240
rect 50264 122200 52880 122228
rect 50264 122188 50270 122200
rect 52874 122188 52880 122200
rect 52932 122188 52938 122240
rect 52782 121916 52788 121968
rect 52840 121956 52846 121968
rect 58302 121956 58308 121968
rect 52840 121928 58308 121956
rect 52840 121916 52846 121928
rect 58302 121916 58308 121928
rect 58360 121916 58366 121968
rect 92802 121916 92808 121968
rect 92860 121956 92866 121968
rect 101818 121956 101824 121968
rect 92860 121928 101824 121956
rect 92860 121916 92866 121928
rect 101818 121916 101824 121928
rect 101876 121916 101882 121968
rect 137698 121916 137704 121968
rect 137756 121956 137762 121968
rect 142758 121956 142764 121968
rect 137756 121928 142764 121956
rect 137756 121916 137762 121928
rect 142758 121916 142764 121928
rect 142816 121916 142822 121968
rect 177626 121916 177632 121968
rect 177684 121956 177690 121968
rect 185722 121956 185728 121968
rect 177684 121928 185728 121956
rect 177684 121916 177690 121928
rect 185722 121916 185728 121928
rect 185780 121916 185786 121968
rect 52690 121848 52696 121900
rect 52748 121888 52754 121900
rect 58210 121888 58216 121900
rect 52748 121860 58216 121888
rect 52748 121848 52754 121860
rect 58210 121848 58216 121860
rect 58268 121848 58274 121900
rect 92710 121848 92716 121900
rect 92768 121888 92774 121900
rect 101910 121888 101916 121900
rect 92768 121860 101916 121888
rect 92768 121848 92774 121860
rect 101910 121848 101916 121860
rect 101968 121848 101974 121900
rect 138158 121848 138164 121900
rect 138216 121888 138222 121900
rect 143034 121888 143040 121900
rect 138216 121860 143040 121888
rect 138216 121848 138222 121860
rect 143034 121848 143040 121860
rect 143092 121848 143098 121900
rect 177718 121848 177724 121900
rect 177776 121888 177782 121900
rect 185906 121888 185912 121900
rect 177776 121860 185912 121888
rect 177776 121848 177782 121860
rect 185906 121848 185912 121860
rect 185964 121848 185970 121900
rect 51218 120896 51224 120948
rect 51276 120936 51282 120948
rect 53058 120936 53064 120948
rect 51276 120908 53064 120936
rect 51276 120896 51282 120908
rect 53058 120896 53064 120908
rect 53116 120896 53122 120948
rect 97862 120760 97868 120812
rect 97920 120800 97926 120812
rect 101726 120800 101732 120812
rect 97920 120772 101732 120800
rect 97920 120760 97926 120772
rect 101726 120760 101732 120772
rect 101784 120760 101790 120812
rect 134478 120760 134484 120812
rect 134536 120800 134542 120812
rect 137422 120800 137428 120812
rect 134536 120772 137428 120800
rect 134536 120760 134542 120772
rect 137422 120760 137428 120772
rect 137480 120760 137486 120812
rect 182042 120760 182048 120812
rect 182100 120800 182106 120812
rect 185354 120800 185360 120812
rect 182100 120772 185360 120800
rect 182100 120760 182106 120772
rect 185354 120760 185360 120772
rect 185412 120760 185418 120812
rect 51218 120692 51224 120744
rect 51276 120732 51282 120744
rect 52690 120732 52696 120744
rect 51276 120704 52696 120732
rect 51276 120692 51282 120704
rect 52690 120692 52696 120704
rect 52748 120692 52754 120744
rect 97954 120692 97960 120744
rect 98012 120732 98018 120744
rect 101082 120732 101088 120744
rect 98012 120704 101088 120732
rect 98012 120692 98018 120704
rect 101082 120692 101088 120704
rect 101140 120692 101146 120744
rect 134662 120692 134668 120744
rect 134720 120732 134726 120744
rect 137514 120732 137520 120744
rect 134720 120704 137520 120732
rect 134720 120692 134726 120704
rect 137514 120692 137520 120704
rect 137572 120692 137578 120744
rect 182318 120692 182324 120744
rect 182376 120732 182382 120744
rect 185262 120732 185268 120744
rect 182376 120704 185268 120732
rect 182376 120692 182382 120704
rect 185262 120692 185268 120704
rect 185320 120692 185326 120744
rect 50206 120624 50212 120676
rect 50264 120664 50270 120676
rect 53150 120664 53156 120676
rect 50264 120636 53156 120664
rect 50264 120624 50270 120636
rect 53150 120624 53156 120636
rect 53208 120624 53214 120676
rect 98138 120624 98144 120676
rect 98196 120664 98202 120676
rect 101542 120664 101548 120676
rect 98196 120636 101548 120664
rect 98196 120624 98202 120636
rect 101542 120624 101548 120636
rect 101600 120624 101606 120676
rect 135398 120624 135404 120676
rect 135456 120664 135462 120676
rect 136870 120664 136876 120676
rect 135456 120636 136876 120664
rect 135456 120624 135462 120636
rect 136870 120624 136876 120636
rect 136928 120624 136934 120676
rect 181766 120624 181772 120676
rect 181824 120664 181830 120676
rect 185170 120664 185176 120676
rect 181824 120636 185176 120664
rect 181824 120624 181830 120636
rect 185170 120624 185176 120636
rect 185228 120624 185234 120676
rect 52966 120556 52972 120608
rect 53024 120596 53030 120608
rect 58210 120596 58216 120608
rect 53024 120568 58216 120596
rect 53024 120556 53030 120568
rect 58210 120556 58216 120568
rect 58268 120556 58274 120608
rect 92710 120556 92716 120608
rect 92768 120596 92774 120608
rect 101634 120596 101640 120608
rect 92768 120568 101640 120596
rect 92768 120556 92774 120568
rect 101634 120556 101640 120568
rect 101692 120556 101698 120608
rect 138066 120556 138072 120608
rect 138124 120596 138130 120608
rect 142942 120596 142948 120608
rect 138124 120568 142948 120596
rect 138124 120556 138130 120568
rect 142942 120556 142948 120568
rect 143000 120556 143006 120608
rect 177718 120556 177724 120608
rect 177776 120596 177782 120608
rect 185814 120596 185820 120608
rect 177776 120568 185820 120596
rect 177776 120556 177782 120568
rect 185814 120556 185820 120568
rect 185872 120556 185878 120608
rect 52874 120488 52880 120540
rect 52932 120528 52938 120540
rect 58302 120528 58308 120540
rect 52932 120500 58308 120528
rect 52932 120488 52938 120500
rect 58302 120488 58308 120500
rect 58360 120488 58366 120540
rect 92802 120488 92808 120540
rect 92860 120528 92866 120540
rect 101450 120528 101456 120540
rect 92860 120500 101456 120528
rect 92860 120488 92866 120500
rect 101450 120488 101456 120500
rect 101508 120488 101514 120540
rect 137238 120488 137244 120540
rect 137296 120528 137302 120540
rect 143586 120528 143592 120540
rect 137296 120500 143592 120528
rect 137296 120488 137302 120500
rect 143586 120488 143592 120500
rect 143644 120488 143650 120540
rect 177626 120488 177632 120540
rect 177684 120528 177690 120540
rect 185538 120528 185544 120540
rect 177684 120500 185544 120528
rect 177684 120488 177690 120500
rect 185538 120488 185544 120500
rect 185596 120488 185602 120540
rect 51218 119536 51224 119588
rect 51276 119576 51282 119588
rect 52874 119576 52880 119588
rect 51276 119548 52880 119576
rect 51276 119536 51282 119548
rect 52874 119536 52880 119548
rect 52932 119536 52938 119588
rect 135398 119536 135404 119588
rect 135456 119576 135462 119588
rect 137606 119576 137612 119588
rect 135456 119548 137612 119576
rect 135456 119536 135462 119548
rect 137606 119536 137612 119548
rect 137664 119536 137670 119588
rect 97678 119332 97684 119384
rect 97736 119372 97742 119384
rect 101266 119372 101272 119384
rect 97736 119344 101272 119372
rect 97736 119332 97742 119344
rect 101266 119332 101272 119344
rect 101324 119332 101330 119384
rect 182134 119332 182140 119384
rect 182192 119372 182198 119384
rect 185262 119372 185268 119384
rect 182192 119344 185268 119372
rect 182192 119332 182198 119344
rect 185262 119332 185268 119344
rect 185320 119332 185326 119384
rect 51218 119264 51224 119316
rect 51276 119304 51282 119316
rect 52782 119304 52788 119316
rect 51276 119276 52788 119304
rect 51276 119264 51282 119276
rect 52782 119264 52788 119276
rect 52840 119264 52846 119316
rect 98046 119264 98052 119316
rect 98104 119304 98110 119316
rect 101358 119304 101364 119316
rect 98104 119276 101364 119304
rect 98104 119264 98110 119276
rect 101358 119264 101364 119276
rect 101416 119264 101422 119316
rect 134478 119264 134484 119316
rect 134536 119304 134542 119316
rect 136962 119304 136968 119316
rect 134536 119276 136968 119304
rect 134536 119264 134542 119276
rect 136962 119264 136968 119276
rect 137020 119264 137026 119316
rect 182226 119264 182232 119316
rect 182284 119304 182290 119316
rect 185170 119304 185176 119316
rect 182284 119276 185176 119304
rect 182284 119264 182290 119276
rect 185170 119264 185176 119276
rect 185228 119264 185234 119316
rect 52690 119196 52696 119248
rect 52748 119236 52754 119248
rect 58394 119236 58400 119248
rect 52748 119208 58400 119236
rect 52748 119196 52754 119208
rect 58394 119196 58400 119208
rect 58452 119196 58458 119248
rect 92894 119196 92900 119248
rect 92952 119236 92958 119248
rect 98138 119236 98144 119248
rect 92952 119208 98144 119236
rect 92952 119196 92958 119208
rect 98138 119196 98144 119208
rect 98196 119196 98202 119248
rect 137422 119196 137428 119248
rect 137480 119236 137486 119248
rect 143586 119236 143592 119248
rect 137480 119208 143592 119236
rect 137480 119196 137486 119208
rect 143586 119196 143592 119208
rect 143644 119196 143650 119248
rect 53150 119128 53156 119180
rect 53208 119168 53214 119180
rect 58210 119168 58216 119180
rect 53208 119140 58216 119168
rect 53208 119128 53214 119140
rect 58210 119128 58216 119140
rect 58268 119128 58274 119180
rect 92802 119128 92808 119180
rect 92860 119168 92866 119180
rect 97954 119168 97960 119180
rect 92860 119140 97960 119168
rect 92860 119128 92866 119140
rect 97954 119128 97960 119140
rect 98012 119128 98018 119180
rect 136870 119128 136876 119180
rect 136928 119168 136934 119180
rect 142574 119168 142580 119180
rect 136928 119140 142580 119168
rect 136928 119128 136934 119140
rect 142574 119128 142580 119140
rect 142632 119128 142638 119180
rect 177718 119128 177724 119180
rect 177776 119168 177782 119180
rect 182042 119168 182048 119180
rect 177776 119140 182048 119168
rect 177776 119128 177782 119140
rect 182042 119128 182048 119140
rect 182100 119128 182106 119180
rect 53058 119060 53064 119112
rect 53116 119100 53122 119112
rect 58302 119100 58308 119112
rect 53116 119072 58308 119100
rect 53116 119060 53122 119072
rect 58302 119060 58308 119072
rect 58360 119060 58366 119112
rect 92710 119060 92716 119112
rect 92768 119100 92774 119112
rect 97862 119100 97868 119112
rect 92768 119072 97868 119100
rect 92768 119060 92774 119072
rect 97862 119060 97868 119072
rect 97920 119060 97926 119112
rect 137514 119060 137520 119112
rect 137572 119100 137578 119112
rect 143586 119100 143592 119112
rect 137572 119072 143592 119100
rect 137572 119060 137578 119072
rect 143586 119060 143592 119072
rect 143644 119060 143650 119112
rect 177718 118924 177724 118976
rect 177776 118964 177782 118976
rect 181766 118964 181772 118976
rect 177776 118936 181772 118964
rect 177776 118924 177782 118936
rect 181766 118924 181772 118936
rect 181824 118924 181830 118976
rect 177626 118788 177632 118840
rect 177684 118828 177690 118840
rect 182318 118828 182324 118840
rect 177684 118800 182324 118828
rect 177684 118788 177690 118800
rect 182318 118788 182324 118800
rect 182376 118788 182382 118840
rect 134662 118448 134668 118500
rect 134720 118488 134726 118500
rect 136870 118488 136876 118500
rect 134720 118460 136876 118488
rect 134720 118448 134726 118460
rect 136870 118448 136876 118460
rect 136928 118448 136934 118500
rect 51218 118176 51224 118228
rect 51276 118216 51282 118228
rect 52966 118216 52972 118228
rect 51276 118188 52972 118216
rect 51276 118176 51282 118188
rect 52966 118176 52972 118188
rect 53024 118176 53030 118228
rect 134662 118176 134668 118228
rect 134720 118216 134726 118228
rect 137514 118216 137520 118228
rect 134720 118188 137520 118216
rect 134720 118176 134726 118188
rect 137514 118176 137520 118188
rect 137572 118176 137578 118228
rect 51218 117904 51224 117956
rect 51276 117944 51282 117956
rect 52690 117944 52696 117956
rect 51276 117916 52696 117944
rect 51276 117904 51282 117916
rect 52690 117904 52696 117916
rect 52748 117904 52754 117956
rect 97954 117904 97960 117956
rect 98012 117944 98018 117956
rect 101358 117944 101364 117956
rect 98012 117916 101364 117944
rect 98012 117904 98018 117916
rect 101358 117904 101364 117916
rect 101416 117904 101422 117956
rect 181398 117904 181404 117956
rect 181456 117944 181462 117956
rect 185262 117944 185268 117956
rect 181456 117916 185268 117944
rect 181456 117904 181462 117916
rect 185262 117904 185268 117916
rect 185320 117904 185326 117956
rect 98138 117836 98144 117888
rect 98196 117876 98202 117888
rect 101726 117876 101732 117888
rect 98196 117848 101732 117876
rect 98196 117836 98202 117848
rect 101726 117836 101732 117848
rect 101784 117836 101790 117888
rect 182318 117836 182324 117888
rect 182376 117876 182382 117888
rect 185170 117876 185176 117888
rect 182376 117848 185176 117876
rect 182376 117836 182382 117848
rect 185170 117836 185176 117848
rect 185228 117836 185234 117888
rect 52874 117768 52880 117820
rect 52932 117808 52938 117820
rect 58210 117808 58216 117820
rect 52932 117780 58216 117808
rect 52932 117768 52938 117780
rect 58210 117768 58216 117780
rect 58268 117768 58274 117820
rect 92710 117768 92716 117820
rect 92768 117808 92774 117820
rect 97678 117808 97684 117820
rect 92768 117780 97684 117808
rect 92768 117768 92774 117780
rect 97678 117768 97684 117780
rect 97736 117768 97742 117820
rect 136962 117768 136968 117820
rect 137020 117808 137026 117820
rect 142574 117808 142580 117820
rect 137020 117780 142580 117808
rect 137020 117768 137026 117780
rect 142574 117768 142580 117780
rect 142632 117768 142638 117820
rect 52782 117700 52788 117752
rect 52840 117740 52846 117752
rect 58302 117740 58308 117752
rect 52840 117712 58308 117740
rect 52840 117700 52846 117712
rect 58302 117700 58308 117712
rect 58360 117700 58366 117752
rect 92802 117700 92808 117752
rect 92860 117740 92866 117752
rect 98046 117740 98052 117752
rect 92860 117712 98052 117740
rect 92860 117700 92866 117712
rect 98046 117700 98052 117712
rect 98104 117700 98110 117752
rect 137606 117700 137612 117752
rect 137664 117740 137670 117752
rect 143218 117740 143224 117752
rect 137664 117712 143224 117740
rect 137664 117700 137670 117712
rect 143218 117700 143224 117712
rect 143276 117700 143282 117752
rect 177718 117700 177724 117752
rect 177776 117740 177782 117752
rect 182134 117740 182140 117752
rect 177776 117712 182140 117740
rect 177776 117700 177782 117712
rect 182134 117700 182140 117712
rect 182192 117700 182198 117752
rect 177626 117564 177632 117616
rect 177684 117604 177690 117616
rect 182226 117604 182232 117616
rect 177684 117576 182232 117604
rect 177684 117564 177690 117576
rect 182226 117564 182232 117576
rect 182284 117564 182290 117616
rect 51218 116680 51224 116732
rect 51276 116720 51282 116732
rect 56462 116720 56468 116732
rect 51276 116692 56468 116720
rect 51276 116680 51282 116692
rect 56462 116680 56468 116692
rect 56520 116680 56526 116732
rect 93998 116544 94004 116596
rect 94056 116584 94062 116596
rect 101082 116584 101088 116596
rect 94056 116556 101088 116584
rect 94056 116544 94062 116556
rect 101082 116544 101088 116556
rect 101140 116544 101146 116596
rect 178178 116544 178184 116596
rect 178236 116584 178242 116596
rect 185262 116584 185268 116596
rect 178236 116556 185268 116584
rect 178236 116544 178242 116556
rect 185262 116544 185268 116556
rect 185320 116544 185326 116596
rect 92618 116476 92624 116528
rect 92676 116516 92682 116528
rect 100990 116516 100996 116528
rect 92676 116488 100996 116516
rect 92676 116476 92682 116488
rect 100990 116476 100996 116488
rect 101048 116476 101054 116528
rect 134846 116476 134852 116528
rect 134904 116516 134910 116528
rect 134904 116488 139676 116516
rect 134904 116476 134910 116488
rect 52966 116408 52972 116460
rect 53024 116448 53030 116460
rect 58210 116448 58216 116460
rect 53024 116420 58216 116448
rect 53024 116408 53030 116420
rect 58210 116408 58216 116420
rect 58268 116408 58274 116460
rect 92894 116408 92900 116460
rect 92952 116448 92958 116460
rect 101174 116448 101180 116460
rect 92952 116420 101180 116448
rect 92952 116408 92958 116420
rect 101174 116408 101180 116420
rect 101232 116408 101238 116460
rect 139648 116448 139676 116488
rect 176798 116476 176804 116528
rect 176856 116516 176862 116528
rect 185170 116516 185176 116528
rect 176856 116488 185176 116516
rect 176856 116476 176862 116488
rect 185170 116476 185176 116488
rect 185228 116476 185234 116528
rect 142758 116448 142764 116460
rect 139648 116420 142764 116448
rect 142758 116408 142764 116420
rect 142816 116408 142822 116460
rect 177074 116408 177080 116460
rect 177132 116448 177138 116460
rect 185354 116448 185360 116460
rect 177132 116420 185360 116448
rect 177132 116408 177138 116420
rect 185354 116408 185360 116420
rect 185412 116408 185418 116460
rect 52690 116340 52696 116392
rect 52748 116380 52754 116392
rect 58302 116380 58308 116392
rect 52748 116352 58308 116380
rect 52748 116340 52754 116352
rect 58302 116340 58308 116352
rect 58360 116340 58366 116392
rect 92710 116340 92716 116392
rect 92768 116380 92774 116392
rect 97954 116380 97960 116392
rect 92768 116352 97960 116380
rect 92768 116340 92774 116352
rect 97954 116340 97960 116352
rect 98012 116340 98018 116392
rect 136870 116340 136876 116392
rect 136928 116380 136934 116392
rect 142942 116380 142948 116392
rect 136928 116352 142948 116380
rect 136928 116340 136934 116352
rect 142942 116340 142948 116352
rect 143000 116340 143006 116392
rect 177718 116340 177724 116392
rect 177776 116380 177782 116392
rect 181398 116380 181404 116392
rect 177776 116352 181404 116380
rect 177776 116340 177782 116352
rect 181398 116340 181404 116352
rect 181456 116340 181462 116392
rect 56462 116272 56468 116324
rect 56520 116312 56526 116324
rect 58394 116312 58400 116324
rect 56520 116284 58400 116312
rect 56520 116272 56526 116284
rect 58394 116272 58400 116284
rect 58452 116272 58458 116324
rect 92802 116272 92808 116324
rect 92860 116312 92866 116324
rect 98138 116312 98144 116324
rect 92860 116284 98144 116312
rect 92860 116272 92866 116284
rect 98138 116272 98144 116284
rect 98196 116272 98202 116324
rect 137514 116272 137520 116324
rect 137572 116312 137578 116324
rect 143586 116312 143592 116324
rect 137572 116284 143592 116312
rect 137572 116272 137578 116284
rect 143586 116272 143592 116284
rect 143644 116272 143650 116324
rect 177718 116068 177724 116120
rect 177776 116108 177782 116120
rect 182318 116108 182324 116120
rect 177776 116080 182324 116108
rect 177776 116068 177782 116080
rect 182318 116068 182324 116080
rect 182376 116068 182382 116120
rect 91238 115184 91244 115236
rect 91296 115224 91302 115236
rect 101082 115224 101088 115236
rect 91296 115196 101088 115224
rect 91296 115184 91302 115196
rect 101082 115184 101088 115196
rect 101140 115184 101146 115236
rect 175418 115184 175424 115236
rect 175476 115224 175482 115236
rect 185262 115224 185268 115236
rect 175476 115196 185268 115224
rect 175476 115184 175482 115196
rect 185262 115184 185268 115196
rect 185320 115184 185326 115236
rect 59314 115156 59320 115168
rect 59275 115128 59320 115156
rect 59314 115116 59320 115128
rect 59372 115116 59378 115168
rect 90594 115116 90600 115168
rect 90652 115156 90658 115168
rect 100990 115156 100996 115168
rect 90652 115128 100996 115156
rect 90652 115116 90658 115128
rect 100990 115116 100996 115128
rect 101048 115116 101054 115168
rect 174774 115116 174780 115168
rect 174832 115156 174838 115168
rect 185170 115156 185176 115168
rect 174832 115128 185176 115156
rect 174832 115116 174838 115128
rect 185170 115116 185176 115128
rect 185228 115116 185234 115168
rect 51218 113824 51224 113876
rect 51276 113864 51282 113876
rect 57566 113864 57572 113876
rect 51276 113836 57572 113864
rect 51276 113824 51282 113836
rect 57566 113824 57572 113836
rect 57624 113824 57630 113876
rect 135398 113688 135404 113740
rect 135456 113728 135462 113740
rect 141562 113728 141568 113740
rect 135456 113700 141568 113728
rect 135456 113688 135462 113700
rect 141562 113688 141568 113700
rect 141620 113688 141626 113740
rect 17822 113280 17828 113332
rect 17880 113320 17886 113332
rect 64098 113320 64104 113332
rect 17880 113292 64104 113320
rect 17880 113280 17886 113292
rect 64098 113280 64104 113292
rect 64156 113280 64162 113332
rect 147266 113280 147272 113332
rect 147324 113320 147330 113332
rect 218382 113320 218388 113332
rect 147324 113292 218388 113320
rect 147324 113280 147330 113292
rect 218382 113280 218388 113292
rect 218440 113280 218446 113332
rect 18006 112940 18012 112992
rect 18064 112980 18070 112992
rect 52598 112980 52604 112992
rect 18064 112952 52604 112980
rect 18064 112940 18070 112952
rect 52598 112940 52604 112952
rect 52656 112940 52662 112992
rect 85718 112328 85724 112380
rect 85776 112368 85782 112380
rect 100990 112368 100996 112380
rect 85776 112340 100996 112368
rect 85776 112328 85782 112340
rect 100990 112328 100996 112340
rect 101048 112328 101054 112380
rect 169898 112328 169904 112380
rect 169956 112368 169962 112380
rect 185170 112368 185176 112380
rect 169956 112340 185176 112368
rect 169956 112328 169962 112340
rect 185170 112328 185176 112340
rect 185228 112328 185234 112380
rect 52598 112260 52604 112312
rect 52656 112300 52662 112312
rect 61890 112300 61896 112312
rect 52656 112272 61896 112300
rect 52656 112260 52662 112272
rect 61890 112260 61896 112272
rect 61948 112260 61954 112312
rect 90410 112192 90416 112244
rect 90468 112232 90474 112244
rect 93354 112232 93360 112244
rect 90468 112204 93360 112232
rect 90468 112192 90474 112204
rect 93354 112192 93360 112204
rect 93412 112192 93418 112244
rect 134018 111648 134024 111700
rect 134076 111688 134082 111700
rect 145334 111688 145340 111700
rect 134076 111660 145340 111688
rect 134076 111648 134082 111660
rect 145334 111648 145340 111660
rect 145392 111648 145398 111700
rect 82314 111580 82320 111632
rect 82372 111620 82378 111632
rect 85442 111620 85448 111632
rect 82372 111592 85448 111620
rect 82372 111580 82378 111592
rect 85442 111580 85448 111592
rect 85500 111580 85506 111632
rect 129970 111580 129976 111632
rect 130028 111620 130034 111632
rect 148094 111620 148100 111632
rect 130028 111592 148100 111620
rect 130028 111580 130034 111592
rect 148094 111580 148100 111592
rect 148152 111580 148158 111632
rect 83694 111512 83700 111564
rect 83752 111552 83758 111564
rect 87190 111552 87196 111564
rect 83752 111524 87196 111552
rect 83752 111512 83758 111524
rect 87190 111512 87196 111524
rect 87248 111512 87254 111564
rect 80934 111444 80940 111496
rect 80992 111484 80998 111496
rect 84062 111484 84068 111496
rect 80992 111456 84068 111484
rect 80992 111444 80998 111456
rect 84062 111444 84068 111456
rect 84120 111444 84126 111496
rect 79646 111104 79652 111156
rect 79704 111144 79710 111156
rect 82590 111144 82596 111156
rect 79704 111116 82596 111144
rect 79704 111104 79710 111116
rect 82590 111104 82596 111116
rect 82648 111104 82654 111156
rect 163826 111104 163832 111156
rect 163884 111144 163890 111156
rect 166586 111144 166592 111156
rect 163884 111116 166592 111144
rect 163884 111104 163890 111116
rect 166586 111104 166592 111116
rect 166644 111104 166650 111156
rect 167874 111104 167880 111156
rect 167932 111144 167938 111156
rect 170910 111144 170916 111156
rect 167932 111116 170916 111144
rect 167932 111104 167938 111116
rect 170910 111104 170916 111116
rect 170968 111104 170974 111156
rect 74034 111036 74040 111088
rect 74092 111076 74098 111088
rect 75506 111076 75512 111088
rect 74092 111048 75512 111076
rect 74092 111036 74098 111048
rect 75506 111036 75512 111048
rect 75564 111036 75570 111088
rect 77438 111036 77444 111088
rect 77496 111076 77502 111088
rect 79738 111076 79744 111088
rect 77496 111048 79744 111076
rect 77496 111036 77502 111048
rect 79738 111036 79744 111048
rect 79796 111036 79802 111088
rect 158858 111036 158864 111088
rect 158916 111076 158922 111088
rect 160882 111076 160888 111088
rect 158916 111048 160888 111076
rect 158916 111036 158922 111048
rect 160882 111036 160888 111048
rect 160940 111036 160946 111088
rect 166494 111036 166500 111088
rect 166552 111076 166558 111088
rect 169438 111076 169444 111088
rect 166552 111048 169444 111076
rect 166552 111036 166558 111048
rect 169438 111036 169444 111048
rect 169496 111036 169502 111088
rect 74678 110968 74684 111020
rect 74736 111008 74742 111020
rect 76886 111008 76892 111020
rect 74736 110980 76892 111008
rect 74736 110968 74742 110980
rect 76886 110968 76892 110980
rect 76944 110968 76950 111020
rect 79554 110968 79560 111020
rect 79612 111008 79618 111020
rect 81210 111008 81216 111020
rect 79612 110980 81216 111008
rect 79612 110968 79618 110980
rect 81210 110968 81216 110980
rect 81268 110968 81274 111020
rect 156834 110968 156840 111020
rect 156892 111008 156898 111020
rect 158030 111008 158036 111020
rect 156892 110980 158036 111008
rect 156892 110968 156898 110980
rect 158030 110968 158036 110980
rect 158088 110968 158094 111020
rect 158306 110968 158312 111020
rect 158364 111008 158370 111020
rect 159502 111008 159508 111020
rect 158364 110980 159508 111008
rect 158364 110968 158370 110980
rect 159502 110968 159508 110980
rect 159560 110968 159566 111020
rect 161618 110968 161624 111020
rect 161676 111008 161682 111020
rect 163734 111008 163740 111020
rect 161676 110980 163740 111008
rect 161676 110968 161682 110980
rect 163734 110968 163740 110980
rect 163792 110968 163798 111020
rect 165114 110968 165120 111020
rect 165172 111008 165178 111020
rect 168058 111008 168064 111020
rect 165172 110980 168064 111008
rect 165172 110968 165178 110980
rect 168058 110968 168064 110980
rect 168116 110968 168122 111020
rect 172658 110968 172664 111020
rect 172716 111008 172722 111020
rect 176154 111008 176160 111020
rect 172716 110980 176160 111008
rect 172716 110968 172722 110980
rect 176154 110968 176160 110980
rect 176212 110968 176218 111020
rect 108994 110900 109000 110952
rect 109052 110940 109058 110952
rect 129970 110940 129976 110952
rect 109052 110912 129976 110940
rect 109052 110900 109058 110912
rect 129970 110900 129976 110912
rect 130028 110900 130034 110952
rect 63270 110832 63276 110884
rect 63328 110872 63334 110884
rect 109546 110872 109552 110884
rect 63328 110844 109552 110872
rect 63328 110832 63334 110844
rect 109546 110832 109552 110844
rect 109604 110832 109610 110884
rect 113226 110560 113232 110612
rect 113284 110600 113290 110612
rect 114514 110600 114520 110612
rect 113284 110572 114520 110600
rect 113284 110560 113290 110572
rect 114514 110560 114520 110572
rect 114572 110560 114578 110612
rect 115802 110560 115808 110612
rect 115860 110600 115866 110612
rect 118286 110600 118292 110612
rect 115860 110572 118292 110600
rect 115860 110560 115866 110572
rect 118286 110560 118292 110572
rect 118344 110560 118350 110612
rect 113134 110492 113140 110544
rect 113192 110532 113198 110544
rect 113962 110532 113968 110544
rect 113192 110504 113968 110532
rect 113192 110492 113198 110504
rect 113962 110492 113968 110504
rect 114020 110492 114026 110544
rect 114606 110492 114612 110544
rect 114664 110532 114670 110544
rect 115618 110532 115624 110544
rect 114664 110504 115624 110532
rect 114664 110492 114670 110504
rect 115618 110492 115624 110504
rect 115676 110492 115682 110544
rect 115894 110492 115900 110544
rect 115952 110532 115958 110544
rect 116722 110532 116728 110544
rect 115952 110504 116728 110532
rect 115952 110492 115958 110504
rect 116722 110492 116728 110504
rect 116780 110492 116786 110544
rect 117458 110492 117464 110544
rect 117516 110532 117522 110544
rect 118838 110532 118844 110544
rect 117516 110504 118844 110532
rect 117516 110492 117522 110504
rect 118838 110492 118844 110504
rect 118896 110492 118902 110544
rect 31070 110424 31076 110476
rect 31128 110464 31134 110476
rect 31898 110464 31904 110476
rect 31128 110436 31904 110464
rect 31128 110424 31134 110436
rect 31898 110424 31904 110436
rect 31956 110424 31962 110476
rect 99518 110424 99524 110476
rect 99576 110464 99582 110476
rect 107338 110464 107344 110476
rect 99576 110436 107344 110464
rect 99576 110424 99582 110436
rect 107338 110424 107344 110436
rect 107396 110424 107402 110476
rect 183606 110356 183612 110408
rect 183664 110396 183670 110408
rect 191610 110396 191616 110408
rect 183664 110368 191616 110396
rect 183664 110356 183670 110368
rect 191610 110356 191616 110368
rect 191668 110356 191674 110408
rect 99426 110288 99432 110340
rect 99484 110328 99490 110340
rect 106786 110328 106792 110340
rect 99484 110300 106792 110328
rect 99484 110288 99490 110300
rect 106786 110288 106792 110300
rect 106844 110288 106850 110340
rect 115986 110288 115992 110340
rect 116044 110328 116050 110340
rect 117274 110328 117280 110340
rect 116044 110300 117280 110328
rect 116044 110288 116050 110300
rect 117274 110288 117280 110300
rect 117332 110288 117338 110340
rect 183698 110288 183704 110340
rect 183756 110328 183762 110340
rect 192162 110328 192168 110340
rect 183756 110300 192168 110328
rect 183756 110288 183762 110300
rect 192162 110288 192168 110300
rect 192220 110288 192226 110340
rect 208262 110288 208268 110340
rect 208320 110328 208326 110340
rect 213230 110328 213236 110340
rect 208320 110300 213236 110328
rect 208320 110288 208326 110300
rect 213230 110288 213236 110300
rect 213288 110288 213294 110340
rect 20214 110220 20220 110272
rect 20272 110260 20278 110272
rect 41742 110260 41748 110272
rect 20272 110232 41748 110260
rect 20272 110220 20278 110232
rect 41742 110220 41748 110232
rect 41800 110220 41806 110272
rect 98782 110220 98788 110272
rect 98840 110260 98846 110272
rect 107890 110260 107896 110272
rect 98840 110232 107896 110260
rect 98840 110220 98846 110232
rect 107890 110220 107896 110232
rect 107948 110220 107954 110272
rect 183514 110220 183520 110272
rect 183572 110260 183578 110272
rect 191058 110260 191064 110272
rect 183572 110232 191064 110260
rect 183572 110220 183578 110232
rect 191058 110220 191064 110232
rect 191116 110220 191122 110272
rect 191978 110220 191984 110272
rect 192036 110260 192042 110272
rect 215530 110260 215536 110272
rect 192036 110232 215536 110260
rect 192036 110220 192042 110232
rect 215530 110220 215536 110232
rect 215588 110220 215594 110272
rect 25918 109948 25924 110000
rect 25976 109988 25982 110000
rect 26286 109988 26292 110000
rect 25976 109960 26292 109988
rect 25976 109948 25982 109960
rect 26286 109948 26292 109960
rect 26344 109948 26350 110000
rect 29046 109948 29052 110000
rect 29104 109988 29110 110000
rect 30886 109988 30892 110000
rect 29104 109960 30892 109988
rect 29104 109948 29110 109960
rect 30886 109948 30892 109960
rect 30944 109948 30950 110000
rect 24906 109880 24912 109932
rect 24964 109920 24970 109932
rect 24964 109892 27528 109920
rect 24964 109880 24970 109892
rect 22882 109812 22888 109864
rect 22940 109852 22946 109864
rect 27298 109852 27304 109864
rect 22940 109824 27304 109852
rect 22940 109812 22946 109824
rect 27298 109812 27304 109824
rect 27356 109812 27362 109864
rect 27500 109852 27528 109892
rect 27666 109880 27672 109932
rect 27724 109920 27730 109932
rect 30058 109920 30064 109932
rect 27724 109892 30064 109920
rect 27724 109880 27730 109892
rect 30058 109880 30064 109892
rect 30116 109880 30122 109932
rect 28494 109852 28500 109864
rect 27500 109824 28500 109852
rect 28494 109812 28500 109824
rect 28552 109812 28558 109864
rect 99242 109812 99248 109864
rect 99300 109852 99306 109864
rect 106234 109852 106240 109864
rect 99300 109824 106240 109852
rect 99300 109812 99306 109824
rect 106234 109812 106240 109824
rect 106292 109812 106298 109864
rect 115710 109812 115716 109864
rect 115768 109852 115774 109864
rect 117826 109852 117832 109864
rect 115768 109824 117832 109852
rect 115768 109812 115774 109824
rect 117826 109812 117832 109824
rect 117884 109812 117890 109864
rect 118930 109812 118936 109864
rect 118988 109852 118994 109864
rect 119942 109852 119948 109864
rect 118988 109824 119948 109852
rect 118988 109812 118994 109824
rect 119942 109812 119948 109824
rect 120000 109812 120006 109864
rect 183330 109812 183336 109864
rect 183388 109852 183394 109864
rect 190414 109852 190420 109864
rect 183388 109824 190420 109852
rect 183388 109812 183394 109824
rect 190414 109812 190420 109824
rect 190472 109812 190478 109864
rect 23618 109744 23624 109796
rect 23676 109784 23682 109796
rect 27666 109784 27672 109796
rect 23676 109756 27672 109784
rect 23676 109744 23682 109756
rect 27666 109744 27672 109756
rect 27724 109744 27730 109796
rect 44410 109744 44416 109796
rect 44468 109784 44474 109796
rect 45054 109784 45060 109796
rect 44468 109756 45060 109784
rect 44468 109744 44474 109756
rect 45054 109744 45060 109756
rect 45112 109744 45118 109796
rect 99150 109744 99156 109796
rect 99208 109784 99214 109796
rect 105130 109784 105136 109796
rect 99208 109756 105136 109784
rect 99208 109744 99214 109756
rect 105130 109744 105136 109756
rect 105188 109744 105194 109796
rect 119574 109744 119580 109796
rect 119632 109784 119638 109796
rect 121046 109784 121052 109796
rect 119632 109756 121052 109784
rect 119632 109744 119638 109756
rect 121046 109744 121052 109756
rect 121104 109744 121110 109796
rect 126658 109744 126664 109796
rect 126716 109784 126722 109796
rect 129326 109784 129332 109796
rect 126716 109756 129332 109784
rect 126716 109744 126722 109756
rect 129326 109744 129332 109756
rect 129384 109744 129390 109796
rect 183238 109744 183244 109796
rect 183296 109784 183302 109796
rect 189310 109784 189316 109796
rect 183296 109756 189316 109784
rect 183296 109744 183302 109756
rect 189310 109744 189316 109756
rect 189368 109744 189374 109796
rect 205226 109744 205232 109796
rect 205284 109784 205290 109796
rect 206974 109784 206980 109796
rect 205284 109756 206980 109784
rect 205284 109744 205290 109756
rect 206974 109744 206980 109756
rect 207032 109744 207038 109796
rect 21502 109676 21508 109728
rect 21560 109716 21566 109728
rect 26470 109716 26476 109728
rect 21560 109688 26476 109716
rect 21560 109676 21566 109688
rect 26470 109676 26476 109688
rect 26528 109676 26534 109728
rect 37510 109676 37516 109728
rect 37568 109716 37574 109728
rect 38246 109716 38252 109728
rect 37568 109688 38252 109716
rect 37568 109676 37574 109688
rect 38246 109676 38252 109688
rect 38304 109676 38310 109728
rect 42938 109676 42944 109728
rect 42996 109716 43002 109728
rect 47446 109716 47452 109728
rect 42996 109688 47452 109716
rect 42996 109676 43002 109688
rect 47446 109676 47452 109688
rect 47504 109676 47510 109728
rect 99058 109676 99064 109728
rect 99116 109716 99122 109728
rect 104578 109716 104584 109728
rect 99116 109688 104584 109716
rect 99116 109676 99122 109688
rect 104578 109676 104584 109688
rect 104636 109676 104642 109728
rect 119942 109676 119948 109728
rect 120000 109716 120006 109728
rect 122150 109716 122156 109728
rect 120000 109688 122156 109716
rect 120000 109676 120006 109688
rect 122150 109676 122156 109688
rect 122208 109676 122214 109728
rect 183146 109676 183152 109728
rect 183204 109716 183210 109728
rect 188758 109716 188764 109728
rect 183204 109688 188764 109716
rect 183204 109676 183210 109688
rect 188758 109676 188764 109688
rect 188816 109676 188822 109728
rect 203754 109676 203760 109728
rect 203812 109716 203818 109728
rect 205318 109716 205324 109728
rect 203812 109688 205324 109716
rect 203812 109676 203818 109688
rect 205318 109676 205324 109688
rect 205376 109676 205382 109728
rect 208170 109676 208176 109728
rect 208228 109716 208234 109728
rect 212126 109716 212132 109728
rect 208228 109688 212132 109716
rect 208228 109676 208234 109688
rect 212126 109676 212132 109688
rect 212184 109676 212190 109728
rect 22238 109608 22244 109660
rect 22296 109648 22302 109660
rect 26838 109648 26844 109660
rect 22296 109620 26844 109648
rect 22296 109608 22302 109620
rect 26838 109608 26844 109620
rect 26896 109608 26902 109660
rect 27022 109608 27028 109660
rect 27080 109648 27086 109660
rect 29690 109648 29696 109660
rect 27080 109620 29696 109648
rect 27080 109608 27086 109620
rect 29690 109608 29696 109620
rect 29748 109608 29754 109660
rect 38154 109608 38160 109660
rect 38212 109648 38218 109660
rect 39994 109648 40000 109660
rect 38212 109620 40000 109648
rect 38212 109608 38218 109620
rect 39994 109608 40000 109620
rect 40052 109608 40058 109660
rect 45054 109608 45060 109660
rect 45112 109648 45118 109660
rect 46802 109648 46808 109660
rect 45112 109620 46808 109648
rect 45112 109608 45118 109620
rect 46802 109608 46808 109620
rect 46860 109608 46866 109660
rect 98966 109608 98972 109660
rect 99024 109648 99030 109660
rect 104118 109648 104124 109660
rect 99024 109620 104124 109648
rect 99024 109608 99030 109620
rect 104118 109608 104124 109620
rect 104176 109608 104182 109660
rect 119850 109608 119856 109660
rect 119908 109648 119914 109660
rect 121598 109648 121604 109660
rect 119908 109620 121604 109648
rect 119908 109608 119914 109620
rect 121598 109608 121604 109620
rect 121656 109608 121662 109660
rect 126474 109608 126480 109660
rect 126532 109648 126538 109660
rect 128774 109648 128780 109660
rect 126532 109620 128780 109648
rect 126532 109608 126538 109620
rect 128774 109608 128780 109620
rect 128832 109608 128838 109660
rect 129326 109608 129332 109660
rect 129384 109648 129390 109660
rect 130982 109648 130988 109660
rect 129384 109620 130988 109648
rect 129384 109608 129390 109620
rect 130982 109608 130988 109620
rect 131040 109608 131046 109660
rect 183054 109608 183060 109660
rect 183112 109648 183118 109660
rect 188206 109648 188212 109660
rect 183112 109620 188212 109648
rect 183112 109608 183118 109620
rect 188206 109608 188212 109620
rect 188264 109608 188270 109660
rect 201454 109608 201460 109660
rect 201512 109648 201518 109660
rect 202466 109648 202472 109660
rect 201512 109620 202472 109648
rect 201512 109608 201518 109620
rect 202466 109608 202472 109620
rect 202524 109608 202530 109660
rect 205134 109608 205140 109660
rect 205192 109648 205198 109660
rect 206422 109648 206428 109660
rect 205192 109620 206428 109648
rect 205192 109608 205198 109620
rect 206422 109608 206428 109620
rect 206480 109608 206486 109660
rect 208354 109608 208360 109660
rect 208412 109648 208418 109660
rect 212678 109648 212684 109660
rect 208412 109620 212684 109648
rect 208412 109608 208418 109620
rect 212678 109608 212684 109620
rect 212736 109608 212742 109660
rect 213506 109608 213512 109660
rect 213564 109648 213570 109660
rect 214978 109648 214984 109660
rect 213564 109620 214984 109648
rect 213564 109608 213570 109620
rect 214978 109608 214984 109620
rect 215036 109608 215042 109660
rect 20858 109540 20864 109592
rect 20916 109580 20922 109592
rect 22974 109580 22980 109592
rect 20916 109552 22980 109580
rect 20916 109540 20922 109552
rect 22974 109540 22980 109552
rect 23032 109540 23038 109592
rect 24262 109540 24268 109592
rect 24320 109580 24326 109592
rect 28126 109580 28132 109592
rect 24320 109552 28132 109580
rect 24320 109540 24326 109552
rect 28126 109540 28132 109552
rect 28184 109540 28190 109592
rect 28310 109540 28316 109592
rect 28368 109580 28374 109592
rect 29138 109580 29144 109592
rect 28368 109552 29144 109580
rect 28368 109540 28374 109552
rect 29138 109540 29144 109552
rect 29196 109540 29202 109592
rect 38246 109540 38252 109592
rect 38304 109580 38310 109592
rect 39258 109580 39264 109592
rect 38304 109552 39264 109580
rect 38304 109540 38310 109552
rect 39258 109540 39264 109552
rect 39316 109540 39322 109592
rect 45146 109540 45152 109592
rect 45204 109580 45210 109592
rect 46066 109580 46072 109592
rect 45204 109552 46072 109580
rect 45204 109540 45210 109552
rect 46066 109540 46072 109552
rect 46124 109540 46130 109592
rect 99334 109540 99340 109592
rect 99392 109580 99398 109592
rect 105682 109580 105688 109592
rect 99392 109552 105688 109580
rect 99392 109540 99398 109552
rect 105682 109540 105688 109552
rect 105740 109540 105746 109592
rect 119758 109540 119764 109592
rect 119816 109580 119822 109592
rect 120494 109580 120500 109592
rect 119816 109552 120500 109580
rect 119816 109540 119822 109552
rect 120494 109540 120500 109552
rect 120552 109540 120558 109592
rect 120954 109540 120960 109592
rect 121012 109580 121018 109592
rect 122702 109580 122708 109592
rect 121012 109552 122708 109580
rect 121012 109540 121018 109552
rect 122702 109540 122708 109552
rect 122760 109540 122766 109592
rect 126566 109540 126572 109592
rect 126624 109580 126630 109592
rect 128222 109580 128228 109592
rect 126624 109552 128228 109580
rect 126624 109540 126630 109552
rect 128222 109540 128228 109552
rect 128280 109540 128286 109592
rect 129234 109540 129240 109592
rect 129292 109580 129298 109592
rect 130430 109580 130436 109592
rect 129292 109552 130436 109580
rect 129292 109540 129298 109552
rect 130430 109540 130436 109552
rect 130488 109540 130494 109592
rect 183422 109540 183428 109592
rect 183480 109580 183486 109592
rect 189862 109580 189868 109592
rect 183480 109552 189868 109580
rect 183480 109540 183486 109552
rect 189862 109540 189868 109552
rect 189920 109540 189926 109592
rect 193910 109540 193916 109592
rect 193968 109580 193974 109592
rect 194738 109580 194744 109592
rect 193968 109552 194744 109580
rect 193968 109540 193974 109552
rect 194738 109540 194744 109552
rect 194796 109540 194802 109592
rect 201638 109540 201644 109592
rect 201696 109580 201702 109592
rect 203018 109580 203024 109592
rect 201696 109552 203024 109580
rect 201696 109540 201702 109552
rect 203018 109540 203024 109552
rect 203076 109540 203082 109592
rect 203846 109540 203852 109592
rect 203904 109580 203910 109592
rect 204674 109580 204680 109592
rect 203904 109552 204680 109580
rect 203904 109540 203910 109552
rect 204674 109540 204680 109552
rect 204732 109540 204738 109592
rect 205410 109540 205416 109592
rect 205468 109580 205474 109592
rect 205870 109580 205876 109592
rect 205468 109552 205876 109580
rect 205468 109540 205474 109552
rect 205870 109540 205876 109552
rect 205928 109540 205934 109592
rect 208538 109540 208544 109592
rect 208596 109580 208602 109592
rect 211574 109580 211580 109592
rect 208596 109552 211580 109580
rect 208596 109540 208602 109552
rect 211574 109540 211580 109552
rect 211632 109540 211638 109592
rect 213414 109540 213420 109592
rect 213472 109580 213478 109592
rect 214426 109580 214432 109592
rect 213472 109552 214432 109580
rect 213472 109540 213478 109552
rect 214426 109540 214432 109552
rect 214484 109540 214490 109592
rect 59314 108180 59320 108232
rect 59372 108180 59378 108232
rect 59332 108152 59360 108180
rect 59406 108152 59412 108164
rect 59332 108124 59412 108152
rect 59406 108112 59412 108124
rect 59464 108112 59470 108164
rect 41650 107500 41656 107552
rect 41708 107540 41714 107552
rect 42294 107540 42300 107552
rect 41708 107512 42300 107540
rect 41708 107500 41714 107512
rect 42294 107500 42300 107512
rect 42352 107500 42358 107552
rect 43030 107500 43036 107552
rect 43088 107540 43094 107552
rect 43766 107540 43772 107552
rect 43088 107512 43772 107540
rect 43088 107500 43094 107512
rect 43766 107500 43772 107512
rect 43824 107500 43830 107552
rect 208630 107500 208636 107552
rect 208688 107540 208694 107552
rect 208998 107540 209004 107552
rect 208688 107512 209004 107540
rect 208688 107500 208694 107512
rect 208998 107500 209004 107512
rect 209056 107500 209062 107552
rect 210010 107500 210016 107552
rect 210068 107540 210074 107552
rect 210654 107540 210660 107552
rect 210068 107512 210660 107540
rect 210068 107500 210074 107512
rect 210654 107500 210660 107512
rect 210712 107500 210718 107552
rect 30242 102604 30248 102656
rect 30300 102644 30306 102656
rect 31254 102644 31260 102656
rect 30300 102616 31260 102644
rect 30300 102604 30306 102616
rect 31254 102604 31260 102616
rect 31312 102604 31318 102656
rect 32082 102604 32088 102656
rect 32140 102644 32146 102656
rect 32818 102644 32824 102656
rect 32140 102616 32824 102644
rect 32140 102604 32146 102616
rect 32818 102604 32824 102616
rect 32876 102604 32882 102656
rect 35302 102604 35308 102656
rect 35360 102644 35366 102656
rect 36130 102644 36136 102656
rect 35360 102616 36136 102644
rect 35360 102604 35366 102616
rect 36130 102604 36136 102616
rect 36188 102604 36194 102656
rect 36866 102604 36872 102656
rect 36924 102644 36930 102656
rect 38246 102644 38252 102656
rect 36924 102616 38252 102644
rect 36924 102604 36930 102616
rect 38246 102604 38252 102616
rect 38304 102604 38310 102656
rect 111294 102604 111300 102656
rect 111352 102644 111358 102656
rect 111754 102644 111760 102656
rect 111352 102616 111760 102644
rect 111352 102604 111358 102616
rect 111754 102604 111760 102616
rect 111812 102604 111818 102656
rect 112490 102604 112496 102656
rect 112548 102644 112554 102656
rect 113318 102644 113324 102656
rect 112548 102616 113324 102644
rect 112548 102604 112554 102616
rect 113318 102604 113324 102616
rect 113376 102604 113382 102656
rect 113686 102604 113692 102656
rect 113744 102644 113750 102656
rect 114698 102644 114704 102656
rect 113744 102616 114704 102644
rect 113744 102604 113750 102616
rect 114698 102604 114704 102616
rect 114756 102604 114762 102656
rect 193266 102604 193272 102656
rect 193324 102644 193330 102656
rect 194094 102644 194100 102656
rect 193324 102616 194100 102644
rect 193324 102604 193330 102616
rect 194094 102604 194100 102616
rect 194152 102604 194158 102656
rect 196302 102604 196308 102656
rect 196360 102644 196366 102656
rect 196854 102644 196860 102656
rect 196360 102616 196860 102644
rect 196360 102604 196366 102616
rect 196854 102604 196860 102616
rect 196912 102604 196918 102656
rect 198418 102604 198424 102656
rect 198476 102644 198482 102656
rect 199154 102644 199160 102656
rect 198476 102616 199160 102644
rect 198476 102604 198482 102616
rect 199154 102604 199160 102616
rect 199212 102604 199218 102656
rect 199614 102604 199620 102656
rect 199672 102644 199678 102656
rect 200350 102644 200356 102656
rect 199672 102616 200356 102644
rect 199672 102604 199678 102616
rect 200350 102604 200356 102616
rect 200408 102604 200414 102656
rect 200810 102604 200816 102656
rect 200868 102644 200874 102656
rect 201362 102644 201368 102656
rect 200868 102616 201368 102644
rect 200868 102604 200874 102616
rect 201362 102604 201368 102616
rect 201420 102604 201426 102656
rect 201454 102604 201460 102656
rect 201512 102644 201518 102656
rect 203110 102644 203116 102656
rect 201512 102616 203116 102644
rect 201512 102604 201518 102616
rect 203110 102604 203116 102616
rect 203168 102604 203174 102656
rect 204858 102604 204864 102656
rect 204916 102644 204922 102656
rect 207342 102644 207348 102656
rect 204916 102616 207348 102644
rect 204916 102604 204922 102616
rect 207342 102604 207348 102616
rect 207400 102604 207406 102656
rect 32726 102536 32732 102588
rect 32784 102576 32790 102588
rect 33278 102576 33284 102588
rect 32784 102548 33284 102576
rect 32784 102536 32790 102548
rect 33278 102536 33284 102548
rect 33336 102536 33342 102588
rect 35670 102536 35676 102588
rect 35728 102576 35734 102588
rect 36774 102576 36780 102588
rect 35728 102548 36780 102576
rect 35728 102536 35734 102548
rect 36774 102536 36780 102548
rect 36832 102536 36838 102588
rect 37694 102536 37700 102588
rect 37752 102576 37758 102588
rect 40270 102576 40276 102588
rect 37752 102548 40276 102576
rect 37752 102536 37758 102548
rect 40270 102536 40276 102548
rect 40328 102536 40334 102588
rect 111662 102536 111668 102588
rect 111720 102576 111726 102588
rect 112306 102576 112312 102588
rect 111720 102548 112312 102576
rect 111720 102536 111726 102548
rect 112306 102536 112312 102548
rect 112364 102536 112370 102588
rect 119666 102536 119672 102588
rect 119724 102576 119730 102588
rect 123254 102576 123260 102588
rect 119724 102548 123260 102576
rect 119724 102536 119730 102548
rect 123254 102536 123260 102548
rect 123312 102536 123318 102588
rect 200074 102536 200080 102588
rect 200132 102576 200138 102588
rect 200626 102576 200632 102588
rect 200132 102548 200632 102576
rect 200132 102536 200138 102548
rect 200626 102536 200632 102548
rect 200684 102536 200690 102588
rect 201270 102536 201276 102588
rect 201328 102576 201334 102588
rect 201638 102576 201644 102588
rect 201328 102548 201644 102576
rect 201328 102536 201334 102548
rect 201638 102536 201644 102548
rect 201696 102536 201702 102588
rect 203294 102536 203300 102588
rect 203352 102576 203358 102588
rect 205410 102576 205416 102588
rect 203352 102548 205416 102576
rect 203352 102536 203358 102548
rect 205410 102536 205416 102548
rect 205468 102536 205474 102588
rect 206422 102536 206428 102588
rect 206480 102576 206486 102588
rect 210102 102576 210108 102588
rect 206480 102548 210108 102576
rect 206480 102536 206486 102548
rect 210102 102536 210108 102548
rect 210160 102536 210166 102588
rect 36038 102468 36044 102520
rect 36096 102508 36102 102520
rect 37602 102508 37608 102520
rect 36096 102480 37608 102508
rect 36096 102468 36102 102480
rect 37602 102468 37608 102480
rect 37660 102468 37666 102520
rect 38062 102468 38068 102520
rect 38120 102508 38126 102520
rect 40822 102508 40828 102520
rect 38120 102480 40828 102508
rect 38120 102468 38126 102480
rect 40822 102468 40828 102480
rect 40880 102468 40886 102520
rect 114054 102468 114060 102520
rect 114112 102508 114118 102520
rect 114606 102508 114612 102520
rect 114112 102480 114612 102508
rect 114112 102468 114118 102480
rect 114606 102468 114612 102480
rect 114664 102468 114670 102520
rect 115250 102468 115256 102520
rect 115308 102508 115314 102520
rect 115986 102508 115992 102520
rect 115308 102480 115992 102508
rect 115308 102468 115314 102480
rect 115986 102468 115992 102480
rect 116044 102468 116050 102520
rect 120862 102468 120868 102520
rect 120920 102508 120926 102520
rect 124910 102508 124916 102520
rect 120920 102480 124916 102508
rect 120920 102468 120926 102480
rect 124910 102468 124916 102480
rect 124968 102468 124974 102520
rect 22974 102400 22980 102452
rect 23032 102440 23038 102452
rect 26102 102440 26108 102452
rect 23032 102412 26108 102440
rect 23032 102400 23038 102412
rect 26102 102400 26108 102412
rect 26160 102400 26166 102452
rect 93354 102400 93360 102452
rect 93412 102440 93418 102452
rect 94182 102440 94188 102452
rect 93412 102412 94188 102440
rect 93412 102400 93418 102412
rect 94182 102400 94188 102412
rect 94240 102400 94246 102452
rect 120034 102400 120040 102452
rect 120092 102440 120098 102452
rect 123806 102440 123812 102452
rect 120092 102412 123812 102440
rect 120092 102400 120098 102412
rect 123806 102400 123812 102412
rect 123864 102400 123870 102452
rect 202466 102400 202472 102452
rect 202524 102440 202530 102452
rect 203846 102440 203852 102452
rect 202524 102412 203852 102440
rect 202524 102400 202530 102412
rect 203846 102400 203852 102412
rect 203904 102400 203910 102452
rect 50942 102332 50948 102384
rect 51000 102372 51006 102384
rect 59774 102372 59780 102384
rect 51000 102344 59780 102372
rect 51000 102332 51006 102344
rect 59774 102332 59780 102344
rect 59832 102332 59838 102384
rect 114422 102332 114428 102384
rect 114480 102372 114486 102384
rect 116170 102372 116176 102384
rect 114480 102344 116176 102372
rect 114480 102332 114486 102344
rect 116170 102332 116176 102344
rect 116228 102332 116234 102384
rect 122426 102332 122432 102384
rect 122484 102372 122490 102384
rect 127118 102372 127124 102384
rect 122484 102344 127124 102372
rect 122484 102332 122490 102344
rect 127118 102332 127124 102344
rect 127176 102332 127182 102384
rect 135122 102332 135128 102384
rect 135180 102372 135186 102384
rect 143770 102372 143776 102384
rect 135180 102344 143776 102372
rect 135180 102332 135186 102344
rect 143770 102332 143776 102344
rect 143828 102332 143834 102384
rect 159318 102332 159324 102384
rect 159376 102372 159382 102384
rect 161710 102372 161716 102384
rect 159376 102344 161716 102372
rect 159376 102332 159382 102344
rect 161710 102332 161716 102344
rect 161768 102332 161774 102384
rect 206054 102332 206060 102384
rect 206112 102372 206118 102384
rect 208814 102372 208820 102384
rect 206112 102344 208820 102372
rect 206112 102332 206118 102344
rect 208814 102332 208820 102344
rect 208872 102332 208878 102384
rect 122058 102264 122064 102316
rect 122116 102304 122122 102316
rect 126106 102304 126112 102316
rect 122116 102276 126112 102304
rect 122116 102264 122122 102276
rect 126106 102264 126112 102276
rect 126164 102264 126170 102316
rect 50666 102196 50672 102248
rect 50724 102236 50730 102248
rect 60878 102236 60884 102248
rect 50724 102208 60884 102236
rect 50724 102196 50730 102208
rect 60878 102196 60884 102208
rect 60936 102196 60942 102248
rect 121690 102196 121696 102248
rect 121748 102236 121754 102248
rect 126014 102236 126020 102248
rect 121748 102208 126020 102236
rect 121748 102196 121754 102208
rect 126014 102196 126020 102208
rect 126072 102196 126078 102248
rect 134846 102196 134852 102248
rect 134904 102236 134910 102248
rect 144874 102236 144880 102248
rect 134904 102208 144880 102236
rect 134904 102196 134910 102208
rect 144874 102196 144880 102208
rect 144932 102196 144938 102248
rect 200442 102196 200448 102248
rect 200500 102236 200506 102248
rect 201546 102236 201552 102248
rect 200500 102208 201552 102236
rect 200500 102196 200506 102208
rect 201546 102196 201552 102208
rect 201604 102196 201610 102248
rect 208814 102196 208820 102248
rect 208872 102236 208878 102248
rect 212862 102236 212868 102248
rect 208872 102208 212868 102236
rect 208872 102196 208878 102208
rect 212862 102196 212868 102208
rect 212920 102196 212926 102248
rect 50850 102128 50856 102180
rect 50908 102168 50914 102180
rect 61982 102168 61988 102180
rect 50908 102140 61988 102168
rect 50908 102128 50914 102140
rect 61982 102128 61988 102140
rect 62040 102128 62046 102180
rect 120494 102128 120500 102180
rect 120552 102168 120558 102180
rect 124358 102168 124364 102180
rect 120552 102140 124364 102168
rect 120552 102128 120558 102140
rect 124358 102128 124364 102140
rect 124416 102128 124422 102180
rect 135030 102128 135036 102180
rect 135088 102168 135094 102180
rect 145978 102168 145984 102180
rect 135088 102140 145984 102168
rect 135088 102128 135094 102140
rect 145978 102128 145984 102140
rect 146036 102128 146042 102180
rect 50758 102060 50764 102112
rect 50816 102100 50822 102112
rect 63086 102100 63092 102112
rect 50816 102072 63092 102100
rect 50816 102060 50822 102072
rect 63086 102060 63092 102072
rect 63144 102060 63150 102112
rect 88662 102060 88668 102112
rect 88720 102100 88726 102112
rect 101818 102100 101824 102112
rect 88720 102072 101824 102100
rect 88720 102060 88726 102072
rect 101818 102060 101824 102072
rect 101876 102060 101882 102112
rect 122886 102060 122892 102112
rect 122944 102100 122950 102112
rect 127670 102100 127676 102112
rect 122944 102072 127676 102100
rect 122944 102060 122950 102072
rect 127670 102060 127676 102072
rect 127728 102060 127734 102112
rect 134754 102060 134760 102112
rect 134812 102100 134818 102112
rect 147082 102100 147088 102112
rect 134812 102072 147088 102100
rect 134812 102060 134818 102072
rect 147082 102060 147088 102072
rect 147140 102060 147146 102112
rect 172658 102060 172664 102112
rect 172716 102100 172722 102112
rect 185814 102100 185820 102112
rect 172716 102072 185820 102100
rect 172716 102060 172722 102072
rect 185814 102060 185820 102072
rect 185872 102060 185878 102112
rect 199246 102060 199252 102112
rect 199304 102100 199310 102112
rect 199706 102100 199712 102112
rect 199304 102072 199712 102100
rect 199304 102060 199310 102072
rect 199706 102060 199712 102072
rect 199764 102060 199770 102112
rect 202098 102060 202104 102112
rect 202156 102100 202162 102112
rect 203202 102100 203208 102112
rect 202156 102072 203208 102100
rect 202156 102060 202162 102072
rect 203202 102060 203208 102072
rect 203260 102060 203266 102112
rect 204030 102060 204036 102112
rect 204088 102100 204094 102112
rect 205226 102100 205232 102112
rect 204088 102072 205232 102100
rect 204088 102060 204094 102072
rect 205226 102060 205232 102072
rect 205284 102060 205290 102112
rect 209274 102060 209280 102112
rect 209332 102100 209338 102112
rect 213414 102100 213420 102112
rect 209332 102072 213420 102100
rect 209332 102060 209338 102072
rect 213414 102060 213420 102072
rect 213472 102060 213478 102112
rect 26286 101992 26292 102044
rect 26344 102032 26350 102044
rect 28862 102032 28868 102044
rect 26344 102004 28868 102032
rect 26344 101992 26350 102004
rect 28862 101992 28868 102004
rect 28920 101992 28926 102044
rect 29138 101992 29144 102044
rect 29196 102032 29202 102044
rect 30426 102032 30432 102044
rect 29196 102004 30432 102032
rect 29196 101992 29202 102004
rect 30426 101992 30432 102004
rect 30484 101992 30490 102044
rect 36498 101992 36504 102044
rect 36556 102032 36562 102044
rect 37510 102032 37516 102044
rect 36556 102004 37516 102032
rect 36556 101992 36562 102004
rect 37510 101992 37516 102004
rect 37568 101992 37574 102044
rect 50574 101992 50580 102044
rect 50632 102032 50638 102044
rect 64190 102032 64196 102044
rect 50632 102004 64196 102032
rect 50632 101992 50638 102004
rect 64190 101992 64196 102004
rect 64248 101992 64254 102044
rect 87558 101992 87564 102044
rect 87616 102032 87622 102044
rect 102002 102032 102008 102044
rect 87616 102004 102008 102032
rect 87616 101992 87622 102004
rect 102002 101992 102008 102004
rect 102060 101992 102066 102044
rect 114882 101992 114888 102044
rect 114940 102032 114946 102044
rect 115894 102032 115900 102044
rect 114940 102004 115900 102032
rect 114940 101992 114946 102004
rect 115894 101992 115900 102004
rect 115952 101992 115958 102044
rect 134938 101992 134944 102044
rect 134996 102032 135002 102044
rect 148186 102032 148192 102044
rect 134996 102004 148192 102032
rect 134996 101992 135002 102004
rect 148186 101992 148192 102004
rect 148244 101992 148250 102044
rect 161526 101992 161532 102044
rect 161584 102032 161590 102044
rect 164470 102032 164476 102044
rect 161584 102004 164476 102032
rect 161584 101992 161590 102004
rect 164470 101992 164476 102004
rect 164528 101992 164534 102044
rect 171554 101992 171560 102044
rect 171612 102032 171618 102044
rect 185998 102032 186004 102044
rect 171612 102004 186004 102032
rect 171612 101992 171618 102004
rect 185998 101992 186004 102004
rect 186056 101992 186062 102044
rect 209642 101992 209648 102044
rect 209700 102032 209706 102044
rect 213506 102032 213512 102044
rect 209700 102004 213512 102032
rect 209700 101992 209706 102004
rect 213506 101992 213512 102004
rect 213564 101992 213570 102044
rect 51126 101924 51132 101976
rect 51184 101964 51190 101976
rect 58670 101964 58676 101976
rect 51184 101936 58676 101964
rect 51184 101924 51190 101936
rect 58670 101924 58676 101936
rect 58728 101924 58734 101976
rect 59406 101924 59412 101976
rect 59464 101964 59470 101976
rect 83142 101964 83148 101976
rect 59464 101936 83148 101964
rect 59464 101924 59470 101936
rect 83142 101924 83148 101936
rect 83200 101924 83206 101976
rect 86454 101924 86460 101976
rect 86512 101964 86518 101976
rect 101634 101964 101640 101976
rect 86512 101936 101640 101964
rect 86512 101924 86518 101936
rect 101634 101924 101640 101936
rect 101692 101924 101698 101976
rect 112030 101924 112036 101976
rect 112088 101964 112094 101976
rect 112858 101964 112864 101976
rect 112088 101936 112864 101964
rect 112088 101924 112094 101936
rect 112858 101924 112864 101936
rect 112916 101924 112922 101976
rect 135306 101924 135312 101976
rect 135364 101964 135370 101976
rect 142666 101964 142672 101976
rect 135364 101936 142672 101964
rect 135364 101924 135370 101936
rect 142666 101924 142672 101936
rect 142724 101924 142730 101976
rect 143678 101924 143684 101976
rect 143736 101964 143742 101976
rect 167138 101964 167144 101976
rect 143736 101936 167144 101964
rect 143736 101924 143742 101936
rect 167138 101924 167144 101936
rect 167196 101924 167202 101976
rect 170450 101924 170456 101976
rect 170508 101964 170514 101976
rect 186182 101964 186188 101976
rect 170508 101936 186188 101964
rect 170508 101924 170514 101936
rect 186182 101924 186188 101936
rect 186240 101924 186246 101976
rect 40086 101856 40092 101908
rect 40144 101896 40150 101908
rect 44502 101896 44508 101908
rect 40144 101868 44508 101896
rect 40144 101856 40150 101868
rect 44502 101856 44508 101868
rect 44560 101856 44566 101908
rect 30518 101788 30524 101840
rect 30576 101828 30582 101840
rect 31622 101828 31628 101840
rect 30576 101800 31628 101828
rect 30576 101788 30582 101800
rect 31622 101788 31628 101800
rect 31680 101788 31686 101840
rect 37234 101788 37240 101840
rect 37292 101828 37298 101840
rect 38154 101828 38160 101840
rect 37292 101800 38160 101828
rect 37292 101788 37298 101800
rect 38154 101788 38160 101800
rect 38212 101788 38218 101840
rect 39258 101788 39264 101840
rect 39316 101828 39322 101840
rect 43122 101828 43128 101840
rect 39316 101800 43128 101828
rect 39316 101788 39322 101800
rect 43122 101788 43128 101800
rect 43180 101788 43186 101840
rect 116446 101788 116452 101840
rect 116504 101828 116510 101840
rect 117458 101828 117464 101840
rect 116504 101800 117464 101828
rect 116504 101788 116510 101800
rect 117458 101788 117464 101800
rect 117516 101788 117522 101840
rect 124450 101788 124456 101840
rect 124508 101828 124514 101840
rect 129878 101828 129884 101840
rect 124508 101800 129884 101828
rect 124508 101788 124514 101800
rect 129878 101788 129884 101800
rect 129936 101788 129942 101840
rect 205226 101788 205232 101840
rect 205284 101828 205290 101840
rect 208722 101828 208728 101840
rect 205284 101800 208728 101828
rect 205284 101788 205290 101800
rect 208722 101788 208728 101800
rect 208780 101788 208786 101840
rect 26378 101720 26384 101772
rect 26436 101760 26442 101772
rect 29230 101760 29236 101772
rect 26436 101732 29236 101760
rect 26436 101720 26442 101732
rect 29230 101720 29236 101732
rect 29288 101720 29294 101772
rect 38430 101720 38436 101772
rect 38488 101760 38494 101772
rect 41834 101760 41840 101772
rect 38488 101732 41840 101760
rect 38488 101720 38494 101732
rect 41834 101720 41840 101732
rect 41892 101720 41898 101772
rect 51034 101720 51040 101772
rect 51092 101760 51098 101772
rect 56462 101760 56468 101772
rect 51092 101732 56468 101760
rect 51092 101720 51098 101732
rect 56462 101720 56468 101732
rect 56520 101720 56526 101772
rect 121230 101720 121236 101772
rect 121288 101760 121294 101772
rect 125462 101760 125468 101772
rect 121288 101732 125468 101760
rect 121288 101720 121294 101732
rect 125462 101720 125468 101732
rect 125520 101720 125526 101772
rect 206882 101720 206888 101772
rect 206940 101760 206946 101772
rect 210010 101760 210016 101772
rect 206940 101732 210016 101760
rect 206940 101720 206946 101732
rect 210010 101720 210016 101732
rect 210068 101720 210074 101772
rect 40822 101652 40828 101704
rect 40880 101692 40886 101704
rect 45146 101692 45152 101704
rect 40880 101664 45152 101692
rect 40880 101652 40886 101664
rect 45146 101652 45152 101664
rect 45204 101652 45210 101704
rect 116814 101652 116820 101704
rect 116872 101692 116878 101704
rect 119390 101692 119396 101704
rect 116872 101664 119396 101692
rect 116872 101652 116878 101664
rect 119390 101652 119396 101664
rect 119448 101652 119454 101704
rect 123254 101652 123260 101704
rect 123312 101692 123318 101704
rect 126566 101692 126572 101704
rect 123312 101664 126572 101692
rect 123312 101652 123318 101664
rect 126566 101652 126572 101664
rect 126624 101652 126630 101704
rect 202834 101652 202840 101704
rect 202892 101692 202898 101704
rect 203754 101692 203760 101704
rect 202892 101664 203760 101692
rect 202892 101652 202898 101664
rect 203754 101652 203760 101664
rect 203812 101652 203818 101704
rect 204490 101652 204496 101704
rect 204548 101692 204554 101704
rect 207250 101692 207256 101704
rect 204548 101664 207256 101692
rect 204548 101652 204554 101664
rect 207250 101652 207256 101664
rect 207308 101652 207314 101704
rect 39626 101584 39632 101636
rect 39684 101624 39690 101636
rect 43030 101624 43036 101636
rect 39684 101596 43036 101624
rect 39684 101584 39690 101596
rect 43030 101584 43036 101596
rect 43088 101584 43094 101636
rect 117642 101584 117648 101636
rect 117700 101624 117706 101636
rect 119758 101624 119764 101636
rect 117700 101596 119764 101624
rect 117700 101584 117706 101596
rect 119758 101584 119764 101596
rect 119816 101584 119822 101636
rect 124818 101584 124824 101636
rect 124876 101624 124882 101636
rect 129234 101624 129240 101636
rect 124876 101596 129240 101624
rect 124876 101584 124882 101596
rect 129234 101584 129240 101596
rect 129292 101584 129298 101636
rect 40454 101516 40460 101568
rect 40512 101556 40518 101568
rect 44410 101556 44416 101568
rect 40512 101528 44416 101556
rect 40512 101516 40518 101528
rect 44410 101516 44416 101528
rect 44468 101516 44474 101568
rect 75322 101516 75328 101568
rect 75380 101556 75386 101568
rect 77530 101556 77536 101568
rect 75380 101528 77536 101556
rect 75380 101516 75386 101528
rect 77530 101516 77536 101528
rect 77588 101516 77594 101568
rect 118470 101516 118476 101568
rect 118528 101556 118534 101568
rect 119850 101556 119856 101568
rect 118528 101528 119856 101556
rect 118528 101516 118534 101528
rect 119850 101516 119856 101528
rect 119908 101516 119914 101568
rect 123622 101516 123628 101568
rect 123680 101556 123686 101568
rect 126474 101556 126480 101568
rect 123680 101528 126480 101556
rect 123680 101516 123686 101528
rect 126474 101516 126480 101528
rect 126532 101516 126538 101568
rect 207618 101516 207624 101568
rect 207676 101556 207682 101568
rect 208170 101556 208176 101568
rect 207676 101528 208176 101556
rect 207676 101516 207682 101528
rect 208170 101516 208176 101528
rect 208228 101516 208234 101568
rect 38890 101448 38896 101500
rect 38948 101488 38954 101500
rect 41650 101488 41656 101500
rect 38948 101460 41656 101488
rect 38948 101448 38954 101460
rect 41650 101448 41656 101460
rect 41708 101448 41714 101500
rect 118838 101448 118844 101500
rect 118896 101488 118902 101500
rect 119942 101488 119948 101500
rect 118896 101460 119948 101488
rect 118896 101448 118902 101460
rect 119942 101448 119948 101460
rect 120000 101448 120006 101500
rect 124082 101448 124088 101500
rect 124140 101488 124146 101500
rect 126658 101488 126664 101500
rect 124140 101460 126664 101488
rect 124140 101448 124146 101460
rect 126658 101448 126664 101460
rect 126716 101448 126722 101500
rect 194646 101448 194652 101500
rect 194704 101488 194710 101500
rect 195290 101488 195296 101500
rect 194704 101460 195296 101488
rect 194704 101448 194710 101460
rect 195290 101448 195296 101460
rect 195348 101448 195354 101500
rect 203662 101448 203668 101500
rect 203720 101488 203726 101500
rect 205134 101488 205140 101500
rect 203720 101460 205140 101488
rect 203720 101448 203726 101460
rect 205134 101448 205140 101460
rect 205192 101448 205198 101500
rect 205686 101448 205692 101500
rect 205744 101488 205750 101500
rect 208630 101488 208636 101500
rect 205744 101460 208636 101488
rect 205744 101448 205750 101460
rect 208630 101448 208636 101460
rect 208688 101448 208694 101500
rect 31806 101380 31812 101432
rect 31864 101420 31870 101432
rect 32450 101420 32456 101432
rect 31864 101392 32456 101420
rect 31864 101380 31870 101392
rect 32450 101380 32456 101392
rect 32508 101380 32514 101432
rect 41282 101380 41288 101432
rect 41340 101420 41346 101432
rect 45054 101420 45060 101432
rect 41340 101392 45060 101420
rect 41340 101380 41346 101392
rect 45054 101380 45060 101392
rect 45112 101380 45118 101432
rect 72378 101380 72384 101432
rect 72436 101420 72442 101432
rect 73482 101420 73488 101432
rect 72436 101392 73488 101420
rect 72436 101380 72442 101392
rect 73482 101380 73488 101392
rect 73540 101380 73546 101432
rect 77530 101380 77536 101432
rect 77588 101420 77594 101432
rect 79554 101420 79560 101432
rect 77588 101392 79560 101420
rect 77588 101380 77594 101392
rect 79554 101380 79560 101392
rect 79612 101380 79618 101432
rect 80842 101380 80848 101432
rect 80900 101420 80906 101432
rect 82314 101420 82320 101432
rect 80900 101392 82320 101420
rect 80900 101380 80906 101392
rect 82314 101380 82320 101392
rect 82372 101380 82378 101432
rect 117274 101380 117280 101432
rect 117332 101420 117338 101432
rect 118930 101420 118936 101432
rect 117332 101392 118936 101420
rect 117332 101380 117338 101392
rect 118930 101380 118936 101392
rect 118988 101380 118994 101432
rect 119298 101380 119304 101432
rect 119356 101420 119362 101432
rect 120954 101420 120960 101432
rect 119356 101392 120960 101420
rect 119356 101380 119362 101392
rect 120954 101380 120960 101392
rect 121012 101380 121018 101432
rect 125646 101380 125652 101432
rect 125704 101420 125710 101432
rect 131534 101420 131540 101432
rect 125704 101392 131540 101420
rect 125704 101380 125710 101392
rect 131534 101380 131540 101392
rect 131592 101380 131598 101432
rect 154902 101380 154908 101432
rect 154960 101420 154966 101432
rect 156190 101420 156196 101432
rect 154960 101392 156196 101420
rect 154960 101380 154966 101392
rect 156190 101380 156196 101392
rect 156248 101380 156254 101432
rect 158214 101380 158220 101432
rect 158272 101420 158278 101432
rect 158858 101420 158864 101432
rect 158272 101392 158864 101420
rect 158272 101380 158278 101392
rect 158858 101380 158864 101392
rect 158916 101380 158922 101432
rect 163734 101380 163740 101432
rect 163792 101420 163798 101432
rect 165114 101420 165120 101432
rect 163792 101392 165120 101420
rect 163792 101380 163798 101392
rect 165114 101380 165120 101392
rect 165172 101380 165178 101432
rect 165942 101380 165948 101432
rect 166000 101420 166006 101432
rect 167874 101420 167880 101432
rect 166000 101392 167880 101420
rect 166000 101380 166006 101392
rect 167874 101380 167880 101392
rect 167932 101380 167938 101432
rect 176154 101380 176160 101432
rect 176212 101420 176218 101432
rect 179282 101420 179288 101432
rect 176212 101392 179288 101420
rect 176212 101380 176218 101392
rect 179282 101380 179288 101392
rect 179340 101380 179346 101432
rect 193358 101380 193364 101432
rect 193416 101420 193422 101432
rect 194462 101420 194468 101432
rect 193416 101392 194468 101420
rect 193416 101380 193422 101392
rect 194462 101380 194468 101392
rect 194520 101380 194526 101432
rect 194738 101380 194744 101432
rect 194796 101420 194802 101432
rect 195014 101420 195020 101432
rect 194796 101392 195020 101420
rect 194796 101380 194802 101392
rect 195014 101380 195020 101392
rect 195072 101380 195078 101432
rect 195106 101380 195112 101432
rect 195164 101420 195170 101432
rect 196026 101420 196032 101432
rect 195164 101392 196032 101420
rect 195164 101380 195170 101392
rect 196026 101380 196032 101392
rect 196084 101380 196090 101432
rect 207250 101380 207256 101432
rect 207308 101420 207314 101432
rect 208538 101420 208544 101432
rect 207308 101392 208544 101420
rect 207308 101380 207314 101392
rect 208538 101380 208544 101392
rect 208596 101380 208602 101432
rect 41650 101312 41656 101364
rect 41708 101352 41714 101364
rect 42938 101352 42944 101364
rect 41708 101324 42944 101352
rect 41708 101312 41714 101324
rect 42938 101312 42944 101324
rect 42996 101312 43002 101364
rect 68606 101312 68612 101364
rect 68664 101352 68670 101364
rect 69250 101352 69256 101364
rect 68664 101324 69256 101352
rect 68664 101312 68670 101324
rect 69250 101312 69256 101324
rect 69308 101312 69314 101364
rect 69802 101312 69808 101364
rect 69860 101352 69866 101364
rect 70630 101352 70636 101364
rect 69860 101324 70636 101352
rect 69860 101312 69866 101324
rect 70630 101312 70636 101324
rect 70688 101312 70694 101364
rect 70906 101312 70912 101364
rect 70964 101352 70970 101364
rect 72010 101352 72016 101364
rect 70964 101324 72016 101352
rect 70964 101312 70970 101324
rect 72010 101312 72016 101324
rect 72068 101312 72074 101364
rect 73114 101312 73120 101364
rect 73172 101352 73178 101364
rect 74034 101352 74040 101364
rect 73172 101324 74040 101352
rect 73172 101312 73178 101324
rect 74034 101312 74040 101324
rect 74092 101312 74098 101364
rect 76426 101312 76432 101364
rect 76484 101352 76490 101364
rect 77438 101352 77444 101364
rect 76484 101324 77444 101352
rect 76484 101312 76490 101324
rect 77438 101312 77444 101324
rect 77496 101312 77502 101364
rect 78634 101312 78640 101364
rect 78692 101352 78698 101364
rect 79646 101352 79652 101364
rect 78692 101324 79652 101352
rect 78692 101312 78698 101324
rect 79646 101312 79652 101324
rect 79704 101312 79710 101364
rect 79738 101312 79744 101364
rect 79796 101352 79802 101364
rect 80934 101352 80940 101364
rect 79796 101324 80940 101352
rect 79796 101312 79802 101324
rect 80934 101312 80940 101324
rect 80992 101312 80998 101364
rect 81946 101312 81952 101364
rect 82004 101352 82010 101364
rect 83694 101352 83700 101364
rect 82004 101324 83700 101352
rect 82004 101312 82010 101324
rect 83694 101312 83700 101324
rect 83752 101312 83758 101364
rect 89766 101312 89772 101364
rect 89824 101352 89830 101364
rect 90594 101352 90600 101364
rect 89824 101324 90600 101352
rect 89824 101312 89830 101324
rect 90594 101312 90600 101324
rect 90652 101312 90658 101364
rect 91974 101312 91980 101364
rect 92032 101352 92038 101364
rect 92618 101352 92624 101364
rect 92032 101324 92624 101352
rect 92032 101312 92038 101324
rect 92618 101312 92624 101324
rect 92676 101312 92682 101364
rect 93078 101312 93084 101364
rect 93136 101352 93142 101364
rect 93998 101352 94004 101364
rect 93136 101324 94004 101352
rect 93136 101312 93142 101324
rect 93998 101312 94004 101324
rect 94056 101312 94062 101364
rect 118102 101312 118108 101364
rect 118160 101352 118166 101364
rect 119574 101352 119580 101364
rect 118160 101324 119580 101352
rect 118160 101312 118166 101324
rect 119574 101312 119580 101324
rect 119632 101312 119638 101364
rect 125278 101312 125284 101364
rect 125336 101352 125342 101364
rect 129326 101352 129332 101364
rect 125336 101324 129332 101352
rect 125336 101312 125342 101324
rect 129326 101312 129332 101324
rect 129384 101312 129390 101364
rect 135214 101312 135220 101364
rect 135272 101352 135278 101364
rect 140458 101352 140464 101364
rect 135272 101324 140464 101352
rect 135272 101312 135278 101324
rect 140458 101312 140464 101324
rect 140516 101312 140522 101364
rect 152602 101312 152608 101364
rect 152660 101352 152666 101364
rect 153430 101352 153436 101364
rect 152660 101324 153436 101352
rect 152660 101312 152666 101324
rect 153430 101312 153436 101324
rect 153488 101312 153494 101364
rect 153798 101312 153804 101364
rect 153856 101352 153862 101364
rect 154810 101352 154816 101364
rect 153856 101324 154816 101352
rect 153856 101312 153862 101324
rect 154810 101312 154816 101324
rect 154868 101312 154874 101364
rect 156006 101312 156012 101364
rect 156064 101352 156070 101364
rect 156834 101352 156840 101364
rect 156064 101324 156840 101352
rect 156064 101312 156070 101324
rect 156834 101312 156840 101324
rect 156892 101312 156898 101364
rect 157110 101312 157116 101364
rect 157168 101352 157174 101364
rect 158306 101352 158312 101364
rect 157168 101324 158312 101352
rect 157168 101312 157174 101324
rect 158306 101312 158312 101324
rect 158364 101312 158370 101364
rect 160422 101312 160428 101364
rect 160480 101352 160486 101364
rect 161618 101352 161624 101364
rect 160480 101324 161624 101352
rect 160480 101312 160486 101324
rect 161618 101312 161624 101324
rect 161676 101312 161682 101364
rect 162630 101312 162636 101364
rect 162688 101352 162694 101364
rect 163826 101352 163832 101364
rect 162688 101324 163832 101352
rect 162688 101312 162694 101324
rect 163826 101312 163832 101324
rect 163884 101312 163890 101364
rect 164838 101312 164844 101364
rect 164896 101352 164902 101364
rect 166494 101352 166500 101364
rect 164896 101324 166500 101352
rect 164896 101312 164902 101324
rect 166494 101312 166500 101324
rect 166552 101312 166558 101364
rect 173762 101312 173768 101364
rect 173820 101352 173826 101364
rect 174774 101352 174780 101364
rect 173820 101324 174780 101352
rect 173820 101312 173826 101324
rect 174774 101312 174780 101324
rect 174832 101312 174838 101364
rect 175970 101312 175976 101364
rect 176028 101352 176034 101364
rect 176798 101352 176804 101364
rect 176028 101324 176804 101352
rect 176028 101312 176034 101324
rect 176798 101312 176804 101324
rect 176856 101312 176862 101364
rect 177074 101312 177080 101364
rect 177132 101352 177138 101364
rect 178178 101352 178184 101364
rect 177132 101324 178184 101352
rect 177132 101312 177138 101324
rect 178178 101312 178184 101324
rect 178236 101312 178242 101364
rect 194922 101312 194928 101364
rect 194980 101352 194986 101364
rect 195658 101352 195664 101364
rect 194980 101324 195664 101352
rect 194980 101312 194986 101324
rect 195658 101312 195664 101324
rect 195716 101312 195722 101364
rect 208078 101312 208084 101364
rect 208136 101352 208142 101364
rect 208354 101352 208360 101364
rect 208136 101324 208360 101352
rect 208136 101312 208142 101324
rect 208354 101312 208360 101324
rect 208412 101312 208418 101364
rect 212034 99884 212040 99936
rect 212092 99924 212098 99936
rect 222338 99924 222344 99936
rect 212092 99896 222344 99924
rect 212092 99884 212098 99896
rect 222338 99884 222344 99896
rect 222396 99884 222402 99936
rect 98782 97164 98788 97216
rect 98840 97204 98846 97216
rect 106786 97204 106792 97216
rect 98840 97176 106792 97204
rect 98840 97164 98846 97176
rect 106786 97164 106792 97176
rect 106844 97164 106850 97216
rect 13314 97096 13320 97148
rect 13372 97136 13378 97148
rect 22330 97136 22336 97148
rect 13372 97108 22336 97136
rect 13372 97096 13378 97108
rect 22330 97096 22336 97108
rect 22388 97096 22394 97148
rect 211758 97096 211764 97148
rect 211816 97136 211822 97148
rect 216174 97136 216180 97148
rect 211816 97108 216180 97136
rect 211816 97096 211822 97108
rect 216174 97096 216180 97108
rect 216232 97096 216238 97148
rect 99518 95804 99524 95856
rect 99576 95844 99582 95856
rect 106786 95844 106792 95856
rect 99576 95816 106792 95844
rect 99576 95804 99582 95816
rect 106786 95804 106792 95816
rect 106844 95804 106850 95856
rect 188574 94376 188580 94428
rect 188632 94416 188638 94428
rect 191978 94416 191984 94428
rect 188632 94388 191984 94416
rect 188632 94376 188638 94388
rect 191978 94376 191984 94388
rect 192036 94376 192042 94428
rect 98690 93016 98696 93068
rect 98748 93056 98754 93068
rect 106510 93056 106516 93068
rect 98748 93028 106516 93056
rect 98748 93016 98754 93028
rect 106510 93016 106516 93028
rect 106568 93016 106574 93068
rect 13314 90228 13320 90280
rect 13372 90268 13378 90280
rect 22330 90268 22336 90280
rect 13372 90240 22336 90268
rect 13372 90228 13378 90240
rect 22330 90228 22336 90240
rect 22388 90228 22394 90280
rect 105038 90228 105044 90280
rect 105096 90268 105102 90280
rect 106786 90268 106792 90280
rect 105096 90240 106792 90268
rect 105096 90228 105102 90240
rect 106786 90228 106792 90240
rect 106844 90228 106850 90280
rect 182870 90160 182876 90212
rect 182928 90200 182934 90212
rect 188574 90200 188580 90212
rect 182928 90172 188580 90200
rect 182928 90160 182934 90172
rect 188574 90160 188580 90172
rect 188632 90160 188638 90212
rect 211850 90160 211856 90212
rect 211908 90200 211914 90212
rect 221694 90200 221700 90212
rect 211908 90172 221700 90200
rect 211908 90160 211914 90172
rect 221694 90160 221700 90172
rect 221752 90160 221758 90212
rect 104946 88868 104952 88920
rect 105004 88908 105010 88920
rect 106786 88908 106792 88920
rect 105004 88880 106792 88908
rect 105004 88868 105010 88880
rect 106786 88868 106792 88880
rect 106844 88868 106850 88920
rect 128498 88868 128504 88920
rect 128556 88908 128562 88920
rect 131994 88908 132000 88920
rect 128556 88880 132000 88908
rect 128556 88868 128562 88880
rect 131994 88868 132000 88880
rect 132052 88868 132058 88920
rect 183514 88800 183520 88852
rect 183572 88840 183578 88852
rect 191150 88840 191156 88852
rect 183572 88812 191156 88840
rect 183572 88800 183578 88812
rect 191150 88800 191156 88812
rect 191208 88800 191214 88852
rect 183698 87440 183704 87492
rect 183756 87480 183762 87492
rect 190782 87480 190788 87492
rect 183756 87452 190788 87480
rect 183756 87440 183762 87452
rect 190782 87440 190788 87452
rect 190840 87440 190846 87492
rect 183698 86012 183704 86064
rect 183756 86052 183762 86064
rect 191702 86052 191708 86064
rect 183756 86024 191708 86052
rect 183756 86012 183762 86024
rect 191702 86012 191708 86024
rect 191760 86012 191766 86064
rect 99518 85196 99524 85248
rect 99576 85236 99582 85248
rect 105038 85236 105044 85248
rect 99576 85208 105044 85236
rect 99576 85196 99582 85208
rect 105038 85196 105044 85208
rect 105096 85196 105102 85248
rect 99426 84652 99432 84704
rect 99484 84692 99490 84704
rect 106786 84692 106792 84704
rect 99484 84664 106792 84692
rect 99484 84652 99490 84664
rect 106786 84652 106792 84664
rect 106844 84652 106850 84704
rect 182502 84652 182508 84704
rect 182560 84692 182566 84704
rect 191978 84692 191984 84704
rect 182560 84664 191984 84692
rect 182560 84652 182566 84664
rect 191978 84652 191984 84664
rect 192036 84652 192042 84704
rect 183698 84584 183704 84636
rect 183756 84624 183762 84636
rect 191610 84624 191616 84636
rect 183756 84596 191616 84624
rect 183756 84584 183762 84596
rect 191610 84584 191616 84596
rect 191668 84584 191674 84636
rect 99518 84448 99524 84500
rect 99576 84488 99582 84500
rect 104946 84488 104952 84500
rect 99576 84460 104952 84488
rect 99576 84448 99582 84460
rect 104946 84448 104952 84460
rect 105004 84448 105010 84500
rect 99518 83292 99524 83344
rect 99576 83332 99582 83344
rect 107798 83332 107804 83344
rect 99576 83304 107804 83332
rect 99576 83292 99582 83304
rect 107798 83292 107804 83304
rect 107856 83292 107862 83344
rect 183698 82612 183704 82664
rect 183756 82652 183762 82664
rect 191978 82652 191984 82664
rect 183756 82624 191984 82652
rect 183756 82612 183762 82624
rect 191978 82612 191984 82624
rect 192036 82612 192042 82664
rect 106786 82108 106792 82120
rect 103768 82080 106792 82108
rect 13314 82000 13320 82052
rect 13372 82040 13378 82052
rect 22330 82040 22336 82052
rect 13372 82012 22336 82040
rect 13372 82000 13378 82012
rect 22330 82000 22336 82012
rect 22388 82000 22394 82052
rect 99518 81932 99524 81984
rect 99576 81972 99582 81984
rect 103768 81972 103796 82080
rect 106786 82068 106792 82080
rect 106844 82068 106850 82120
rect 99576 81944 103796 81972
rect 99576 81932 99582 81944
rect 183238 81252 183244 81304
rect 183296 81292 183302 81304
rect 191886 81292 191892 81304
rect 183296 81264 191892 81292
rect 183296 81252 183302 81264
rect 191886 81252 191892 81264
rect 191944 81252 191950 81304
rect 131994 80504 132000 80556
rect 132052 80544 132058 80556
rect 136870 80544 136876 80556
rect 132052 80516 136876 80544
rect 132052 80504 132058 80516
rect 136870 80504 136876 80516
rect 136928 80504 136934 80556
rect 99518 79824 99524 79876
rect 99576 79864 99582 79876
rect 106786 79864 106792 79876
rect 99576 79836 106792 79864
rect 99576 79824 99582 79836
rect 106786 79824 106792 79836
rect 106844 79824 106850 79876
rect 183698 79212 183704 79264
rect 183756 79252 183762 79264
rect 183756 79224 187976 79252
rect 183756 79212 183762 79224
rect 187948 79184 187976 79224
rect 191978 79184 191984 79196
rect 187948 79156 191984 79184
rect 191978 79144 191984 79156
rect 192036 79144 192042 79196
rect 99518 77852 99524 77904
rect 99576 77892 99582 77904
rect 106510 77892 106516 77904
rect 99576 77864 106516 77892
rect 99576 77852 99582 77864
rect 106510 77852 106516 77864
rect 106568 77852 106574 77904
rect 183514 77852 183520 77904
rect 183572 77892 183578 77904
rect 191978 77892 191984 77904
rect 183572 77864 191984 77892
rect 183572 77852 183578 77864
rect 191978 77852 191984 77864
rect 192036 77852 192042 77904
rect 99518 76424 99524 76476
rect 99576 76464 99582 76476
rect 100990 76464 100996 76476
rect 99576 76436 100996 76464
rect 99576 76424 99582 76436
rect 100990 76424 100996 76436
rect 101048 76424 101054 76476
rect 183054 76424 183060 76476
rect 183112 76464 183118 76476
rect 185170 76464 185176 76476
rect 183112 76436 185176 76464
rect 183112 76424 183118 76436
rect 185170 76424 185176 76436
rect 185228 76424 185234 76476
rect 98230 75064 98236 75116
rect 98288 75104 98294 75116
rect 98288 75076 100944 75104
rect 98288 75064 98294 75076
rect 44410 74996 44416 75048
rect 44468 75036 44474 75048
rect 52598 75036 52604 75048
rect 44468 75008 52604 75036
rect 44468 74996 44474 75008
rect 52598 74996 52604 75008
rect 52656 74996 52662 75048
rect 100916 74900 100944 75076
rect 183238 75064 183244 75116
rect 183296 75104 183302 75116
rect 185998 75104 186004 75116
rect 183296 75076 186004 75104
rect 183296 75064 183302 75076
rect 185998 75064 186004 75076
rect 186056 75064 186062 75116
rect 100990 74996 100996 75048
rect 101048 75036 101054 75048
rect 106786 75036 106792 75048
rect 101048 75008 106792 75036
rect 101048 74996 101054 75008
rect 106786 74996 106792 75008
rect 106844 74996 106850 75048
rect 185170 74996 185176 75048
rect 185228 75036 185234 75048
rect 191518 75036 191524 75048
rect 185228 75008 191524 75036
rect 185228 74996 185234 75008
rect 191518 74996 191524 75008
rect 191576 74996 191582 75048
rect 100990 74900 100996 74912
rect 100916 74872 100996 74900
rect 100990 74860 100996 74872
rect 101048 74860 101054 74912
rect 52598 74656 52604 74708
rect 52656 74696 52662 74708
rect 53426 74696 53432 74708
rect 52656 74668 53432 74696
rect 52656 74656 52662 74668
rect 53426 74656 53432 74668
rect 53484 74656 53490 74708
rect 183698 73840 183704 73892
rect 183756 73880 183762 73892
rect 183756 73852 188620 73880
rect 183756 73840 183762 73852
rect 99518 73772 99524 73824
rect 99576 73812 99582 73824
rect 105130 73812 105136 73824
rect 99576 73784 105136 73812
rect 99576 73772 99582 73784
rect 105130 73772 105136 73784
rect 105188 73772 105194 73824
rect 99426 73704 99432 73756
rect 99484 73744 99490 73756
rect 106694 73744 106700 73756
rect 99484 73716 106700 73744
rect 99484 73704 99490 73716
rect 106694 73704 106700 73716
rect 106752 73704 106758 73756
rect 183698 73704 183704 73756
rect 183756 73744 183762 73756
rect 188482 73744 188488 73756
rect 183756 73716 188488 73744
rect 183756 73704 183762 73716
rect 188482 73704 188488 73716
rect 188540 73704 188546 73756
rect 188592 73744 188620 73852
rect 217554 73772 217560 73824
rect 217612 73812 217618 73824
rect 222338 73812 222344 73824
rect 217612 73784 222344 73812
rect 217612 73772 217618 73784
rect 222338 73772 222344 73784
rect 222396 73772 222402 73824
rect 190782 73744 190788 73756
rect 188592 73716 190788 73744
rect 190782 73704 190788 73716
rect 190840 73704 190846 73756
rect 100990 73636 100996 73688
rect 101048 73676 101054 73688
rect 106786 73676 106792 73688
rect 101048 73648 106792 73676
rect 101048 73636 101054 73648
rect 106786 73636 106792 73648
rect 106844 73636 106850 73688
rect 185998 73636 186004 73688
rect 186056 73676 186062 73688
rect 191978 73676 191984 73688
rect 186056 73648 191984 73676
rect 186056 73636 186062 73648
rect 191978 73636 191984 73648
rect 192036 73636 192042 73688
rect 99518 72344 99524 72396
rect 99576 72384 99582 72396
rect 106510 72384 106516 72396
rect 99576 72356 106516 72384
rect 99576 72344 99582 72356
rect 106510 72344 106516 72356
rect 106568 72344 106574 72396
rect 99518 70984 99524 71036
rect 99576 71024 99582 71036
rect 104486 71024 104492 71036
rect 99576 70996 104492 71024
rect 99576 70984 99582 70996
rect 104486 70984 104492 70996
rect 104544 70984 104550 71036
rect 183698 70916 183704 70968
rect 183756 70956 183762 70968
rect 191518 70956 191524 70968
rect 183756 70928 191524 70956
rect 183756 70916 183762 70928
rect 191518 70916 191524 70928
rect 191576 70916 191582 70968
rect 128498 70168 128504 70220
rect 128556 70208 128562 70220
rect 134018 70208 134024 70220
rect 128556 70180 134024 70208
rect 128556 70168 128562 70180
rect 134018 70168 134024 70180
rect 134076 70208 134082 70220
rect 136870 70208 136876 70220
rect 134076 70180 136876 70208
rect 134076 70168 134082 70180
rect 136870 70168 136876 70180
rect 136928 70168 136934 70220
rect 182870 69896 182876 69948
rect 182928 69936 182934 69948
rect 189954 69936 189960 69948
rect 182928 69908 189960 69936
rect 182928 69896 182934 69908
rect 189954 69896 189960 69908
rect 190012 69896 190018 69948
rect 99518 69556 99524 69608
rect 99576 69596 99582 69608
rect 104394 69596 104400 69608
rect 99576 69568 104400 69596
rect 99576 69556 99582 69568
rect 104394 69556 104400 69568
rect 104452 69556 104458 69608
rect 188482 69488 188488 69540
rect 188540 69528 188546 69540
rect 190966 69528 190972 69540
rect 188540 69500 190972 69528
rect 188540 69488 188546 69500
rect 190966 69488 190972 69500
rect 191024 69488 191030 69540
rect 105130 68128 105136 68180
rect 105188 68168 105194 68180
rect 106602 68168 106608 68180
rect 105188 68140 106608 68168
rect 105188 68128 105194 68140
rect 106602 68128 106608 68140
rect 106660 68128 106666 68180
rect 183790 68128 183796 68180
rect 183848 68168 183854 68180
rect 191334 68168 191340 68180
rect 183848 68140 191340 68168
rect 183848 68128 183854 68140
rect 191334 68128 191340 68140
rect 191392 68128 191398 68180
rect 104486 63640 104492 63692
rect 104544 63680 104550 63692
rect 106602 63680 106608 63692
rect 104544 63652 106608 63680
rect 104544 63640 104550 63652
rect 106602 63640 106608 63652
rect 106660 63640 106666 63692
rect 18098 63572 18104 63624
rect 18156 63612 18162 63624
rect 22330 63612 22336 63624
rect 18156 63584 22336 63612
rect 18156 63572 18162 63584
rect 22330 63572 22336 63584
rect 22388 63572 22394 63624
rect 212678 63164 212684 63216
rect 212736 63204 212742 63216
rect 217554 63204 217560 63216
rect 212736 63176 217560 63204
rect 212736 63164 212742 63176
rect 217554 63164 217560 63176
rect 217612 63164 217618 63216
rect 183698 61464 183704 61516
rect 183756 61504 183762 61516
rect 188022 61504 188028 61516
rect 183756 61476 188028 61504
rect 183756 61464 183762 61476
rect 188022 61464 188028 61476
rect 188080 61464 188086 61516
rect 99518 61260 99524 61312
rect 99576 61300 99582 61312
rect 103014 61300 103020 61312
rect 99576 61272 103020 61300
rect 99576 61260 99582 61272
rect 103014 61260 103020 61272
rect 103072 61260 103078 61312
rect 104394 61192 104400 61244
rect 104452 61232 104458 61244
rect 107154 61232 107160 61244
rect 104452 61204 107160 61232
rect 104452 61192 104458 61204
rect 107154 61192 107160 61204
rect 107212 61192 107218 61244
rect 182686 60376 182692 60428
rect 182744 60416 182750 60428
rect 184434 60416 184440 60428
rect 182744 60388 184440 60416
rect 182744 60376 182750 60388
rect 184434 60376 184440 60388
rect 184492 60376 184498 60428
rect 99518 59900 99524 59952
rect 99576 59940 99582 59952
rect 100346 59940 100352 59952
rect 99576 59912 100352 59940
rect 99576 59900 99582 59912
rect 100346 59900 100352 59912
rect 100404 59900 100410 59952
rect 36130 58472 36136 58524
rect 36188 58512 36194 58524
rect 37510 58512 37516 58524
rect 36188 58484 37516 58512
rect 36188 58472 36194 58484
rect 37510 58472 37516 58484
rect 37568 58472 37574 58524
rect 84341 58515 84399 58521
rect 84341 58481 84353 58515
rect 84387 58512 84399 58515
rect 84433 58515 84491 58521
rect 84433 58512 84445 58515
rect 84387 58484 84445 58512
rect 84387 58481 84399 58484
rect 84341 58475 84399 58481
rect 84433 58481 84445 58484
rect 84479 58481 84491 58515
rect 84433 58475 84491 58481
rect 96853 58515 96911 58521
rect 96853 58481 96865 58515
rect 96899 58512 96911 58515
rect 98874 58512 98880 58524
rect 96899 58484 98880 58512
rect 96899 58481 96911 58484
rect 96853 58475 96911 58481
rect 98874 58472 98880 58484
rect 98932 58512 98938 58524
rect 163182 58512 163188 58524
rect 98932 58484 163188 58512
rect 98932 58472 98938 58484
rect 163182 58472 163188 58484
rect 163240 58472 163246 58524
rect 208078 58472 208084 58524
rect 208136 58512 208142 58524
rect 210654 58512 210660 58524
rect 208136 58484 210660 58512
rect 208136 58472 208142 58484
rect 210654 58472 210660 58484
rect 210712 58472 210718 58524
rect 99521 58447 99579 58453
rect 99521 58413 99533 58447
rect 99567 58444 99579 58447
rect 128593 58447 128651 58453
rect 128593 58444 128605 58447
rect 99567 58416 109132 58444
rect 99567 58413 99579 58416
rect 99521 58407 99579 58413
rect 72562 58336 72568 58388
rect 72620 58376 72626 58388
rect 72620 58348 77944 58376
rect 72620 58336 72626 58348
rect 77916 58308 77944 58348
rect 79186 58336 79192 58388
rect 79244 58376 79250 58388
rect 88481 58379 88539 58385
rect 88481 58376 88493 58379
rect 79244 58348 88493 58376
rect 79244 58336 79250 58348
rect 88481 58345 88493 58348
rect 88527 58345 88539 58379
rect 88481 58339 88539 58345
rect 84341 58311 84399 58317
rect 84341 58308 84353 58311
rect 77916 58280 84353 58308
rect 84341 58277 84353 58280
rect 84387 58277 84399 58311
rect 84341 58271 84399 58277
rect 84433 58311 84491 58317
rect 84433 58277 84445 58311
rect 84479 58308 84491 58311
rect 95378 58308 95384 58320
rect 84479 58280 95384 58308
rect 84479 58277 84491 58280
rect 84433 58271 84491 58277
rect 95378 58268 95384 58280
rect 95436 58308 95442 58320
rect 99521 58311 99579 58317
rect 99521 58308 99533 58311
rect 95436 58280 99533 58308
rect 95436 58268 95442 58280
rect 99521 58277 99533 58280
rect 99567 58277 99579 58311
rect 109104 58308 109132 58416
rect 120328 58416 128605 58444
rect 109641 58311 109699 58317
rect 109641 58308 109653 58311
rect 109104 58280 109653 58308
rect 99521 58271 99579 58277
rect 109641 58277 109653 58280
rect 109687 58277 109699 58311
rect 109641 58271 109699 58277
rect 109733 58311 109791 58317
rect 109733 58277 109745 58311
rect 109779 58308 109791 58311
rect 120328 58308 120356 58416
rect 128593 58413 128605 58416
rect 128639 58413 128651 58447
rect 128593 58407 128651 58413
rect 209642 58404 209648 58456
rect 209700 58444 209706 58456
rect 212034 58444 212040 58456
rect 209700 58416 212040 58444
rect 209700 58404 209706 58416
rect 212034 58404 212040 58416
rect 212092 58404 212098 58456
rect 145061 58379 145119 58385
rect 145061 58345 145073 58379
rect 145107 58376 145119 58379
rect 147821 58379 147879 58385
rect 147821 58376 147833 58379
rect 145107 58348 147833 58376
rect 145107 58345 145119 58348
rect 145061 58339 145119 58345
rect 147821 58345 147833 58348
rect 147867 58345 147879 58379
rect 147821 58339 147879 58345
rect 147913 58379 147971 58385
rect 147913 58345 147925 58379
rect 147959 58376 147971 58379
rect 147959 58348 149152 58376
rect 147959 58345 147971 58348
rect 147913 58339 147971 58345
rect 109779 58280 120356 58308
rect 109779 58277 109791 58280
rect 109733 58271 109791 58277
rect 122058 58268 122064 58320
rect 122116 58308 122122 58320
rect 124542 58308 124548 58320
rect 122116 58280 124548 58308
rect 122116 58268 122122 58280
rect 124542 58268 124548 58280
rect 124600 58268 124606 58320
rect 128593 58311 128651 58317
rect 128593 58277 128605 58311
rect 128639 58308 128651 58311
rect 135493 58311 135551 58317
rect 135493 58308 135505 58311
rect 128639 58280 135505 58308
rect 128639 58277 128651 58280
rect 128593 58271 128651 58277
rect 135493 58277 135505 58280
rect 135539 58277 135551 58311
rect 149124 58308 149152 58348
rect 209274 58336 209280 58388
rect 209332 58376 209338 58388
rect 212126 58376 212132 58388
rect 209332 58348 212132 58376
rect 209332 58336 209338 58348
rect 212126 58336 212132 58348
rect 212184 58336 212190 58388
rect 156558 58308 156564 58320
rect 149124 58280 156564 58308
rect 135493 58271 135551 58277
rect 156558 58268 156564 58280
rect 156616 58268 156622 58320
rect 207618 58268 207624 58320
rect 207676 58308 207682 58320
rect 210746 58308 210752 58320
rect 207676 58280 210752 58308
rect 207676 58268 207682 58280
rect 210746 58268 210752 58280
rect 210804 58268 210810 58320
rect 41650 58200 41656 58252
rect 41708 58240 41714 58252
rect 46434 58240 46440 58252
rect 41708 58212 46440 58240
rect 41708 58200 41714 58212
rect 46434 58200 46440 58212
rect 46492 58200 46498 58252
rect 206882 58200 206888 58252
rect 206940 58240 206946 58252
rect 210010 58240 210016 58252
rect 206940 58212 210016 58240
rect 206940 58200 206946 58212
rect 210010 58200 210016 58212
rect 210068 58200 210074 58252
rect 119298 58132 119304 58184
rect 119356 58172 119362 58184
rect 121138 58172 121144 58184
rect 119356 58144 121144 58172
rect 119356 58132 119362 58144
rect 121138 58132 121144 58144
rect 121196 58132 121202 58184
rect 135493 58175 135551 58181
rect 135493 58141 135505 58175
rect 135539 58172 135551 58175
rect 145061 58175 145119 58181
rect 145061 58172 145073 58175
rect 135539 58144 145073 58172
rect 135539 58141 135551 58144
rect 135493 58135 135551 58141
rect 145061 58141 145073 58144
rect 145107 58141 145119 58175
rect 145061 58135 145119 58141
rect 207250 58132 207256 58184
rect 207308 58172 207314 58184
rect 210838 58172 210844 58184
rect 207308 58144 210844 58172
rect 207308 58132 207314 58144
rect 210838 58132 210844 58144
rect 210896 58132 210902 58184
rect 88481 58107 88539 58113
rect 88481 58073 88493 58107
rect 88527 58104 88539 58107
rect 96853 58107 96911 58113
rect 96853 58104 96865 58107
rect 88527 58076 96865 58104
rect 88527 58073 88539 58076
rect 88481 58067 88539 58073
rect 96853 58073 96865 58076
rect 96899 58073 96911 58107
rect 96853 58067 96911 58073
rect 116446 58064 116452 58116
rect 116504 58104 116510 58116
rect 117642 58104 117648 58116
rect 116504 58076 117648 58104
rect 116504 58064 116510 58076
rect 117642 58064 117648 58076
rect 117700 58064 117706 58116
rect 208814 58064 208820 58116
rect 208872 58104 208878 58116
rect 212218 58104 212224 58116
rect 208872 58076 212224 58104
rect 208872 58064 208878 58076
rect 212218 58064 212224 58076
rect 212276 58064 212282 58116
rect 122426 57996 122432 58048
rect 122484 58036 122490 58048
rect 125186 58036 125192 58048
rect 122484 58008 125192 58036
rect 122484 57996 122490 58008
rect 125186 57996 125192 58008
rect 125244 57996 125250 58048
rect 206422 57996 206428 58048
rect 206480 58036 206486 58048
rect 210102 58036 210108 58048
rect 206480 58008 210108 58036
rect 206480 57996 206486 58008
rect 210102 57996 210108 58008
rect 210160 57996 210166 58048
rect 70538 57928 70544 57980
rect 70596 57968 70602 57980
rect 92526 57968 92532 57980
rect 70596 57940 92532 57968
rect 70596 57928 70602 57940
rect 92526 57928 92532 57940
rect 92584 57928 92590 57980
rect 124450 57928 124456 57980
rect 124508 57968 124514 57980
rect 128590 57968 128596 57980
rect 124508 57940 128596 57968
rect 124508 57928 124514 57940
rect 128590 57928 128596 57940
rect 128648 57928 128654 57980
rect 13314 57860 13320 57912
rect 13372 57900 13378 57912
rect 72562 57900 72568 57912
rect 13372 57872 72568 57900
rect 13372 57860 13378 57872
rect 72562 57860 72568 57872
rect 72620 57860 72626 57912
rect 201546 57860 201552 57912
rect 201604 57900 201610 57912
rect 202742 57900 202748 57912
rect 201604 57872 202748 57900
rect 201604 57860 201610 57872
rect 202742 57860 202748 57872
rect 202800 57860 202806 57912
rect 13406 57792 13412 57844
rect 13464 57832 13470 57844
rect 79186 57832 79192 57844
rect 13464 57804 79192 57832
rect 13464 57792 13470 57804
rect 79186 57792 79192 57804
rect 79244 57792 79250 57844
rect 123622 57792 123628 57844
rect 123680 57832 123686 57844
rect 127210 57832 127216 57844
rect 123680 57804 127216 57832
rect 123680 57792 123686 57804
rect 127210 57792 127216 57804
rect 127268 57792 127274 57844
rect 156098 57792 156104 57844
rect 156156 57832 156162 57844
rect 169898 57832 169904 57844
rect 156156 57804 169904 57832
rect 156156 57792 156162 57804
rect 169898 57792 169904 57804
rect 169956 57792 169962 57844
rect 208446 57792 208452 57844
rect 208504 57832 208510 57844
rect 212862 57832 212868 57844
rect 208504 57804 212868 57832
rect 208504 57792 208510 57804
rect 212862 57792 212868 57804
rect 212920 57792 212926 57844
rect 120494 57656 120500 57708
rect 120552 57696 120558 57708
rect 123162 57696 123168 57708
rect 120552 57668 123168 57696
rect 120552 57656 120558 57668
rect 123162 57656 123168 57668
rect 123220 57656 123226 57708
rect 39258 57588 39264 57640
rect 39316 57628 39322 57640
rect 43030 57628 43036 57640
rect 39316 57600 43036 57628
rect 39316 57588 39322 57600
rect 43030 57588 43036 57600
rect 43088 57588 43094 57640
rect 117274 57588 117280 57640
rect 117332 57628 117338 57640
rect 118286 57628 118292 57640
rect 117332 57600 118292 57628
rect 117332 57588 117338 57600
rect 118286 57588 118292 57600
rect 118344 57588 118350 57640
rect 200810 57588 200816 57640
rect 200868 57628 200874 57640
rect 202190 57628 202196 57640
rect 200868 57600 202196 57628
rect 200868 57588 200874 57600
rect 202190 57588 202196 57600
rect 202248 57588 202254 57640
rect 40086 57520 40092 57572
rect 40144 57560 40150 57572
rect 43674 57560 43680 57572
rect 40144 57532 43680 57560
rect 40144 57520 40150 57532
rect 43674 57520 43680 57532
rect 43732 57520 43738 57572
rect 199614 57520 199620 57572
rect 199672 57560 199678 57572
rect 200442 57560 200448 57572
rect 199672 57532 200448 57560
rect 199672 57520 199678 57532
rect 200442 57520 200448 57532
rect 200500 57520 200506 57572
rect 205226 57520 205232 57572
rect 205284 57560 205290 57572
rect 207986 57560 207992 57572
rect 205284 57532 207992 57560
rect 205284 57520 205290 57532
rect 207986 57520 207992 57532
rect 208044 57520 208050 57572
rect 39626 57452 39632 57504
rect 39684 57492 39690 57504
rect 43122 57492 43128 57504
rect 39684 57464 43128 57492
rect 39684 57452 39690 57464
rect 43122 57452 43128 57464
rect 43180 57452 43186 57504
rect 123254 57452 123260 57504
rect 123312 57492 123318 57504
rect 126106 57492 126112 57504
rect 123312 57464 126112 57492
rect 123312 57452 123318 57464
rect 126106 57452 126112 57464
rect 126164 57452 126170 57504
rect 204490 57452 204496 57504
rect 204548 57492 204554 57504
rect 207342 57492 207348 57504
rect 204548 57464 207348 57492
rect 204548 57452 204554 57464
rect 207342 57452 207348 57464
rect 207400 57452 207406 57504
rect 38890 57384 38896 57436
rect 38948 57424 38954 57436
rect 41834 57424 41840 57436
rect 38948 57396 41840 57424
rect 38948 57384 38954 57396
rect 41834 57384 41840 57396
rect 41892 57384 41898 57436
rect 109086 57384 109092 57436
rect 109144 57424 109150 57436
rect 110466 57424 110472 57436
rect 109144 57396 110472 57424
rect 109144 57384 109150 57396
rect 110466 57384 110472 57396
rect 110524 57384 110530 57436
rect 203662 57384 203668 57436
rect 203720 57424 203726 57436
rect 205226 57424 205232 57436
rect 203720 57396 205232 57424
rect 203720 57384 203726 57396
rect 205226 57384 205232 57396
rect 205284 57384 205290 57436
rect 29138 57316 29144 57368
rect 29196 57356 29202 57368
rect 30426 57356 30432 57368
rect 29196 57328 30432 57356
rect 29196 57316 29202 57328
rect 30426 57316 30432 57328
rect 30484 57316 30490 57368
rect 37694 57316 37700 57368
rect 37752 57356 37758 57368
rect 40270 57356 40276 57368
rect 37752 57328 40276 57356
rect 37752 57316 37758 57328
rect 40270 57316 40276 57328
rect 40328 57316 40334 57368
rect 40822 57316 40828 57368
rect 40880 57356 40886 57368
rect 45146 57356 45152 57368
rect 40880 57328 45152 57356
rect 40880 57316 40886 57328
rect 45146 57316 45152 57328
rect 45204 57316 45210 57368
rect 118470 57316 118476 57368
rect 118528 57356 118534 57368
rect 120494 57356 120500 57368
rect 118528 57328 120500 57356
rect 118528 57316 118534 57328
rect 120494 57316 120500 57328
rect 120552 57316 120558 57368
rect 120862 57316 120868 57368
rect 120920 57356 120926 57368
rect 123346 57356 123352 57368
rect 120920 57328 123352 57356
rect 120920 57316 120926 57328
rect 123346 57316 123352 57328
rect 123404 57316 123410 57368
rect 124082 57316 124088 57368
rect 124140 57356 124146 57368
rect 127302 57356 127308 57368
rect 124140 57328 127308 57356
rect 124140 57316 124146 57328
rect 127302 57316 127308 57328
rect 127360 57316 127366 57368
rect 204030 57316 204036 57368
rect 204088 57356 204094 57368
rect 205318 57356 205324 57368
rect 204088 57328 205324 57356
rect 204088 57316 204094 57328
rect 205318 57316 205324 57328
rect 205376 57316 205382 57368
rect 36866 57248 36872 57300
rect 36924 57288 36930 57300
rect 38154 57288 38160 57300
rect 36924 57260 38160 57288
rect 36924 57248 36930 57260
rect 38154 57248 38160 57260
rect 38212 57248 38218 57300
rect 40454 57248 40460 57300
rect 40512 57288 40518 57300
rect 44594 57288 44600 57300
rect 40512 57260 44600 57288
rect 40512 57248 40518 57260
rect 44594 57248 44600 57260
rect 44652 57248 44658 57300
rect 118838 57248 118844 57300
rect 118896 57288 118902 57300
rect 120770 57288 120776 57300
rect 118896 57260 120776 57288
rect 118896 57248 118902 57260
rect 120770 57248 120776 57260
rect 120828 57248 120834 57300
rect 121690 57248 121696 57300
rect 121748 57288 121754 57300
rect 124450 57288 124456 57300
rect 121748 57260 124456 57288
rect 121748 57248 121754 57260
rect 124450 57248 124456 57260
rect 124508 57248 124514 57300
rect 124818 57248 124824 57300
rect 124876 57288 124882 57300
rect 128866 57288 128872 57300
rect 124876 57260 128872 57288
rect 124876 57248 124882 57260
rect 128866 57248 128872 57260
rect 128924 57248 128930 57300
rect 194922 57248 194928 57300
rect 194980 57288 194986 57300
rect 195658 57288 195664 57300
rect 194980 57260 195664 57288
rect 194980 57248 194986 57260
rect 195658 57248 195664 57260
rect 195716 57248 195722 57300
rect 199062 57248 199068 57300
rect 199120 57288 199126 57300
rect 199798 57288 199804 57300
rect 199120 57260 199804 57288
rect 199120 57248 199126 57260
rect 199798 57248 199804 57260
rect 199856 57248 199862 57300
rect 202466 57248 202472 57300
rect 202524 57288 202530 57300
rect 204490 57288 204496 57300
rect 202524 57260 204496 57288
rect 202524 57248 202530 57260
rect 204490 57248 204496 57260
rect 204548 57248 204554 57300
rect 204858 57248 204864 57300
rect 204916 57288 204922 57300
rect 207250 57288 207256 57300
rect 204916 57260 207256 57288
rect 204916 57248 204922 57260
rect 207250 57248 207256 57260
rect 207308 57248 207314 57300
rect 30426 57180 30432 57232
rect 30484 57220 30490 57232
rect 31254 57220 31260 57232
rect 30484 57192 31260 57220
rect 30484 57180 30490 57192
rect 31254 57180 31260 57192
rect 31312 57180 31318 57232
rect 32450 57220 32456 57232
rect 31916 57192 32456 57220
rect 26470 57112 26476 57164
rect 26528 57152 26534 57164
rect 27390 57152 27396 57164
rect 26528 57124 27396 57152
rect 26528 57112 26534 57124
rect 27390 57112 27396 57124
rect 27448 57112 27454 57164
rect 29414 57112 29420 57164
rect 29472 57152 29478 57164
rect 29782 57152 29788 57164
rect 29472 57124 29788 57152
rect 29472 57112 29478 57124
rect 29782 57112 29788 57124
rect 29840 57112 29846 57164
rect 30518 57112 30524 57164
rect 30576 57152 30582 57164
rect 31622 57152 31628 57164
rect 30576 57124 31628 57152
rect 30576 57112 30582 57124
rect 31622 57112 31628 57124
rect 31680 57112 31686 57164
rect 31916 57096 31944 57192
rect 32450 57180 32456 57192
rect 32508 57180 32514 57232
rect 37234 57180 37240 57232
rect 37292 57220 37298 57232
rect 38246 57220 38252 57232
rect 37292 57192 38252 57220
rect 37292 57180 37298 57192
rect 38246 57180 38252 57192
rect 38304 57180 38310 57232
rect 38430 57180 38436 57232
rect 38488 57220 38494 57232
rect 40914 57220 40920 57232
rect 38488 57192 40920 57220
rect 38488 57180 38494 57192
rect 40914 57180 40920 57192
rect 40972 57180 40978 57232
rect 112858 57220 112864 57232
rect 112600 57192 112864 57220
rect 112600 57164 112628 57192
rect 112858 57180 112864 57192
rect 112916 57180 112922 57232
rect 116078 57180 116084 57232
rect 116136 57220 116142 57232
rect 116630 57220 116636 57232
rect 116136 57192 116636 57220
rect 116136 57180 116142 57192
rect 116630 57180 116636 57192
rect 116688 57180 116694 57232
rect 118010 57180 118016 57232
rect 118068 57220 118074 57232
rect 118068 57192 118884 57220
rect 118068 57180 118074 57192
rect 118856 57164 118884 57192
rect 119666 57180 119672 57232
rect 119724 57220 119730 57232
rect 120954 57220 120960 57232
rect 119724 57192 120960 57220
rect 119724 57180 119730 57192
rect 120954 57180 120960 57192
rect 121012 57180 121018 57232
rect 122886 57180 122892 57232
rect 122944 57220 122950 57232
rect 125094 57220 125100 57232
rect 122944 57192 125100 57220
rect 122944 57180 122950 57192
rect 125094 57180 125100 57192
rect 125152 57180 125158 57232
rect 125646 57180 125652 57232
rect 125704 57220 125710 57232
rect 130062 57220 130068 57232
rect 125704 57192 130068 57220
rect 125704 57180 125710 57192
rect 130062 57180 130068 57192
rect 130120 57180 130126 57232
rect 193266 57180 193272 57232
rect 193324 57220 193330 57232
rect 194462 57220 194468 57232
rect 193324 57192 194468 57220
rect 193324 57180 193330 57192
rect 194462 57180 194468 57192
rect 194520 57180 194526 57232
rect 200718 57180 200724 57232
rect 200776 57220 200782 57232
rect 201822 57220 201828 57232
rect 200776 57192 201828 57220
rect 200776 57180 200782 57192
rect 201822 57180 201828 57192
rect 201880 57180 201886 57232
rect 202098 57180 202104 57232
rect 202156 57220 202162 57232
rect 203018 57220 203024 57232
rect 202156 57192 203024 57220
rect 202156 57180 202162 57192
rect 203018 57180 203024 57192
rect 203076 57180 203082 57232
rect 203294 57180 203300 57232
rect 203352 57220 203358 57232
rect 205134 57220 205140 57232
rect 203352 57192 205140 57220
rect 203352 57180 203358 57192
rect 205134 57180 205140 57192
rect 205192 57180 205198 57232
rect 205686 57180 205692 57232
rect 205744 57220 205750 57232
rect 207894 57220 207900 57232
rect 205744 57192 207900 57220
rect 205744 57180 205750 57192
rect 207894 57180 207900 57192
rect 207952 57180 207958 57232
rect 32082 57112 32088 57164
rect 32140 57152 32146 57164
rect 32818 57152 32824 57164
rect 32140 57124 32824 57152
rect 32140 57112 32146 57124
rect 32818 57112 32824 57124
rect 32876 57112 32882 57164
rect 33278 57152 33284 57164
rect 32928 57124 33284 57152
rect 31898 57044 31904 57096
rect 31956 57044 31962 57096
rect 31990 57044 31996 57096
rect 32048 57084 32054 57096
rect 32928 57084 32956 57124
rect 33278 57112 33284 57124
rect 33336 57112 33342 57164
rect 33370 57112 33376 57164
rect 33428 57152 33434 57164
rect 34106 57152 34112 57164
rect 33428 57124 34112 57152
rect 33428 57112 33434 57124
rect 34106 57112 34112 57124
rect 34164 57112 34170 57164
rect 35302 57112 35308 57164
rect 35360 57152 35366 57164
rect 36038 57152 36044 57164
rect 35360 57124 36044 57152
rect 35360 57112 35366 57124
rect 36038 57112 36044 57124
rect 36096 57112 36102 57164
rect 36498 57112 36504 57164
rect 36556 57152 36562 57164
rect 37602 57152 37608 57164
rect 36556 57124 37608 57152
rect 36556 57112 36562 57124
rect 37602 57112 37608 57124
rect 37660 57112 37666 57164
rect 38062 57112 38068 57164
rect 38120 57152 38126 57164
rect 40362 57152 40368 57164
rect 38120 57124 40368 57152
rect 38120 57112 38126 57124
rect 40362 57112 40368 57124
rect 40420 57112 40426 57164
rect 41282 57112 41288 57164
rect 41340 57152 41346 57164
rect 45054 57152 45060 57164
rect 41340 57124 45060 57152
rect 41340 57112 41346 57124
rect 45054 57112 45060 57124
rect 45112 57112 45118 57164
rect 109178 57112 109184 57164
rect 109236 57152 109242 57164
rect 110098 57152 110104 57164
rect 109236 57124 110104 57152
rect 109236 57112 109242 57124
rect 110098 57112 110104 57124
rect 110156 57112 110162 57164
rect 111662 57152 111668 57164
rect 110668 57124 111668 57152
rect 110668 57096 110696 57124
rect 111662 57112 111668 57124
rect 111720 57112 111726 57164
rect 112582 57112 112588 57164
rect 112640 57112 112646 57164
rect 112766 57112 112772 57164
rect 112824 57152 112830 57164
rect 113226 57152 113232 57164
rect 112824 57124 113232 57152
rect 112824 57112 112830 57124
rect 113226 57112 113232 57124
rect 113284 57112 113290 57164
rect 113502 57112 113508 57164
rect 113560 57152 113566 57164
rect 114054 57152 114060 57164
rect 113560 57124 114060 57152
rect 113560 57112 113566 57124
rect 114054 57112 114060 57124
rect 114112 57112 114118 57164
rect 114422 57112 114428 57164
rect 114480 57152 114486 57164
rect 114974 57152 114980 57164
rect 114480 57124 114980 57152
rect 114480 57112 114486 57124
rect 114974 57112 114980 57124
rect 115032 57112 115038 57164
rect 115618 57112 115624 57164
rect 115676 57152 115682 57164
rect 116262 57152 116268 57164
rect 115676 57124 116268 57152
rect 115676 57112 115682 57124
rect 116262 57112 116268 57124
rect 116320 57112 116326 57164
rect 116814 57112 116820 57164
rect 116872 57152 116878 57164
rect 117734 57152 117740 57164
rect 116872 57124 117740 57152
rect 116872 57112 116878 57124
rect 117734 57112 117740 57124
rect 117792 57112 117798 57164
rect 118102 57112 118108 57164
rect 118160 57152 118166 57164
rect 118654 57152 118660 57164
rect 118160 57124 118660 57152
rect 118160 57112 118166 57124
rect 118654 57112 118660 57124
rect 118712 57112 118718 57164
rect 118838 57112 118844 57164
rect 118896 57112 118902 57164
rect 120034 57112 120040 57164
rect 120092 57152 120098 57164
rect 121046 57152 121052 57164
rect 120092 57124 121052 57152
rect 120092 57112 120098 57124
rect 121046 57112 121052 57124
rect 121104 57112 121110 57164
rect 121230 57112 121236 57164
rect 121288 57152 121294 57164
rect 123990 57152 123996 57164
rect 121288 57124 123996 57152
rect 121288 57112 121294 57124
rect 123990 57112 123996 57124
rect 124048 57112 124054 57164
rect 125278 57112 125284 57164
rect 125336 57152 125342 57164
rect 128958 57152 128964 57164
rect 125336 57124 128964 57152
rect 125336 57112 125342 57124
rect 128958 57112 128964 57124
rect 129016 57112 129022 57164
rect 193358 57112 193364 57164
rect 193416 57152 193422 57164
rect 194094 57152 194100 57164
rect 193416 57124 194100 57152
rect 193416 57112 193422 57124
rect 194094 57112 194100 57124
rect 194152 57112 194158 57164
rect 194738 57112 194744 57164
rect 194796 57152 194802 57164
rect 195014 57152 195020 57164
rect 194796 57124 195020 57152
rect 194796 57112 194802 57124
rect 195014 57112 195020 57124
rect 195072 57112 195078 57164
rect 195106 57112 195112 57164
rect 195164 57152 195170 57164
rect 196026 57152 196032 57164
rect 195164 57124 196032 57152
rect 195164 57112 195170 57124
rect 196026 57112 196032 57124
rect 196084 57112 196090 57164
rect 196302 57112 196308 57164
rect 196360 57152 196366 57164
rect 196854 57152 196860 57164
rect 196360 57124 196860 57152
rect 196360 57112 196366 57124
rect 196854 57112 196860 57124
rect 196912 57112 196918 57164
rect 198786 57112 198792 57164
rect 198844 57152 198850 57164
rect 198844 57124 199108 57152
rect 198844 57112 198850 57124
rect 32048 57056 32956 57084
rect 32048 57044 32054 57056
rect 110650 57044 110656 57096
rect 110708 57044 110714 57096
rect 198050 57084 198056 57096
rect 198011 57056 198056 57084
rect 198050 57044 198056 57056
rect 198108 57044 198114 57096
rect 199080 57028 199108 57124
rect 200166 57112 200172 57164
rect 200224 57152 200230 57164
rect 200902 57152 200908 57164
rect 200224 57124 200908 57152
rect 200224 57112 200230 57124
rect 200902 57112 200908 57124
rect 200960 57112 200966 57164
rect 201638 57112 201644 57164
rect 201696 57152 201702 57164
rect 202374 57152 202380 57164
rect 201696 57124 202380 57152
rect 201696 57112 201702 57124
rect 202374 57112 202380 57124
rect 202432 57112 202438 57164
rect 202834 57112 202840 57164
rect 202892 57152 202898 57164
rect 204582 57152 204588 57164
rect 202892 57124 204588 57152
rect 202892 57112 202898 57124
rect 204582 57112 204588 57124
rect 204640 57112 204646 57164
rect 206054 57112 206060 57164
rect 206112 57152 206118 57164
rect 207158 57152 207164 57164
rect 206112 57124 207164 57152
rect 206112 57112 206118 57124
rect 207158 57112 207164 57124
rect 207216 57112 207222 57164
rect 199062 56976 199068 57028
rect 199120 56976 199126 57028
rect 98782 55004 98788 55056
rect 98840 55044 98846 55056
rect 99518 55044 99524 55056
rect 98840 55016 99524 55044
rect 98840 55004 98846 55016
rect 99518 55004 99524 55016
rect 99576 55004 99582 55056
rect 26654 54392 26660 54444
rect 26712 54432 26718 54444
rect 26838 54432 26844 54444
rect 26712 54404 26844 54432
rect 26712 54392 26718 54404
rect 26838 54392 26844 54404
rect 26896 54392 26902 54444
rect 210654 50516 210660 50568
rect 210712 50556 210718 50568
rect 210930 50556 210936 50568
rect 210712 50528 210936 50556
rect 210712 50516 210718 50528
rect 210930 50516 210936 50528
rect 210988 50516 210994 50568
rect 210010 50380 210016 50432
rect 210068 50420 210074 50432
rect 210654 50420 210660 50432
rect 210068 50392 210660 50420
rect 210068 50380 210074 50392
rect 210654 50380 210660 50392
rect 210712 50380 210718 50432
rect 114882 50312 114888 50364
rect 114940 50352 114946 50364
rect 114940 50324 115112 50352
rect 114940 50312 114946 50324
rect 31990 50244 31996 50296
rect 32048 50284 32054 50296
rect 32726 50284 32732 50296
rect 32048 50256 32732 50284
rect 32048 50244 32054 50256
rect 32726 50244 32732 50256
rect 32784 50244 32790 50296
rect 33370 50244 33376 50296
rect 33428 50284 33434 50296
rect 34198 50284 34204 50296
rect 33428 50256 34204 50284
rect 33428 50244 33434 50256
rect 34198 50244 34204 50256
rect 34256 50244 34262 50296
rect 41834 50244 41840 50296
rect 41892 50284 41898 50296
rect 42294 50284 42300 50296
rect 41892 50256 42300 50284
rect 41892 50244 41898 50256
rect 42294 50244 42300 50256
rect 42352 50244 42358 50296
rect 114974 50244 114980 50296
rect 115032 50244 115038 50296
rect 22882 50176 22888 50228
rect 22940 50216 22946 50228
rect 26746 50216 26752 50228
rect 22940 50188 26752 50216
rect 22940 50176 22946 50188
rect 26746 50176 26752 50188
rect 26804 50176 26810 50228
rect 28310 50176 28316 50228
rect 28368 50216 28374 50228
rect 29138 50216 29144 50228
rect 28368 50188 29144 50216
rect 28368 50176 28374 50188
rect 29138 50176 29144 50188
rect 29196 50176 29202 50228
rect 29690 50176 29696 50228
rect 29748 50216 29754 50228
rect 30426 50216 30432 50228
rect 29748 50188 30432 50216
rect 29748 50176 29754 50188
rect 30426 50176 30432 50188
rect 30484 50176 30490 50228
rect 31070 50176 31076 50228
rect 31128 50216 31134 50228
rect 31806 50216 31812 50228
rect 31128 50188 31812 50216
rect 31128 50176 31134 50188
rect 31806 50176 31812 50188
rect 31864 50176 31870 50228
rect 40914 50176 40920 50228
rect 40972 50216 40978 50228
rect 42018 50216 42024 50228
rect 40972 50188 42024 50216
rect 40972 50176 40978 50188
rect 42018 50176 42024 50188
rect 42076 50176 42082 50228
rect 114992 50160 115020 50244
rect 115084 50160 115112 50324
rect 118654 50176 118660 50228
rect 118712 50216 118718 50228
rect 119850 50216 119856 50228
rect 118712 50188 119856 50216
rect 118712 50176 118718 50188
rect 119850 50176 119856 50188
rect 119908 50176 119914 50228
rect 120954 50176 120960 50228
rect 121012 50216 121018 50228
rect 122058 50216 122064 50228
rect 121012 50188 122064 50216
rect 121012 50176 121018 50188
rect 122058 50176 122064 50188
rect 122116 50176 122122 50228
rect 125186 50176 125192 50228
rect 125244 50216 125250 50228
rect 126014 50216 126020 50228
rect 125244 50188 126020 50216
rect 125244 50176 125250 50188
rect 126014 50176 126020 50188
rect 126072 50176 126078 50228
rect 184434 50176 184440 50228
rect 184492 50216 184498 50228
rect 188206 50216 188212 50228
rect 184492 50188 188212 50216
rect 184492 50176 184498 50188
rect 188206 50176 188212 50188
rect 188264 50176 188270 50228
rect 193910 50176 193916 50228
rect 193968 50216 193974 50228
rect 194646 50216 194652 50228
rect 193968 50188 194652 50216
rect 193968 50176 193974 50188
rect 194646 50176 194652 50188
rect 194704 50176 194710 50228
rect 202374 50176 202380 50228
rect 202432 50216 202438 50228
rect 203570 50216 203576 50228
rect 202432 50188 203576 50216
rect 202432 50176 202438 50188
rect 203570 50176 203576 50188
rect 203628 50176 203634 50228
rect 205134 50176 205140 50228
rect 205192 50216 205198 50228
rect 205870 50216 205876 50228
rect 205192 50188 205876 50216
rect 205192 50176 205198 50188
rect 205870 50176 205876 50188
rect 205928 50176 205934 50228
rect 207986 50176 207992 50228
rect 208044 50216 208050 50228
rect 208722 50216 208728 50228
rect 208044 50188 208728 50216
rect 208044 50176 208050 50188
rect 208722 50176 208728 50188
rect 208780 50176 208786 50228
rect 212034 50176 212040 50228
rect 212092 50216 212098 50228
rect 214978 50216 214984 50228
rect 212092 50188 214984 50216
rect 212092 50176 212098 50188
rect 214978 50176 214984 50188
rect 215036 50176 215042 50228
rect 24906 50108 24912 50160
rect 24964 50148 24970 50160
rect 27942 50148 27948 50160
rect 24964 50120 27948 50148
rect 24964 50108 24970 50120
rect 27942 50108 27948 50120
rect 28000 50108 28006 50160
rect 114974 50108 114980 50160
rect 115032 50108 115038 50160
rect 115066 50108 115072 50160
rect 115124 50108 115130 50160
rect 205226 50108 205232 50160
rect 205284 50148 205290 50160
rect 206422 50148 206428 50160
rect 205284 50120 206428 50148
rect 205284 50108 205290 50120
rect 206422 50108 206428 50120
rect 206480 50108 206486 50160
rect 207894 50108 207900 50160
rect 207952 50148 207958 50160
rect 209274 50148 209280 50160
rect 207952 50120 209280 50148
rect 207952 50108 207958 50120
rect 209274 50108 209280 50120
rect 209332 50108 209338 50160
rect 210930 50108 210936 50160
rect 210988 50148 210994 50160
rect 212678 50148 212684 50160
rect 210988 50120 212684 50148
rect 210988 50108 210994 50120
rect 212678 50108 212684 50120
rect 212736 50108 212742 50160
rect 24262 50040 24268 50092
rect 24320 50080 24326 50092
rect 27850 50080 27856 50092
rect 24320 50052 27856 50080
rect 24320 50040 24326 50052
rect 27850 50040 27856 50052
rect 27908 50040 27914 50092
rect 29046 50040 29052 50092
rect 29104 50080 29110 50092
rect 30702 50080 30708 50092
rect 29104 50052 30708 50080
rect 29104 50040 29110 50052
rect 30702 50040 30708 50052
rect 30760 50040 30766 50092
rect 99518 50040 99524 50092
rect 99576 50080 99582 50092
rect 105314 50080 105320 50092
rect 99576 50052 105320 50080
rect 99576 50040 99582 50052
rect 105314 50040 105320 50052
rect 105372 50040 105378 50092
rect 205318 50040 205324 50092
rect 205376 50080 205382 50092
rect 206974 50080 206980 50092
rect 205376 50052 206980 50080
rect 205376 50040 205382 50052
rect 206974 50040 206980 50052
rect 207032 50040 207038 50092
rect 22238 49972 22244 50024
rect 22296 50012 22302 50024
rect 26838 50012 26844 50024
rect 22296 49984 26844 50012
rect 22296 49972 22302 49984
rect 26838 49972 26844 49984
rect 26896 49972 26902 50024
rect 27666 49972 27672 50024
rect 27724 50012 27730 50024
rect 29414 50012 29420 50024
rect 27724 49984 29420 50012
rect 27724 49972 27730 49984
rect 29414 49972 29420 49984
rect 29472 49972 29478 50024
rect 99242 49972 99248 50024
rect 99300 50012 99306 50024
rect 106418 50012 106424 50024
rect 99300 49984 106424 50012
rect 99300 49972 99306 49984
rect 106418 49972 106424 49984
rect 106476 49972 106482 50024
rect 183606 49972 183612 50024
rect 183664 50012 183670 50024
rect 189310 50012 189316 50024
rect 183664 49984 189316 50012
rect 183664 49972 183670 49984
rect 189310 49972 189316 49984
rect 189368 49972 189374 50024
rect 207250 49972 207256 50024
rect 207308 50012 207314 50024
rect 207894 50012 207900 50024
rect 207308 49984 207900 50012
rect 207308 49972 207314 49984
rect 207894 49972 207900 49984
rect 207952 49972 207958 50024
rect 23618 49904 23624 49956
rect 23676 49944 23682 49956
rect 26470 49944 26476 49956
rect 23676 49916 26476 49944
rect 23676 49904 23682 49916
rect 26470 49904 26476 49916
rect 26528 49904 26534 49956
rect 99334 49904 99340 49956
rect 99392 49944 99398 49956
rect 105866 49944 105872 49956
rect 99392 49916 105872 49944
rect 99392 49904 99398 49916
rect 105866 49904 105872 49916
rect 105924 49904 105930 49956
rect 121046 49904 121052 49956
rect 121104 49944 121110 49956
rect 122610 49944 122616 49956
rect 121104 49916 122616 49944
rect 121104 49904 121110 49916
rect 122610 49904 122616 49916
rect 122668 49904 122674 49956
rect 99150 49700 99156 49752
rect 99208 49740 99214 49752
rect 106970 49740 106976 49752
rect 99208 49712 106976 49740
rect 99208 49700 99214 49712
rect 106970 49700 106976 49712
rect 107028 49700 107034 49752
rect 26286 49632 26292 49684
rect 26344 49672 26350 49684
rect 29322 49672 29328 49684
rect 26344 49644 29328 49672
rect 26344 49632 26350 49644
rect 29322 49632 29328 49644
rect 29380 49632 29386 49684
rect 183238 49632 183244 49684
rect 183296 49672 183302 49684
rect 191058 49672 191064 49684
rect 183296 49644 191064 49672
rect 183296 49632 183302 49644
rect 191058 49632 191064 49644
rect 191116 49632 191122 49684
rect 99058 49564 99064 49616
rect 99116 49604 99122 49616
rect 107522 49604 107528 49616
rect 99116 49576 107528 49604
rect 99116 49564 99122 49576
rect 107522 49564 107528 49576
rect 107580 49564 107586 49616
rect 125094 49564 125100 49616
rect 125152 49604 125158 49616
rect 126566 49604 126572 49616
rect 125152 49576 126572 49604
rect 125152 49564 125158 49576
rect 126566 49564 126572 49576
rect 126624 49564 126630 49616
rect 183054 49564 183060 49616
rect 183112 49604 183118 49616
rect 192162 49604 192168 49616
rect 183112 49576 192168 49604
rect 183112 49564 183118 49576
rect 192162 49564 192168 49576
rect 192220 49564 192226 49616
rect 215530 49604 215536 49616
rect 210764 49576 215536 49604
rect 20214 49496 20220 49548
rect 20272 49536 20278 49548
rect 44502 49536 44508 49548
rect 20272 49508 44508 49536
rect 20272 49496 20278 49508
rect 44502 49496 44508 49508
rect 44560 49496 44566 49548
rect 98966 49496 98972 49548
rect 99024 49536 99030 49548
rect 108074 49536 108080 49548
rect 99024 49508 108080 49536
rect 99024 49496 99030 49508
rect 108074 49496 108080 49508
rect 108132 49496 108138 49548
rect 183146 49496 183152 49548
rect 183204 49536 183210 49548
rect 191610 49536 191616 49548
rect 183204 49508 191616 49536
rect 183204 49496 183210 49508
rect 191610 49496 191616 49508
rect 191668 49496 191674 49548
rect 191978 49496 191984 49548
rect 192036 49536 192042 49548
rect 210764 49536 210792 49576
rect 215530 49564 215536 49576
rect 215588 49564 215594 49616
rect 192036 49508 210792 49536
rect 192036 49496 192042 49508
rect 210838 49496 210844 49548
rect 210896 49536 210902 49548
rect 211574 49536 211580 49548
rect 210896 49508 211580 49536
rect 210896 49496 210902 49508
rect 211574 49496 211580 49508
rect 211632 49496 211638 49548
rect 212218 49496 212224 49548
rect 212276 49536 212282 49548
rect 213874 49536 213880 49548
rect 212276 49508 213880 49536
rect 212276 49496 212282 49508
rect 213874 49496 213880 49508
rect 213932 49496 213938 49548
rect 21502 49428 21508 49480
rect 21560 49468 21566 49480
rect 26562 49468 26568 49480
rect 21560 49440 26568 49468
rect 21560 49428 21566 49440
rect 26562 49428 26568 49440
rect 26620 49428 26626 49480
rect 183422 49224 183428 49276
rect 183480 49264 183486 49276
rect 189862 49264 189868 49276
rect 183480 49236 189868 49264
rect 183480 49224 183486 49236
rect 189862 49224 189868 49236
rect 189920 49224 189926 49276
rect 212126 49224 212132 49276
rect 212184 49264 212190 49276
rect 214426 49264 214432 49276
rect 212184 49236 214432 49264
rect 212184 49224 212190 49236
rect 214426 49224 214432 49236
rect 214484 49224 214490 49276
rect 28034 49196 28040 49208
rect 26948 49168 28040 49196
rect 25642 49088 25648 49140
rect 25700 49128 25706 49140
rect 26948 49128 26976 49168
rect 28034 49156 28040 49168
rect 28092 49156 28098 49208
rect 207158 49156 207164 49208
rect 207216 49196 207222 49208
rect 209826 49196 209832 49208
rect 207216 49168 209832 49196
rect 207216 49156 207222 49168
rect 209826 49156 209832 49168
rect 209884 49156 209890 49208
rect 25700 49100 26976 49128
rect 25700 49088 25706 49100
rect 27022 49088 27028 49140
rect 27080 49128 27086 49140
rect 29506 49128 29512 49140
rect 27080 49100 29512 49128
rect 27080 49088 27086 49100
rect 29506 49088 29512 49100
rect 29564 49088 29570 49140
rect 38154 49088 38160 49140
rect 38212 49128 38218 49140
rect 39258 49128 39264 49140
rect 38212 49100 39264 49128
rect 38212 49088 38218 49100
rect 39258 49088 39264 49100
rect 39316 49088 39322 49140
rect 183330 49088 183336 49140
rect 183388 49128 183394 49140
rect 190414 49128 190420 49140
rect 183388 49100 190420 49128
rect 183388 49088 183394 49100
rect 190414 49088 190420 49100
rect 190472 49088 190478 49140
rect 203018 49088 203024 49140
rect 203076 49128 203082 49140
rect 204122 49128 204128 49140
rect 203076 49100 204128 49128
rect 203076 49088 203082 49100
rect 204122 49088 204128 49100
rect 204180 49088 204186 49140
rect 210746 49088 210752 49140
rect 210804 49128 210810 49140
rect 212126 49128 212132 49140
rect 210804 49100 212132 49128
rect 210804 49088 210810 49100
rect 212126 49088 212132 49100
rect 212184 49088 212190 49140
rect 20858 49020 20864 49072
rect 20916 49060 20922 49072
rect 25090 49060 25096 49072
rect 20916 49032 25096 49060
rect 20916 49020 20922 49032
rect 25090 49020 25096 49032
rect 25148 49020 25154 49072
rect 38246 49020 38252 49072
rect 38304 49060 38310 49072
rect 39994 49060 40000 49072
rect 38304 49032 40000 49060
rect 38304 49020 38310 49032
rect 39994 49020 40000 49032
rect 40052 49020 40058 49072
rect 100254 49020 100260 49072
rect 100312 49060 100318 49072
rect 100312 49032 104900 49060
rect 100312 49020 100318 49032
rect 45054 48952 45060 49004
rect 45112 48992 45118 49004
rect 46802 48992 46808 49004
rect 45112 48964 46808 48992
rect 45112 48952 45118 48964
rect 46802 48952 46808 48964
rect 46860 48952 46866 49004
rect 100346 48952 100352 49004
rect 100404 48992 100410 49004
rect 104210 48992 104216 49004
rect 100404 48964 104216 48992
rect 100404 48952 100410 48964
rect 104210 48952 104216 48964
rect 104268 48952 104274 49004
rect 36130 48884 36136 48936
rect 36188 48924 36194 48936
rect 37234 48924 37240 48936
rect 36188 48896 37240 48924
rect 36188 48884 36194 48896
rect 37234 48884 37240 48896
rect 37292 48884 37298 48936
rect 43674 48884 43680 48936
rect 43732 48924 43738 48936
rect 44686 48924 44692 48936
rect 43732 48896 44692 48924
rect 43732 48884 43738 48896
rect 44686 48884 44692 48896
rect 44744 48884 44750 48936
rect 45146 48884 45152 48936
rect 45204 48924 45210 48936
rect 46066 48924 46072 48936
rect 45204 48896 46072 48924
rect 45204 48884 45210 48896
rect 46066 48884 46072 48896
rect 46124 48884 46130 48936
rect 46434 48884 46440 48936
rect 46492 48924 46498 48936
rect 47446 48924 47452 48936
rect 46492 48896 47452 48924
rect 46492 48884 46498 48896
rect 47446 48884 47452 48896
rect 47504 48884 47510 48936
rect 103014 48884 103020 48936
rect 103072 48924 103078 48936
rect 104762 48924 104768 48936
rect 103072 48896 104768 48924
rect 103072 48884 103078 48896
rect 104762 48884 104768 48896
rect 104820 48884 104826 48936
rect 104872 48924 104900 49032
rect 108626 48952 108632 49004
rect 108684 48992 108690 49004
rect 109178 48992 109184 49004
rect 108684 48964 109184 48992
rect 108684 48952 108690 48964
rect 109178 48952 109184 48964
rect 109236 48952 109242 49004
rect 109730 48952 109736 49004
rect 109788 48992 109794 49004
rect 110466 48992 110472 49004
rect 109788 48964 110472 48992
rect 109788 48952 109794 48964
rect 110466 48952 110472 48964
rect 110524 48952 110530 49004
rect 130982 48924 130988 48936
rect 104872 48896 130988 48924
rect 130982 48884 130988 48896
rect 131040 48884 131046 48936
rect 192714 48884 192720 48936
rect 192772 48924 192778 48936
rect 193358 48924 193364 48936
rect 192772 48896 193364 48924
rect 192772 48884 192778 48896
rect 193358 48884 193364 48896
rect 193416 48884 193422 48936
rect 96114 48816 96120 48868
rect 96172 48856 96178 48868
rect 222246 48856 222252 48868
rect 96172 48828 222252 48856
rect 96172 48816 96178 48828
rect 222246 48816 222252 48828
rect 222304 48816 222310 48868
rect 112490 47456 112496 47508
rect 112548 47496 112554 47508
rect 112582 47496 112588 47508
rect 112548 47468 112588 47496
rect 112548 47456 112554 47468
rect 112582 47456 112588 47468
rect 112640 47456 112646 47508
rect 197038 47456 197044 47508
rect 197096 47496 197102 47508
rect 197222 47496 197228 47508
rect 197096 47468 197228 47496
rect 197096 47456 197102 47468
rect 197222 47456 197228 47468
rect 197280 47456 197286 47508
rect 198053 47499 198111 47505
rect 198053 47465 198065 47499
rect 198099 47496 198111 47499
rect 198142 47496 198148 47508
rect 198099 47468 198148 47496
rect 198099 47465 198111 47468
rect 198053 47459 198111 47465
rect 198142 47456 198148 47468
rect 198200 47456 198206 47508
rect 50758 46504 50764 46556
rect 50816 46544 50822 46556
rect 61338 46544 61344 46556
rect 50816 46516 61344 46544
rect 50816 46504 50822 46516
rect 61338 46504 61344 46516
rect 61396 46504 61402 46556
rect 135122 46504 135128 46556
rect 135180 46544 135186 46556
rect 151314 46544 151320 46556
rect 135180 46516 151320 46544
rect 135180 46504 135186 46516
rect 151314 46504 151320 46516
rect 151372 46504 151378 46556
rect 49930 46436 49936 46488
rect 49988 46476 49994 46488
rect 58946 46476 58952 46488
rect 49988 46448 58952 46476
rect 49988 46436 49994 46448
rect 58946 46436 58952 46448
rect 59004 46436 59010 46488
rect 134754 46436 134760 46488
rect 134812 46476 134818 46488
rect 145334 46476 145340 46488
rect 134812 46448 145340 46476
rect 134812 46436 134818 46448
rect 145334 46436 145340 46448
rect 145392 46436 145398 46488
rect 50574 46368 50580 46420
rect 50632 46408 50638 46420
rect 62810 46408 62816 46420
rect 50632 46380 62816 46408
rect 50632 46368 50638 46380
rect 62810 46368 62816 46380
rect 62868 46368 62874 46420
rect 134938 46368 134944 46420
rect 134996 46408 135002 46420
rect 146806 46408 146812 46420
rect 134996 46380 146812 46408
rect 134996 46368 135002 46380
rect 146806 46368 146812 46380
rect 146864 46368 146870 46420
rect 51034 46300 51040 46352
rect 51092 46340 51098 46352
rect 64282 46340 64288 46352
rect 51092 46312 64288 46340
rect 51092 46300 51098 46312
rect 64282 46300 64288 46312
rect 64340 46300 64346 46352
rect 93354 46340 93360 46352
rect 84448 46312 93360 46340
rect 50850 46232 50856 46284
rect 50908 46272 50914 46284
rect 65754 46272 65760 46284
rect 50908 46244 65760 46272
rect 50908 46232 50914 46244
rect 65754 46232 65760 46244
rect 65812 46232 65818 46284
rect 50666 46164 50672 46216
rect 50724 46204 50730 46216
rect 67318 46204 67324 46216
rect 50724 46176 67324 46204
rect 50724 46164 50730 46176
rect 67318 46164 67324 46176
rect 67376 46164 67382 46216
rect 82958 46164 82964 46216
rect 83016 46204 83022 46216
rect 84448 46204 84476 46312
rect 93354 46300 93360 46312
rect 93412 46300 93418 46352
rect 134846 46300 134852 46352
rect 134904 46340 134910 46352
rect 148278 46340 148284 46352
rect 134904 46312 148284 46340
rect 134904 46300 134910 46312
rect 148278 46300 148284 46312
rect 148336 46300 148342 46352
rect 135030 46232 135036 46284
rect 135088 46272 135094 46284
rect 149750 46272 149756 46284
rect 135088 46244 149756 46272
rect 135088 46232 135094 46244
rect 149750 46232 149756 46244
rect 149808 46232 149814 46284
rect 94734 46204 94740 46216
rect 83016 46176 84476 46204
rect 88864 46176 94740 46204
rect 83016 46164 83022 46176
rect 50942 46096 50948 46148
rect 51000 46136 51006 46148
rect 68790 46136 68796 46148
rect 51000 46108 68796 46136
rect 51000 46096 51006 46108
rect 68790 46096 68796 46108
rect 68848 46096 68854 46148
rect 84062 46096 84068 46148
rect 84120 46136 84126 46148
rect 88864 46136 88892 46176
rect 94734 46164 94740 46176
rect 94792 46164 94798 46216
rect 135398 46164 135404 46216
rect 135456 46204 135462 46216
rect 140182 46204 140188 46216
rect 135456 46176 140188 46204
rect 135456 46164 135462 46176
rect 140182 46164 140188 46176
rect 140240 46164 140246 46216
rect 166954 46164 166960 46216
rect 167012 46204 167018 46216
rect 176154 46204 176160 46216
rect 167012 46176 176160 46204
rect 167012 46164 167018 46176
rect 176154 46164 176160 46176
rect 176212 46164 176218 46216
rect 84120 46108 88892 46136
rect 84120 46096 84126 46108
rect 88938 46096 88944 46148
rect 88996 46136 89002 46148
rect 96114 46136 96120 46148
rect 88996 46108 96120 46136
rect 88996 46096 89002 46108
rect 96114 46096 96120 46108
rect 96172 46096 96178 46148
rect 135306 46096 135312 46148
rect 135364 46136 135370 46148
rect 152786 46136 152792 46148
rect 135364 46108 152792 46136
rect 135364 46096 135370 46108
rect 152786 46096 152792 46108
rect 152844 46096 152850 46148
rect 168426 46096 168432 46148
rect 168484 46136 168490 46148
rect 177534 46136 177540 46148
rect 168484 46108 177540 46136
rect 168484 46096 168490 46108
rect 177534 46096 177540 46108
rect 177592 46096 177598 46148
rect 135398 45280 135404 45332
rect 135456 45320 135462 45332
rect 140274 45320 140280 45332
rect 135456 45292 140280 45320
rect 135456 45280 135462 45292
rect 140274 45280 140280 45292
rect 140332 45280 140338 45332
rect 181030 45280 181036 45332
rect 181088 45320 181094 45332
rect 185170 45320 185176 45332
rect 181088 45292 185176 45320
rect 181088 45280 181094 45292
rect 185170 45280 185176 45292
rect 185228 45280 185234 45332
rect 135398 45008 135404 45060
rect 135456 45048 135462 45060
rect 142298 45048 142304 45060
rect 135456 45020 142304 45048
rect 135456 45008 135462 45020
rect 142298 45008 142304 45020
rect 142356 45008 142362 45060
rect 53242 44736 53248 44788
rect 53300 44776 53306 44788
rect 59038 44776 59044 44788
rect 53300 44748 59044 44776
rect 53300 44736 53306 44748
rect 59038 44736 59044 44748
rect 59096 44736 59102 44788
rect 135398 44736 135404 44788
rect 135456 44776 135462 44788
rect 142206 44776 142212 44788
rect 135456 44748 142212 44776
rect 135456 44736 135462 44748
rect 142206 44736 142212 44748
rect 142264 44736 142270 44788
rect 53334 44668 53340 44720
rect 53392 44708 53398 44720
rect 58210 44708 58216 44720
rect 53392 44680 58216 44708
rect 53392 44668 53398 44680
rect 58210 44668 58216 44680
rect 58268 44668 58274 44720
rect 92802 44668 92808 44720
rect 92860 44708 92866 44720
rect 101726 44708 101732 44720
rect 92860 44680 101732 44708
rect 92860 44668 92866 44680
rect 101726 44668 101732 44680
rect 101784 44668 101790 44720
rect 140182 44668 140188 44720
rect 140240 44708 140246 44720
rect 143678 44708 143684 44720
rect 140240 44680 143684 44708
rect 140240 44668 140246 44680
rect 143678 44668 143684 44680
rect 143736 44668 143742 44720
rect 177718 44668 177724 44720
rect 177776 44708 177782 44720
rect 185906 44708 185912 44720
rect 177776 44680 185912 44708
rect 177776 44668 177782 44680
rect 185906 44668 185912 44680
rect 185964 44668 185970 44720
rect 92710 44600 92716 44652
rect 92768 44640 92774 44652
rect 101358 44640 101364 44652
rect 92768 44612 101364 44640
rect 92768 44600 92774 44612
rect 101358 44600 101364 44612
rect 101416 44600 101422 44652
rect 140274 44396 140280 44448
rect 140332 44436 140338 44448
rect 143494 44436 143500 44448
rect 140332 44408 143500 44436
rect 140332 44396 140338 44408
rect 143494 44396 143500 44408
rect 143552 44396 143558 44448
rect 177718 43852 177724 43904
rect 177776 43892 177782 43904
rect 181030 43892 181036 43904
rect 177776 43864 181036 43892
rect 177776 43852 177782 43864
rect 181030 43852 181036 43864
rect 181088 43852 181094 43904
rect 50022 43512 50028 43564
rect 50080 43552 50086 43564
rect 50080 43524 56784 43552
rect 50080 43512 50086 43524
rect 49930 43308 49936 43360
rect 49988 43348 49994 43360
rect 49988 43320 56692 43348
rect 49988 43308 49994 43320
rect 56664 43212 56692 43320
rect 56756 43280 56784 43524
rect 98138 43444 98144 43496
rect 98196 43484 98202 43496
rect 101634 43484 101640 43496
rect 98196 43456 101640 43484
rect 98196 43444 98202 43456
rect 101634 43444 101640 43456
rect 101692 43444 101698 43496
rect 135214 43376 135220 43428
rect 135272 43416 135278 43428
rect 136962 43416 136968 43428
rect 135272 43388 136968 43416
rect 135272 43376 135278 43388
rect 136962 43376 136968 43388
rect 137020 43376 137026 43428
rect 135398 43308 135404 43360
rect 135456 43348 135462 43360
rect 135456 43320 139676 43348
rect 135456 43308 135462 43320
rect 58210 43280 58216 43292
rect 56756 43252 58216 43280
rect 58210 43240 58216 43252
rect 58268 43240 58274 43292
rect 92710 43240 92716 43292
rect 92768 43280 92774 43292
rect 101818 43280 101824 43292
rect 92768 43252 101824 43280
rect 92768 43240 92774 43252
rect 101818 43240 101824 43252
rect 101876 43240 101882 43292
rect 139648 43280 139676 43320
rect 181858 43308 181864 43360
rect 181916 43348 181922 43360
rect 185170 43348 185176 43360
rect 181916 43320 185176 43348
rect 181916 43308 181922 43320
rect 185170 43308 185176 43320
rect 185228 43308 185234 43360
rect 142758 43280 142764 43292
rect 139648 43252 142764 43280
rect 142758 43240 142764 43252
rect 142816 43240 142822 43292
rect 177810 43240 177816 43292
rect 177868 43280 177874 43292
rect 185446 43280 185452 43292
rect 177868 43252 185452 43280
rect 177868 43240 177874 43252
rect 185446 43240 185452 43252
rect 185504 43240 185510 43292
rect 58302 43212 58308 43224
rect 56664 43184 58308 43212
rect 58302 43172 58308 43184
rect 58360 43172 58366 43224
rect 92894 43172 92900 43224
rect 92952 43212 92958 43224
rect 101266 43212 101272 43224
rect 92952 43184 101272 43212
rect 92952 43172 92958 43184
rect 101266 43172 101272 43184
rect 101324 43172 101330 43224
rect 177718 43172 177724 43224
rect 177776 43212 177782 43224
rect 185814 43212 185820 43224
rect 177776 43184 185820 43212
rect 177776 43172 177782 43184
rect 185814 43172 185820 43184
rect 185872 43172 185878 43224
rect 92802 43104 92808 43156
rect 92860 43144 92866 43156
rect 98138 43144 98144 43156
rect 92860 43116 98144 43144
rect 92860 43104 92866 43116
rect 98138 43104 98144 43116
rect 98196 43104 98202 43156
rect 49930 42424 49936 42476
rect 49988 42464 49994 42476
rect 56278 42464 56284 42476
rect 49988 42436 56284 42464
rect 49988 42424 49994 42436
rect 56278 42424 56284 42436
rect 56336 42424 56342 42476
rect 177718 42356 177724 42408
rect 177776 42396 177782 42408
rect 181858 42396 181864 42408
rect 177776 42368 181864 42396
rect 177776 42356 177782 42368
rect 181858 42356 181864 42368
rect 181916 42356 181922 42408
rect 50022 42288 50028 42340
rect 50080 42328 50086 42340
rect 56646 42328 56652 42340
rect 50080 42300 56652 42328
rect 50080 42288 50086 42300
rect 56646 42288 56652 42300
rect 56704 42288 56710 42340
rect 135214 42152 135220 42204
rect 135272 42192 135278 42204
rect 136870 42192 136876 42204
rect 135272 42164 136876 42192
rect 135272 42152 135278 42164
rect 136870 42152 136876 42164
rect 136928 42152 136934 42204
rect 49930 41948 49936 42000
rect 49988 41988 49994 42000
rect 58394 41988 58400 42000
rect 49988 41960 58400 41988
rect 49988 41948 49994 41960
rect 58394 41948 58400 41960
rect 58452 41948 58458 42000
rect 135398 41948 135404 42000
rect 135456 41988 135462 42000
rect 135456 41960 139676 41988
rect 135456 41948 135462 41960
rect 14694 41880 14700 41932
rect 14752 41920 14758 41932
rect 18098 41920 18104 41932
rect 14752 41892 18104 41920
rect 14752 41880 14758 41892
rect 18098 41880 18104 41892
rect 18156 41880 18162 41932
rect 56646 41880 56652 41932
rect 56704 41920 56710 41932
rect 58210 41920 58216 41932
rect 56704 41892 58216 41920
rect 56704 41880 56710 41892
rect 58210 41880 58216 41892
rect 58268 41880 58274 41932
rect 92802 41880 92808 41932
rect 92860 41920 92866 41932
rect 101726 41920 101732 41932
rect 92860 41892 101732 41920
rect 92860 41880 92866 41892
rect 101726 41880 101732 41892
rect 101784 41880 101790 41932
rect 139648 41920 139676 41960
rect 143310 41920 143316 41932
rect 139648 41892 143316 41920
rect 143310 41880 143316 41892
rect 143368 41880 143374 41932
rect 177626 41880 177632 41932
rect 177684 41920 177690 41932
rect 185170 41920 185176 41932
rect 177684 41892 185176 41920
rect 177684 41880 177690 41892
rect 185170 41880 185176 41892
rect 185228 41880 185234 41932
rect 92710 41812 92716 41864
rect 92768 41852 92774 41864
rect 100806 41852 100812 41864
rect 92768 41824 100812 41852
rect 92768 41812 92774 41824
rect 100806 41812 100812 41824
rect 100864 41812 100870 41864
rect 136962 41812 136968 41864
rect 137020 41852 137026 41864
rect 143402 41852 143408 41864
rect 137020 41824 143408 41852
rect 137020 41812 137026 41824
rect 143402 41812 143408 41824
rect 143460 41812 143466 41864
rect 177718 41812 177724 41864
rect 177776 41852 177782 41864
rect 184986 41852 184992 41864
rect 177776 41824 184992 41852
rect 177776 41812 177782 41824
rect 184986 41812 184992 41824
rect 185044 41812 185050 41864
rect 56278 41608 56284 41660
rect 56336 41648 56342 41660
rect 58302 41648 58308 41660
rect 56336 41620 58308 41648
rect 56336 41608 56342 41620
rect 58302 41608 58308 41620
rect 58360 41608 58366 41660
rect 135214 40792 135220 40844
rect 135272 40832 135278 40844
rect 136962 40832 136968 40844
rect 135272 40804 136968 40832
rect 135272 40792 135278 40804
rect 136962 40792 136968 40804
rect 137020 40792 137026 40844
rect 49930 40656 49936 40708
rect 49988 40696 49994 40708
rect 56646 40696 56652 40708
rect 49988 40668 56652 40696
rect 49988 40656 49994 40668
rect 56646 40656 56652 40668
rect 56704 40656 56710 40708
rect 50022 40588 50028 40640
rect 50080 40628 50086 40640
rect 56554 40628 56560 40640
rect 50080 40600 56560 40628
rect 50080 40588 50086 40600
rect 56554 40588 56560 40600
rect 56612 40588 56618 40640
rect 135398 40588 135404 40640
rect 135456 40628 135462 40640
rect 135456 40600 139676 40628
rect 135456 40588 135462 40600
rect 92802 40520 92808 40572
rect 92860 40560 92866 40572
rect 100990 40560 100996 40572
rect 92860 40532 100996 40560
rect 92860 40520 92866 40532
rect 100990 40520 100996 40532
rect 101048 40520 101054 40572
rect 139648 40560 139676 40600
rect 142482 40560 142488 40572
rect 139648 40532 142488 40560
rect 142482 40520 142488 40532
rect 142540 40520 142546 40572
rect 177258 40520 177264 40572
rect 177316 40560 177322 40572
rect 185170 40560 185176 40572
rect 177316 40532 185176 40560
rect 177316 40520 177322 40532
rect 185170 40520 185176 40532
rect 185228 40520 185234 40572
rect 92710 40452 92716 40504
rect 92768 40492 92774 40504
rect 100898 40492 100904 40504
rect 92768 40464 100904 40492
rect 92768 40452 92774 40464
rect 100898 40452 100904 40464
rect 100956 40452 100962 40504
rect 136870 40452 136876 40504
rect 136928 40492 136934 40504
rect 143678 40492 143684 40504
rect 136928 40464 143684 40492
rect 136928 40452 136934 40464
rect 143678 40452 143684 40464
rect 143736 40452 143742 40504
rect 177718 40452 177724 40504
rect 177776 40492 177782 40504
rect 185078 40492 185084 40504
rect 177776 40464 185084 40492
rect 177776 40452 177782 40464
rect 185078 40452 185084 40464
rect 185136 40452 185142 40504
rect 56554 40112 56560 40164
rect 56612 40152 56618 40164
rect 58210 40152 58216 40164
rect 56612 40124 58216 40152
rect 56612 40112 56618 40124
rect 58210 40112 58216 40124
rect 58268 40112 58274 40164
rect 51218 39228 51224 39280
rect 51276 39268 51282 39280
rect 56738 39268 56744 39280
rect 51276 39240 56744 39268
rect 51276 39228 51282 39240
rect 56738 39228 56744 39240
rect 56796 39228 56802 39280
rect 135214 39228 135220 39280
rect 135272 39268 135278 39280
rect 135272 39240 139860 39268
rect 135272 39228 135278 39240
rect 51126 39160 51132 39212
rect 51184 39200 51190 39212
rect 51184 39172 56140 39200
rect 51184 39160 51190 39172
rect 56112 38996 56140 39172
rect 135398 39160 135404 39212
rect 135456 39200 135462 39212
rect 135456 39172 139768 39200
rect 135456 39160 135462 39172
rect 92894 39092 92900 39144
rect 92952 39132 92958 39144
rect 100990 39132 100996 39144
rect 92952 39104 100996 39132
rect 92952 39092 92958 39104
rect 100990 39092 100996 39104
rect 101048 39092 101054 39144
rect 56646 39024 56652 39076
rect 56704 39064 56710 39076
rect 58302 39064 58308 39076
rect 56704 39036 58308 39064
rect 56704 39024 56710 39036
rect 58302 39024 58308 39036
rect 58360 39024 58366 39076
rect 92802 39024 92808 39076
rect 92860 39064 92866 39076
rect 101082 39064 101088 39076
rect 92860 39036 101088 39064
rect 92860 39024 92866 39036
rect 101082 39024 101088 39036
rect 101140 39024 101146 39076
rect 139740 39064 139768 39172
rect 139832 39132 139860 39240
rect 142850 39132 142856 39144
rect 139832 39104 142856 39132
rect 142850 39092 142856 39104
rect 142908 39092 142914 39144
rect 177718 39092 177724 39144
rect 177776 39132 177782 39144
rect 185170 39132 185176 39144
rect 177776 39104 185176 39132
rect 177776 39092 177782 39104
rect 185170 39092 185176 39104
rect 185228 39092 185234 39144
rect 143402 39064 143408 39076
rect 139740 39036 143408 39064
rect 143402 39024 143408 39036
rect 143460 39024 143466 39076
rect 177350 39024 177356 39076
rect 177408 39064 177414 39076
rect 185262 39064 185268 39076
rect 177408 39036 185268 39064
rect 177408 39024 177414 39036
rect 185262 39024 185268 39036
rect 185320 39024 185326 39076
rect 58210 38996 58216 39008
rect 56112 38968 58216 38996
rect 58210 38956 58216 38968
rect 58268 38956 58274 39008
rect 92710 38956 92716 39008
rect 92768 38996 92774 39008
rect 100806 38996 100812 39008
rect 92768 38968 100812 38996
rect 92768 38956 92774 38968
rect 100806 38956 100812 38968
rect 100864 38956 100870 39008
rect 136962 38956 136968 39008
rect 137020 38996 137026 39008
rect 143678 38996 143684 39008
rect 137020 38968 143684 38996
rect 137020 38956 137026 38968
rect 143678 38956 143684 38968
rect 143736 38956 143742 39008
rect 177258 38956 177264 39008
rect 177316 38996 177322 39008
rect 184986 38996 184992 39008
rect 177316 38968 184992 38996
rect 177316 38956 177322 38968
rect 184986 38956 184992 38968
rect 185044 38956 185050 39008
rect 56738 38616 56744 38668
rect 56796 38656 56802 38668
rect 58394 38656 58400 38668
rect 56796 38628 58400 38656
rect 56796 38616 56802 38628
rect 58394 38616 58400 38628
rect 58452 38616 58458 38668
rect 98966 38344 98972 38396
rect 99024 38384 99030 38396
rect 101174 38384 101180 38396
rect 99024 38356 101180 38384
rect 99024 38344 99030 38356
rect 101174 38344 101180 38356
rect 101232 38344 101238 38396
rect 98874 38208 98880 38260
rect 98932 38248 98938 38260
rect 100990 38248 100996 38260
rect 98932 38220 100996 38248
rect 98932 38208 98938 38220
rect 100990 38208 100996 38220
rect 101048 38208 101054 38260
rect 135398 38208 135404 38260
rect 135456 38248 135462 38260
rect 139630 38248 139636 38260
rect 135456 38220 139636 38248
rect 135456 38208 135462 38220
rect 139630 38208 139636 38220
rect 139688 38208 139694 38260
rect 183238 38072 183244 38124
rect 183296 38112 183302 38124
rect 185262 38112 185268 38124
rect 183296 38084 185268 38112
rect 183296 38072 183302 38084
rect 185262 38072 185268 38084
rect 185320 38072 185326 38124
rect 51218 37868 51224 37920
rect 51276 37908 51282 37920
rect 58302 37908 58308 37920
rect 51276 37880 58308 37908
rect 51276 37868 51282 37880
rect 58302 37868 58308 37880
rect 58360 37868 58366 37920
rect 135398 37868 135404 37920
rect 135456 37908 135462 37920
rect 136870 37908 136876 37920
rect 135456 37880 136876 37908
rect 135456 37868 135462 37880
rect 136870 37868 136876 37880
rect 136928 37868 136934 37920
rect 51126 37800 51132 37852
rect 51184 37840 51190 37852
rect 58210 37840 58216 37852
rect 51184 37812 58216 37840
rect 51184 37800 51190 37812
rect 58210 37800 58216 37812
rect 58268 37800 58274 37852
rect 135214 37800 135220 37852
rect 135272 37840 135278 37852
rect 135272 37812 139768 37840
rect 135272 37800 135278 37812
rect 92802 37732 92808 37784
rect 92860 37772 92866 37784
rect 98874 37772 98880 37784
rect 92860 37744 98880 37772
rect 92860 37732 92866 37744
rect 98874 37732 98880 37744
rect 98932 37732 98938 37784
rect 92710 37664 92716 37716
rect 92768 37704 92774 37716
rect 98966 37704 98972 37716
rect 92768 37676 98972 37704
rect 92768 37664 92774 37676
rect 98966 37664 98972 37676
rect 99024 37664 99030 37716
rect 139740 37500 139768 37812
rect 183698 37800 183704 37852
rect 183756 37840 183762 37852
rect 185170 37840 185176 37852
rect 183756 37812 185176 37840
rect 183756 37800 183762 37812
rect 185170 37800 185176 37812
rect 185228 37800 185234 37852
rect 143678 37500 143684 37512
rect 139740 37472 143684 37500
rect 143678 37460 143684 37472
rect 143736 37460 143742 37512
rect 177718 37324 177724 37376
rect 177776 37364 177782 37376
rect 183238 37364 183244 37376
rect 177776 37336 183244 37364
rect 177776 37324 177782 37336
rect 183238 37324 183244 37336
rect 183296 37324 183302 37376
rect 139630 37188 139636 37240
rect 139688 37228 139694 37240
rect 143494 37228 143500 37240
rect 139688 37200 143500 37228
rect 139688 37188 139694 37200
rect 143494 37188 143500 37200
rect 143552 37188 143558 37240
rect 177442 36848 177448 36900
rect 177500 36888 177506 36900
rect 183698 36888 183704 36900
rect 177500 36860 183704 36888
rect 177500 36848 177506 36860
rect 183698 36848 183704 36860
rect 183756 36848 183762 36900
rect 51126 36576 51132 36628
rect 51184 36616 51190 36628
rect 55542 36616 55548 36628
rect 51184 36588 55548 36616
rect 51184 36576 51190 36588
rect 55542 36576 55548 36588
rect 55600 36576 55606 36628
rect 134662 36576 134668 36628
rect 134720 36616 134726 36628
rect 136778 36616 136784 36628
rect 134720 36588 136784 36616
rect 134720 36576 134726 36588
rect 136778 36576 136784 36588
rect 136836 36576 136842 36628
rect 51218 36508 51224 36560
rect 51276 36548 51282 36560
rect 58302 36548 58308 36560
rect 51276 36520 58308 36548
rect 51276 36508 51282 36520
rect 58302 36508 58308 36520
rect 58360 36508 58366 36560
rect 50206 36440 50212 36492
rect 50264 36480 50270 36492
rect 58210 36480 58216 36492
rect 50264 36452 58216 36480
rect 50264 36440 50270 36452
rect 58210 36440 58216 36452
rect 58268 36440 58274 36492
rect 135398 36440 135404 36492
rect 135456 36480 135462 36492
rect 135456 36452 139676 36480
rect 135456 36440 135462 36452
rect 92802 36372 92808 36424
rect 92860 36412 92866 36424
rect 100990 36412 100996 36424
rect 92860 36384 100996 36412
rect 92860 36372 92866 36384
rect 100990 36372 100996 36384
rect 101048 36372 101054 36424
rect 139648 36412 139676 36452
rect 143034 36412 143040 36424
rect 139648 36384 143040 36412
rect 143034 36372 143040 36384
rect 143092 36372 143098 36424
rect 177350 36372 177356 36424
rect 177408 36412 177414 36424
rect 185170 36412 185176 36424
rect 177408 36384 185176 36412
rect 177408 36372 177414 36384
rect 185170 36372 185176 36384
rect 185228 36372 185234 36424
rect 92710 36304 92716 36356
rect 92768 36344 92774 36356
rect 100530 36344 100536 36356
rect 92768 36316 100536 36344
rect 92768 36304 92774 36316
rect 100530 36304 100536 36316
rect 100588 36304 100594 36356
rect 177442 36304 177448 36356
rect 177500 36344 177506 36356
rect 184986 36344 184992 36356
rect 177500 36316 184992 36344
rect 177500 36304 177506 36316
rect 184986 36304 184992 36316
rect 185044 36304 185050 36356
rect 136870 36236 136876 36288
rect 136928 36276 136934 36288
rect 143678 36276 143684 36288
rect 136928 36248 143684 36276
rect 136928 36236 136934 36248
rect 143678 36236 143684 36248
rect 143736 36236 143742 36288
rect 51218 35352 51224 35404
rect 51276 35392 51282 35404
rect 55450 35392 55456 35404
rect 51276 35364 55456 35392
rect 51276 35352 51282 35364
rect 55450 35352 55456 35364
rect 55508 35352 55514 35404
rect 135214 35216 135220 35268
rect 135272 35256 135278 35268
rect 138158 35256 138164 35268
rect 135272 35228 138164 35256
rect 135272 35216 135278 35228
rect 138158 35216 138164 35228
rect 138216 35216 138222 35268
rect 51218 35080 51224 35132
rect 51276 35120 51282 35132
rect 59222 35120 59228 35132
rect 51276 35092 59228 35120
rect 51276 35080 51282 35092
rect 59222 35080 59228 35092
rect 59280 35080 59286 35132
rect 135398 35080 135404 35132
rect 135456 35120 135462 35132
rect 142390 35120 142396 35132
rect 135456 35092 142396 35120
rect 135456 35080 135462 35092
rect 142390 35080 142396 35092
rect 142448 35080 142454 35132
rect 92802 35012 92808 35064
rect 92860 35052 92866 35064
rect 100990 35052 100996 35064
rect 92860 35024 100996 35052
rect 92860 35012 92866 35024
rect 100990 35012 100996 35024
rect 101048 35012 101054 35064
rect 136778 35012 136784 35064
rect 136836 35052 136842 35064
rect 143678 35052 143684 35064
rect 136836 35024 143684 35052
rect 136836 35012 136842 35024
rect 143678 35012 143684 35024
rect 143736 35012 143742 35064
rect 177718 35012 177724 35064
rect 177776 35052 177782 35064
rect 185446 35052 185452 35064
rect 177776 35024 185452 35052
rect 177776 35012 177782 35024
rect 185446 35012 185452 35024
rect 185504 35012 185510 35064
rect 55542 34944 55548 34996
rect 55600 34984 55606 34996
rect 58302 34984 58308 34996
rect 55600 34956 58308 34984
rect 55600 34944 55606 34956
rect 58302 34944 58308 34956
rect 58360 34944 58366 34996
rect 92710 34944 92716 34996
rect 92768 34984 92774 34996
rect 100898 34984 100904 34996
rect 92768 34956 100904 34984
rect 92768 34944 92774 34956
rect 100898 34944 100904 34956
rect 100956 34944 100962 34996
rect 177258 34944 177264 34996
rect 177316 34984 177322 34996
rect 185078 34984 185084 34996
rect 177316 34956 185084 34984
rect 177316 34944 177322 34956
rect 185078 34944 185084 34956
rect 185136 34944 185142 34996
rect 55450 34740 55456 34792
rect 55508 34780 55514 34792
rect 58210 34780 58216 34792
rect 55508 34752 58216 34780
rect 55508 34740 55514 34752
rect 58210 34740 58216 34752
rect 58268 34740 58274 34792
rect 134662 33788 134668 33840
rect 134720 33828 134726 33840
rect 136962 33828 136968 33840
rect 134720 33800 136968 33828
rect 134720 33788 134726 33800
rect 136962 33788 136968 33800
rect 137020 33788 137026 33840
rect 51218 33720 51224 33772
rect 51276 33760 51282 33772
rect 56462 33760 56468 33772
rect 51276 33732 56468 33760
rect 51276 33720 51282 33732
rect 56462 33720 56468 33732
rect 56520 33720 56526 33772
rect 135214 33720 135220 33772
rect 135272 33760 135278 33772
rect 135272 33732 139768 33760
rect 135272 33720 135278 33732
rect 51126 33652 51132 33704
rect 51184 33692 51190 33704
rect 56738 33692 56744 33704
rect 51184 33664 56744 33692
rect 51184 33652 51190 33664
rect 56738 33652 56744 33664
rect 56796 33652 56802 33704
rect 135398 33652 135404 33704
rect 135456 33692 135462 33704
rect 135456 33664 139676 33692
rect 135456 33652 135462 33664
rect 92802 33584 92808 33636
rect 92860 33624 92866 33636
rect 101082 33624 101088 33636
rect 92860 33596 101088 33624
rect 92860 33584 92866 33596
rect 101082 33584 101088 33596
rect 101140 33584 101146 33636
rect 92894 33516 92900 33568
rect 92952 33556 92958 33568
rect 100990 33556 100996 33568
rect 92952 33528 100996 33556
rect 92952 33516 92958 33528
rect 100990 33516 100996 33528
rect 101048 33516 101054 33568
rect 139648 33556 139676 33664
rect 139740 33624 139768 33732
rect 143310 33624 143316 33636
rect 139740 33596 143316 33624
rect 143310 33584 143316 33596
rect 143368 33584 143374 33636
rect 177810 33584 177816 33636
rect 177868 33624 177874 33636
rect 185170 33624 185176 33636
rect 177868 33596 185176 33624
rect 177868 33584 177874 33596
rect 185170 33584 185176 33596
rect 185228 33584 185234 33636
rect 142758 33556 142764 33568
rect 139648 33528 142764 33556
rect 142758 33516 142764 33528
rect 142816 33516 142822 33568
rect 177718 33516 177724 33568
rect 177776 33556 177782 33568
rect 185262 33556 185268 33568
rect 177776 33528 185268 33556
rect 177776 33516 177782 33528
rect 185262 33516 185268 33528
rect 185320 33516 185326 33568
rect 92710 33448 92716 33500
rect 92768 33488 92774 33500
rect 100714 33488 100720 33500
rect 92768 33460 100720 33488
rect 92768 33448 92774 33460
rect 100714 33448 100720 33460
rect 100772 33448 100778 33500
rect 138158 33448 138164 33500
rect 138216 33488 138222 33500
rect 143678 33488 143684 33500
rect 138216 33460 143684 33488
rect 138216 33448 138222 33460
rect 143678 33448 143684 33460
rect 143736 33448 143742 33500
rect 177626 33448 177632 33500
rect 177684 33488 177690 33500
rect 184894 33488 184900 33500
rect 177684 33460 184900 33488
rect 177684 33448 177690 33460
rect 184894 33448 184900 33460
rect 184952 33448 184958 33500
rect 56738 33380 56744 33432
rect 56796 33420 56802 33432
rect 58210 33420 58216 33432
rect 56796 33392 58216 33420
rect 56796 33380 56802 33392
rect 58210 33380 58216 33392
rect 58268 33380 58274 33432
rect 56462 33040 56468 33092
rect 56520 33080 56526 33092
rect 58302 33080 58308 33092
rect 56520 33052 58308 33080
rect 56520 33040 56526 33052
rect 58302 33040 58308 33052
rect 58360 33040 58366 33092
rect 50022 32496 50028 32548
rect 50080 32536 50086 32548
rect 50080 32508 56784 32536
rect 50080 32496 50086 32508
rect 51218 32292 51224 32344
rect 51276 32332 51282 32344
rect 51276 32304 56692 32332
rect 51276 32292 51282 32304
rect 56664 32196 56692 32304
rect 56756 32264 56784 32508
rect 135214 32360 135220 32412
rect 135272 32400 135278 32412
rect 136870 32400 136876 32412
rect 135272 32372 136876 32400
rect 135272 32360 135278 32372
rect 136870 32360 136876 32372
rect 136928 32360 136934 32412
rect 135398 32292 135404 32344
rect 135456 32332 135462 32344
rect 135456 32304 139676 32332
rect 135456 32292 135462 32304
rect 58210 32264 58216 32276
rect 56756 32236 58216 32264
rect 58210 32224 58216 32236
rect 58268 32224 58274 32276
rect 92802 32224 92808 32276
rect 92860 32264 92866 32276
rect 100990 32264 100996 32276
rect 92860 32236 100996 32264
rect 92860 32224 92866 32236
rect 100990 32224 100996 32236
rect 101048 32224 101054 32276
rect 139648 32264 139676 32304
rect 142574 32264 142580 32276
rect 139648 32236 142580 32264
rect 142574 32224 142580 32236
rect 142632 32224 142638 32276
rect 177626 32224 177632 32276
rect 177684 32264 177690 32276
rect 185170 32264 185176 32276
rect 177684 32236 185176 32264
rect 177684 32224 177690 32236
rect 185170 32224 185176 32236
rect 185228 32224 185234 32276
rect 58302 32196 58308 32208
rect 56664 32168 58308 32196
rect 58302 32156 58308 32168
rect 58360 32156 58366 32208
rect 92710 32156 92716 32208
rect 92768 32196 92774 32208
rect 100806 32196 100812 32208
rect 92768 32168 100812 32196
rect 92768 32156 92774 32168
rect 100806 32156 100812 32168
rect 100864 32156 100870 32208
rect 136962 32156 136968 32208
rect 137020 32196 137026 32208
rect 143678 32196 143684 32208
rect 137020 32168 143684 32196
rect 137020 32156 137026 32168
rect 143678 32156 143684 32168
rect 143736 32156 143742 32208
rect 177718 32156 177724 32208
rect 177776 32196 177782 32208
rect 184986 32196 184992 32208
rect 177776 32168 184992 32196
rect 177776 32156 177782 32168
rect 184986 32156 184992 32168
rect 185044 32156 185050 32208
rect 50022 31272 50028 31324
rect 50080 31312 50086 31324
rect 56738 31312 56744 31324
rect 50080 31284 56744 31312
rect 50080 31272 50086 31284
rect 56738 31272 56744 31284
rect 56796 31272 56802 31324
rect 51218 31136 51224 31188
rect 51276 31176 51282 31188
rect 56646 31176 56652 31188
rect 51276 31148 56652 31176
rect 51276 31136 51282 31148
rect 56646 31136 56652 31148
rect 56704 31136 56710 31188
rect 135214 31136 135220 31188
rect 135272 31176 135278 31188
rect 136962 31176 136968 31188
rect 135272 31148 136968 31176
rect 135272 31136 135278 31148
rect 136962 31136 136968 31148
rect 137020 31136 137026 31188
rect 51218 30932 51224 30984
rect 51276 30972 51282 30984
rect 58394 30972 58400 30984
rect 51276 30944 58400 30972
rect 51276 30932 51282 30944
rect 58394 30932 58400 30944
rect 58452 30932 58458 30984
rect 135398 30932 135404 30984
rect 135456 30972 135462 30984
rect 135456 30944 139676 30972
rect 135456 30932 135462 30944
rect 56646 30864 56652 30916
rect 56704 30904 56710 30916
rect 58210 30904 58216 30916
rect 56704 30876 58216 30904
rect 56704 30864 56710 30876
rect 58210 30864 58216 30876
rect 58268 30864 58274 30916
rect 92802 30864 92808 30916
rect 92860 30904 92866 30916
rect 100990 30904 100996 30916
rect 92860 30876 100996 30904
rect 92860 30864 92866 30876
rect 100990 30864 100996 30876
rect 101048 30864 101054 30916
rect 139648 30904 139676 30944
rect 142758 30904 142764 30916
rect 139648 30876 142764 30904
rect 142758 30864 142764 30876
rect 142816 30864 142822 30916
rect 177718 30864 177724 30916
rect 177776 30904 177782 30916
rect 185170 30904 185176 30916
rect 177776 30876 185176 30904
rect 177776 30864 177782 30876
rect 185170 30864 185176 30876
rect 185228 30864 185234 30916
rect 56738 30796 56744 30848
rect 56796 30836 56802 30848
rect 58302 30836 58308 30848
rect 56796 30808 58308 30836
rect 56796 30796 56802 30808
rect 58302 30796 58308 30808
rect 58360 30796 58366 30848
rect 92710 30796 92716 30848
rect 92768 30836 92774 30848
rect 100898 30836 100904 30848
rect 92768 30808 100904 30836
rect 92768 30796 92774 30808
rect 100898 30796 100904 30808
rect 100956 30796 100962 30848
rect 136870 30796 136876 30848
rect 136928 30836 136934 30848
rect 143678 30836 143684 30848
rect 136928 30808 143684 30836
rect 136928 30796 136934 30808
rect 143678 30796 143684 30808
rect 143736 30796 143742 30848
rect 177442 30796 177448 30848
rect 177500 30836 177506 30848
rect 185078 30836 185084 30848
rect 177500 30808 185084 30836
rect 177500 30796 177506 30808
rect 185078 30796 185084 30808
rect 185136 30796 185142 30848
rect 51218 29640 51224 29692
rect 51276 29680 51282 29692
rect 56002 29680 56008 29692
rect 51276 29652 56008 29680
rect 51276 29640 51282 29652
rect 56002 29640 56008 29652
rect 56060 29640 56066 29692
rect 135214 29572 135220 29624
rect 135272 29612 135278 29624
rect 135272 29584 139860 29612
rect 135272 29572 135278 29584
rect 51126 29504 51132 29556
rect 51184 29544 51190 29556
rect 51184 29516 56784 29544
rect 51184 29504 51190 29516
rect 56756 29408 56784 29516
rect 135398 29504 135404 29556
rect 135456 29544 135462 29556
rect 135456 29516 139768 29544
rect 135456 29504 135462 29516
rect 92894 29436 92900 29488
rect 92952 29476 92958 29488
rect 101082 29476 101088 29488
rect 92952 29448 101088 29476
rect 92952 29436 92958 29448
rect 101082 29436 101088 29448
rect 101140 29436 101146 29488
rect 58210 29408 58216 29420
rect 56756 29380 58216 29408
rect 58210 29368 58216 29380
rect 58268 29368 58274 29420
rect 92802 29368 92808 29420
rect 92860 29408 92866 29420
rect 100990 29408 100996 29420
rect 92860 29380 100996 29408
rect 92860 29368 92866 29380
rect 100990 29368 100996 29380
rect 101048 29368 101054 29420
rect 139740 29408 139768 29516
rect 139832 29476 139860 29584
rect 143586 29476 143592 29488
rect 139832 29448 143592 29476
rect 143586 29436 143592 29448
rect 143644 29436 143650 29488
rect 177718 29436 177724 29488
rect 177776 29476 177782 29488
rect 185262 29476 185268 29488
rect 177776 29448 185268 29476
rect 177776 29436 177782 29448
rect 185262 29436 185268 29448
rect 185320 29436 185326 29488
rect 142758 29408 142764 29420
rect 139740 29380 142764 29408
rect 142758 29368 142764 29380
rect 142816 29368 142822 29420
rect 177442 29368 177448 29420
rect 177500 29408 177506 29420
rect 185170 29408 185176 29420
rect 177500 29380 185176 29408
rect 177500 29368 177506 29380
rect 185170 29368 185176 29380
rect 185228 29368 185234 29420
rect 92710 29300 92716 29352
rect 92768 29340 92774 29352
rect 100806 29340 100812 29352
rect 92768 29312 100812 29340
rect 92768 29300 92774 29312
rect 100806 29300 100812 29312
rect 100864 29300 100870 29352
rect 136962 29300 136968 29352
rect 137020 29340 137026 29352
rect 143678 29340 143684 29352
rect 137020 29312 143684 29340
rect 137020 29300 137026 29312
rect 143678 29300 143684 29312
rect 143736 29300 143742 29352
rect 177258 29300 177264 29352
rect 177316 29340 177322 29352
rect 184986 29340 184992 29352
rect 177316 29312 184992 29340
rect 177316 29300 177322 29312
rect 184986 29300 184992 29312
rect 185044 29300 185050 29352
rect 56002 28892 56008 28944
rect 56060 28932 56066 28944
rect 58302 28932 58308 28944
rect 56060 28904 58308 28932
rect 56060 28892 56066 28904
rect 58302 28892 58308 28904
rect 58360 28892 58366 28944
rect 135398 28416 135404 28468
rect 135456 28456 135462 28468
rect 139630 28456 139636 28468
rect 135456 28428 139636 28456
rect 135456 28416 135462 28428
rect 139630 28416 139636 28428
rect 139688 28416 139694 28468
rect 51126 28280 51132 28332
rect 51184 28320 51190 28332
rect 56370 28320 56376 28332
rect 51184 28292 56376 28320
rect 51184 28280 51190 28292
rect 56370 28280 56376 28292
rect 56428 28280 56434 28332
rect 135398 28280 135404 28332
rect 135456 28320 135462 28332
rect 137330 28320 137336 28332
rect 135456 28292 137336 28320
rect 135456 28280 135462 28292
rect 137330 28280 137336 28292
rect 137388 28280 137394 28332
rect 51218 28144 51224 28196
rect 51276 28184 51282 28196
rect 51276 28156 56324 28184
rect 51276 28144 51282 28156
rect 56296 27980 56324 28156
rect 92894 28144 92900 28196
rect 92952 28184 92958 28196
rect 100990 28184 100996 28196
rect 92952 28156 100996 28184
rect 92952 28144 92958 28156
rect 100990 28144 100996 28156
rect 101048 28144 101054 28196
rect 135214 28144 135220 28196
rect 135272 28184 135278 28196
rect 135272 28156 139768 28184
rect 135272 28144 135278 28156
rect 92802 28076 92808 28128
rect 92860 28116 92866 28128
rect 101910 28116 101916 28128
rect 92860 28088 101916 28116
rect 92860 28076 92866 28088
rect 101910 28076 101916 28088
rect 101968 28076 101974 28128
rect 56370 28008 56376 28060
rect 56428 28048 56434 28060
rect 58302 28048 58308 28060
rect 56428 28020 58308 28048
rect 56428 28008 56434 28020
rect 58302 28008 58308 28020
rect 58360 28008 58366 28060
rect 92710 28008 92716 28060
rect 92768 28048 92774 28060
rect 101726 28048 101732 28060
rect 92768 28020 101732 28048
rect 92768 28008 92774 28020
rect 101726 28008 101732 28020
rect 101784 28008 101790 28060
rect 58210 27980 58216 27992
rect 56296 27952 58216 27980
rect 58210 27940 58216 27952
rect 58268 27940 58274 27992
rect 139740 27980 139768 28156
rect 177626 28144 177632 28196
rect 177684 28184 177690 28196
rect 185170 28184 185176 28196
rect 177684 28156 185176 28184
rect 177684 28144 177690 28156
rect 185170 28144 185176 28156
rect 185228 28144 185234 28196
rect 177350 28076 177356 28128
rect 177408 28116 177414 28128
rect 185262 28116 185268 28128
rect 177408 28088 185268 28116
rect 177408 28076 177414 28088
rect 185262 28076 185268 28088
rect 185320 28076 185326 28128
rect 177718 28008 177724 28060
rect 177776 28048 177782 28060
rect 185354 28048 185360 28060
rect 177776 28020 185360 28048
rect 177776 28008 177782 28020
rect 185354 28008 185360 28020
rect 185412 28008 185418 28060
rect 143678 27980 143684 27992
rect 139740 27952 143684 27980
rect 143678 27940 143684 27952
rect 143736 27940 143742 27992
rect 139630 27532 139636 27584
rect 139688 27572 139694 27584
rect 143402 27572 143408 27584
rect 139688 27544 143408 27572
rect 139688 27532 139694 27544
rect 143402 27532 143408 27544
rect 143460 27532 143466 27584
rect 51126 26920 51132 26972
rect 51184 26960 51190 26972
rect 59038 26960 59044 26972
rect 51184 26932 59044 26960
rect 51184 26920 51190 26932
rect 59038 26920 59044 26932
rect 59096 26920 59102 26972
rect 135214 26920 135220 26972
rect 135272 26960 135278 26972
rect 138158 26960 138164 26972
rect 135272 26932 138164 26960
rect 135272 26920 135278 26932
rect 138158 26920 138164 26932
rect 138216 26920 138222 26972
rect 51218 26852 51224 26904
rect 51276 26892 51282 26904
rect 58302 26892 58308 26904
rect 51276 26864 58308 26892
rect 51276 26852 51282 26864
rect 58302 26852 58308 26864
rect 58360 26852 58366 26904
rect 50022 26784 50028 26836
rect 50080 26824 50086 26836
rect 58210 26824 58216 26836
rect 50080 26796 58216 26824
rect 50080 26784 50086 26796
rect 58210 26784 58216 26796
rect 58268 26784 58274 26836
rect 100990 26824 100996 26836
rect 98616 26796 100996 26824
rect 92710 26716 92716 26768
rect 92768 26756 92774 26768
rect 98616 26756 98644 26796
rect 100990 26784 100996 26796
rect 101048 26784 101054 26836
rect 135398 26784 135404 26836
rect 135456 26824 135462 26836
rect 185170 26824 185176 26836
rect 135456 26796 139676 26824
rect 135456 26784 135462 26796
rect 92768 26728 98644 26756
rect 139648 26756 139676 26796
rect 183716 26796 185176 26824
rect 143586 26756 143592 26768
rect 139648 26728 143592 26756
rect 92768 26716 92774 26728
rect 143586 26716 143592 26728
rect 143644 26716 143650 26768
rect 177718 26716 177724 26768
rect 177776 26756 177782 26768
rect 183716 26756 183744 26796
rect 185170 26784 185176 26796
rect 185228 26784 185234 26836
rect 177776 26728 183744 26756
rect 177776 26716 177782 26728
rect 137330 26580 137336 26632
rect 137388 26620 137394 26632
rect 143678 26620 143684 26632
rect 137388 26592 143684 26620
rect 137388 26580 137394 26592
rect 143678 26580 143684 26592
rect 143736 26580 143742 26632
rect 51218 25492 51224 25544
rect 51276 25532 51282 25544
rect 59406 25532 59412 25544
rect 51276 25504 59412 25532
rect 51276 25492 51282 25504
rect 59406 25492 59412 25504
rect 59464 25492 59470 25544
rect 135214 25492 135220 25544
rect 135272 25532 135278 25544
rect 135272 25504 140228 25532
rect 135272 25492 135278 25504
rect 51126 25424 51132 25476
rect 51184 25464 51190 25476
rect 59498 25464 59504 25476
rect 51184 25436 59504 25464
rect 51184 25424 51190 25436
rect 59498 25424 59504 25436
rect 59556 25424 59562 25476
rect 135398 25424 135404 25476
rect 135456 25464 135462 25476
rect 135456 25436 140136 25464
rect 135456 25424 135462 25436
rect 50298 25356 50304 25408
rect 50356 25396 50362 25408
rect 50666 25396 50672 25408
rect 50356 25368 50672 25396
rect 50356 25356 50362 25368
rect 50666 25356 50672 25368
rect 50724 25356 50730 25408
rect 92894 25356 92900 25408
rect 92952 25396 92958 25408
rect 101174 25396 101180 25408
rect 92952 25368 101180 25396
rect 92952 25356 92958 25368
rect 101174 25356 101180 25368
rect 101232 25356 101238 25408
rect 92802 25288 92808 25340
rect 92860 25328 92866 25340
rect 101082 25328 101088 25340
rect 92860 25300 101088 25328
rect 92860 25288 92866 25300
rect 101082 25288 101088 25300
rect 101140 25288 101146 25340
rect 140108 25328 140136 25436
rect 140200 25396 140228 25504
rect 143678 25396 143684 25408
rect 140200 25368 143684 25396
rect 143678 25356 143684 25368
rect 143736 25356 143742 25408
rect 177350 25356 177356 25408
rect 177408 25396 177414 25408
rect 185722 25396 185728 25408
rect 177408 25368 185728 25396
rect 177408 25356 177414 25368
rect 185722 25356 185728 25368
rect 185780 25356 185786 25408
rect 143494 25328 143500 25340
rect 140108 25300 143500 25328
rect 143494 25288 143500 25300
rect 143552 25288 143558 25340
rect 177810 25288 177816 25340
rect 177868 25328 177874 25340
rect 185262 25328 185268 25340
rect 177868 25300 185268 25328
rect 177868 25288 177874 25300
rect 185262 25288 185268 25300
rect 185320 25288 185326 25340
rect 92710 25220 92716 25272
rect 92768 25260 92774 25272
rect 100990 25260 100996 25272
rect 92768 25232 100996 25260
rect 92768 25220 92774 25232
rect 100990 25220 100996 25232
rect 101048 25220 101054 25272
rect 138158 25220 138164 25272
rect 138216 25260 138222 25272
rect 143126 25260 143132 25272
rect 138216 25232 143132 25260
rect 138216 25220 138222 25232
rect 143126 25220 143132 25232
rect 143184 25220 143190 25272
rect 177718 25220 177724 25272
rect 177776 25260 177782 25272
rect 185814 25260 185820 25272
rect 177776 25232 185820 25260
rect 177776 25220 177782 25232
rect 185814 25220 185820 25232
rect 185872 25220 185878 25272
rect 134662 25016 134668 25068
rect 134720 25056 134726 25068
rect 134938 25056 134944 25068
rect 134720 25028 134944 25056
rect 134720 25016 134726 25028
rect 134938 25016 134944 25028
rect 134996 25016 135002 25068
rect 51218 24064 51224 24116
rect 51276 24104 51282 24116
rect 56094 24104 56100 24116
rect 51276 24076 56100 24104
rect 51276 24064 51282 24076
rect 56094 24064 56100 24076
rect 56152 24064 56158 24116
rect 135398 24064 135404 24116
rect 135456 24104 135462 24116
rect 143586 24104 143592 24116
rect 135456 24076 143592 24104
rect 135456 24064 135462 24076
rect 143586 24064 143592 24076
rect 143644 24064 143650 24116
rect 51126 23996 51132 24048
rect 51184 24036 51190 24048
rect 51184 24008 56784 24036
rect 51184 23996 51190 24008
rect 56756 23968 56784 24008
rect 135030 23996 135036 24048
rect 135088 24036 135094 24048
rect 143678 24036 143684 24048
rect 135088 24008 143684 24036
rect 135088 23996 135094 24008
rect 143678 23996 143684 24008
rect 143736 23996 143742 24048
rect 58210 23968 58216 23980
rect 56756 23940 58216 23968
rect 58210 23928 58216 23940
rect 58268 23928 58274 23980
rect 92802 23928 92808 23980
rect 92860 23968 92866 23980
rect 100990 23968 100996 23980
rect 92860 23940 100996 23968
rect 92860 23928 92866 23940
rect 100990 23928 100996 23940
rect 101048 23928 101054 23980
rect 177626 23928 177632 23980
rect 177684 23968 177690 23980
rect 185170 23968 185176 23980
rect 177684 23940 185176 23968
rect 177684 23928 177690 23940
rect 185170 23928 185176 23940
rect 185228 23928 185234 23980
rect 92710 23860 92716 23912
rect 92768 23900 92774 23912
rect 101082 23900 101088 23912
rect 92768 23872 101088 23900
rect 92768 23860 92774 23872
rect 101082 23860 101088 23872
rect 101140 23860 101146 23912
rect 177350 23860 177356 23912
rect 177408 23900 177414 23912
rect 185262 23900 185268 23912
rect 177408 23872 185268 23900
rect 177408 23860 177414 23872
rect 185262 23860 185268 23872
rect 185320 23860 185326 23912
rect 56094 23452 56100 23504
rect 56152 23492 56158 23504
rect 58302 23492 58308 23504
rect 56152 23464 58308 23492
rect 56152 23452 56158 23464
rect 58302 23452 58308 23464
rect 58360 23452 58366 23504
rect 97678 23112 97684 23164
rect 97736 23152 97742 23164
rect 100990 23152 100996 23164
rect 97736 23124 100996 23152
rect 97736 23112 97742 23124
rect 100990 23112 100996 23124
rect 101048 23112 101054 23164
rect 135030 22908 135036 22960
rect 135088 22948 135094 22960
rect 135306 22948 135312 22960
rect 135088 22920 135312 22948
rect 135088 22908 135094 22920
rect 135306 22908 135312 22920
rect 135364 22908 135370 22960
rect 135306 22772 135312 22824
rect 135364 22812 135370 22824
rect 136870 22812 136876 22824
rect 135364 22784 136876 22812
rect 135364 22772 135370 22784
rect 136870 22772 136876 22784
rect 136928 22772 136934 22824
rect 185262 22812 185268 22824
rect 182244 22784 185268 22812
rect 51218 22704 51224 22756
rect 51276 22744 51282 22756
rect 55726 22744 55732 22756
rect 51276 22716 55732 22744
rect 51276 22704 51282 22716
rect 55726 22704 55732 22716
rect 55784 22704 55790 22756
rect 134478 22704 134484 22756
rect 134536 22744 134542 22756
rect 134536 22716 139768 22744
rect 134536 22704 134542 22716
rect 50390 22636 50396 22688
rect 50448 22676 50454 22688
rect 50448 22648 56784 22676
rect 50448 22636 50454 22648
rect 56756 22608 56784 22648
rect 98138 22636 98144 22688
rect 98196 22676 98202 22688
rect 101082 22676 101088 22688
rect 98196 22648 101088 22676
rect 98196 22636 98202 22648
rect 101082 22636 101088 22648
rect 101140 22636 101146 22688
rect 135398 22636 135404 22688
rect 135456 22676 135462 22688
rect 135456 22648 139676 22676
rect 135456 22636 135462 22648
rect 58210 22608 58216 22620
rect 56756 22580 58216 22608
rect 58210 22568 58216 22580
rect 58268 22568 58274 22620
rect 90410 22568 90416 22620
rect 90468 22608 90474 22620
rect 100990 22608 100996 22620
rect 90468 22580 100996 22608
rect 90468 22568 90474 22580
rect 100990 22568 100996 22580
rect 101048 22568 101054 22620
rect 96114 22500 96120 22552
rect 96172 22540 96178 22552
rect 101082 22540 101088 22552
rect 96172 22512 101088 22540
rect 96172 22500 96178 22512
rect 101082 22500 101088 22512
rect 101140 22500 101146 22552
rect 139648 22540 139676 22648
rect 139740 22608 139768 22716
rect 142758 22608 142764 22620
rect 139740 22580 142764 22608
rect 142758 22568 142764 22580
rect 142816 22568 142822 22620
rect 177626 22568 177632 22620
rect 177684 22608 177690 22620
rect 182244 22608 182272 22784
rect 185262 22772 185268 22784
rect 185320 22772 185326 22824
rect 185170 22676 185176 22688
rect 177684 22580 182272 22608
rect 182336 22648 185176 22676
rect 177684 22568 177690 22580
rect 143310 22540 143316 22552
rect 139648 22512 143316 22540
rect 143310 22500 143316 22512
rect 143368 22500 143374 22552
rect 177718 22500 177724 22552
rect 177776 22540 177782 22552
rect 182336 22540 182364 22648
rect 185170 22636 185176 22648
rect 185228 22636 185234 22688
rect 177776 22512 182364 22540
rect 177776 22500 177782 22512
rect 92802 22432 92808 22484
rect 92860 22472 92866 22484
rect 98138 22472 98144 22484
rect 92860 22444 98144 22472
rect 92860 22432 92866 22444
rect 98138 22432 98144 22444
rect 98196 22432 98202 22484
rect 174406 22432 174412 22484
rect 174464 22472 174470 22484
rect 185170 22472 185176 22484
rect 174464 22444 185176 22472
rect 174464 22432 174470 22444
rect 185170 22432 185176 22444
rect 185228 22432 185234 22484
rect 92710 22364 92716 22416
rect 92768 22404 92774 22416
rect 97678 22404 97684 22416
rect 92768 22376 97684 22404
rect 92768 22364 92774 22376
rect 97678 22364 97684 22376
rect 97736 22364 97742 22416
rect 55726 22160 55732 22212
rect 55784 22200 55790 22212
rect 58302 22200 58308 22212
rect 55784 22172 58308 22200
rect 55784 22160 55790 22172
rect 58302 22160 58308 22172
rect 58360 22160 58366 22212
rect 50574 21276 50580 21328
rect 50632 21316 50638 21328
rect 50632 21288 56784 21316
rect 50632 21276 50638 21288
rect 56756 21248 56784 21288
rect 58210 21248 58216 21260
rect 56756 21220 58216 21248
rect 58210 21208 58216 21220
rect 58268 21208 58274 21260
rect 92710 21208 92716 21260
rect 92768 21248 92774 21260
rect 101174 21248 101180 21260
rect 92768 21220 101180 21248
rect 92768 21208 92774 21220
rect 101174 21208 101180 21220
rect 101232 21208 101238 21260
rect 136870 21208 136876 21260
rect 136928 21248 136934 21260
rect 143678 21248 143684 21260
rect 136928 21220 143684 21248
rect 136928 21208 136934 21220
rect 143678 21208 143684 21220
rect 143736 21208 143742 21260
rect 177718 21208 177724 21260
rect 177776 21248 177782 21260
rect 185262 21248 185268 21260
rect 177776 21220 185268 21248
rect 177776 21208 177782 21220
rect 185262 21208 185268 21220
rect 185320 21208 185326 21260
rect 93354 19780 93360 19832
rect 93412 19820 93418 19832
rect 101082 19820 101088 19832
rect 93412 19792 101088 19820
rect 93412 19780 93418 19792
rect 101082 19780 101088 19792
rect 101140 19780 101146 19832
rect 176154 19780 176160 19832
rect 176212 19820 176218 19832
rect 185262 19820 185268 19832
rect 176212 19792 185268 19820
rect 176212 19780 176218 19792
rect 185262 19780 185268 19792
rect 185320 19780 185326 19832
rect 94734 19712 94740 19764
rect 94792 19752 94798 19764
rect 100990 19752 100996 19764
rect 94792 19724 100996 19752
rect 94792 19712 94798 19724
rect 100990 19712 100996 19724
rect 101048 19712 101054 19764
rect 177534 19712 177540 19764
rect 177592 19752 177598 19764
rect 185170 19752 185176 19764
rect 177592 19724 185176 19752
rect 177592 19712 177598 19724
rect 185170 19712 185176 19724
rect 185228 19712 185234 19764
rect 18098 18420 18104 18472
rect 18156 18460 18162 18472
rect 68238 18460 68244 18472
rect 18156 18432 68244 18460
rect 18156 18420 18162 18432
rect 68238 18420 68244 18432
rect 68296 18420 68302 18472
rect 69802 18420 69808 18472
rect 69860 18460 69866 18472
rect 106694 18460 106700 18472
rect 69860 18432 106700 18460
rect 69860 18420 69866 18432
rect 106694 18420 106700 18432
rect 106752 18460 106758 18472
rect 153522 18460 153528 18472
rect 106752 18432 153528 18460
rect 106752 18420 106758 18432
rect 153522 18420 153528 18432
rect 153580 18460 153586 18472
rect 192530 18460 192536 18472
rect 153580 18432 192536 18460
rect 153580 18420 153586 18432
rect 192530 18420 192536 18432
rect 192588 18460 192594 18472
rect 211390 18460 211396 18472
rect 192588 18432 211396 18460
rect 192588 18420 192594 18432
rect 211390 18420 211396 18432
rect 211448 18420 211454 18472
rect 53978 18352 53984 18404
rect 54036 18392 54042 18404
rect 69820 18392 69848 18420
rect 54036 18364 69848 18392
rect 54036 18352 54042 18364
rect 71918 18352 71924 18404
rect 71976 18392 71982 18404
rect 100254 18392 100260 18404
rect 71976 18364 100260 18392
rect 71976 18352 71982 18364
rect 100254 18352 100260 18364
rect 100312 18352 100318 18404
rect 112214 18352 112220 18404
rect 112272 18392 112278 18404
rect 152234 18392 152240 18404
rect 112272 18364 152240 18392
rect 112272 18352 112278 18364
rect 152234 18352 152240 18364
rect 152292 18352 152298 18404
rect 60786 18284 60792 18336
rect 60844 18324 60850 18336
rect 60844 18296 76104 18324
rect 60844 18284 60850 18296
rect 54806 18216 54812 18268
rect 54864 18256 54870 18268
rect 75969 18259 76027 18265
rect 75969 18256 75981 18259
rect 54864 18228 75981 18256
rect 54864 18216 54870 18228
rect 75969 18225 75981 18228
rect 76015 18225 76027 18259
rect 76076 18256 76104 18296
rect 76150 18284 76156 18336
rect 76208 18324 76214 18336
rect 80658 18324 80664 18336
rect 76208 18296 80664 18324
rect 76208 18284 76214 18296
rect 80658 18284 80664 18296
rect 80716 18284 80722 18336
rect 88478 18284 88484 18336
rect 88536 18324 88542 18336
rect 92710 18324 92716 18336
rect 88536 18296 92716 18324
rect 88536 18284 88542 18296
rect 92710 18284 92716 18296
rect 92768 18284 92774 18336
rect 156006 18284 156012 18336
rect 156064 18324 156070 18336
rect 157570 18324 157576 18336
rect 156064 18296 157576 18324
rect 156064 18284 156070 18296
rect 157570 18284 157576 18296
rect 157628 18284 157634 18336
rect 161894 18284 161900 18336
rect 161952 18324 161958 18336
rect 162630 18324 162636 18336
rect 161952 18296 162636 18324
rect 161952 18284 161958 18296
rect 162630 18284 162636 18296
rect 162688 18284 162694 18336
rect 163090 18284 163096 18336
rect 163148 18324 163154 18336
rect 163642 18324 163648 18336
rect 163148 18296 163648 18324
rect 163148 18284 163154 18296
rect 163642 18284 163648 18296
rect 163700 18284 163706 18336
rect 167138 18284 167144 18336
rect 167196 18324 167202 18336
rect 167782 18324 167788 18336
rect 167196 18296 167788 18324
rect 167196 18284 167202 18296
rect 167782 18284 167788 18296
rect 167840 18284 167846 18336
rect 171370 18284 171376 18336
rect 171428 18324 171434 18336
rect 171922 18324 171928 18336
rect 171428 18296 171928 18324
rect 171428 18284 171434 18296
rect 171922 18284 171928 18296
rect 171980 18284 171986 18336
rect 81670 18256 81676 18268
rect 76076 18228 81676 18256
rect 75969 18219 76027 18225
rect 81670 18216 81676 18228
rect 81728 18216 81734 18268
rect 166310 18216 166316 18268
rect 166368 18256 166374 18268
rect 168518 18256 168524 18268
rect 166368 18228 168524 18256
rect 166368 18216 166374 18228
rect 168518 18216 168524 18228
rect 168576 18216 168582 18268
rect 42846 18148 42852 18200
rect 42904 18188 42910 18200
rect 72378 18188 72384 18200
rect 42904 18160 72384 18188
rect 42904 18148 42910 18160
rect 72378 18148 72384 18160
rect 72436 18148 72442 18200
rect 48826 18080 48832 18132
rect 48884 18120 48890 18132
rect 83786 18120 83792 18132
rect 48884 18092 83792 18120
rect 48884 18080 48890 18092
rect 83786 18080 83792 18092
rect 83844 18080 83850 18132
rect 30794 18012 30800 18064
rect 30852 18052 30858 18064
rect 74770 18052 74776 18064
rect 30852 18024 74776 18052
rect 30852 18012 30858 18024
rect 74770 18012 74776 18024
rect 74828 18012 74834 18064
rect 75969 18055 76027 18061
rect 75969 18021 75981 18055
rect 76015 18052 76027 18055
rect 83050 18052 83056 18064
rect 76015 18024 83056 18052
rect 76015 18021 76027 18024
rect 75969 18015 76027 18021
rect 83050 18012 83056 18024
rect 83108 18012 83114 18064
rect 36774 17944 36780 17996
rect 36832 17984 36838 17996
rect 73390 17984 73396 17996
rect 36832 17956 73396 17984
rect 36832 17944 36838 17956
rect 73390 17944 73396 17956
rect 73448 17944 73454 17996
rect 138802 17944 138808 17996
rect 138860 17984 138866 17996
rect 158490 17984 158496 17996
rect 138860 17956 158496 17984
rect 138860 17944 138866 17956
rect 158490 17944 158496 17956
rect 158548 17944 158554 17996
rect 165298 17944 165304 17996
rect 165356 17984 165362 17996
rect 168978 17984 168984 17996
rect 165356 17956 168984 17984
rect 165356 17944 165362 17956
rect 168978 17944 168984 17956
rect 169036 17944 169042 17996
rect 24814 17876 24820 17928
rect 24872 17916 24878 17928
rect 75506 17916 75512 17928
rect 24872 17888 75512 17916
rect 24872 17876 24878 17888
rect 75506 17876 75512 17888
rect 75564 17876 75570 17928
rect 132822 17876 132828 17928
rect 132880 17916 132886 17928
rect 159502 17916 159508 17928
rect 132880 17888 159508 17916
rect 132880 17876 132886 17888
rect 159502 17876 159508 17888
rect 159560 17876 159566 17928
rect 18834 17808 18840 17860
rect 18892 17848 18898 17860
rect 76518 17848 76524 17860
rect 18892 17820 76524 17848
rect 18892 17808 18898 17820
rect 76518 17808 76524 17820
rect 76576 17808 76582 17860
rect 126842 17808 126848 17860
rect 126900 17848 126906 17860
rect 160514 17848 160520 17860
rect 126900 17820 160520 17848
rect 126900 17808 126906 17820
rect 160514 17808 160520 17820
rect 160572 17808 160578 17860
rect 12854 17740 12860 17792
rect 12912 17780 12918 17792
rect 77530 17780 77536 17792
rect 12912 17752 77536 17780
rect 12912 17740 12918 17752
rect 77530 17740 77536 17752
rect 77588 17740 77594 17792
rect 120862 17740 120868 17792
rect 120920 17780 120926 17792
rect 161710 17780 161716 17792
rect 120920 17752 161716 17780
rect 120920 17740 120926 17752
rect 161710 17740 161716 17752
rect 161768 17740 161774 17792
rect 89582 17536 89588 17588
rect 89640 17576 89646 17588
rect 90778 17576 90784 17588
rect 89640 17548 90784 17576
rect 89640 17536 89646 17548
rect 90778 17536 90784 17548
rect 90836 17536 90842 17588
rect 169990 17536 169996 17588
rect 170048 17576 170054 17588
rect 170910 17576 170916 17588
rect 170048 17548 170916 17576
rect 170048 17536 170054 17548
rect 170910 17536 170916 17548
rect 170968 17536 170974 17588
rect 67778 17060 67784 17112
rect 67836 17100 67842 17112
rect 117826 17100 117832 17112
rect 67836 17072 117832 17100
rect 67836 17060 67842 17072
rect 117826 17060 117832 17072
rect 117884 17060 117890 17112
rect 151866 17060 151872 17112
rect 151924 17100 151930 17112
rect 211114 17100 211120 17112
rect 151924 17072 211120 17100
rect 151924 17060 151930 17072
rect 211114 17060 211120 17072
rect 211172 17060 211178 17112
rect 180846 12884 180852 12896
rect 173044 12856 180852 12884
rect 163090 12708 163096 12760
rect 163148 12748 163154 12760
rect 173044 12748 173072 12856
rect 180846 12844 180852 12856
rect 180904 12844 180910 12896
rect 174866 12748 174872 12760
rect 163148 12720 173072 12748
rect 173136 12720 174872 12748
rect 163148 12708 163154 12720
rect 168978 12640 168984 12692
rect 169036 12680 169042 12692
rect 173136 12680 173164 12720
rect 174866 12708 174872 12720
rect 174924 12708 174930 12760
rect 169036 12652 173164 12680
rect 169036 12640 169042 12652
rect 174130 12640 174136 12692
rect 174188 12680 174194 12692
rect 192806 12680 192812 12692
rect 174188 12652 192812 12680
rect 174188 12640 174194 12652
rect 192806 12640 192812 12652
rect 192864 12640 192870 12692
rect 172750 12572 172756 12624
rect 172808 12612 172814 12624
rect 198786 12612 198792 12624
rect 172808 12584 198792 12612
rect 172808 12572 172814 12584
rect 198786 12572 198792 12584
rect 198844 12572 198850 12624
rect 161894 12504 161900 12556
rect 161952 12544 161958 12556
rect 186826 12544 186832 12556
rect 161952 12516 186832 12544
rect 161952 12504 161958 12516
rect 186826 12504 186832 12516
rect 186884 12504 186890 12556
rect 92710 12436 92716 12488
rect 92768 12476 92774 12488
rect 96850 12476 96856 12488
rect 92768 12448 96856 12476
rect 92768 12436 92774 12448
rect 96850 12436 96856 12448
rect 96908 12436 96914 12488
rect 171370 12436 171376 12488
rect 171428 12476 171434 12488
rect 204858 12476 204864 12488
rect 171428 12448 204864 12476
rect 171428 12436 171434 12448
rect 204858 12436 204864 12448
rect 204916 12436 204922 12488
rect 87282 12368 87288 12420
rect 87340 12408 87346 12420
rect 102830 12408 102836 12420
rect 87340 12380 102836 12408
rect 87340 12368 87346 12380
rect 102830 12368 102836 12380
rect 102888 12368 102894 12420
rect 168610 12368 168616 12420
rect 168668 12408 168674 12420
rect 168668 12380 168748 12408
rect 168668 12368 168674 12380
rect 72838 12300 72844 12352
rect 72896 12340 72902 12352
rect 79094 12340 79100 12352
rect 72896 12312 79100 12340
rect 72896 12300 72902 12312
rect 79094 12300 79100 12312
rect 79152 12300 79158 12352
rect 85810 12300 85816 12352
rect 85868 12340 85874 12352
rect 108810 12340 108816 12352
rect 85868 12312 108816 12340
rect 85868 12300 85874 12312
rect 108810 12300 108816 12312
rect 108868 12300 108874 12352
rect 150854 12300 150860 12352
rect 150912 12340 150918 12352
rect 156098 12340 156104 12352
rect 150912 12312 156104 12340
rect 150912 12300 150918 12312
rect 156098 12300 156104 12312
rect 156156 12300 156162 12352
rect 162814 12300 162820 12352
rect 162872 12340 162878 12352
rect 165850 12340 165856 12352
rect 162872 12312 165856 12340
rect 162872 12300 162878 12312
rect 165850 12300 165856 12312
rect 165908 12300 165914 12352
rect 66858 12232 66864 12284
rect 66916 12272 66922 12284
rect 76150 12272 76156 12284
rect 66916 12244 76156 12272
rect 66916 12232 66922 12244
rect 76150 12232 76156 12244
rect 76208 12232 76214 12284
rect 84430 12232 84436 12284
rect 84488 12272 84494 12284
rect 114790 12272 114796 12284
rect 84488 12244 114796 12272
rect 84488 12232 84494 12244
rect 114790 12232 114796 12244
rect 114848 12232 114854 12284
rect 144782 12232 144788 12284
rect 144840 12272 144846 12284
rect 156006 12272 156012 12284
rect 144840 12244 156012 12272
rect 144840 12232 144846 12244
rect 156006 12232 156012 12244
rect 156064 12232 156070 12284
rect 156834 12232 156840 12284
rect 156892 12272 156898 12284
rect 167138 12272 167144 12284
rect 156892 12244 167144 12272
rect 156892 12232 156898 12244
rect 167138 12232 167144 12244
rect 167196 12232 167202 12284
rect 168720 12272 168748 12380
rect 169990 12368 169996 12420
rect 170048 12408 170054 12420
rect 210838 12408 210844 12420
rect 170048 12380 210844 12408
rect 170048 12368 170054 12380
rect 210838 12368 210844 12380
rect 210896 12368 210902 12420
rect 170082 12300 170088 12352
rect 170140 12340 170146 12352
rect 216818 12340 216824 12352
rect 170140 12312 216824 12340
rect 170140 12300 170146 12312
rect 216818 12300 216824 12312
rect 216876 12300 216882 12352
rect 222798 12272 222804 12284
rect 168720 12244 222804 12272
rect 222798 12232 222804 12244
rect 222856 12232 222862 12284
rect 84798 11824 84804 11876
rect 84856 11864 84862 11876
rect 89858 11864 89864 11876
rect 84856 11836 89864 11864
rect 84856 11824 84862 11836
rect 89858 11824 89864 11836
rect 89916 11824 89922 11876
<< via1 >>
rect 99616 244248 99668 244300
rect 99800 244248 99852 244300
rect 89864 241324 89916 241376
rect 171836 241324 171888 241376
rect 174044 241324 174096 241376
rect 207808 241324 207860 241376
rect 27856 241120 27908 241172
rect 29144 241120 29196 241172
rect 63828 241120 63880 241172
rect 65024 241120 65076 241172
rect 22704 236632 22756 236684
rect 49844 236632 49896 236684
rect 72844 236632 72896 236684
rect 121420 236632 121472 236684
rect 39448 236564 39500 236616
rect 96120 236564 96172 236616
rect 29144 235884 29196 235936
rect 82228 235884 82280 235936
rect 86184 235884 86236 235936
rect 99616 235884 99668 235936
rect 135864 235884 135916 235936
rect 169536 235884 169588 235936
rect 65024 235816 65076 235868
rect 166224 235816 166276 235868
rect 47268 235272 47320 235324
rect 65576 235272 65628 235324
rect 49844 235204 49896 235256
rect 62540 235204 62592 235256
rect 107436 235340 107488 235392
rect 139452 235340 139504 235392
rect 114428 235204 114480 235256
rect 159508 235204 159560 235256
rect 173492 235204 173544 235256
rect 174044 235204 174096 235256
rect 28224 235136 28276 235188
rect 75512 235136 75564 235188
rect 146536 235136 146588 235188
rect 156840 235136 156892 235188
rect 215628 235136 215680 235188
rect 107436 235000 107488 235052
rect 134760 234499 134812 234508
rect 134760 234465 134769 234499
rect 134769 234465 134803 234499
rect 134803 234465 134812 234499
rect 134760 234456 134812 234465
rect 51224 233912 51276 233964
rect 58124 233912 58176 233964
rect 90232 233844 90284 233896
rect 101180 233844 101232 233896
rect 134760 233844 134812 233896
rect 142304 233844 142356 233896
rect 180300 233844 180352 233896
rect 185176 233844 185228 233896
rect 13320 233776 13372 233828
rect 185268 233776 185320 233828
rect 92716 233028 92768 233080
rect 101364 233028 101416 233080
rect 177724 233028 177776 233080
rect 185176 233028 185228 233080
rect 134760 232688 134812 232740
rect 142212 232688 142264 232740
rect 134852 232620 134904 232672
rect 142304 232620 142356 232672
rect 51224 232552 51276 232604
rect 58032 232552 58084 232604
rect 50028 232416 50080 232468
rect 58124 232416 58176 232468
rect 94004 232348 94056 232400
rect 101732 232416 101784 232468
rect 177724 232348 177776 232400
rect 185176 232416 185228 232468
rect 92716 231668 92768 231720
rect 101272 231668 101324 231720
rect 177724 231668 177776 231720
rect 185176 231668 185228 231720
rect 134760 231464 134812 231516
rect 139636 231464 139688 231516
rect 50120 231124 50172 231176
rect 56468 231124 56520 231176
rect 50764 231056 50816 231108
rect 51224 230988 51276 231040
rect 52696 230988 52748 231040
rect 98880 231056 98932 231108
rect 101456 231056 101508 231108
rect 134760 231056 134812 231108
rect 136876 231056 136928 231108
rect 58216 230920 58268 230972
rect 92716 230920 92768 230972
rect 101732 230988 101784 231040
rect 134852 230988 134904 231040
rect 93728 230852 93780 230904
rect 98880 230852 98932 230904
rect 143684 230852 143736 230904
rect 177724 230852 177776 230904
rect 185268 231056 185320 231108
rect 217560 231056 217612 231108
rect 222344 231056 222396 231108
rect 183704 230988 183756 231040
rect 185176 230988 185228 231040
rect 56468 230580 56520 230632
rect 58216 230580 58268 230632
rect 139636 230580 139688 230632
rect 142948 230580 143000 230632
rect 177724 230580 177776 230632
rect 183704 230580 183756 230632
rect 134300 229968 134352 230020
rect 139636 229968 139688 230020
rect 51224 229832 51276 229884
rect 56468 229832 56520 229884
rect 51132 229696 51184 229748
rect 56192 229696 56244 229748
rect 134392 229628 134444 229680
rect 52696 229560 52748 229612
rect 58216 229560 58268 229612
rect 92716 229560 92768 229612
rect 101732 229560 101784 229612
rect 143592 229560 143644 229612
rect 177632 229560 177684 229612
rect 185176 229560 185228 229612
rect 92808 229492 92860 229544
rect 101548 229492 101600 229544
rect 136876 229492 136928 229544
rect 143684 229492 143736 229544
rect 177724 229492 177776 229544
rect 185268 229492 185320 229544
rect 139636 229424 139688 229476
rect 143500 229424 143552 229476
rect 56192 229288 56244 229340
rect 58216 229288 58268 229340
rect 56468 229016 56520 229068
rect 58308 229016 58360 229068
rect 92716 228880 92768 228932
rect 101732 228880 101784 228932
rect 176988 228880 177040 228932
rect 185176 228880 185228 228932
rect 51040 228404 51092 228456
rect 52696 228404 52748 228456
rect 134392 228404 134444 228456
rect 51224 228336 51276 228388
rect 55456 228336 55508 228388
rect 51132 228268 51184 228320
rect 58216 228200 58268 228252
rect 93176 228200 93228 228252
rect 101456 228336 101508 228388
rect 134760 228336 134812 228388
rect 92716 228132 92768 228184
rect 101732 228268 101784 228320
rect 134852 228268 134904 228320
rect 136876 228268 136928 228320
rect 143684 228200 143736 228252
rect 177724 228200 177776 228252
rect 185268 228336 185320 228388
rect 143316 228132 143368 228184
rect 177632 228132 177684 228184
rect 185176 228268 185228 228320
rect 55456 227860 55508 227912
rect 58308 227860 58360 227912
rect 50764 226840 50816 226892
rect 55916 226840 55968 226892
rect 134760 226840 134812 226892
rect 52696 226772 52748 226824
rect 58216 226772 58268 226824
rect 92716 226772 92768 226824
rect 101364 226772 101416 226824
rect 143316 226772 143368 226824
rect 177172 226772 177224 226824
rect 185176 226772 185228 226824
rect 92808 226704 92860 226756
rect 101456 226704 101508 226756
rect 136876 226704 136928 226756
rect 143684 226704 143736 226756
rect 177724 226704 177776 226756
rect 185268 226704 185320 226756
rect 55916 226364 55968 226416
rect 58216 226364 58268 226416
rect 51224 225548 51276 225600
rect 58308 225548 58360 225600
rect 134392 225548 134444 225600
rect 143316 225548 143368 225600
rect 50028 225480 50080 225532
rect 58400 225480 58452 225532
rect 134760 225480 134812 225532
rect 142580 225480 142632 225532
rect 51316 225412 51368 225464
rect 58216 225412 58268 225464
rect 93728 225412 93780 225464
rect 101548 225412 101600 225464
rect 135496 225412 135548 225464
rect 143684 225412 143736 225464
rect 177724 225412 177776 225464
rect 185360 225412 185412 225464
rect 92808 225344 92860 225396
rect 101824 225344 101876 225396
rect 177172 225344 177224 225396
rect 185176 225344 185228 225396
rect 92716 225276 92768 225328
rect 101640 225276 101692 225328
rect 177724 225276 177776 225328
rect 185268 225276 185320 225328
rect 51132 224392 51184 224444
rect 56744 224392 56796 224444
rect 51132 224256 51184 224308
rect 52696 224256 52748 224308
rect 134668 224256 134720 224308
rect 135404 224188 135456 224240
rect 136876 224188 136928 224240
rect 51224 224120 51276 224172
rect 134300 224120 134352 224172
rect 58216 224052 58268 224104
rect 93912 224052 93964 224104
rect 100996 224052 101048 224104
rect 56744 223984 56796 224036
rect 58308 223984 58360 224036
rect 93728 223984 93780 224036
rect 101088 223984 101140 224036
rect 134760 224027 134812 224036
rect 134760 223993 134769 224027
rect 134769 223993 134803 224027
rect 134803 223993 134812 224027
rect 134760 223984 134812 223993
rect 143684 224052 143736 224104
rect 177724 224052 177776 224104
rect 185268 224052 185320 224104
rect 143316 223984 143368 224036
rect 177632 223984 177684 224036
rect 185176 223984 185228 224036
rect 51132 223032 51184 223084
rect 52788 223032 52840 223084
rect 134484 223032 134536 223084
rect 136968 223032 137020 223084
rect 51224 222896 51276 222948
rect 55824 222896 55876 222948
rect 135404 222760 135456 222812
rect 52696 222692 52748 222744
rect 58216 222692 58268 222744
rect 92716 222692 92768 222744
rect 101456 222692 101508 222744
rect 143316 222692 143368 222744
rect 177632 222692 177684 222744
rect 185176 222692 185228 222744
rect 92992 222624 93044 222676
rect 101364 222624 101416 222676
rect 136876 222624 136928 222676
rect 143684 222624 143736 222676
rect 177724 222624 177776 222676
rect 185268 222624 185320 222676
rect 55824 222284 55876 222336
rect 58308 222284 58360 222336
rect 51224 221672 51276 221724
rect 56008 221672 56060 221724
rect 134852 221672 134904 221724
rect 139636 221672 139688 221724
rect 51132 221400 51184 221452
rect 56468 221400 56520 221452
rect 134668 221400 134720 221452
rect 139728 221400 139780 221452
rect 51224 221332 51276 221384
rect 52696 221332 52748 221384
rect 135404 221332 135456 221384
rect 136876 221332 136928 221384
rect 52788 221264 52840 221316
rect 58216 221264 58268 221316
rect 92808 221264 92860 221316
rect 101548 221264 101600 221316
rect 136968 221264 137020 221316
rect 143684 221264 143736 221316
rect 177172 221264 177224 221316
rect 185176 221264 185228 221316
rect 93728 221196 93780 221248
rect 101640 221196 101692 221248
rect 177632 221196 177684 221248
rect 185268 221196 185320 221248
rect 92716 221128 92768 221180
rect 100904 221128 100956 221180
rect 177724 221128 177776 221180
rect 185084 221128 185136 221180
rect 56008 221060 56060 221112
rect 58216 221060 58268 221112
rect 139636 220924 139688 220976
rect 143316 220924 143368 220976
rect 56468 220652 56520 220704
rect 58308 220652 58360 220704
rect 139728 220584 139780 220636
rect 143684 220584 143736 220636
rect 135312 220108 135364 220160
rect 138164 220108 138216 220160
rect 51132 220040 51184 220092
rect 52788 220040 52840 220092
rect 51224 219972 51276 220024
rect 55824 219972 55876 220024
rect 135404 219972 135456 220024
rect 52696 219904 52748 219956
rect 58216 219904 58268 219956
rect 93728 219904 93780 219956
rect 101824 219904 101876 219956
rect 143132 219904 143184 219956
rect 177172 219904 177224 219956
rect 185176 219904 185228 219956
rect 93912 219836 93964 219888
rect 101272 219836 101324 219888
rect 136876 219836 136928 219888
rect 143684 219836 143736 219888
rect 177724 219836 177776 219888
rect 185360 219836 185412 219888
rect 55824 219292 55876 219344
rect 58308 219292 58360 219344
rect 51224 218816 51276 218868
rect 53340 218816 53392 218868
rect 135036 218816 135088 218868
rect 137520 218816 137572 218868
rect 51224 218680 51276 218732
rect 52788 218680 52840 218732
rect 135404 218680 135456 218732
rect 50856 218612 50908 218664
rect 55456 218612 55508 218664
rect 93544 218612 93596 218664
rect 101732 218612 101784 218664
rect 135312 218612 135364 218664
rect 137980 218612 138032 218664
rect 52696 218544 52748 218596
rect 58216 218544 58268 218596
rect 93728 218544 93780 218596
rect 101364 218544 101416 218596
rect 178000 218612 178052 218664
rect 185176 218612 185228 218664
rect 143500 218544 143552 218596
rect 177172 218544 177224 218596
rect 185820 218544 185872 218596
rect 93176 218476 93228 218528
rect 100904 218476 100956 218528
rect 138164 218476 138216 218528
rect 143684 218476 143736 218528
rect 177724 218476 177776 218528
rect 185084 218476 185136 218528
rect 55456 218000 55508 218052
rect 58216 218000 58268 218052
rect 51224 217320 51276 217372
rect 52880 217320 52932 217372
rect 134484 217320 134536 217372
rect 137612 217320 137664 217372
rect 135404 217252 135456 217304
rect 137704 217252 137756 217304
rect 50764 217184 50816 217236
rect 52696 217184 52748 217236
rect 53340 217116 53392 217168
rect 58216 217116 58268 217168
rect 92716 217116 92768 217168
rect 101180 217184 101232 217236
rect 137520 217116 137572 217168
rect 143684 217116 143736 217168
rect 177724 217116 177776 217168
rect 185176 217184 185228 217236
rect 52788 217048 52840 217100
rect 58308 217048 58360 217100
rect 137980 217048 138032 217100
rect 143132 217048 143184 217100
rect 51132 215824 51184 215876
rect 56468 215824 56520 215876
rect 135404 215824 135456 215876
rect 52696 215756 52748 215808
rect 58216 215756 58268 215808
rect 93544 215756 93596 215808
rect 101364 215756 101416 215808
rect 143500 215756 143552 215808
rect 177172 215756 177224 215808
rect 185176 215756 185228 215808
rect 52880 215688 52932 215740
rect 58308 215688 58360 215740
rect 92716 215688 92768 215740
rect 100812 215688 100864 215740
rect 137704 215688 137756 215740
rect 143132 215688 143184 215740
rect 177724 215688 177776 215740
rect 184992 215688 185044 215740
rect 92808 215620 92860 215672
rect 100904 215620 100956 215672
rect 137612 215620 137664 215672
rect 142948 215620 143000 215672
rect 177632 215620 177684 215672
rect 185084 215620 185136 215672
rect 56468 215144 56520 215196
rect 58216 215144 58268 215196
rect 50396 214872 50448 214924
rect 52788 214872 52840 214924
rect 134852 214872 134904 214924
rect 137612 214872 137664 214924
rect 51132 214532 51184 214584
rect 52696 214532 52748 214584
rect 135312 214532 135364 214584
rect 136876 214532 136928 214584
rect 51224 214464 51276 214516
rect 58308 214464 58360 214516
rect 135404 214464 135456 214516
rect 143684 214464 143736 214516
rect 51316 214396 51368 214448
rect 58216 214396 58268 214448
rect 93360 214396 93412 214448
rect 100996 214396 101048 214448
rect 134760 214396 134812 214448
rect 135312 214396 135364 214448
rect 135496 214396 135548 214448
rect 142948 214396 143000 214448
rect 177632 214396 177684 214448
rect 185176 214396 185228 214448
rect 92716 214328 92768 214380
rect 100720 214328 100772 214380
rect 177724 214328 177776 214380
rect 184808 214328 184860 214380
rect 134484 213512 134536 213564
rect 137060 213512 137112 213564
rect 51224 213376 51276 213428
rect 52880 213376 52932 213428
rect 50396 213104 50448 213156
rect 52972 213104 53024 213156
rect 134484 213104 134536 213156
rect 136968 213104 137020 213156
rect 52788 213036 52840 213088
rect 58216 213036 58268 213088
rect 93360 213036 93412 213088
rect 100996 213036 101048 213088
rect 137612 213036 137664 213088
rect 143684 213036 143736 213088
rect 177172 213036 177224 213088
rect 185268 213036 185320 213088
rect 52696 212968 52748 213020
rect 58308 212968 58360 213020
rect 92716 212968 92768 213020
rect 100812 212968 100864 213020
rect 136876 212968 136928 213020
rect 143500 212968 143552 213020
rect 177724 212968 177776 213020
rect 184900 212968 184952 213020
rect 51132 212016 51184 212068
rect 52696 212016 52748 212068
rect 97500 211948 97552 212000
rect 100996 211948 101048 212000
rect 134484 211880 134536 211932
rect 139636 211880 139688 211932
rect 51224 211744 51276 211796
rect 56284 211744 56336 211796
rect 134668 211744 134720 211796
rect 136876 211744 136928 211796
rect 181772 211676 181824 211728
rect 185176 211676 185228 211728
rect 52972 211608 53024 211660
rect 58216 211608 58268 211660
rect 92808 211608 92860 211660
rect 100904 211608 100956 211660
rect 137060 211608 137112 211660
rect 143684 211608 143736 211660
rect 177724 211608 177776 211660
rect 184992 211608 185044 211660
rect 52880 211540 52932 211592
rect 58308 211540 58360 211592
rect 92716 211540 92768 211592
rect 100720 211540 100772 211592
rect 177172 211540 177224 211592
rect 185084 211540 185136 211592
rect 92900 211472 92952 211524
rect 97500 211472 97552 211524
rect 136968 211336 137020 211388
rect 143684 211336 143736 211388
rect 56284 210996 56336 211048
rect 58400 210996 58452 211048
rect 139636 210928 139688 210980
rect 143592 210928 143644 210980
rect 177724 210792 177776 210844
rect 181772 210792 181824 210844
rect 51224 210520 51276 210572
rect 56100 210520 56152 210572
rect 94004 210384 94056 210436
rect 101088 210384 101140 210436
rect 178184 210384 178236 210436
rect 185268 210384 185320 210436
rect 92624 210316 92676 210368
rect 100996 210316 101048 210368
rect 134576 210316 134628 210368
rect 52696 210248 52748 210300
rect 58216 210248 58268 210300
rect 93176 210248 93228 210300
rect 101272 210248 101324 210300
rect 176804 210316 176856 210368
rect 185176 210316 185228 210368
rect 143684 210248 143736 210300
rect 177172 210248 177224 210300
rect 185452 210248 185504 210300
rect 92716 210180 92768 210232
rect 101180 210180 101232 210232
rect 136876 210180 136928 210232
rect 142948 210180 143000 210232
rect 177724 210180 177776 210232
rect 185360 210180 185412 210232
rect 56100 209840 56152 209892
rect 58308 209840 58360 209892
rect 83056 208956 83108 209008
rect 84252 208956 84304 209008
rect 91244 208956 91296 209008
rect 100996 208956 101048 209008
rect 175424 208956 175476 209008
rect 185176 208956 185228 209008
rect 134208 207664 134260 207716
rect 140280 207664 140332 207716
rect 50580 207460 50632 207512
rect 61252 207460 61304 207512
rect 135312 207460 135364 207512
rect 145340 207460 145392 207512
rect 174044 207460 174096 207512
rect 180300 207460 180352 207512
rect 76800 206304 76852 206356
rect 78364 206304 78416 206356
rect 73212 206236 73264 206288
rect 75512 206236 75564 206288
rect 78180 206236 78232 206288
rect 79744 206236 79796 206288
rect 157484 206236 157536 206288
rect 159508 206236 159560 206288
rect 160980 206236 161032 206288
rect 162452 206236 162504 206288
rect 73304 206168 73356 206220
rect 74040 206168 74092 206220
rect 74684 206168 74736 206220
rect 76892 206168 76944 206220
rect 79560 206168 79612 206220
rect 81216 206168 81268 206220
rect 85724 206168 85776 206220
rect 100996 206168 101048 206220
rect 147272 206168 147324 206220
rect 147824 206168 147876 206220
rect 156840 206168 156892 206220
rect 158036 206168 158088 206220
rect 158864 206168 158916 206220
rect 160888 206168 160940 206220
rect 162360 206168 162412 206220
rect 163740 206168 163792 206220
rect 169904 206168 169956 206220
rect 185176 206168 185228 206220
rect 216180 204808 216232 204860
rect 222344 204808 222396 204860
rect 148744 204740 148796 204792
rect 215536 204740 215588 204792
rect 24084 204672 24136 204724
rect 28132 204672 28184 204724
rect 21508 204604 21560 204656
rect 26936 204604 26988 204656
rect 22796 204536 22848 204588
rect 26844 204536 26896 204588
rect 121420 204536 121472 204588
rect 123168 204536 123220 204588
rect 208544 204536 208596 204588
rect 211120 204536 211172 204588
rect 23440 204468 23492 204520
rect 26752 204468 26804 204520
rect 45060 204400 45112 204452
rect 45888 204400 45940 204452
rect 98972 204400 99024 204452
rect 104768 204400 104820 204452
rect 121604 204400 121656 204452
rect 123720 204400 123772 204452
rect 207900 204400 207952 204452
rect 210568 204400 210620 204452
rect 24728 204332 24780 204384
rect 28040 204332 28092 204384
rect 120132 204332 120184 204384
rect 121512 204332 121564 204384
rect 200264 204332 200316 204384
rect 201000 204332 201052 204384
rect 22152 204264 22204 204316
rect 26660 204264 26712 204316
rect 99432 204264 99484 204316
rect 107528 204264 107580 204316
rect 208084 204264 208136 204316
rect 210016 204264 210068 204316
rect 121512 204196 121564 204248
rect 124272 204196 124324 204248
rect 183612 204196 183664 204248
rect 191524 204196 191576 204248
rect 208452 204196 208504 204248
rect 211672 204196 211724 204248
rect 99248 204128 99300 204180
rect 106976 204128 107028 204180
rect 183704 204128 183756 204180
rect 192076 204128 192128 204180
rect 208360 204128 208412 204180
rect 212224 204128 212276 204180
rect 20220 204060 20272 204112
rect 41748 204060 41800 204112
rect 99524 204060 99576 204112
rect 108080 204060 108132 204112
rect 183428 204060 183480 204112
rect 190972 204060 191024 204112
rect 191984 204060 192036 204112
rect 214984 204060 215036 204112
rect 99156 203788 99208 203840
rect 106424 203788 106476 203840
rect 117464 203788 117516 203840
rect 118752 203788 118804 203840
rect 124272 203788 124324 203840
rect 128228 203788 128280 203840
rect 123720 203720 123772 203772
rect 125468 203720 125520 203772
rect 205692 203720 205744 203772
rect 208820 203720 208872 203772
rect 110288 203652 110340 203704
rect 111024 203652 111076 203704
rect 118752 203652 118804 203704
rect 120960 203652 121012 203704
rect 123904 203652 123956 203704
rect 126572 203652 126624 203704
rect 183336 203652 183388 203704
rect 189868 203652 189920 203704
rect 204312 203652 204364 203704
rect 206612 203652 206664 203704
rect 99340 203584 99392 203636
rect 105872 203584 105924 203636
rect 124180 203584 124232 203636
rect 127124 203584 127176 203636
rect 127952 203584 128004 203636
rect 130436 203584 130488 203636
rect 183244 203584 183296 203636
rect 189316 203584 189368 203636
rect 201460 203584 201512 203636
rect 203300 203584 203352 203636
rect 204220 203584 204272 203636
rect 206060 203584 206112 203636
rect 40920 203516 40972 203568
rect 43036 203516 43088 203568
rect 99064 203516 99116 203568
rect 105320 203516 105372 203568
rect 109276 203516 109328 203568
rect 110288 203516 110340 203568
rect 116360 203516 116412 203568
rect 117556 203516 117608 203568
rect 118844 203516 118896 203568
rect 120408 203516 120460 203568
rect 123996 203516 124048 203568
rect 126020 203516 126072 203568
rect 127860 203516 127912 203568
rect 128780 203516 128832 203568
rect 183152 203516 183204 203568
rect 188764 203516 188816 203568
rect 202932 203516 202984 203568
rect 204404 203516 204456 203568
rect 205784 203516 205836 203568
rect 208268 203516 208320 203568
rect 20864 203448 20916 203500
rect 25464 203448 25516 203500
rect 41104 203448 41156 203500
rect 42300 203448 42352 203500
rect 43772 203448 43824 203500
rect 44876 203448 44928 203500
rect 98880 203448 98932 203500
rect 104216 203448 104268 203500
rect 116084 203448 116136 203500
rect 117004 203448 117056 203500
rect 117648 203448 117700 203500
rect 25372 203380 25424 203432
rect 26108 203380 26160 203432
rect 27212 203380 27264 203432
rect 27672 203380 27724 203432
rect 28592 203380 28644 203432
rect 29144 203380 29196 203432
rect 29972 203380 30024 203432
rect 30524 203380 30576 203432
rect 31260 203380 31312 203432
rect 31812 203380 31864 203432
rect 37424 203380 37476 203432
rect 38436 203380 38488 203432
rect 39540 203380 39592 203432
rect 40368 203380 40420 203432
rect 41012 203380 41064 203432
rect 41656 203380 41708 203432
rect 43680 203380 43732 203432
rect 44416 203380 44468 203432
rect 108632 203380 108684 203432
rect 109276 203380 109328 203432
rect 109736 203380 109788 203432
rect 110748 203380 110800 203432
rect 111484 203380 111536 203432
rect 112312 203380 112364 203432
rect 114612 203380 114664 203432
rect 114796 203380 114848 203432
rect 115992 203380 116044 203432
rect 116452 203380 116504 203432
rect 117372 203380 117424 203432
rect 118200 203380 118252 203432
rect 118660 203448 118712 203500
rect 119856 203448 119908 203500
rect 120040 203448 120092 203500
rect 122064 203448 122116 203500
rect 123812 203448 123864 203500
rect 124824 203448 124876 203500
rect 128136 203448 128188 203500
rect 129884 203448 129936 203500
rect 183060 203448 183112 203500
rect 188212 203448 188264 203500
rect 203024 203448 203076 203500
rect 204956 203448 205008 203500
rect 205416 203448 205468 203500
rect 207164 203448 207216 203500
rect 119304 203380 119356 203432
rect 120224 203380 120276 203432
rect 122616 203380 122668 203432
rect 124364 203380 124416 203432
rect 127676 203380 127728 203432
rect 128044 203380 128096 203432
rect 129332 203380 129384 203432
rect 183520 203380 183572 203432
rect 190420 203380 190472 203432
rect 192628 203380 192680 203432
rect 193364 203380 193416 203432
rect 193732 203380 193784 203432
rect 194744 203380 194796 203432
rect 201552 203380 201604 203432
rect 202748 203380 202800 203432
rect 202840 203380 202892 203432
rect 203852 203380 203904 203432
rect 204404 203380 204456 203432
rect 205508 203380 205560 203432
rect 205600 203380 205652 203432
rect 207716 203380 207768 203432
rect 207992 203380 208044 203432
rect 209464 203380 209516 203432
rect 213420 203380 213472 203432
rect 214432 203380 214484 203432
rect 33376 203040 33428 203092
rect 33836 203040 33888 203092
rect 212868 203040 212920 203092
rect 213052 203040 213104 203092
rect 197504 202836 197556 202888
rect 197780 202836 197832 202888
rect 196216 201408 196268 201460
rect 196860 201408 196912 201460
rect 50488 196444 50540 196496
rect 57572 196444 57624 196496
rect 110840 196444 110892 196496
rect 111668 196444 111720 196496
rect 112036 196444 112088 196496
rect 112496 196444 112548 196496
rect 114888 196444 114940 196496
rect 115348 196444 115400 196496
rect 123628 196444 123680 196496
rect 124364 196444 124416 196496
rect 26752 196376 26804 196428
rect 27396 196376 27448 196428
rect 27764 196376 27816 196428
rect 30156 196376 30208 196428
rect 72016 196376 72068 196428
rect 73304 196376 73356 196428
rect 115256 196376 115308 196428
rect 115900 196376 115952 196428
rect 120868 196376 120920 196428
rect 121604 196376 121656 196428
rect 121696 196376 121748 196428
rect 123812 196376 123864 196428
rect 135312 196376 135364 196428
rect 140464 196376 140516 196428
rect 196308 196376 196360 196428
rect 196860 196376 196912 196428
rect 200816 196376 200868 196428
rect 201644 196376 201696 196428
rect 203668 196376 203720 196428
rect 204220 196376 204272 196428
rect 204496 196376 204548 196428
rect 205508 196376 205560 196428
rect 26568 196308 26620 196360
rect 26936 196308 26988 196360
rect 28040 196308 28092 196360
rect 28224 196308 28276 196360
rect 38436 196308 38488 196360
rect 39540 196308 39592 196360
rect 40092 196308 40144 196360
rect 40920 196308 40972 196360
rect 41656 196308 41708 196360
rect 45060 196308 45112 196360
rect 69808 196308 69860 196360
rect 70636 196308 70688 196360
rect 70912 196308 70964 196360
rect 72200 196308 72252 196360
rect 75328 196308 75380 196360
rect 76800 196308 76852 196360
rect 78640 196308 78692 196360
rect 81676 196308 81728 196360
rect 93084 196308 93136 196360
rect 94004 196308 94056 196360
rect 119672 196308 119724 196360
rect 120040 196308 120092 196360
rect 120500 196308 120552 196360
rect 121420 196308 121472 196360
rect 123260 196308 123312 196360
rect 124180 196308 124232 196360
rect 140280 196308 140332 196360
rect 141568 196308 141620 196360
rect 152608 196308 152660 196360
rect 153436 196308 153488 196360
rect 153804 196308 153856 196360
rect 154816 196308 154868 196360
rect 156012 196308 156064 196360
rect 156840 196308 156892 196360
rect 162636 196308 162688 196360
rect 165856 196308 165908 196360
rect 165948 196308 166000 196360
rect 169996 196308 170048 196360
rect 175976 196308 176028 196360
rect 176804 196308 176856 196360
rect 177080 196308 177132 196360
rect 178184 196308 178236 196360
rect 195112 196308 195164 196360
rect 196032 196308 196084 196360
rect 196216 196308 196268 196360
rect 197228 196308 197280 196360
rect 203300 196308 203352 196360
rect 204404 196308 204456 196360
rect 204864 196308 204916 196360
rect 205600 196308 205652 196360
rect 207624 196308 207676 196360
rect 208452 196308 208504 196360
rect 27672 196240 27724 196292
rect 30064 196240 30116 196292
rect 80848 196240 80900 196292
rect 84528 196240 84580 196292
rect 122432 196240 122484 196292
rect 123996 196240 124048 196292
rect 201460 196240 201512 196292
rect 201644 196240 201696 196292
rect 205232 196240 205284 196292
rect 205784 196240 205836 196292
rect 39632 196172 39684 196224
rect 41104 196172 41156 196224
rect 30524 196104 30576 196156
rect 31628 196104 31680 196156
rect 51040 196104 51092 196156
rect 59780 196104 59832 196156
rect 135404 196104 135456 196156
rect 143776 196104 143828 196156
rect 154908 196104 154960 196156
rect 156196 196104 156248 196156
rect 160428 196104 160480 196156
rect 162360 196104 162412 196156
rect 206428 196104 206480 196156
rect 208084 196104 208136 196156
rect 51224 196036 51276 196088
rect 58676 196036 58728 196088
rect 89772 196036 89824 196088
rect 101640 196036 101692 196088
rect 135220 196036 135272 196088
rect 142672 196036 142724 196088
rect 173768 196036 173820 196088
rect 185820 196036 185872 196088
rect 39264 195968 39316 196020
rect 41012 195968 41064 196020
rect 50948 195968 51000 196020
rect 60884 195968 60936 196020
rect 88668 195968 88720 196020
rect 101732 195968 101784 196020
rect 124456 195968 124508 196020
rect 127860 195968 127912 196020
rect 134944 195968 134996 196020
rect 144880 195968 144932 196020
rect 161532 195968 161584 196020
rect 164476 195968 164528 196020
rect 164844 195968 164896 196020
rect 168616 195968 168668 196020
rect 172664 195968 172716 196020
rect 185912 195968 185964 196020
rect 193272 195968 193324 196020
rect 194468 195968 194520 196020
rect 202104 195968 202156 196020
rect 202840 195968 202892 196020
rect 209280 195968 209332 196020
rect 213052 195968 213104 196020
rect 50764 195900 50816 195952
rect 61988 195900 62040 195952
rect 81952 195900 82004 195952
rect 87196 195900 87248 195952
rect 87564 195900 87616 195952
rect 102100 195900 102152 195952
rect 135128 195900 135180 195952
rect 145984 195900 146036 195952
rect 171560 195900 171612 195952
rect 186280 195900 186332 195952
rect 208820 195900 208872 195952
rect 212868 195900 212920 195952
rect 26384 195832 26436 195884
rect 29696 195832 29748 195884
rect 31904 195832 31956 195884
rect 32824 195832 32876 195884
rect 36872 195832 36924 195884
rect 37332 195832 37384 195884
rect 41288 195832 41340 195884
rect 43772 195832 43824 195884
rect 50672 195832 50724 195884
rect 63092 195832 63144 195884
rect 86460 195832 86512 195884
rect 101916 195832 101968 195884
rect 122064 195832 122116 195884
rect 123720 195832 123772 195884
rect 135036 195832 135088 195884
rect 148192 195832 148244 195884
rect 163740 195832 163792 195884
rect 167236 195832 167288 195884
rect 170456 195832 170508 195884
rect 186096 195832 186148 195884
rect 209648 195832 209700 195884
rect 213420 195832 213472 195884
rect 26292 195764 26344 195816
rect 29236 195764 29288 195816
rect 50856 195764 50908 195816
rect 64196 195764 64248 195816
rect 65024 195764 65076 195816
rect 94188 195764 94240 195816
rect 125652 195764 125704 195816
rect 127952 195764 128004 195816
rect 134852 195764 134904 195816
rect 147088 195764 147140 195816
rect 147824 195764 147876 195816
rect 179288 195764 179340 195816
rect 208452 195764 208504 195816
rect 212960 195764 213012 195816
rect 26200 195696 26252 195748
rect 28868 195696 28920 195748
rect 31996 195696 32048 195748
rect 32916 195696 32968 195748
rect 33376 195696 33428 195748
rect 34480 195696 34532 195748
rect 79744 195696 79796 195748
rect 83056 195696 83108 195748
rect 91980 195696 92032 195748
rect 92624 195696 92676 195748
rect 122892 195696 122944 195748
rect 123904 195696 123956 195748
rect 194928 195696 194980 195748
rect 195664 195696 195716 195748
rect 206060 195696 206112 195748
rect 207992 195696 208044 195748
rect 38068 195628 38120 195680
rect 38988 195628 39040 195680
rect 40460 195628 40512 195680
rect 43128 195628 43180 195680
rect 125284 195628 125336 195680
rect 128136 195628 128188 195680
rect 207256 195628 207308 195680
rect 208544 195628 208596 195680
rect 124824 195560 124876 195612
rect 128044 195560 128096 195612
rect 206888 195560 206940 195612
rect 207900 195560 207952 195612
rect 33468 195492 33520 195544
rect 34112 195492 34164 195544
rect 77536 195492 77588 195544
rect 79560 195492 79612 195544
rect 29144 195424 29196 195476
rect 30892 195424 30944 195476
rect 37700 195424 37752 195476
rect 38896 195424 38948 195476
rect 51132 195424 51184 195476
rect 56468 195424 56520 195476
rect 76432 195424 76484 195476
rect 78180 195424 78232 195476
rect 119304 195424 119356 195476
rect 120132 195424 120184 195476
rect 197596 195356 197648 195408
rect 198056 195356 198108 195408
rect 38896 195288 38948 195340
rect 40828 195288 40880 195340
rect 159324 195288 159376 195340
rect 160980 195288 161032 195340
rect 29052 195220 29104 195272
rect 31260 195220 31312 195272
rect 194652 195220 194704 195272
rect 195296 195220 195348 195272
rect 30432 195152 30484 195204
rect 40828 195152 40880 195204
rect 43680 195152 43732 195204
rect 32088 195084 32140 195136
rect 118660 194132 118712 194184
rect 118844 194132 118896 194184
rect 211948 190596 212000 190648
rect 217560 190596 217612 190648
rect 187936 188216 187988 188268
rect 191984 188216 192036 188268
rect 99432 186856 99484 186908
rect 106792 186856 106844 186908
rect 13320 186788 13372 186840
rect 22796 186788 22848 186840
rect 104400 184068 104452 184120
rect 106792 184068 106844 184120
rect 99524 184000 99576 184052
rect 105780 184000 105832 184052
rect 182876 184000 182928 184052
rect 187936 184000 187988 184052
rect 13412 182708 13464 182760
rect 22336 182708 22388 182760
rect 104492 182708 104544 182760
rect 107160 182708 107212 182760
rect 128504 182708 128556 182760
rect 137520 182708 137572 182760
rect 212500 182708 212552 182760
rect 220412 182708 220464 182760
rect 98604 182640 98656 182692
rect 106976 182640 107028 182692
rect 183152 182640 183204 182692
rect 191156 182640 191208 182692
rect 183704 181280 183756 181332
rect 191984 181280 192036 181332
rect 105136 180328 105188 180380
rect 106976 180328 107028 180380
rect 98420 179852 98472 179904
rect 104492 179852 104544 179904
rect 182508 179852 182560 179904
rect 190696 179852 190748 179904
rect 183704 179784 183756 179836
rect 190604 179784 190656 179836
rect 99524 179512 99576 179564
rect 104400 179512 104452 179564
rect 182508 178492 182560 178544
rect 191984 178492 192036 178544
rect 99524 177336 99576 177388
rect 105136 177336 105188 177388
rect 98604 177132 98656 177184
rect 106792 177132 106844 177184
rect 183244 176452 183296 176504
rect 191984 176452 192036 176504
rect 211764 176316 211816 176368
rect 216272 176316 216324 176368
rect 13320 175840 13372 175892
rect 22336 175840 22388 175892
rect 98236 175772 98288 175824
rect 106608 175772 106660 175824
rect 183704 175092 183756 175144
rect 191524 175092 191576 175144
rect 99524 173664 99576 173716
rect 106792 173664 106844 173716
rect 183336 173052 183388 173104
rect 191984 173052 192036 173104
rect 99524 171692 99576 171744
rect 106792 171692 106844 171744
rect 183520 171692 183572 171744
rect 191156 171692 191208 171744
rect 182692 171216 182744 171268
rect 185084 171216 185136 171268
rect 99432 170264 99484 170316
rect 106792 170196 106844 170248
rect 99524 168904 99576 168956
rect 106700 168904 106752 168956
rect 182508 168904 182560 168956
rect 191892 168904 191944 168956
rect 44416 168836 44468 168888
rect 49844 168836 49896 168888
rect 185084 168836 185136 168888
rect 191984 168836 192036 168888
rect 99524 167612 99576 167664
rect 106884 167612 106936 167664
rect 49844 167544 49896 167596
rect 53432 167544 53484 167596
rect 99432 167544 99484 167596
rect 106792 167544 106844 167596
rect 183704 167544 183756 167596
rect 191340 167544 191392 167596
rect 182876 166456 182928 166508
rect 187936 166456 187988 166508
rect 99524 166184 99576 166236
rect 107252 166184 107304 166236
rect 212684 165232 212736 165284
rect 218296 165232 218348 165284
rect 183704 164960 183756 165012
rect 190052 164960 190104 165012
rect 99524 164756 99576 164808
rect 107160 164756 107212 164808
rect 211764 163600 211816 163652
rect 218296 163600 218348 163652
rect 99524 163396 99576 163448
rect 104400 163396 104452 163448
rect 128504 163396 128556 163448
rect 138164 163396 138216 163448
rect 183060 163396 183112 163448
rect 189960 163396 190012 163448
rect 183796 162988 183848 163040
rect 191984 162988 192036 163040
rect 187936 161968 187988 162020
rect 191340 161968 191392 162020
rect 211948 156460 212000 156512
rect 212684 156460 212736 156512
rect 216916 156460 216968 156512
rect 182692 155440 182744 155492
rect 188028 155440 188080 155492
rect 104400 155032 104452 155084
rect 106516 155032 106568 155084
rect 27764 152312 27816 152364
rect 29696 152312 29748 152364
rect 30524 152312 30576 152364
rect 31260 152312 31312 152364
rect 32088 152312 32140 152364
rect 32824 152312 32876 152364
rect 37240 152312 37292 152364
rect 38988 152312 39040 152364
rect 39264 152312 39316 152364
rect 40184 152312 40236 152364
rect 41656 152312 41708 152364
rect 43680 152312 43732 152364
rect 109184 152312 109236 152364
rect 110104 152312 110156 152364
rect 119672 152312 119724 152364
rect 121972 152312 122024 152364
rect 124824 152312 124876 152364
rect 129240 152312 129292 152364
rect 193272 152312 193324 152364
rect 194468 152312 194520 152364
rect 194928 152312 194980 152364
rect 195664 152312 195716 152364
rect 196584 152312 196636 152364
rect 197228 152312 197280 152364
rect 197596 152312 197648 152364
rect 198056 152312 198108 152364
rect 202104 152312 202156 152364
rect 202932 152312 202984 152364
rect 203668 152312 203720 152364
rect 205968 152312 206020 152364
rect 30432 152244 30484 152296
rect 31628 152244 31680 152296
rect 38896 152244 38948 152296
rect 39908 152244 39960 152296
rect 118476 152244 118528 152296
rect 120592 152244 120644 152296
rect 124456 152244 124508 152296
rect 128780 152244 128832 152296
rect 193364 152244 193416 152296
rect 194100 152244 194152 152296
rect 203300 152244 203352 152296
rect 206060 152244 206112 152296
rect 29144 152176 29196 152228
rect 30892 152176 30944 152228
rect 38436 152176 38488 152228
rect 41840 152176 41892 152228
rect 120500 152176 120552 152228
rect 123168 152176 123220 152228
rect 123628 152176 123680 152228
rect 127952 152176 128004 152228
rect 204864 152176 204916 152228
rect 207348 152176 207400 152228
rect 36872 152108 36924 152160
rect 38896 152108 38948 152160
rect 120040 152108 120092 152160
rect 123076 152108 123128 152160
rect 204496 152108 204548 152160
rect 207256 152108 207308 152160
rect 118844 152040 118896 152092
rect 120960 152040 121012 152092
rect 205232 152040 205284 152092
rect 207992 152040 208044 152092
rect 208820 152040 208872 152092
rect 212868 152040 212920 152092
rect 119304 151972 119356 152024
rect 121788 151972 121840 152024
rect 31812 151836 31864 151888
rect 32456 151836 32508 151888
rect 40460 151836 40512 151888
rect 44968 151836 45020 151888
rect 122892 151836 122944 151888
rect 127308 151904 127360 151956
rect 206428 151904 206480 151956
rect 210016 151904 210068 151956
rect 123260 151836 123312 151888
rect 127216 151836 127268 151888
rect 206336 151836 206388 151888
rect 208820 151836 208872 151888
rect 79192 151768 79244 151820
rect 98236 151768 98288 151820
rect 207624 151768 207676 151820
rect 210936 151768 210988 151820
rect 26292 151700 26344 151752
rect 29236 151700 29288 151752
rect 38068 151700 38120 151752
rect 40920 151700 40972 151752
rect 69164 151700 69216 151752
rect 92532 151700 92584 151752
rect 41288 151632 41340 151684
rect 45152 151632 45204 151684
rect 37700 151564 37752 151616
rect 40276 151564 40328 151616
rect 72568 151564 72620 151616
rect 36044 151428 36096 151480
rect 37608 151428 37660 151480
rect 95384 151700 95436 151752
rect 156564 151700 156616 151752
rect 209648 151700 209700 151752
rect 214248 151700 214300 151752
rect 98236 151632 98288 151684
rect 98880 151632 98932 151684
rect 163188 151632 163240 151684
rect 200448 151632 200500 151684
rect 201184 151632 201236 151684
rect 205692 151632 205744 151684
rect 207900 151632 207952 151684
rect 209280 151632 209332 151684
rect 214156 151632 214208 151684
rect 124088 151496 124140 151548
rect 127860 151496 127912 151548
rect 195112 151496 195164 151548
rect 196032 151496 196084 151548
rect 122432 151428 122484 151480
rect 125100 151428 125152 151480
rect 25004 151360 25056 151412
rect 28500 151360 28552 151412
rect 29052 151360 29104 151412
rect 30156 151360 30208 151412
rect 24912 151292 24964 151344
rect 28040 151292 28092 151344
rect 121696 151292 121748 151344
rect 124640 151292 124692 151344
rect 125652 151292 125704 151344
rect 131356 151292 131408 151344
rect 208084 151292 208136 151344
rect 210752 151292 210804 151344
rect 26384 151224 26436 151276
rect 28868 151224 28920 151276
rect 31996 151224 32048 151276
rect 33284 151224 33336 151276
rect 118108 151224 118160 151276
rect 120316 151224 120368 151276
rect 121236 151224 121288 151276
rect 123720 151224 123772 151276
rect 194652 151224 194704 151276
rect 195296 151224 195348 151276
rect 25740 151156 25792 151208
rect 27672 151156 27724 151208
rect 36504 151156 36556 151208
rect 37424 151156 37476 151208
rect 206888 151156 206940 151208
rect 210108 151156 210160 151208
rect 26016 151088 26068 151140
rect 27304 151088 27356 151140
rect 35308 151088 35360 151140
rect 36044 151088 36096 151140
rect 199620 151088 199672 151140
rect 200172 151088 200224 151140
rect 25924 151020 25976 151072
rect 26844 151020 26896 151072
rect 27672 151020 27724 151072
rect 30064 151020 30116 151072
rect 40828 151020 40880 151072
rect 45060 151020 45112 151072
rect 25832 150952 25884 151004
rect 26476 150952 26528 151004
rect 33468 150952 33520 151004
rect 34112 150952 34164 151004
rect 109552 150952 109604 151004
rect 110472 150952 110524 151004
rect 110472 150816 110524 150868
rect 111300 151020 111352 151072
rect 111668 150952 111720 151004
rect 112496 151020 112548 151072
rect 120868 151020 120920 151072
rect 123812 151020 123864 151072
rect 125284 151020 125336 151072
rect 129332 151020 129384 151072
rect 112128 150952 112180 151004
rect 112864 150952 112916 151004
rect 115624 150952 115676 151004
rect 115992 150952 116044 151004
rect 116452 150952 116504 151004
rect 117464 150952 117516 151004
rect 117648 150952 117700 151004
rect 118844 150952 118896 151004
rect 122064 150952 122116 151004
rect 125192 150952 125244 151004
rect 194744 150952 194796 151004
rect 195020 150952 195072 151004
rect 196860 151020 196912 151072
rect 208452 151020 208504 151072
rect 210660 151020 210712 151072
rect 204036 150952 204088 151004
rect 206244 150952 206296 151004
rect 207532 150952 207584 151004
rect 210844 150952 210896 151004
rect 110656 150884 110708 150936
rect 112036 150884 112088 150936
rect 196216 150884 196268 150936
rect 59228 146804 59280 146856
rect 59412 146736 59464 146788
rect 127216 146124 127268 146176
rect 127676 146124 127728 146176
rect 197596 146124 197648 146176
rect 198148 146124 198200 146176
rect 40184 144016 40236 144068
rect 43036 144016 43088 144068
rect 59412 144059 59464 144068
rect 59412 144025 59421 144059
rect 59421 144025 59455 144059
rect 59455 144025 59464 144059
rect 59412 144016 59464 144025
rect 118844 144016 118896 144068
rect 119580 144016 119632 144068
rect 120960 144016 121012 144068
rect 121696 144016 121748 144068
rect 123812 144016 123864 144068
rect 124456 144016 124508 144068
rect 125192 144016 125244 144068
rect 126020 144016 126072 144068
rect 127952 144016 128004 144068
rect 128596 144016 128648 144068
rect 129240 144016 129292 144068
rect 130068 144016 130120 144068
rect 183612 144016 183664 144068
rect 187936 144016 187988 144068
rect 193088 144016 193140 144068
rect 193364 144016 193416 144068
rect 198424 144016 198476 144068
rect 199068 144016 199120 144068
rect 201184 144016 201236 144068
rect 201736 144016 201788 144068
rect 202932 144016 202984 144068
rect 203852 144016 203904 144068
rect 39908 143948 39960 144000
rect 42300 143948 42352 144000
rect 123720 143948 123772 144000
rect 124548 143948 124600 144000
rect 125100 143948 125152 144000
rect 126572 143948 126624 144000
rect 127860 143948 127912 144000
rect 128688 143948 128740 144000
rect 129332 143948 129384 144000
rect 130620 143948 130672 144000
rect 183428 143948 183480 144000
rect 189408 143948 189460 144000
rect 198884 143948 198936 144000
rect 199252 143948 199304 144000
rect 201276 143948 201328 144000
rect 202748 143948 202800 144000
rect 203024 143948 203076 144000
rect 204956 143948 205008 144000
rect 40092 143880 40144 143932
rect 44416 143880 44468 143932
rect 117280 143880 117332 143932
rect 119028 143880 119080 143932
rect 183520 143880 183572 143932
rect 189500 143880 189552 143932
rect 200816 143880 200868 143932
rect 202288 143880 202340 143932
rect 202472 143880 202524 143932
rect 204496 143880 204548 143932
rect 23256 143812 23308 143864
rect 26016 143812 26068 143864
rect 39632 143812 39684 143864
rect 43772 143812 43824 143864
rect 183336 143812 183388 143864
rect 190052 143812 190104 143864
rect 201644 143812 201696 143864
rect 203300 143812 203352 143864
rect 22152 143744 22204 143796
rect 25924 143744 25976 143796
rect 24452 143676 24504 143728
rect 24912 143676 24964 143728
rect 20772 143608 20824 143660
rect 25096 143608 25148 143660
rect 26016 143608 26068 143660
rect 26384 143608 26436 143660
rect 27304 143608 27356 143660
rect 27764 143608 27816 143660
rect 28592 143608 28644 143660
rect 29052 143608 29104 143660
rect 30064 143608 30116 143660
rect 30524 143608 30576 143660
rect 31996 143608 32048 143660
rect 32732 143608 32784 143660
rect 34480 143608 34532 143660
rect 34940 143608 34992 143660
rect 43680 143608 43732 143660
rect 47176 143608 47228 143660
rect 114428 143608 114480 143660
rect 114980 143608 115032 143660
rect 115992 143608 116044 143660
rect 116636 143608 116688 143660
rect 117464 143608 117516 143660
rect 117924 143608 117976 143660
rect 205968 143608 206020 143660
rect 206152 143608 206204 143660
rect 207992 143608 208044 143660
rect 208636 143608 208688 143660
rect 208820 143608 208872 143660
rect 209556 143608 209608 143660
rect 210844 143608 210896 143660
rect 211396 143608 211448 143660
rect 214248 143608 214300 143660
rect 214708 143608 214760 143660
rect 23532 143540 23584 143592
rect 25740 143540 25792 143592
rect 34848 143540 34900 143592
rect 35492 143540 35544 143592
rect 99248 143540 99300 143592
rect 106608 143540 106660 143592
rect 114888 143540 114940 143592
rect 115532 143540 115584 143592
rect 115900 143540 115952 143592
rect 117648 143540 117700 143592
rect 207900 143540 207952 143592
rect 209004 143540 209056 143592
rect 35676 143472 35728 143524
rect 36964 143472 37016 143524
rect 99156 143472 99208 143524
rect 106792 143472 106844 143524
rect 183244 143472 183296 143524
rect 190788 143472 190840 143524
rect 99064 143404 99116 143456
rect 107436 143404 107488 143456
rect 183060 143404 183112 143456
rect 192076 143404 192128 143456
rect 194192 143404 194244 143456
rect 194744 143404 194796 143456
rect 20496 143336 20548 143388
rect 44508 143336 44560 143388
rect 98972 143336 99024 143388
rect 107988 143336 108040 143388
rect 183152 143336 183204 143388
rect 191340 143336 191392 143388
rect 191984 143336 192036 143388
rect 215628 143336 215680 143388
rect 45152 143200 45204 143252
rect 46532 143200 46584 143252
rect 110288 143200 110340 143252
rect 110564 143200 110616 143252
rect 116820 143064 116872 143116
rect 118476 143064 118528 143116
rect 210936 143064 210988 143116
rect 211764 143064 211816 143116
rect 45060 142928 45112 142980
rect 45796 142928 45848 142980
rect 98788 142928 98840 142980
rect 103940 142928 103992 142980
rect 210660 142928 210712 142980
rect 212868 142928 212920 142980
rect 99432 142860 99484 142912
rect 105596 142860 105648 142912
rect 200264 142860 200316 142912
rect 200908 142860 200960 142912
rect 21784 142792 21836 142844
rect 25832 142792 25884 142844
rect 31352 142792 31404 142844
rect 31904 142792 31956 142844
rect 37424 142792 37476 142844
rect 38252 142792 38304 142844
rect 99340 142792 99392 142844
rect 105136 142792 105188 142844
rect 210752 142792 210804 142844
rect 212316 142792 212368 142844
rect 99524 142724 99576 142776
rect 104584 142724 104636 142776
rect 68704 142656 68756 142708
rect 69164 142656 69216 142708
rect 167696 142452 167748 142504
rect 169904 142452 169956 142504
rect 134852 140004 134904 140056
rect 143592 140004 143644 140056
rect 49936 139936 49988 139988
rect 56192 139936 56244 139988
rect 135404 139936 135456 139988
rect 143316 139936 143368 139988
rect 135404 138712 135456 138764
rect 139820 138712 139872 138764
rect 49936 138644 49988 138696
rect 58492 138644 58544 138696
rect 50028 138576 50080 138628
rect 58400 138576 58452 138628
rect 134668 138576 134720 138628
rect 139636 138576 139688 138628
rect 51408 138508 51460 138560
rect 59228 138508 59280 138560
rect 92716 138508 92768 138560
rect 100812 138508 100864 138560
rect 177632 138508 177684 138560
rect 185084 138508 185136 138560
rect 56192 138440 56244 138492
rect 58676 138440 58728 138492
rect 92808 138440 92860 138492
rect 100904 138440 100956 138492
rect 177724 138440 177776 138492
rect 184992 138440 185044 138492
rect 134668 137352 134720 137404
rect 139728 137352 139780 137404
rect 97868 137284 97920 137336
rect 100996 137284 101048 137336
rect 49936 137216 49988 137268
rect 58308 137216 58360 137268
rect 97960 137216 98012 137268
rect 101272 137216 101324 137268
rect 181588 137216 181640 137268
rect 185176 137216 185228 137268
rect 50028 137148 50080 137200
rect 135404 137148 135456 137200
rect 143408 137148 143460 137200
rect 182232 137148 182284 137200
rect 185452 137148 185504 137200
rect 58216 137080 58268 137132
rect 92716 137080 92768 137132
rect 101180 137080 101232 137132
rect 177632 137080 177684 137132
rect 185268 137080 185320 137132
rect 92808 137012 92860 137064
rect 101088 137012 101140 137064
rect 139636 137012 139688 137064
rect 143592 137012 143644 137064
rect 177724 137012 177776 137064
rect 185360 137012 185412 137064
rect 92716 136944 92768 136996
rect 97868 136944 97920 136996
rect 139820 136944 139872 136996
rect 143132 136944 143184 136996
rect 139728 136604 139780 136656
rect 143500 136604 143552 136656
rect 177724 136604 177776 136656
rect 181588 136604 181640 136656
rect 51224 136128 51276 136180
rect 52788 136128 52840 136180
rect 51224 135992 51276 136044
rect 52696 135992 52748 136044
rect 135036 135924 135088 135976
rect 143316 135924 143368 135976
rect 98052 135856 98104 135908
rect 101456 135856 101508 135908
rect 135312 135856 135364 135908
rect 143592 135856 143644 135908
rect 182324 135856 182376 135908
rect 185360 135856 185412 135908
rect 50396 135788 50448 135840
rect 98144 135788 98196 135840
rect 101732 135788 101784 135840
rect 135404 135788 135456 135840
rect 143224 135788 143276 135840
rect 181956 135788 182008 135840
rect 185268 135788 185320 135840
rect 58216 135720 58268 135772
rect 92808 135720 92860 135772
rect 101824 135720 101876 135772
rect 177632 135720 177684 135772
rect 185176 135720 185228 135772
rect 92716 135652 92768 135704
rect 97960 135652 98012 135704
rect 177724 135652 177776 135704
rect 182232 135652 182284 135704
rect 51224 134564 51276 134616
rect 56744 134564 56796 134616
rect 134668 134564 134720 134616
rect 136876 134564 136928 134616
rect 51132 134496 51184 134548
rect 52880 134496 52932 134548
rect 59412 134539 59464 134548
rect 59412 134505 59421 134539
rect 59421 134505 59455 134539
rect 59455 134505 59464 134539
rect 59412 134496 59464 134505
rect 134852 134496 134904 134548
rect 139636 134496 139688 134548
rect 52788 134360 52840 134412
rect 58216 134360 58268 134412
rect 92900 134360 92952 134412
rect 101456 134360 101508 134412
rect 177632 134360 177684 134412
rect 185176 134360 185228 134412
rect 52696 134292 52748 134344
rect 58308 134292 58360 134344
rect 92716 134292 92768 134344
rect 98052 134292 98104 134344
rect 177724 134292 177776 134344
rect 181956 134292 182008 134344
rect 92808 134224 92860 134276
rect 98144 134224 98196 134276
rect 177724 134020 177776 134072
rect 182324 134020 182376 134072
rect 56744 133816 56796 133868
rect 58216 133816 58268 133868
rect 139636 133748 139688 133800
rect 142948 133748 143000 133800
rect 50948 133068 51000 133120
rect 52696 133068 52748 133120
rect 134116 133068 134168 133120
rect 138164 133068 138216 133120
rect 50212 133000 50264 133052
rect 56100 133000 56152 133052
rect 135404 133000 135456 133052
rect 52880 132932 52932 132984
rect 58216 132932 58268 132984
rect 59412 132932 59464 132984
rect 92808 132932 92860 132984
rect 101824 132932 101876 132984
rect 143224 132932 143276 132984
rect 177632 132932 177684 132984
rect 185176 132932 185228 132984
rect 92716 132864 92768 132916
rect 100904 132864 100956 132916
rect 177724 132864 177776 132916
rect 185084 132864 185136 132916
rect 136876 132796 136928 132848
rect 143592 132796 143644 132848
rect 56100 132388 56152 132440
rect 58308 132388 58360 132440
rect 50396 131980 50448 132032
rect 53432 131980 53484 132032
rect 51224 131912 51276 131964
rect 55456 131912 55508 131964
rect 134484 131912 134536 131964
rect 137152 131912 137204 131964
rect 135312 131708 135364 131760
rect 137980 131708 138032 131760
rect 51224 131640 51276 131692
rect 52788 131640 52840 131692
rect 135128 131640 135180 131692
rect 52696 131572 52748 131624
rect 58216 131572 58268 131624
rect 92716 131572 92768 131624
rect 101732 131572 101784 131624
rect 142488 131572 142540 131624
rect 177632 131572 177684 131624
rect 185912 131572 185964 131624
rect 92808 131504 92860 131556
rect 101824 131504 101876 131556
rect 138164 131504 138216 131556
rect 143592 131504 143644 131556
rect 177724 131504 177776 131556
rect 185820 131504 185872 131556
rect 55456 131300 55508 131352
rect 58308 131300 58360 131352
rect 51224 130688 51276 130740
rect 52972 130688 53024 130740
rect 134668 130552 134720 130604
rect 137612 130552 137664 130604
rect 51224 130280 51276 130332
rect 52696 130280 52748 130332
rect 134852 130280 134904 130332
rect 137428 130280 137480 130332
rect 53432 130212 53484 130264
rect 58216 130212 58268 130264
rect 92716 130212 92768 130264
rect 101180 130212 101232 130264
rect 137152 130212 137204 130264
rect 143592 130212 143644 130264
rect 177632 130212 177684 130264
rect 185544 130212 185596 130264
rect 52788 130144 52840 130196
rect 58308 130144 58360 130196
rect 92808 130144 92860 130196
rect 101548 130144 101600 130196
rect 137980 130144 138032 130196
rect 143040 130144 143092 130196
rect 177724 130144 177776 130196
rect 185728 130144 185780 130196
rect 134668 129328 134720 129380
rect 137520 129328 137572 129380
rect 50396 129056 50448 129108
rect 56468 129056 56520 129108
rect 51224 128920 51276 128972
rect 52880 128920 52932 128972
rect 135404 128920 135456 128972
rect 52696 128852 52748 128904
rect 58308 128852 58360 128904
rect 92716 128852 92768 128904
rect 101824 128852 101876 128904
rect 143132 128852 143184 128904
rect 177356 128852 177408 128904
rect 185176 128852 185228 128904
rect 52972 128784 53024 128836
rect 58216 128784 58268 128836
rect 92808 128784 92860 128836
rect 101364 128784 101416 128836
rect 137428 128784 137480 128836
rect 142764 128784 142816 128836
rect 177632 128784 177684 128836
rect 185268 128784 185320 128836
rect 92716 128716 92768 128768
rect 101732 128716 101784 128768
rect 137612 128716 137664 128768
rect 143592 128716 143644 128768
rect 177724 128716 177776 128768
rect 185360 128716 185412 128768
rect 56468 128308 56520 128360
rect 58216 128308 58268 128360
rect 50948 127832 51000 127884
rect 56744 127832 56796 127884
rect 134668 127832 134720 127884
rect 137612 127832 137664 127884
rect 51224 127764 51276 127816
rect 52788 127764 52840 127816
rect 134668 127696 134720 127748
rect 136876 127696 136928 127748
rect 51224 127560 51276 127612
rect 52696 127560 52748 127612
rect 135404 127492 135456 127544
rect 52880 127424 52932 127476
rect 58216 127424 58268 127476
rect 92808 127424 92860 127476
rect 100996 127424 101048 127476
rect 143316 127424 143368 127476
rect 177724 127424 177776 127476
rect 185176 127424 185228 127476
rect 216272 127424 216324 127476
rect 222344 127424 222396 127476
rect 92716 127356 92768 127408
rect 101272 127356 101324 127408
rect 137520 127356 137572 127408
rect 142488 127356 142540 127408
rect 177172 127356 177224 127408
rect 185452 127356 185504 127408
rect 56744 127152 56796 127204
rect 58308 127152 58360 127204
rect 98052 126200 98104 126252
rect 101824 126200 101876 126252
rect 182232 126200 182284 126252
rect 185452 126200 185504 126252
rect 98144 126132 98196 126184
rect 101732 126132 101784 126184
rect 182324 126132 182376 126184
rect 185176 126132 185228 126184
rect 52696 126064 52748 126116
rect 58308 126064 58360 126116
rect 92808 126064 92860 126116
rect 101088 126064 101140 126116
rect 137612 126064 137664 126116
rect 143592 126064 143644 126116
rect 177632 126064 177684 126116
rect 185268 126064 185320 126116
rect 52788 125996 52840 126048
rect 58216 125996 58268 126048
rect 92716 125996 92768 126048
rect 101180 125996 101232 126048
rect 136876 125996 136928 126048
rect 143040 125996 143092 126048
rect 177724 125996 177776 126048
rect 185360 125996 185412 126048
rect 135036 125248 135088 125300
rect 137612 125248 137664 125300
rect 51224 124976 51276 125028
rect 52972 124976 53024 125028
rect 51224 124840 51276 124892
rect 52880 124840 52932 124892
rect 135404 124840 135456 124892
rect 136876 124840 136928 124892
rect 50212 124772 50264 124824
rect 58400 124772 58452 124824
rect 135220 124772 135272 124824
rect 142764 124772 142816 124824
rect 51316 124704 51368 124756
rect 58308 124704 58360 124756
rect 92900 124704 92952 124756
rect 101456 124704 101508 124756
rect 135588 124704 135640 124756
rect 143592 124704 143644 124756
rect 177632 124704 177684 124756
rect 185176 124704 185228 124756
rect 51408 124636 51460 124688
rect 58216 124636 58268 124688
rect 92716 124636 92768 124688
rect 98052 124636 98104 124688
rect 177724 124636 177776 124688
rect 182232 124636 182284 124688
rect 92808 124568 92860 124620
rect 98144 124568 98196 124620
rect 135496 124364 135548 124416
rect 142488 124364 142540 124416
rect 177172 124364 177224 124416
rect 182324 124364 182376 124416
rect 134484 123480 134536 123532
rect 137704 123480 137756 123532
rect 50580 123412 50632 123464
rect 52696 123412 52748 123464
rect 51132 123344 51184 123396
rect 52788 123344 52840 123396
rect 134116 123344 134168 123396
rect 138164 123344 138216 123396
rect 52972 123276 53024 123328
rect 58216 123276 58268 123328
rect 92716 123276 92768 123328
rect 101640 123276 101692 123328
rect 137612 123276 137664 123328
rect 143592 123276 143644 123328
rect 177632 123276 177684 123328
rect 185268 123276 185320 123328
rect 52880 123208 52932 123260
rect 58308 123208 58360 123260
rect 92808 123208 92860 123260
rect 101732 123208 101784 123260
rect 177724 123208 177776 123260
rect 185360 123208 185412 123260
rect 136876 122868 136928 122920
rect 142856 122868 142908 122920
rect 134484 122392 134536 122444
rect 138072 122392 138124 122444
rect 50856 122324 50908 122376
rect 52972 122324 53024 122376
rect 134944 122256 134996 122308
rect 137244 122256 137296 122308
rect 50212 122188 50264 122240
rect 52880 122188 52932 122240
rect 52788 121916 52840 121968
rect 58308 121916 58360 121968
rect 92808 121916 92860 121968
rect 101824 121916 101876 121968
rect 137704 121916 137756 121968
rect 142764 121916 142816 121968
rect 177632 121916 177684 121968
rect 185728 121916 185780 121968
rect 52696 121848 52748 121900
rect 58216 121848 58268 121900
rect 92716 121848 92768 121900
rect 101916 121848 101968 121900
rect 138164 121848 138216 121900
rect 143040 121848 143092 121900
rect 177724 121848 177776 121900
rect 185912 121848 185964 121900
rect 51224 120896 51276 120948
rect 53064 120896 53116 120948
rect 97868 120760 97920 120812
rect 101732 120760 101784 120812
rect 134484 120760 134536 120812
rect 137428 120760 137480 120812
rect 182048 120760 182100 120812
rect 185360 120760 185412 120812
rect 51224 120692 51276 120744
rect 52696 120692 52748 120744
rect 97960 120692 98012 120744
rect 101088 120692 101140 120744
rect 134668 120692 134720 120744
rect 137520 120692 137572 120744
rect 182324 120692 182376 120744
rect 185268 120692 185320 120744
rect 50212 120624 50264 120676
rect 53156 120624 53208 120676
rect 98144 120624 98196 120676
rect 101548 120624 101600 120676
rect 135404 120624 135456 120676
rect 136876 120624 136928 120676
rect 181772 120624 181824 120676
rect 185176 120624 185228 120676
rect 52972 120556 53024 120608
rect 58216 120556 58268 120608
rect 92716 120556 92768 120608
rect 101640 120556 101692 120608
rect 138072 120556 138124 120608
rect 142948 120556 143000 120608
rect 177724 120556 177776 120608
rect 185820 120556 185872 120608
rect 52880 120488 52932 120540
rect 58308 120488 58360 120540
rect 92808 120488 92860 120540
rect 101456 120488 101508 120540
rect 137244 120488 137296 120540
rect 143592 120488 143644 120540
rect 177632 120488 177684 120540
rect 185544 120488 185596 120540
rect 51224 119536 51276 119588
rect 52880 119536 52932 119588
rect 135404 119536 135456 119588
rect 137612 119536 137664 119588
rect 97684 119332 97736 119384
rect 101272 119332 101324 119384
rect 182140 119332 182192 119384
rect 185268 119332 185320 119384
rect 51224 119264 51276 119316
rect 52788 119264 52840 119316
rect 98052 119264 98104 119316
rect 101364 119264 101416 119316
rect 134484 119264 134536 119316
rect 136968 119264 137020 119316
rect 182232 119264 182284 119316
rect 185176 119264 185228 119316
rect 52696 119196 52748 119248
rect 58400 119196 58452 119248
rect 92900 119196 92952 119248
rect 98144 119196 98196 119248
rect 137428 119196 137480 119248
rect 143592 119196 143644 119248
rect 53156 119128 53208 119180
rect 58216 119128 58268 119180
rect 92808 119128 92860 119180
rect 97960 119128 98012 119180
rect 136876 119128 136928 119180
rect 142580 119128 142632 119180
rect 177724 119128 177776 119180
rect 182048 119128 182100 119180
rect 53064 119060 53116 119112
rect 58308 119060 58360 119112
rect 92716 119060 92768 119112
rect 97868 119060 97920 119112
rect 137520 119060 137572 119112
rect 143592 119060 143644 119112
rect 177724 118924 177776 118976
rect 181772 118924 181824 118976
rect 177632 118788 177684 118840
rect 182324 118788 182376 118840
rect 134668 118448 134720 118500
rect 136876 118448 136928 118500
rect 51224 118176 51276 118228
rect 52972 118176 53024 118228
rect 134668 118176 134720 118228
rect 137520 118176 137572 118228
rect 51224 117904 51276 117956
rect 52696 117904 52748 117956
rect 97960 117904 98012 117956
rect 101364 117904 101416 117956
rect 181404 117904 181456 117956
rect 185268 117904 185320 117956
rect 98144 117836 98196 117888
rect 101732 117836 101784 117888
rect 182324 117836 182376 117888
rect 185176 117836 185228 117888
rect 52880 117768 52932 117820
rect 58216 117768 58268 117820
rect 92716 117768 92768 117820
rect 97684 117768 97736 117820
rect 136968 117768 137020 117820
rect 142580 117768 142632 117820
rect 52788 117700 52840 117752
rect 58308 117700 58360 117752
rect 92808 117700 92860 117752
rect 98052 117700 98104 117752
rect 137612 117700 137664 117752
rect 143224 117700 143276 117752
rect 177724 117700 177776 117752
rect 182140 117700 182192 117752
rect 177632 117564 177684 117616
rect 182232 117564 182284 117616
rect 51224 116680 51276 116732
rect 56468 116680 56520 116732
rect 94004 116544 94056 116596
rect 101088 116544 101140 116596
rect 178184 116544 178236 116596
rect 185268 116544 185320 116596
rect 92624 116476 92676 116528
rect 100996 116476 101048 116528
rect 134852 116476 134904 116528
rect 52972 116408 53024 116460
rect 58216 116408 58268 116460
rect 92900 116408 92952 116460
rect 101180 116408 101232 116460
rect 176804 116476 176856 116528
rect 185176 116476 185228 116528
rect 142764 116408 142816 116460
rect 177080 116408 177132 116460
rect 185360 116408 185412 116460
rect 52696 116340 52748 116392
rect 58308 116340 58360 116392
rect 92716 116340 92768 116392
rect 97960 116340 98012 116392
rect 136876 116340 136928 116392
rect 142948 116340 143000 116392
rect 177724 116340 177776 116392
rect 181404 116340 181456 116392
rect 56468 116272 56520 116324
rect 58400 116272 58452 116324
rect 92808 116272 92860 116324
rect 98144 116272 98196 116324
rect 137520 116272 137572 116324
rect 143592 116272 143644 116324
rect 177724 116068 177776 116120
rect 182324 116068 182376 116120
rect 91244 115184 91296 115236
rect 101088 115184 101140 115236
rect 175424 115184 175476 115236
rect 185268 115184 185320 115236
rect 59320 115159 59372 115168
rect 59320 115125 59329 115159
rect 59329 115125 59363 115159
rect 59363 115125 59372 115159
rect 59320 115116 59372 115125
rect 90600 115116 90652 115168
rect 100996 115116 101048 115168
rect 174780 115116 174832 115168
rect 185176 115116 185228 115168
rect 51224 113824 51276 113876
rect 57572 113824 57624 113876
rect 135404 113688 135456 113740
rect 141568 113688 141620 113740
rect 17828 113280 17880 113332
rect 64104 113280 64156 113332
rect 147272 113280 147324 113332
rect 218388 113280 218440 113332
rect 18012 112940 18064 112992
rect 52604 112940 52656 112992
rect 85724 112328 85776 112380
rect 100996 112328 101048 112380
rect 169904 112328 169956 112380
rect 185176 112328 185228 112380
rect 52604 112260 52656 112312
rect 61896 112260 61948 112312
rect 90416 112192 90468 112244
rect 93360 112192 93412 112244
rect 134024 111648 134076 111700
rect 145340 111648 145392 111700
rect 82320 111580 82372 111632
rect 85448 111580 85500 111632
rect 129976 111580 130028 111632
rect 148100 111580 148152 111632
rect 83700 111512 83752 111564
rect 87196 111512 87248 111564
rect 80940 111444 80992 111496
rect 84068 111444 84120 111496
rect 79652 111104 79704 111156
rect 82596 111104 82648 111156
rect 163832 111104 163884 111156
rect 166592 111104 166644 111156
rect 167880 111104 167932 111156
rect 170916 111104 170968 111156
rect 74040 111036 74092 111088
rect 75512 111036 75564 111088
rect 77444 111036 77496 111088
rect 79744 111036 79796 111088
rect 158864 111036 158916 111088
rect 160888 111036 160940 111088
rect 166500 111036 166552 111088
rect 169444 111036 169496 111088
rect 74684 110968 74736 111020
rect 76892 110968 76944 111020
rect 79560 110968 79612 111020
rect 81216 110968 81268 111020
rect 156840 110968 156892 111020
rect 158036 110968 158088 111020
rect 158312 110968 158364 111020
rect 159508 110968 159560 111020
rect 161624 110968 161676 111020
rect 163740 110968 163792 111020
rect 165120 110968 165172 111020
rect 168064 110968 168116 111020
rect 172664 110968 172716 111020
rect 176160 110968 176212 111020
rect 109000 110900 109052 110952
rect 129976 110900 130028 110952
rect 63276 110832 63328 110884
rect 109552 110832 109604 110884
rect 113232 110560 113284 110612
rect 114520 110560 114572 110612
rect 115808 110560 115860 110612
rect 118292 110560 118344 110612
rect 113140 110492 113192 110544
rect 113968 110492 114020 110544
rect 114612 110492 114664 110544
rect 115624 110492 115676 110544
rect 115900 110492 115952 110544
rect 116728 110492 116780 110544
rect 117464 110492 117516 110544
rect 118844 110492 118896 110544
rect 31076 110424 31128 110476
rect 31904 110424 31956 110476
rect 99524 110424 99576 110476
rect 107344 110424 107396 110476
rect 183612 110356 183664 110408
rect 191616 110356 191668 110408
rect 99432 110288 99484 110340
rect 106792 110288 106844 110340
rect 115992 110288 116044 110340
rect 117280 110288 117332 110340
rect 183704 110288 183756 110340
rect 192168 110288 192220 110340
rect 208268 110288 208320 110340
rect 213236 110288 213288 110340
rect 20220 110220 20272 110272
rect 41748 110220 41800 110272
rect 98788 110220 98840 110272
rect 107896 110220 107948 110272
rect 183520 110220 183572 110272
rect 191064 110220 191116 110272
rect 191984 110220 192036 110272
rect 215536 110220 215588 110272
rect 25924 109948 25976 110000
rect 26292 109948 26344 110000
rect 29052 109948 29104 110000
rect 30892 109948 30944 110000
rect 24912 109880 24964 109932
rect 22888 109812 22940 109864
rect 27304 109812 27356 109864
rect 27672 109880 27724 109932
rect 30064 109880 30116 109932
rect 28500 109812 28552 109864
rect 99248 109812 99300 109864
rect 106240 109812 106292 109864
rect 115716 109812 115768 109864
rect 117832 109812 117884 109864
rect 118936 109812 118988 109864
rect 119948 109812 120000 109864
rect 183336 109812 183388 109864
rect 190420 109812 190472 109864
rect 23624 109744 23676 109796
rect 27672 109744 27724 109796
rect 44416 109744 44468 109796
rect 45060 109744 45112 109796
rect 99156 109744 99208 109796
rect 105136 109744 105188 109796
rect 119580 109744 119632 109796
rect 121052 109744 121104 109796
rect 126664 109744 126716 109796
rect 129332 109744 129384 109796
rect 183244 109744 183296 109796
rect 189316 109744 189368 109796
rect 205232 109744 205284 109796
rect 206980 109744 207032 109796
rect 21508 109676 21560 109728
rect 26476 109676 26528 109728
rect 37516 109676 37568 109728
rect 38252 109676 38304 109728
rect 42944 109676 42996 109728
rect 47452 109676 47504 109728
rect 99064 109676 99116 109728
rect 104584 109676 104636 109728
rect 119948 109676 120000 109728
rect 122156 109676 122208 109728
rect 183152 109676 183204 109728
rect 188764 109676 188816 109728
rect 203760 109676 203812 109728
rect 205324 109676 205376 109728
rect 208176 109676 208228 109728
rect 212132 109676 212184 109728
rect 22244 109608 22296 109660
rect 26844 109608 26896 109660
rect 27028 109608 27080 109660
rect 29696 109608 29748 109660
rect 38160 109608 38212 109660
rect 40000 109608 40052 109660
rect 45060 109608 45112 109660
rect 46808 109608 46860 109660
rect 98972 109608 99024 109660
rect 104124 109608 104176 109660
rect 119856 109608 119908 109660
rect 121604 109608 121656 109660
rect 126480 109608 126532 109660
rect 128780 109608 128832 109660
rect 129332 109608 129384 109660
rect 130988 109608 131040 109660
rect 183060 109608 183112 109660
rect 188212 109608 188264 109660
rect 201460 109608 201512 109660
rect 202472 109608 202524 109660
rect 205140 109608 205192 109660
rect 206428 109608 206480 109660
rect 208360 109608 208412 109660
rect 212684 109608 212736 109660
rect 213512 109608 213564 109660
rect 214984 109608 215036 109660
rect 20864 109540 20916 109592
rect 22980 109540 23032 109592
rect 24268 109540 24320 109592
rect 28132 109540 28184 109592
rect 28316 109540 28368 109592
rect 29144 109540 29196 109592
rect 38252 109540 38304 109592
rect 39264 109540 39316 109592
rect 45152 109540 45204 109592
rect 46072 109540 46124 109592
rect 99340 109540 99392 109592
rect 105688 109540 105740 109592
rect 119764 109540 119816 109592
rect 120500 109540 120552 109592
rect 120960 109540 121012 109592
rect 122708 109540 122760 109592
rect 126572 109540 126624 109592
rect 128228 109540 128280 109592
rect 129240 109540 129292 109592
rect 130436 109540 130488 109592
rect 183428 109540 183480 109592
rect 189868 109540 189920 109592
rect 193916 109540 193968 109592
rect 194744 109540 194796 109592
rect 201644 109540 201696 109592
rect 203024 109540 203076 109592
rect 203852 109540 203904 109592
rect 204680 109540 204732 109592
rect 205416 109540 205468 109592
rect 205876 109540 205928 109592
rect 208544 109540 208596 109592
rect 211580 109540 211632 109592
rect 213420 109540 213472 109592
rect 214432 109540 214484 109592
rect 59320 108180 59372 108232
rect 59412 108112 59464 108164
rect 41656 107500 41708 107552
rect 42300 107500 42352 107552
rect 43036 107500 43088 107552
rect 43772 107500 43824 107552
rect 208636 107500 208688 107552
rect 209004 107500 209056 107552
rect 210016 107500 210068 107552
rect 210660 107500 210712 107552
rect 30248 102604 30300 102656
rect 31260 102604 31312 102656
rect 32088 102604 32140 102656
rect 32824 102604 32876 102656
rect 35308 102604 35360 102656
rect 36136 102604 36188 102656
rect 36872 102604 36924 102656
rect 38252 102604 38304 102656
rect 111300 102604 111352 102656
rect 111760 102604 111812 102656
rect 112496 102604 112548 102656
rect 113324 102604 113376 102656
rect 113692 102604 113744 102656
rect 114704 102604 114756 102656
rect 193272 102604 193324 102656
rect 194100 102604 194152 102656
rect 196308 102604 196360 102656
rect 196860 102604 196912 102656
rect 198424 102604 198476 102656
rect 199160 102604 199212 102656
rect 199620 102604 199672 102656
rect 200356 102604 200408 102656
rect 200816 102604 200868 102656
rect 201368 102604 201420 102656
rect 201460 102604 201512 102656
rect 203116 102604 203168 102656
rect 204864 102604 204916 102656
rect 207348 102604 207400 102656
rect 32732 102536 32784 102588
rect 33284 102536 33336 102588
rect 35676 102536 35728 102588
rect 36780 102536 36832 102588
rect 37700 102536 37752 102588
rect 40276 102536 40328 102588
rect 111668 102536 111720 102588
rect 112312 102536 112364 102588
rect 119672 102536 119724 102588
rect 123260 102536 123312 102588
rect 200080 102536 200132 102588
rect 200632 102536 200684 102588
rect 201276 102536 201328 102588
rect 201644 102536 201696 102588
rect 203300 102536 203352 102588
rect 205416 102536 205468 102588
rect 206428 102536 206480 102588
rect 210108 102536 210160 102588
rect 36044 102468 36096 102520
rect 37608 102468 37660 102520
rect 38068 102468 38120 102520
rect 40828 102468 40880 102520
rect 114060 102468 114112 102520
rect 114612 102468 114664 102520
rect 115256 102468 115308 102520
rect 115992 102468 116044 102520
rect 120868 102468 120920 102520
rect 124916 102468 124968 102520
rect 22980 102400 23032 102452
rect 26108 102400 26160 102452
rect 93360 102400 93412 102452
rect 94188 102400 94240 102452
rect 120040 102400 120092 102452
rect 123812 102400 123864 102452
rect 202472 102400 202524 102452
rect 203852 102400 203904 102452
rect 50948 102332 51000 102384
rect 59780 102332 59832 102384
rect 114428 102332 114480 102384
rect 116176 102332 116228 102384
rect 122432 102332 122484 102384
rect 127124 102332 127176 102384
rect 135128 102332 135180 102384
rect 143776 102332 143828 102384
rect 159324 102332 159376 102384
rect 161716 102332 161768 102384
rect 206060 102332 206112 102384
rect 208820 102332 208872 102384
rect 122064 102264 122116 102316
rect 126112 102264 126164 102316
rect 50672 102196 50724 102248
rect 60884 102196 60936 102248
rect 121696 102196 121748 102248
rect 126020 102196 126072 102248
rect 134852 102196 134904 102248
rect 144880 102196 144932 102248
rect 200448 102196 200500 102248
rect 201552 102196 201604 102248
rect 208820 102196 208872 102248
rect 212868 102196 212920 102248
rect 50856 102128 50908 102180
rect 61988 102128 62040 102180
rect 120500 102128 120552 102180
rect 124364 102128 124416 102180
rect 135036 102128 135088 102180
rect 145984 102128 146036 102180
rect 50764 102060 50816 102112
rect 63092 102060 63144 102112
rect 88668 102060 88720 102112
rect 101824 102060 101876 102112
rect 122892 102060 122944 102112
rect 127676 102060 127728 102112
rect 134760 102060 134812 102112
rect 147088 102060 147140 102112
rect 172664 102060 172716 102112
rect 185820 102060 185872 102112
rect 199252 102060 199304 102112
rect 199712 102060 199764 102112
rect 202104 102060 202156 102112
rect 203208 102060 203260 102112
rect 204036 102060 204088 102112
rect 205232 102060 205284 102112
rect 209280 102060 209332 102112
rect 213420 102060 213472 102112
rect 26292 101992 26344 102044
rect 28868 101992 28920 102044
rect 29144 101992 29196 102044
rect 30432 101992 30484 102044
rect 36504 101992 36556 102044
rect 37516 101992 37568 102044
rect 50580 101992 50632 102044
rect 64196 101992 64248 102044
rect 87564 101992 87616 102044
rect 102008 101992 102060 102044
rect 114888 101992 114940 102044
rect 115900 101992 115952 102044
rect 134944 101992 134996 102044
rect 148192 101992 148244 102044
rect 161532 101992 161584 102044
rect 164476 101992 164528 102044
rect 171560 101992 171612 102044
rect 186004 101992 186056 102044
rect 209648 101992 209700 102044
rect 213512 101992 213564 102044
rect 51132 101924 51184 101976
rect 58676 101924 58728 101976
rect 59412 101924 59464 101976
rect 83148 101924 83200 101976
rect 86460 101924 86512 101976
rect 101640 101924 101692 101976
rect 112036 101924 112088 101976
rect 112864 101924 112916 101976
rect 135312 101924 135364 101976
rect 142672 101924 142724 101976
rect 143684 101924 143736 101976
rect 167144 101924 167196 101976
rect 170456 101924 170508 101976
rect 186188 101924 186240 101976
rect 40092 101856 40144 101908
rect 44508 101856 44560 101908
rect 30524 101788 30576 101840
rect 31628 101788 31680 101840
rect 37240 101788 37292 101840
rect 38160 101788 38212 101840
rect 39264 101788 39316 101840
rect 43128 101788 43180 101840
rect 116452 101788 116504 101840
rect 117464 101788 117516 101840
rect 124456 101788 124508 101840
rect 129884 101788 129936 101840
rect 205232 101788 205284 101840
rect 208728 101788 208780 101840
rect 26384 101720 26436 101772
rect 29236 101720 29288 101772
rect 38436 101720 38488 101772
rect 41840 101720 41892 101772
rect 51040 101720 51092 101772
rect 56468 101720 56520 101772
rect 121236 101720 121288 101772
rect 125468 101720 125520 101772
rect 206888 101720 206940 101772
rect 210016 101720 210068 101772
rect 40828 101652 40880 101704
rect 45152 101652 45204 101704
rect 116820 101652 116872 101704
rect 119396 101652 119448 101704
rect 123260 101652 123312 101704
rect 126572 101652 126624 101704
rect 202840 101652 202892 101704
rect 203760 101652 203812 101704
rect 204496 101652 204548 101704
rect 207256 101652 207308 101704
rect 39632 101584 39684 101636
rect 43036 101584 43088 101636
rect 117648 101584 117700 101636
rect 119764 101584 119816 101636
rect 124824 101584 124876 101636
rect 129240 101584 129292 101636
rect 40460 101516 40512 101568
rect 44416 101516 44468 101568
rect 75328 101516 75380 101568
rect 77536 101516 77588 101568
rect 118476 101516 118528 101568
rect 119856 101516 119908 101568
rect 123628 101516 123680 101568
rect 126480 101516 126532 101568
rect 207624 101516 207676 101568
rect 208176 101516 208228 101568
rect 38896 101448 38948 101500
rect 41656 101448 41708 101500
rect 118844 101448 118896 101500
rect 119948 101448 120000 101500
rect 124088 101448 124140 101500
rect 126664 101448 126716 101500
rect 194652 101448 194704 101500
rect 195296 101448 195348 101500
rect 203668 101448 203720 101500
rect 205140 101448 205192 101500
rect 205692 101448 205744 101500
rect 208636 101448 208688 101500
rect 31812 101380 31864 101432
rect 32456 101380 32508 101432
rect 41288 101380 41340 101432
rect 45060 101380 45112 101432
rect 72384 101380 72436 101432
rect 73488 101380 73540 101432
rect 77536 101380 77588 101432
rect 79560 101380 79612 101432
rect 80848 101380 80900 101432
rect 82320 101380 82372 101432
rect 117280 101380 117332 101432
rect 118936 101380 118988 101432
rect 119304 101380 119356 101432
rect 120960 101380 121012 101432
rect 125652 101380 125704 101432
rect 131540 101380 131592 101432
rect 154908 101380 154960 101432
rect 156196 101380 156248 101432
rect 158220 101380 158272 101432
rect 158864 101380 158916 101432
rect 163740 101380 163792 101432
rect 165120 101380 165172 101432
rect 165948 101380 166000 101432
rect 167880 101380 167932 101432
rect 176160 101380 176212 101432
rect 179288 101380 179340 101432
rect 193364 101380 193416 101432
rect 194468 101380 194520 101432
rect 194744 101380 194796 101432
rect 195020 101380 195072 101432
rect 195112 101380 195164 101432
rect 196032 101380 196084 101432
rect 207256 101380 207308 101432
rect 208544 101380 208596 101432
rect 41656 101312 41708 101364
rect 42944 101312 42996 101364
rect 68612 101312 68664 101364
rect 69256 101312 69308 101364
rect 69808 101312 69860 101364
rect 70636 101312 70688 101364
rect 70912 101312 70964 101364
rect 72016 101312 72068 101364
rect 73120 101312 73172 101364
rect 74040 101312 74092 101364
rect 76432 101312 76484 101364
rect 77444 101312 77496 101364
rect 78640 101312 78692 101364
rect 79652 101312 79704 101364
rect 79744 101312 79796 101364
rect 80940 101312 80992 101364
rect 81952 101312 82004 101364
rect 83700 101312 83752 101364
rect 89772 101312 89824 101364
rect 90600 101312 90652 101364
rect 91980 101312 92032 101364
rect 92624 101312 92676 101364
rect 93084 101312 93136 101364
rect 94004 101312 94056 101364
rect 118108 101312 118160 101364
rect 119580 101312 119632 101364
rect 125284 101312 125336 101364
rect 129332 101312 129384 101364
rect 135220 101312 135272 101364
rect 140464 101312 140516 101364
rect 152608 101312 152660 101364
rect 153436 101312 153488 101364
rect 153804 101312 153856 101364
rect 154816 101312 154868 101364
rect 156012 101312 156064 101364
rect 156840 101312 156892 101364
rect 157116 101312 157168 101364
rect 158312 101312 158364 101364
rect 160428 101312 160480 101364
rect 161624 101312 161676 101364
rect 162636 101312 162688 101364
rect 163832 101312 163884 101364
rect 164844 101312 164896 101364
rect 166500 101312 166552 101364
rect 173768 101312 173820 101364
rect 174780 101312 174832 101364
rect 175976 101312 176028 101364
rect 176804 101312 176856 101364
rect 177080 101312 177132 101364
rect 178184 101312 178236 101364
rect 194928 101312 194980 101364
rect 195664 101312 195716 101364
rect 208084 101312 208136 101364
rect 208360 101312 208412 101364
rect 212040 99884 212092 99936
rect 222344 99884 222396 99936
rect 98788 97164 98840 97216
rect 106792 97164 106844 97216
rect 13320 97096 13372 97148
rect 22336 97096 22388 97148
rect 211764 97096 211816 97148
rect 216180 97096 216232 97148
rect 99524 95804 99576 95856
rect 106792 95804 106844 95856
rect 188580 94376 188632 94428
rect 191984 94376 192036 94428
rect 98696 93016 98748 93068
rect 106516 93016 106568 93068
rect 13320 90228 13372 90280
rect 22336 90228 22388 90280
rect 105044 90228 105096 90280
rect 106792 90228 106844 90280
rect 182876 90160 182928 90212
rect 188580 90160 188632 90212
rect 211856 90160 211908 90212
rect 221700 90160 221752 90212
rect 104952 88868 105004 88920
rect 106792 88868 106844 88920
rect 128504 88868 128556 88920
rect 132000 88868 132052 88920
rect 183520 88800 183572 88852
rect 191156 88800 191208 88852
rect 183704 87440 183756 87492
rect 190788 87440 190840 87492
rect 183704 86012 183756 86064
rect 191708 86012 191760 86064
rect 99524 85196 99576 85248
rect 105044 85196 105096 85248
rect 99432 84652 99484 84704
rect 106792 84652 106844 84704
rect 182508 84652 182560 84704
rect 191984 84652 192036 84704
rect 183704 84584 183756 84636
rect 191616 84584 191668 84636
rect 99524 84448 99576 84500
rect 104952 84448 105004 84500
rect 99524 83292 99576 83344
rect 107804 83292 107856 83344
rect 183704 82612 183756 82664
rect 191984 82612 192036 82664
rect 13320 82000 13372 82052
rect 22336 82000 22388 82052
rect 99524 81932 99576 81984
rect 106792 82068 106844 82120
rect 183244 81252 183296 81304
rect 191892 81252 191944 81304
rect 132000 80504 132052 80556
rect 136876 80504 136928 80556
rect 99524 79824 99576 79876
rect 106792 79824 106844 79876
rect 183704 79212 183756 79264
rect 191984 79144 192036 79196
rect 99524 77852 99576 77904
rect 106516 77852 106568 77904
rect 183520 77852 183572 77904
rect 191984 77852 192036 77904
rect 99524 76424 99576 76476
rect 100996 76424 101048 76476
rect 183060 76424 183112 76476
rect 185176 76424 185228 76476
rect 98236 75064 98288 75116
rect 44416 74996 44468 75048
rect 52604 74996 52656 75048
rect 183244 75064 183296 75116
rect 186004 75064 186056 75116
rect 100996 74996 101048 75048
rect 106792 74996 106844 75048
rect 185176 74996 185228 75048
rect 191524 74996 191576 75048
rect 100996 74860 101048 74912
rect 52604 74656 52656 74708
rect 53432 74656 53484 74708
rect 183704 73840 183756 73892
rect 99524 73772 99576 73824
rect 105136 73772 105188 73824
rect 99432 73704 99484 73756
rect 106700 73704 106752 73756
rect 183704 73704 183756 73756
rect 188488 73704 188540 73756
rect 217560 73772 217612 73824
rect 222344 73772 222396 73824
rect 190788 73704 190840 73756
rect 100996 73636 101048 73688
rect 106792 73636 106844 73688
rect 186004 73636 186056 73688
rect 191984 73636 192036 73688
rect 99524 72344 99576 72396
rect 106516 72344 106568 72396
rect 99524 70984 99576 71036
rect 104492 70984 104544 71036
rect 183704 70916 183756 70968
rect 191524 70916 191576 70968
rect 128504 70168 128556 70220
rect 134024 70168 134076 70220
rect 136876 70168 136928 70220
rect 182876 69896 182928 69948
rect 189960 69896 190012 69948
rect 99524 69556 99576 69608
rect 104400 69556 104452 69608
rect 188488 69488 188540 69540
rect 190972 69488 191024 69540
rect 105136 68128 105188 68180
rect 106608 68128 106660 68180
rect 183796 68128 183848 68180
rect 191340 68128 191392 68180
rect 104492 63640 104544 63692
rect 106608 63640 106660 63692
rect 18104 63572 18156 63624
rect 22336 63572 22388 63624
rect 212684 63164 212736 63216
rect 217560 63164 217612 63216
rect 183704 61464 183756 61516
rect 188028 61464 188080 61516
rect 99524 61260 99576 61312
rect 103020 61260 103072 61312
rect 104400 61192 104452 61244
rect 107160 61192 107212 61244
rect 182692 60376 182744 60428
rect 184440 60376 184492 60428
rect 99524 59900 99576 59952
rect 100352 59900 100404 59952
rect 36136 58472 36188 58524
rect 37516 58472 37568 58524
rect 98880 58472 98932 58524
rect 163188 58472 163240 58524
rect 208084 58472 208136 58524
rect 210660 58472 210712 58524
rect 72568 58336 72620 58388
rect 79192 58336 79244 58388
rect 95384 58268 95436 58320
rect 209648 58404 209700 58456
rect 212040 58404 212092 58456
rect 122064 58268 122116 58320
rect 124548 58268 124600 58320
rect 209280 58336 209332 58388
rect 212132 58336 212184 58388
rect 156564 58268 156616 58320
rect 207624 58268 207676 58320
rect 210752 58268 210804 58320
rect 41656 58200 41708 58252
rect 46440 58200 46492 58252
rect 206888 58200 206940 58252
rect 210016 58200 210068 58252
rect 119304 58132 119356 58184
rect 121144 58132 121196 58184
rect 207256 58132 207308 58184
rect 210844 58132 210896 58184
rect 116452 58064 116504 58116
rect 117648 58064 117700 58116
rect 208820 58064 208872 58116
rect 212224 58064 212276 58116
rect 122432 57996 122484 58048
rect 125192 57996 125244 58048
rect 206428 57996 206480 58048
rect 210108 57996 210160 58048
rect 70544 57928 70596 57980
rect 92532 57928 92584 57980
rect 124456 57928 124508 57980
rect 128596 57928 128648 57980
rect 13320 57860 13372 57912
rect 72568 57860 72620 57912
rect 201552 57860 201604 57912
rect 202748 57860 202800 57912
rect 13412 57792 13464 57844
rect 79192 57792 79244 57844
rect 123628 57792 123680 57844
rect 127216 57792 127268 57844
rect 156104 57792 156156 57844
rect 169904 57792 169956 57844
rect 208452 57792 208504 57844
rect 212868 57792 212920 57844
rect 120500 57656 120552 57708
rect 123168 57656 123220 57708
rect 39264 57588 39316 57640
rect 43036 57588 43088 57640
rect 117280 57588 117332 57640
rect 118292 57588 118344 57640
rect 200816 57588 200868 57640
rect 202196 57588 202248 57640
rect 40092 57520 40144 57572
rect 43680 57520 43732 57572
rect 199620 57520 199672 57572
rect 200448 57520 200500 57572
rect 205232 57520 205284 57572
rect 207992 57520 208044 57572
rect 39632 57452 39684 57504
rect 43128 57452 43180 57504
rect 123260 57452 123312 57504
rect 126112 57452 126164 57504
rect 204496 57452 204548 57504
rect 207348 57452 207400 57504
rect 38896 57384 38948 57436
rect 41840 57384 41892 57436
rect 109092 57384 109144 57436
rect 110472 57384 110524 57436
rect 203668 57384 203720 57436
rect 205232 57384 205284 57436
rect 29144 57316 29196 57368
rect 30432 57316 30484 57368
rect 37700 57316 37752 57368
rect 40276 57316 40328 57368
rect 40828 57316 40880 57368
rect 45152 57316 45204 57368
rect 118476 57316 118528 57368
rect 120500 57316 120552 57368
rect 120868 57316 120920 57368
rect 123352 57316 123404 57368
rect 124088 57316 124140 57368
rect 127308 57316 127360 57368
rect 204036 57316 204088 57368
rect 205324 57316 205376 57368
rect 36872 57248 36924 57300
rect 38160 57248 38212 57300
rect 40460 57248 40512 57300
rect 44600 57248 44652 57300
rect 118844 57248 118896 57300
rect 120776 57248 120828 57300
rect 121696 57248 121748 57300
rect 124456 57248 124508 57300
rect 124824 57248 124876 57300
rect 128872 57248 128924 57300
rect 194928 57248 194980 57300
rect 195664 57248 195716 57300
rect 199068 57248 199120 57300
rect 199804 57248 199856 57300
rect 202472 57248 202524 57300
rect 204496 57248 204548 57300
rect 204864 57248 204916 57300
rect 207256 57248 207308 57300
rect 30432 57180 30484 57232
rect 31260 57180 31312 57232
rect 26476 57112 26528 57164
rect 27396 57112 27448 57164
rect 29420 57112 29472 57164
rect 29788 57112 29840 57164
rect 30524 57112 30576 57164
rect 31628 57112 31680 57164
rect 32456 57180 32508 57232
rect 37240 57180 37292 57232
rect 38252 57180 38304 57232
rect 38436 57180 38488 57232
rect 40920 57180 40972 57232
rect 112864 57180 112916 57232
rect 116084 57180 116136 57232
rect 116636 57180 116688 57232
rect 118016 57180 118068 57232
rect 119672 57180 119724 57232
rect 120960 57180 121012 57232
rect 122892 57180 122944 57232
rect 125100 57180 125152 57232
rect 125652 57180 125704 57232
rect 130068 57180 130120 57232
rect 193272 57180 193324 57232
rect 194468 57180 194520 57232
rect 200724 57180 200776 57232
rect 201828 57180 201880 57232
rect 202104 57180 202156 57232
rect 203024 57180 203076 57232
rect 203300 57180 203352 57232
rect 205140 57180 205192 57232
rect 205692 57180 205744 57232
rect 207900 57180 207952 57232
rect 32088 57112 32140 57164
rect 32824 57112 32876 57164
rect 31904 57044 31956 57096
rect 31996 57044 32048 57096
rect 33284 57112 33336 57164
rect 33376 57112 33428 57164
rect 34112 57112 34164 57164
rect 35308 57112 35360 57164
rect 36044 57112 36096 57164
rect 36504 57112 36556 57164
rect 37608 57112 37660 57164
rect 38068 57112 38120 57164
rect 40368 57112 40420 57164
rect 41288 57112 41340 57164
rect 45060 57112 45112 57164
rect 109184 57112 109236 57164
rect 110104 57112 110156 57164
rect 111668 57112 111720 57164
rect 112588 57112 112640 57164
rect 112772 57112 112824 57164
rect 113232 57112 113284 57164
rect 113508 57112 113560 57164
rect 114060 57112 114112 57164
rect 114428 57112 114480 57164
rect 114980 57112 115032 57164
rect 115624 57112 115676 57164
rect 116268 57112 116320 57164
rect 116820 57112 116872 57164
rect 117740 57112 117792 57164
rect 118108 57112 118160 57164
rect 118660 57112 118712 57164
rect 118844 57112 118896 57164
rect 120040 57112 120092 57164
rect 121052 57112 121104 57164
rect 121236 57112 121288 57164
rect 123996 57112 124048 57164
rect 125284 57112 125336 57164
rect 128964 57112 129016 57164
rect 193364 57112 193416 57164
rect 194100 57112 194152 57164
rect 194744 57112 194796 57164
rect 195020 57112 195072 57164
rect 195112 57112 195164 57164
rect 196032 57112 196084 57164
rect 196308 57112 196360 57164
rect 196860 57112 196912 57164
rect 198792 57112 198844 57164
rect 110656 57044 110708 57096
rect 198056 57087 198108 57096
rect 198056 57053 198065 57087
rect 198065 57053 198099 57087
rect 198099 57053 198108 57087
rect 198056 57044 198108 57053
rect 200172 57112 200224 57164
rect 200908 57112 200960 57164
rect 201644 57112 201696 57164
rect 202380 57112 202432 57164
rect 202840 57112 202892 57164
rect 204588 57112 204640 57164
rect 206060 57112 206112 57164
rect 207164 57112 207216 57164
rect 199068 56976 199120 57028
rect 98788 55004 98840 55056
rect 99524 55004 99576 55056
rect 26660 54392 26712 54444
rect 26844 54392 26896 54444
rect 210660 50516 210712 50568
rect 210936 50516 210988 50568
rect 210016 50380 210068 50432
rect 210660 50380 210712 50432
rect 114888 50312 114940 50364
rect 31996 50244 32048 50296
rect 32732 50244 32784 50296
rect 33376 50244 33428 50296
rect 34204 50244 34256 50296
rect 41840 50244 41892 50296
rect 42300 50244 42352 50296
rect 114980 50244 115032 50296
rect 22888 50176 22940 50228
rect 26752 50176 26804 50228
rect 28316 50176 28368 50228
rect 29144 50176 29196 50228
rect 29696 50176 29748 50228
rect 30432 50176 30484 50228
rect 31076 50176 31128 50228
rect 31812 50176 31864 50228
rect 40920 50176 40972 50228
rect 42024 50176 42076 50228
rect 118660 50176 118712 50228
rect 119856 50176 119908 50228
rect 120960 50176 121012 50228
rect 122064 50176 122116 50228
rect 125192 50176 125244 50228
rect 126020 50176 126072 50228
rect 184440 50176 184492 50228
rect 188212 50176 188264 50228
rect 193916 50176 193968 50228
rect 194652 50176 194704 50228
rect 202380 50176 202432 50228
rect 203576 50176 203628 50228
rect 205140 50176 205192 50228
rect 205876 50176 205928 50228
rect 207992 50176 208044 50228
rect 208728 50176 208780 50228
rect 212040 50176 212092 50228
rect 214984 50176 215036 50228
rect 24912 50108 24964 50160
rect 27948 50108 28000 50160
rect 114980 50108 115032 50160
rect 115072 50108 115124 50160
rect 205232 50108 205284 50160
rect 206428 50108 206480 50160
rect 207900 50108 207952 50160
rect 209280 50108 209332 50160
rect 210936 50108 210988 50160
rect 212684 50108 212736 50160
rect 24268 50040 24320 50092
rect 27856 50040 27908 50092
rect 29052 50040 29104 50092
rect 30708 50040 30760 50092
rect 99524 50040 99576 50092
rect 105320 50040 105372 50092
rect 205324 50040 205376 50092
rect 206980 50040 207032 50092
rect 22244 49972 22296 50024
rect 26844 49972 26896 50024
rect 27672 49972 27724 50024
rect 29420 49972 29472 50024
rect 99248 49972 99300 50024
rect 106424 49972 106476 50024
rect 183612 49972 183664 50024
rect 189316 49972 189368 50024
rect 207256 49972 207308 50024
rect 207900 49972 207952 50024
rect 23624 49904 23676 49956
rect 26476 49904 26528 49956
rect 99340 49904 99392 49956
rect 105872 49904 105924 49956
rect 121052 49904 121104 49956
rect 122616 49904 122668 49956
rect 99156 49700 99208 49752
rect 106976 49700 107028 49752
rect 26292 49632 26344 49684
rect 29328 49632 29380 49684
rect 183244 49632 183296 49684
rect 191064 49632 191116 49684
rect 99064 49564 99116 49616
rect 107528 49564 107580 49616
rect 125100 49564 125152 49616
rect 126572 49564 126624 49616
rect 183060 49564 183112 49616
rect 192168 49564 192220 49616
rect 20220 49496 20272 49548
rect 44508 49496 44560 49548
rect 98972 49496 99024 49548
rect 108080 49496 108132 49548
rect 183152 49496 183204 49548
rect 191616 49496 191668 49548
rect 191984 49496 192036 49548
rect 215536 49564 215588 49616
rect 210844 49496 210896 49548
rect 211580 49496 211632 49548
rect 212224 49496 212276 49548
rect 213880 49496 213932 49548
rect 21508 49428 21560 49480
rect 26568 49428 26620 49480
rect 183428 49224 183480 49276
rect 189868 49224 189920 49276
rect 212132 49224 212184 49276
rect 214432 49224 214484 49276
rect 25648 49088 25700 49140
rect 28040 49156 28092 49208
rect 207164 49156 207216 49208
rect 209832 49156 209884 49208
rect 27028 49088 27080 49140
rect 29512 49088 29564 49140
rect 38160 49088 38212 49140
rect 39264 49088 39316 49140
rect 183336 49088 183388 49140
rect 190420 49088 190472 49140
rect 203024 49088 203076 49140
rect 204128 49088 204180 49140
rect 210752 49088 210804 49140
rect 212132 49088 212184 49140
rect 20864 49020 20916 49072
rect 25096 49020 25148 49072
rect 38252 49020 38304 49072
rect 40000 49020 40052 49072
rect 100260 49020 100312 49072
rect 45060 48952 45112 49004
rect 46808 48952 46860 49004
rect 100352 48952 100404 49004
rect 104216 48952 104268 49004
rect 36136 48884 36188 48936
rect 37240 48884 37292 48936
rect 43680 48884 43732 48936
rect 44692 48884 44744 48936
rect 45152 48884 45204 48936
rect 46072 48884 46124 48936
rect 46440 48884 46492 48936
rect 47452 48884 47504 48936
rect 103020 48884 103072 48936
rect 104768 48884 104820 48936
rect 108632 48952 108684 49004
rect 109184 48952 109236 49004
rect 109736 48952 109788 49004
rect 110472 48952 110524 49004
rect 130988 48884 131040 48936
rect 192720 48884 192772 48936
rect 193364 48884 193416 48936
rect 96120 48816 96172 48868
rect 222252 48816 222304 48868
rect 112496 47456 112548 47508
rect 112588 47456 112640 47508
rect 197044 47456 197096 47508
rect 197228 47456 197280 47508
rect 198148 47456 198200 47508
rect 50764 46504 50816 46556
rect 61344 46504 61396 46556
rect 135128 46504 135180 46556
rect 151320 46504 151372 46556
rect 49936 46436 49988 46488
rect 58952 46436 59004 46488
rect 134760 46436 134812 46488
rect 145340 46436 145392 46488
rect 50580 46368 50632 46420
rect 62816 46368 62868 46420
rect 134944 46368 134996 46420
rect 146812 46368 146864 46420
rect 51040 46300 51092 46352
rect 64288 46300 64340 46352
rect 50856 46232 50908 46284
rect 65760 46232 65812 46284
rect 50672 46164 50724 46216
rect 67324 46164 67376 46216
rect 82964 46164 83016 46216
rect 93360 46300 93412 46352
rect 134852 46300 134904 46352
rect 148284 46300 148336 46352
rect 135036 46232 135088 46284
rect 149756 46232 149808 46284
rect 50948 46096 51000 46148
rect 68796 46096 68848 46148
rect 84068 46096 84120 46148
rect 94740 46164 94792 46216
rect 135404 46164 135456 46216
rect 140188 46164 140240 46216
rect 166960 46164 167012 46216
rect 176160 46164 176212 46216
rect 88944 46096 88996 46148
rect 96120 46096 96172 46148
rect 135312 46096 135364 46148
rect 152792 46096 152844 46148
rect 168432 46096 168484 46148
rect 177540 46096 177592 46148
rect 135404 45280 135456 45332
rect 140280 45280 140332 45332
rect 181036 45280 181088 45332
rect 185176 45280 185228 45332
rect 135404 45008 135456 45060
rect 142304 45008 142356 45060
rect 53248 44736 53300 44788
rect 59044 44736 59096 44788
rect 135404 44736 135456 44788
rect 142212 44736 142264 44788
rect 53340 44668 53392 44720
rect 58216 44668 58268 44720
rect 92808 44668 92860 44720
rect 101732 44668 101784 44720
rect 140188 44668 140240 44720
rect 143684 44668 143736 44720
rect 177724 44668 177776 44720
rect 185912 44668 185964 44720
rect 92716 44600 92768 44652
rect 101364 44600 101416 44652
rect 140280 44396 140332 44448
rect 143500 44396 143552 44448
rect 177724 43852 177776 43904
rect 181036 43852 181088 43904
rect 50028 43512 50080 43564
rect 49936 43308 49988 43360
rect 98144 43444 98196 43496
rect 101640 43444 101692 43496
rect 135220 43376 135272 43428
rect 136968 43376 137020 43428
rect 135404 43308 135456 43360
rect 58216 43240 58268 43292
rect 92716 43240 92768 43292
rect 101824 43240 101876 43292
rect 181864 43308 181916 43360
rect 185176 43308 185228 43360
rect 142764 43240 142816 43292
rect 177816 43240 177868 43292
rect 185452 43240 185504 43292
rect 58308 43172 58360 43224
rect 92900 43172 92952 43224
rect 101272 43172 101324 43224
rect 177724 43172 177776 43224
rect 185820 43172 185872 43224
rect 92808 43104 92860 43156
rect 98144 43104 98196 43156
rect 49936 42424 49988 42476
rect 56284 42424 56336 42476
rect 177724 42356 177776 42408
rect 181864 42356 181916 42408
rect 50028 42288 50080 42340
rect 56652 42288 56704 42340
rect 135220 42152 135272 42204
rect 136876 42152 136928 42204
rect 49936 41948 49988 42000
rect 58400 41948 58452 42000
rect 135404 41948 135456 42000
rect 14700 41880 14752 41932
rect 18104 41880 18156 41932
rect 56652 41880 56704 41932
rect 58216 41880 58268 41932
rect 92808 41880 92860 41932
rect 101732 41880 101784 41932
rect 143316 41880 143368 41932
rect 177632 41880 177684 41932
rect 185176 41880 185228 41932
rect 92716 41812 92768 41864
rect 100812 41812 100864 41864
rect 136968 41812 137020 41864
rect 143408 41812 143460 41864
rect 177724 41812 177776 41864
rect 184992 41812 185044 41864
rect 56284 41608 56336 41660
rect 58308 41608 58360 41660
rect 135220 40792 135272 40844
rect 136968 40792 137020 40844
rect 49936 40656 49988 40708
rect 56652 40656 56704 40708
rect 50028 40588 50080 40640
rect 56560 40588 56612 40640
rect 135404 40588 135456 40640
rect 92808 40520 92860 40572
rect 100996 40520 101048 40572
rect 142488 40520 142540 40572
rect 177264 40520 177316 40572
rect 185176 40520 185228 40572
rect 92716 40452 92768 40504
rect 100904 40452 100956 40504
rect 136876 40452 136928 40504
rect 143684 40452 143736 40504
rect 177724 40452 177776 40504
rect 185084 40452 185136 40504
rect 56560 40112 56612 40164
rect 58216 40112 58268 40164
rect 51224 39228 51276 39280
rect 56744 39228 56796 39280
rect 135220 39228 135272 39280
rect 51132 39160 51184 39212
rect 135404 39160 135456 39212
rect 92900 39092 92952 39144
rect 100996 39092 101048 39144
rect 56652 39024 56704 39076
rect 58308 39024 58360 39076
rect 92808 39024 92860 39076
rect 101088 39024 101140 39076
rect 142856 39092 142908 39144
rect 177724 39092 177776 39144
rect 185176 39092 185228 39144
rect 143408 39024 143460 39076
rect 177356 39024 177408 39076
rect 185268 39024 185320 39076
rect 58216 38956 58268 39008
rect 92716 38956 92768 39008
rect 100812 38956 100864 39008
rect 136968 38956 137020 39008
rect 143684 38956 143736 39008
rect 177264 38956 177316 39008
rect 184992 38956 185044 39008
rect 56744 38616 56796 38668
rect 58400 38616 58452 38668
rect 98972 38344 99024 38396
rect 101180 38344 101232 38396
rect 98880 38208 98932 38260
rect 100996 38208 101048 38260
rect 135404 38208 135456 38260
rect 139636 38208 139688 38260
rect 183244 38072 183296 38124
rect 185268 38072 185320 38124
rect 51224 37868 51276 37920
rect 58308 37868 58360 37920
rect 135404 37868 135456 37920
rect 136876 37868 136928 37920
rect 51132 37800 51184 37852
rect 58216 37800 58268 37852
rect 135220 37800 135272 37852
rect 92808 37732 92860 37784
rect 98880 37732 98932 37784
rect 92716 37664 92768 37716
rect 98972 37664 99024 37716
rect 183704 37800 183756 37852
rect 185176 37800 185228 37852
rect 143684 37460 143736 37512
rect 177724 37324 177776 37376
rect 183244 37324 183296 37376
rect 139636 37188 139688 37240
rect 143500 37188 143552 37240
rect 177448 36848 177500 36900
rect 183704 36848 183756 36900
rect 51132 36576 51184 36628
rect 55548 36576 55600 36628
rect 134668 36576 134720 36628
rect 136784 36576 136836 36628
rect 51224 36508 51276 36560
rect 58308 36508 58360 36560
rect 50212 36440 50264 36492
rect 58216 36440 58268 36492
rect 135404 36440 135456 36492
rect 92808 36372 92860 36424
rect 100996 36372 101048 36424
rect 143040 36372 143092 36424
rect 177356 36372 177408 36424
rect 185176 36372 185228 36424
rect 92716 36304 92768 36356
rect 100536 36304 100588 36356
rect 177448 36304 177500 36356
rect 184992 36304 185044 36356
rect 136876 36236 136928 36288
rect 143684 36236 143736 36288
rect 51224 35352 51276 35404
rect 55456 35352 55508 35404
rect 135220 35216 135272 35268
rect 138164 35216 138216 35268
rect 51224 35080 51276 35132
rect 59228 35080 59280 35132
rect 135404 35080 135456 35132
rect 142396 35080 142448 35132
rect 92808 35012 92860 35064
rect 100996 35012 101048 35064
rect 136784 35012 136836 35064
rect 143684 35012 143736 35064
rect 177724 35012 177776 35064
rect 185452 35012 185504 35064
rect 55548 34944 55600 34996
rect 58308 34944 58360 34996
rect 92716 34944 92768 34996
rect 100904 34944 100956 34996
rect 177264 34944 177316 34996
rect 185084 34944 185136 34996
rect 55456 34740 55508 34792
rect 58216 34740 58268 34792
rect 134668 33788 134720 33840
rect 136968 33788 137020 33840
rect 51224 33720 51276 33772
rect 56468 33720 56520 33772
rect 135220 33720 135272 33772
rect 51132 33652 51184 33704
rect 56744 33652 56796 33704
rect 135404 33652 135456 33704
rect 92808 33584 92860 33636
rect 101088 33584 101140 33636
rect 92900 33516 92952 33568
rect 100996 33516 101048 33568
rect 143316 33584 143368 33636
rect 177816 33584 177868 33636
rect 185176 33584 185228 33636
rect 142764 33516 142816 33568
rect 177724 33516 177776 33568
rect 185268 33516 185320 33568
rect 92716 33448 92768 33500
rect 100720 33448 100772 33500
rect 138164 33448 138216 33500
rect 143684 33448 143736 33500
rect 177632 33448 177684 33500
rect 184900 33448 184952 33500
rect 56744 33380 56796 33432
rect 58216 33380 58268 33432
rect 56468 33040 56520 33092
rect 58308 33040 58360 33092
rect 50028 32496 50080 32548
rect 51224 32292 51276 32344
rect 135220 32360 135272 32412
rect 136876 32360 136928 32412
rect 135404 32292 135456 32344
rect 58216 32224 58268 32276
rect 92808 32224 92860 32276
rect 100996 32224 101048 32276
rect 142580 32224 142632 32276
rect 177632 32224 177684 32276
rect 185176 32224 185228 32276
rect 58308 32156 58360 32208
rect 92716 32156 92768 32208
rect 100812 32156 100864 32208
rect 136968 32156 137020 32208
rect 143684 32156 143736 32208
rect 177724 32156 177776 32208
rect 184992 32156 185044 32208
rect 50028 31272 50080 31324
rect 56744 31272 56796 31324
rect 51224 31136 51276 31188
rect 56652 31136 56704 31188
rect 135220 31136 135272 31188
rect 136968 31136 137020 31188
rect 51224 30932 51276 30984
rect 58400 30932 58452 30984
rect 135404 30932 135456 30984
rect 56652 30864 56704 30916
rect 58216 30864 58268 30916
rect 92808 30864 92860 30916
rect 100996 30864 101048 30916
rect 142764 30864 142816 30916
rect 177724 30864 177776 30916
rect 185176 30864 185228 30916
rect 56744 30796 56796 30848
rect 58308 30796 58360 30848
rect 92716 30796 92768 30848
rect 100904 30796 100956 30848
rect 136876 30796 136928 30848
rect 143684 30796 143736 30848
rect 177448 30796 177500 30848
rect 185084 30796 185136 30848
rect 51224 29640 51276 29692
rect 56008 29640 56060 29692
rect 135220 29572 135272 29624
rect 51132 29504 51184 29556
rect 135404 29504 135456 29556
rect 92900 29436 92952 29488
rect 101088 29436 101140 29488
rect 58216 29368 58268 29420
rect 92808 29368 92860 29420
rect 100996 29368 101048 29420
rect 143592 29436 143644 29488
rect 177724 29436 177776 29488
rect 185268 29436 185320 29488
rect 142764 29368 142816 29420
rect 177448 29368 177500 29420
rect 185176 29368 185228 29420
rect 92716 29300 92768 29352
rect 100812 29300 100864 29352
rect 136968 29300 137020 29352
rect 143684 29300 143736 29352
rect 177264 29300 177316 29352
rect 184992 29300 185044 29352
rect 56008 28892 56060 28944
rect 58308 28892 58360 28944
rect 135404 28416 135456 28468
rect 139636 28416 139688 28468
rect 51132 28280 51184 28332
rect 56376 28280 56428 28332
rect 135404 28280 135456 28332
rect 137336 28280 137388 28332
rect 51224 28144 51276 28196
rect 92900 28144 92952 28196
rect 100996 28144 101048 28196
rect 135220 28144 135272 28196
rect 92808 28076 92860 28128
rect 101916 28076 101968 28128
rect 56376 28008 56428 28060
rect 58308 28008 58360 28060
rect 92716 28008 92768 28060
rect 101732 28008 101784 28060
rect 58216 27940 58268 27992
rect 177632 28144 177684 28196
rect 185176 28144 185228 28196
rect 177356 28076 177408 28128
rect 185268 28076 185320 28128
rect 177724 28008 177776 28060
rect 185360 28008 185412 28060
rect 143684 27940 143736 27992
rect 139636 27532 139688 27584
rect 143408 27532 143460 27584
rect 51132 26920 51184 26972
rect 59044 26920 59096 26972
rect 135220 26920 135272 26972
rect 138164 26920 138216 26972
rect 51224 26852 51276 26904
rect 58308 26852 58360 26904
rect 50028 26784 50080 26836
rect 58216 26784 58268 26836
rect 92716 26716 92768 26768
rect 100996 26784 101048 26836
rect 135404 26784 135456 26836
rect 143592 26716 143644 26768
rect 177724 26716 177776 26768
rect 185176 26784 185228 26836
rect 137336 26580 137388 26632
rect 143684 26580 143736 26632
rect 51224 25492 51276 25544
rect 59412 25492 59464 25544
rect 135220 25492 135272 25544
rect 51132 25424 51184 25476
rect 59504 25424 59556 25476
rect 135404 25424 135456 25476
rect 50304 25356 50356 25408
rect 50672 25356 50724 25408
rect 92900 25356 92952 25408
rect 101180 25356 101232 25408
rect 92808 25288 92860 25340
rect 101088 25288 101140 25340
rect 143684 25356 143736 25408
rect 177356 25356 177408 25408
rect 185728 25356 185780 25408
rect 143500 25288 143552 25340
rect 177816 25288 177868 25340
rect 185268 25288 185320 25340
rect 92716 25220 92768 25272
rect 100996 25220 101048 25272
rect 138164 25220 138216 25272
rect 143132 25220 143184 25272
rect 177724 25220 177776 25272
rect 185820 25220 185872 25272
rect 134668 25016 134720 25068
rect 134944 25016 134996 25068
rect 51224 24064 51276 24116
rect 56100 24064 56152 24116
rect 135404 24064 135456 24116
rect 143592 24064 143644 24116
rect 51132 23996 51184 24048
rect 135036 23996 135088 24048
rect 143684 23996 143736 24048
rect 58216 23928 58268 23980
rect 92808 23928 92860 23980
rect 100996 23928 101048 23980
rect 177632 23928 177684 23980
rect 185176 23928 185228 23980
rect 92716 23860 92768 23912
rect 101088 23860 101140 23912
rect 177356 23860 177408 23912
rect 185268 23860 185320 23912
rect 56100 23452 56152 23504
rect 58308 23452 58360 23504
rect 97684 23112 97736 23164
rect 100996 23112 101048 23164
rect 135036 22908 135088 22960
rect 135312 22908 135364 22960
rect 135312 22772 135364 22824
rect 136876 22772 136928 22824
rect 51224 22704 51276 22756
rect 55732 22704 55784 22756
rect 134484 22704 134536 22756
rect 50396 22636 50448 22688
rect 98144 22636 98196 22688
rect 101088 22636 101140 22688
rect 135404 22636 135456 22688
rect 58216 22568 58268 22620
rect 90416 22568 90468 22620
rect 100996 22568 101048 22620
rect 96120 22500 96172 22552
rect 101088 22500 101140 22552
rect 142764 22568 142816 22620
rect 177632 22568 177684 22620
rect 185268 22772 185320 22824
rect 143316 22500 143368 22552
rect 177724 22500 177776 22552
rect 185176 22636 185228 22688
rect 92808 22432 92860 22484
rect 98144 22432 98196 22484
rect 174412 22432 174464 22484
rect 185176 22432 185228 22484
rect 92716 22364 92768 22416
rect 97684 22364 97736 22416
rect 55732 22160 55784 22212
rect 58308 22160 58360 22212
rect 50580 21276 50632 21328
rect 58216 21208 58268 21260
rect 92716 21208 92768 21260
rect 101180 21208 101232 21260
rect 136876 21208 136928 21260
rect 143684 21208 143736 21260
rect 177724 21208 177776 21260
rect 185268 21208 185320 21260
rect 93360 19780 93412 19832
rect 101088 19780 101140 19832
rect 176160 19780 176212 19832
rect 185268 19780 185320 19832
rect 94740 19712 94792 19764
rect 100996 19712 101048 19764
rect 177540 19712 177592 19764
rect 185176 19712 185228 19764
rect 18104 18420 18156 18472
rect 68244 18420 68296 18472
rect 69808 18420 69860 18472
rect 106700 18420 106752 18472
rect 153528 18420 153580 18472
rect 192536 18420 192588 18472
rect 211396 18420 211448 18472
rect 53984 18352 54036 18404
rect 71924 18352 71976 18404
rect 100260 18352 100312 18404
rect 112220 18352 112272 18404
rect 152240 18352 152292 18404
rect 60792 18284 60844 18336
rect 54812 18216 54864 18268
rect 76156 18284 76208 18336
rect 80664 18284 80716 18336
rect 88484 18284 88536 18336
rect 92716 18284 92768 18336
rect 156012 18284 156064 18336
rect 157576 18284 157628 18336
rect 161900 18284 161952 18336
rect 162636 18284 162688 18336
rect 163096 18284 163148 18336
rect 163648 18284 163700 18336
rect 167144 18284 167196 18336
rect 167788 18284 167840 18336
rect 171376 18284 171428 18336
rect 171928 18284 171980 18336
rect 81676 18216 81728 18268
rect 166316 18216 166368 18268
rect 168524 18216 168576 18268
rect 42852 18148 42904 18200
rect 72384 18148 72436 18200
rect 48832 18080 48884 18132
rect 83792 18080 83844 18132
rect 30800 18012 30852 18064
rect 74776 18012 74828 18064
rect 83056 18012 83108 18064
rect 36780 17944 36832 17996
rect 73396 17944 73448 17996
rect 138808 17944 138860 17996
rect 158496 17944 158548 17996
rect 165304 17944 165356 17996
rect 168984 17944 169036 17996
rect 24820 17876 24872 17928
rect 75512 17876 75564 17928
rect 132828 17876 132880 17928
rect 159508 17876 159560 17928
rect 18840 17808 18892 17860
rect 76524 17808 76576 17860
rect 126848 17808 126900 17860
rect 160520 17808 160572 17860
rect 12860 17740 12912 17792
rect 77536 17740 77588 17792
rect 120868 17740 120920 17792
rect 161716 17740 161768 17792
rect 89588 17536 89640 17588
rect 90784 17536 90836 17588
rect 169996 17536 170048 17588
rect 170916 17536 170968 17588
rect 67784 17060 67836 17112
rect 117832 17060 117884 17112
rect 151872 17060 151924 17112
rect 211120 17060 211172 17112
rect 163096 12708 163148 12760
rect 180852 12844 180904 12896
rect 168984 12640 169036 12692
rect 174872 12708 174924 12760
rect 174136 12640 174188 12692
rect 192812 12640 192864 12692
rect 172756 12572 172808 12624
rect 198792 12572 198844 12624
rect 161900 12504 161952 12556
rect 186832 12504 186884 12556
rect 92716 12436 92768 12488
rect 96856 12436 96908 12488
rect 171376 12436 171428 12488
rect 204864 12436 204916 12488
rect 87288 12368 87340 12420
rect 102836 12368 102888 12420
rect 168616 12368 168668 12420
rect 72844 12300 72896 12352
rect 79100 12300 79152 12352
rect 85816 12300 85868 12352
rect 108816 12300 108868 12352
rect 150860 12300 150912 12352
rect 156104 12300 156156 12352
rect 162820 12300 162872 12352
rect 165856 12300 165908 12352
rect 66864 12232 66916 12284
rect 76156 12232 76208 12284
rect 84436 12232 84488 12284
rect 114796 12232 114848 12284
rect 144788 12232 144840 12284
rect 156012 12232 156064 12284
rect 156840 12232 156892 12284
rect 167144 12232 167196 12284
rect 169996 12368 170048 12420
rect 210844 12368 210896 12420
rect 170088 12300 170140 12352
rect 216824 12300 216876 12352
rect 222804 12232 222856 12284
rect 84804 11824 84856 11876
rect 89864 11824 89916 11876
<< metal2 >>
rect 27854 244344 27910 244824
rect 63826 244344 63882 244824
rect 99798 244344 99854 244824
rect 135862 244344 135918 244824
rect 171834 244344 171890 244824
rect 207806 244344 207862 244824
rect 27868 241178 27896 244344
rect 63840 241178 63868 244344
rect 99812 244306 99840 244344
rect 99616 244300 99668 244306
rect 99616 244242 99668 244248
rect 99800 244300 99852 244306
rect 99800 244242 99852 244248
rect 89864 241376 89916 241382
rect 89864 241318 89916 241324
rect 27856 241172 27908 241178
rect 27856 241114 27908 241120
rect 29144 241172 29196 241178
rect 29144 241114 29196 241120
rect 63828 241172 63880 241178
rect 63828 241114 63880 241120
rect 65024 241172 65076 241178
rect 65024 241114 65076 241120
rect 22704 236684 22756 236690
rect 22704 236626 22756 236632
rect 22716 234802 22744 236626
rect 29156 235942 29184 241114
rect 49844 236684 49896 236690
rect 49844 236626 49896 236632
rect 39448 236616 39500 236622
rect 33374 236584 33430 236593
rect 39448 236558 39500 236564
rect 33374 236519 33430 236528
rect 29144 235936 29196 235942
rect 29144 235878 29196 235884
rect 28224 235188 28276 235194
rect 28224 235130 28276 235136
rect 28236 234802 28264 235130
rect 22408 234774 22744 234802
rect 27928 234774 28264 234802
rect 33388 234802 33416 236519
rect 39460 234802 39488 236558
rect 47268 235324 47320 235330
rect 47268 235266 47320 235272
rect 33388 234774 33540 234802
rect 39152 234774 39488 234802
rect 13320 233828 13372 233834
rect 13320 233770 13372 233776
rect 13332 232921 13360 233770
rect 13318 232912 13374 232921
rect 13318 232847 13374 232856
rect 14698 209384 14754 209393
rect 14698 209319 14754 209328
rect 13320 186840 13372 186846
rect 13320 186782 13372 186788
rect 13332 185729 13360 186782
rect 13318 185720 13374 185729
rect 13318 185655 13374 185664
rect 13412 182760 13464 182766
rect 13412 182702 13464 182708
rect 13320 175892 13372 175898
rect 13320 175834 13372 175840
rect 13332 138537 13360 175834
rect 13424 162201 13452 182702
rect 13410 162192 13466 162201
rect 13410 162127 13466 162136
rect 13318 138528 13374 138537
rect 13318 138463 13374 138472
rect 13318 115000 13374 115009
rect 13318 114935 13374 114944
rect 13332 97154 13360 114935
rect 13320 97148 13372 97154
rect 13320 97090 13372 97096
rect 13318 91336 13374 91345
rect 13318 91271 13374 91280
rect 13332 90286 13360 91271
rect 13320 90280 13372 90286
rect 13320 90222 13372 90228
rect 13320 82052 13372 82058
rect 13320 81994 13372 82000
rect 13332 67817 13360 81994
rect 13318 67808 13374 67817
rect 13318 67743 13374 67752
rect 13320 57912 13372 57918
rect 13320 57854 13372 57860
rect 13332 20625 13360 57854
rect 13412 57844 13464 57850
rect 13412 57786 13464 57792
rect 13424 44153 13452 57786
rect 13410 44144 13466 44153
rect 13410 44079 13466 44088
rect 14712 41938 14740 209319
rect 47280 207194 47308 235266
rect 49856 235262 49884 236626
rect 65036 235874 65064 241114
rect 72844 236684 72896 236690
rect 72844 236626 72896 236632
rect 65024 235868 65076 235874
rect 65024 235810 65076 235816
rect 65576 235324 65628 235330
rect 65576 235266 65628 235272
rect 49844 235256 49896 235262
rect 49844 235198 49896 235204
rect 62540 235256 62592 235262
rect 62540 235198 62592 235204
rect 47156 207166 47308 207194
rect 43416 207030 43936 207058
rect 19924 206894 20260 206922
rect 20568 206894 20904 206922
rect 21212 206894 21548 206922
rect 21856 206894 22192 206922
rect 22500 206894 22836 206922
rect 23144 206894 23480 206922
rect 23788 206894 24124 206922
rect 24432 206894 24768 206922
rect 25076 206894 25412 206922
rect 25720 206894 26240 206922
rect 26364 206894 26424 206922
rect 27008 206894 27252 206922
rect 27652 206894 27804 206922
rect 28296 206894 28632 206922
rect 28940 206894 29092 206922
rect 29676 206894 30012 206922
rect 30320 206894 30472 206922
rect 30964 206894 31300 206922
rect 31608 206894 31944 206922
rect 20232 204118 20260 206894
rect 20220 204112 20272 204118
rect 20220 204054 20272 204060
rect 20876 203506 20904 206894
rect 21520 204662 21548 206894
rect 21508 204656 21560 204662
rect 21508 204598 21560 204604
rect 22164 204322 22192 206894
rect 22808 204594 22836 206894
rect 22796 204588 22848 204594
rect 22796 204530 22848 204536
rect 23452 204526 23480 206894
rect 24096 204730 24124 206894
rect 24084 204724 24136 204730
rect 24084 204666 24136 204672
rect 23440 204520 23492 204526
rect 23440 204462 23492 204468
rect 24740 204390 24768 206894
rect 24728 204384 24780 204390
rect 24728 204326 24780 204332
rect 22152 204316 22204 204322
rect 22152 204258 22204 204264
rect 20864 203500 20916 203506
rect 20864 203442 20916 203448
rect 25384 203438 25412 206894
rect 25464 203500 25516 203506
rect 25464 203442 25516 203448
rect 25372 203432 25424 203438
rect 25372 203374 25424 203380
rect 25476 203114 25504 203442
rect 26108 203432 26160 203438
rect 26108 203374 26160 203380
rect 25384 203086 25504 203114
rect 25384 193594 25412 203086
rect 26120 202978 26148 203374
rect 26212 203114 26240 206894
rect 26212 203086 26332 203114
rect 26120 202950 26240 202978
rect 26212 195754 26240 202950
rect 26304 195822 26332 203086
rect 26396 195890 26424 206894
rect 26936 204656 26988 204662
rect 26936 204598 26988 204604
rect 26844 204588 26896 204594
rect 26844 204530 26896 204536
rect 26752 204520 26804 204526
rect 26752 204462 26804 204468
rect 26660 204316 26712 204322
rect 26660 204258 26712 204264
rect 26568 196360 26620 196366
rect 26568 196302 26620 196308
rect 26384 195884 26436 195890
rect 26384 195826 26436 195832
rect 26292 195816 26344 195822
rect 26292 195758 26344 195764
rect 26200 195748 26252 195754
rect 26200 195690 26252 195696
rect 26580 193730 26608 196302
rect 26502 193702 26608 193730
rect 26672 193730 26700 204258
rect 26764 196434 26792 204462
rect 26752 196428 26804 196434
rect 26752 196370 26804 196376
rect 26856 194138 26884 204530
rect 26948 196366 26976 204598
rect 27224 203438 27252 206894
rect 27212 203432 27264 203438
rect 27212 203374 27264 203380
rect 27672 203432 27724 203438
rect 27672 203374 27724 203380
rect 27396 196428 27448 196434
rect 27396 196370 27448 196376
rect 26936 196360 26988 196366
rect 26936 196302 26988 196308
rect 26856 194110 26976 194138
rect 26948 193730 26976 194110
rect 27408 193730 27436 196370
rect 27684 196298 27712 203374
rect 27776 196434 27804 206894
rect 28132 204724 28184 204730
rect 28132 204666 28184 204672
rect 28040 204384 28092 204390
rect 28040 204326 28092 204332
rect 27764 196428 27816 196434
rect 27764 196370 27816 196376
rect 28052 196366 28080 204326
rect 28040 196360 28092 196366
rect 28040 196302 28092 196308
rect 27672 196292 27724 196298
rect 27672 196234 27724 196240
rect 28144 193730 28172 204666
rect 28604 203438 28632 206894
rect 28592 203432 28644 203438
rect 28592 203374 28644 203380
rect 28224 196360 28276 196366
rect 28224 196302 28276 196308
rect 26672 193702 26870 193730
rect 26948 193702 27330 193730
rect 27408 193702 27698 193730
rect 28066 193702 28172 193730
rect 28236 193730 28264 196302
rect 28868 195748 28920 195754
rect 28868 195690 28920 195696
rect 28236 193702 28526 193730
rect 28880 193716 28908 195690
rect 29064 195278 29092 206894
rect 29984 203438 30012 206894
rect 29144 203432 29196 203438
rect 29144 203374 29196 203380
rect 29972 203432 30024 203438
rect 29972 203374 30024 203380
rect 29156 195482 29184 203374
rect 30156 196428 30208 196434
rect 30156 196370 30208 196376
rect 30064 196292 30116 196298
rect 30064 196234 30116 196240
rect 29696 195884 29748 195890
rect 29696 195826 29748 195832
rect 29236 195816 29288 195822
rect 29236 195758 29288 195764
rect 29144 195476 29196 195482
rect 29144 195418 29196 195424
rect 29052 195272 29104 195278
rect 29052 195214 29104 195220
rect 29248 193716 29276 195758
rect 29708 193716 29736 195826
rect 30076 193716 30104 196234
rect 30168 193730 30196 196370
rect 30444 195210 30472 206894
rect 31272 203438 31300 206894
rect 30524 203432 30576 203438
rect 30524 203374 30576 203380
rect 31260 203432 31312 203438
rect 31260 203374 31312 203380
rect 31812 203432 31864 203438
rect 31812 203374 31864 203380
rect 30536 196162 30564 203374
rect 30524 196156 30576 196162
rect 30524 196098 30576 196104
rect 31628 196156 31680 196162
rect 31628 196098 31680 196104
rect 30892 195476 30944 195482
rect 30892 195418 30944 195424
rect 30432 195204 30484 195210
rect 30432 195146 30484 195152
rect 30168 193702 30458 193730
rect 30904 193716 30932 195418
rect 31260 195272 31312 195278
rect 31260 195214 31312 195220
rect 31272 193716 31300 195214
rect 31640 193716 31668 196098
rect 31824 195226 31852 203374
rect 31916 195890 31944 206894
rect 32008 206894 32252 206922
rect 32896 206894 33324 206922
rect 31904 195884 31956 195890
rect 31904 195826 31956 195832
rect 32008 195754 32036 206894
rect 32824 195884 32876 195890
rect 32824 195826 32876 195832
rect 31996 195748 32048 195754
rect 31996 195690 32048 195696
rect 31824 195198 32220 195226
rect 32088 195136 32140 195142
rect 32088 195078 32140 195084
rect 32100 193716 32128 195078
rect 32192 193730 32220 195198
rect 32192 193702 32482 193730
rect 32836 193716 32864 195826
rect 32916 195748 32968 195754
rect 32916 195690 32968 195696
rect 32928 193730 32956 195690
rect 33296 195226 33324 206894
rect 33526 206650 33554 206908
rect 33480 206622 33554 206650
rect 33848 206894 34184 206922
rect 33376 203092 33428 203098
rect 33376 203034 33428 203040
rect 33388 195754 33416 203034
rect 33376 195748 33428 195754
rect 33376 195690 33428 195696
rect 33480 195550 33508 206622
rect 33848 203098 33876 206894
rect 34814 206650 34842 206908
rect 34768 206622 34842 206650
rect 35136 206894 35472 206922
rect 36116 206894 36176 206922
rect 33836 203092 33888 203098
rect 33836 203034 33888 203040
rect 34480 195748 34532 195754
rect 34480 195690 34532 195696
rect 33468 195544 33520 195550
rect 33468 195486 33520 195492
rect 34112 195544 34164 195550
rect 34112 195486 34164 195492
rect 33296 195198 33416 195226
rect 33388 193730 33416 195198
rect 32928 193702 33310 193730
rect 33388 193702 33678 193730
rect 34124 193716 34152 195486
rect 34492 193716 34520 195690
rect 34768 193730 34796 206622
rect 35136 193730 35164 206894
rect 36148 204474 36176 206894
rect 35964 204446 36176 204474
rect 36240 206894 36760 206922
rect 37068 206894 37404 206922
rect 37528 206894 38048 206922
rect 38448 206894 38784 206922
rect 38908 206894 39428 206922
rect 39644 206894 40072 206922
rect 40380 206894 40716 206922
rect 40840 206894 41360 206922
rect 41668 206894 42004 206922
rect 42312 206894 42648 206922
rect 43048 206894 43292 206922
rect 35964 193730 35992 204446
rect 36240 204338 36268 206894
rect 34768 193702 34874 193730
rect 35136 193702 35334 193730
rect 35702 193702 35992 193730
rect 36056 204310 36268 204338
rect 36056 193716 36084 204310
rect 37068 203114 37096 206894
rect 37528 203522 37556 206894
rect 36332 203086 37096 203114
rect 37344 203494 37556 203522
rect 36332 193730 36360 203086
rect 37344 195890 37372 203494
rect 38448 203438 38476 206894
rect 37424 203432 37476 203438
rect 37424 203374 37476 203380
rect 38436 203432 38488 203438
rect 38436 203374 38488 203380
rect 36872 195884 36924 195890
rect 36872 195826 36924 195832
rect 37332 195884 37384 195890
rect 37332 195826 37384 195832
rect 36332 193702 36530 193730
rect 36884 193716 36912 195826
rect 37436 193730 37464 203374
rect 38436 196360 38488 196366
rect 38436 196302 38488 196308
rect 38068 195680 38120 195686
rect 38068 195622 38120 195628
rect 37700 195476 37752 195482
rect 37700 195418 37752 195424
rect 37266 193702 37464 193730
rect 37712 193716 37740 195418
rect 38080 193716 38108 195622
rect 38448 193716 38476 196302
rect 38908 195482 38936 206894
rect 39644 203522 39672 206894
rect 39000 203494 39672 203522
rect 39000 195686 39028 203494
rect 40380 203438 40408 206894
rect 39540 203432 39592 203438
rect 39540 203374 39592 203380
rect 40368 203432 40420 203438
rect 40368 203374 40420 203380
rect 39552 196366 39580 203374
rect 39540 196360 39592 196366
rect 39540 196302 39592 196308
rect 40092 196360 40144 196366
rect 40092 196302 40144 196308
rect 39632 196224 39684 196230
rect 39632 196166 39684 196172
rect 39264 196020 39316 196026
rect 39264 195962 39316 195968
rect 38988 195680 39040 195686
rect 38988 195622 39040 195628
rect 38896 195476 38948 195482
rect 38896 195418 38948 195424
rect 38896 195340 38948 195346
rect 38896 195282 38948 195288
rect 38908 193716 38936 195282
rect 39276 193716 39304 195962
rect 39644 193716 39672 196166
rect 40104 193716 40132 196302
rect 40460 195680 40512 195686
rect 40460 195622 40512 195628
rect 40472 193716 40500 195622
rect 40840 195346 40868 206894
rect 40920 203568 40972 203574
rect 40920 203510 40972 203516
rect 40932 196366 40960 203510
rect 41104 203500 41156 203506
rect 41104 203442 41156 203448
rect 41012 203432 41064 203438
rect 41012 203374 41064 203380
rect 40920 196360 40972 196366
rect 40920 196302 40972 196308
rect 41024 196026 41052 203374
rect 41116 196230 41144 203442
rect 41668 203438 41696 206894
rect 41748 204112 41800 204118
rect 41748 204054 41800 204060
rect 41656 203432 41708 203438
rect 41656 203374 41708 203380
rect 41656 196360 41708 196366
rect 41656 196302 41708 196308
rect 41104 196224 41156 196230
rect 41104 196166 41156 196172
rect 41012 196020 41064 196026
rect 41012 195962 41064 195968
rect 41288 195884 41340 195890
rect 41288 195826 41340 195832
rect 40828 195340 40880 195346
rect 40828 195282 40880 195288
rect 40828 195204 40880 195210
rect 40828 195146 40880 195152
rect 40840 193716 40868 195146
rect 41300 193716 41328 195826
rect 41668 193716 41696 196302
rect 25384 193566 26134 193594
rect 22794 190480 22850 190489
rect 22794 190415 22850 190424
rect 22808 186846 22836 190415
rect 41760 189242 41788 204054
rect 42312 203506 42340 206894
rect 43048 203574 43076 206894
rect 43036 203568 43088 203574
rect 43036 203510 43088 203516
rect 42300 203500 42352 203506
rect 42300 203442 42352 203448
rect 43416 199306 43444 207030
rect 44428 206894 44580 206922
rect 44888 206894 45224 206922
rect 45868 206894 45928 206922
rect 43772 203500 43824 203506
rect 43772 203442 43824 203448
rect 43680 203432 43732 203438
rect 43680 203374 43732 203380
rect 43140 199278 43444 199306
rect 43140 195686 43168 199278
rect 43128 195680 43180 195686
rect 43128 195622 43180 195628
rect 43692 195210 43720 203374
rect 43784 195890 43812 203442
rect 44428 203438 44456 206894
rect 44888 203506 44916 206894
rect 45900 204458 45928 206894
rect 45060 204452 45112 204458
rect 45060 204394 45112 204400
rect 45888 204452 45940 204458
rect 45888 204394 45940 204400
rect 44876 203500 44928 203506
rect 44876 203442 44928 203448
rect 44416 203432 44468 203438
rect 44416 203374 44468 203380
rect 45072 196366 45100 204394
rect 45060 196360 45112 196366
rect 45060 196302 45112 196308
rect 43772 195884 43824 195890
rect 43772 195826 43824 195832
rect 43680 195204 43732 195210
rect 43680 195146 43732 195152
rect 41838 189256 41894 189265
rect 41760 189214 41838 189242
rect 41838 189191 41894 189200
rect 22796 186840 22848 186846
rect 22796 186782 22848 186788
rect 22334 183816 22390 183825
rect 22334 183751 22390 183760
rect 22348 182766 22376 183751
rect 22336 182760 22388 182766
rect 22336 182702 22388 182708
rect 23622 178784 23678 178793
rect 23622 178719 23678 178728
rect 22334 177152 22390 177161
rect 22334 177087 22390 177096
rect 22348 175898 22376 177087
rect 22336 175892 22388 175898
rect 22336 175834 22388 175840
rect 23636 170497 23664 178719
rect 23622 170488 23678 170497
rect 23622 170423 23678 170432
rect 49856 168894 49884 235198
rect 50578 234544 50634 234553
rect 50578 234479 50634 234488
rect 50026 232912 50082 232921
rect 50026 232847 50082 232856
rect 50040 232474 50068 232847
rect 50028 232468 50080 232474
rect 50028 232410 50080 232416
rect 50118 231688 50174 231697
rect 50118 231623 50174 231632
rect 50132 231182 50160 231623
rect 50120 231176 50172 231182
rect 50120 231118 50172 231124
rect 50026 225976 50082 225985
rect 50026 225911 50082 225920
rect 50040 225538 50068 225911
rect 50028 225532 50080 225538
rect 50028 225474 50080 225480
rect 50394 215096 50450 215105
rect 50394 215031 50450 215040
rect 50408 214930 50436 215031
rect 50396 214924 50448 214930
rect 50396 214866 50448 214872
rect 50394 214008 50450 214017
rect 50394 213943 50450 213952
rect 50408 213162 50436 213943
rect 50396 213156 50448 213162
rect 50396 213098 50448 213104
rect 50486 207752 50542 207761
rect 50486 207687 50542 207696
rect 50500 196502 50528 207687
rect 50592 207518 50620 234479
rect 51222 234000 51278 234009
rect 51222 233935 51224 233944
rect 51276 233935 51278 233944
rect 58124 233964 58176 233970
rect 51224 233906 51276 233912
rect 58124 233906 58176 233912
rect 51222 233456 51278 233465
rect 51222 233391 51278 233400
rect 51236 232610 51264 233391
rect 58136 233057 58164 233906
rect 58122 233048 58178 233057
rect 58122 232983 58178 232992
rect 62552 232762 62580 235198
rect 65588 232762 65616 235266
rect 72856 232762 72884 236626
rect 82228 235936 82280 235942
rect 82228 235878 82280 235884
rect 86184 235936 86236 235942
rect 86184 235878 86236 235884
rect 79558 235224 79614 235233
rect 75512 235188 75564 235194
rect 79558 235159 79614 235168
rect 75512 235130 75564 235136
rect 62552 232734 62612 232762
rect 65588 232734 65924 232762
rect 72548 232734 72884 232762
rect 75524 232762 75552 235130
rect 79572 232762 79600 235159
rect 75524 232734 75860 232762
rect 79264 232734 79600 232762
rect 82240 232762 82268 235878
rect 86196 232762 86224 235878
rect 89876 232762 89904 241318
rect 96120 236616 96172 236622
rect 96120 236558 96172 236564
rect 90232 233896 90284 233902
rect 90232 233838 90284 233844
rect 82240 232734 82576 232762
rect 85888 232734 86224 232762
rect 89200 232734 89904 232762
rect 51224 232604 51276 232610
rect 51224 232546 51276 232552
rect 58032 232604 58084 232610
rect 58032 232546 58084 232552
rect 50762 232232 50818 232241
rect 50762 232167 50818 232176
rect 50776 231114 50804 232167
rect 58044 231969 58072 232546
rect 58124 232468 58176 232474
rect 58124 232410 58176 232416
rect 58030 231960 58086 231969
rect 58030 231895 58086 231904
rect 58136 231289 58164 232410
rect 58122 231280 58178 231289
rect 58122 231215 58178 231224
rect 56468 231176 56520 231182
rect 51222 231144 51278 231153
rect 50764 231108 50816 231114
rect 56468 231118 56520 231124
rect 51222 231079 51278 231088
rect 50764 231050 50816 231056
rect 51236 231046 51264 231079
rect 51224 231040 51276 231046
rect 51224 230982 51276 230988
rect 52696 231040 52748 231046
rect 52696 230982 52748 230988
rect 51130 230600 51186 230609
rect 51130 230535 51186 230544
rect 51144 229754 51172 230535
rect 51222 230056 51278 230065
rect 51222 229991 51278 230000
rect 51236 229890 51264 229991
rect 51224 229884 51276 229890
rect 51224 229826 51276 229832
rect 51132 229748 51184 229754
rect 51132 229690 51184 229696
rect 52708 229618 52736 230982
rect 56480 230638 56508 231118
rect 58216 230972 58268 230978
rect 58216 230914 58268 230920
rect 58228 230745 58256 230914
rect 58214 230736 58270 230745
rect 58214 230671 58270 230680
rect 56468 230632 56520 230638
rect 56468 230574 56520 230580
rect 58216 230632 58268 230638
rect 58216 230574 58268 230580
rect 58228 230201 58256 230574
rect 58214 230192 58270 230201
rect 58214 230127 58270 230136
rect 56468 229884 56520 229890
rect 56468 229826 56520 229832
rect 56192 229748 56244 229754
rect 56192 229690 56244 229696
rect 52696 229612 52748 229618
rect 52696 229554 52748 229560
rect 51130 229376 51186 229385
rect 56204 229346 56232 229690
rect 51130 229311 51186 229320
rect 56192 229340 56244 229346
rect 51040 228456 51092 228462
rect 51040 228398 51092 228404
rect 51052 228297 51080 228398
rect 51144 228326 51172 229311
rect 56192 229282 56244 229288
rect 56480 229074 56508 229826
rect 58216 229612 58268 229618
rect 58216 229554 58268 229560
rect 58228 229521 58256 229554
rect 58214 229512 58270 229521
rect 58214 229447 58270 229456
rect 58216 229340 58268 229346
rect 58216 229282 58268 229288
rect 56468 229068 56520 229074
rect 56468 229010 56520 229016
rect 58228 228977 58256 229282
rect 58308 229068 58360 229074
rect 58308 229010 58360 229016
rect 58214 228968 58270 228977
rect 58214 228903 58270 228912
rect 51222 228832 51278 228841
rect 51222 228767 51278 228776
rect 51236 228394 51264 228767
rect 52696 228456 52748 228462
rect 52696 228398 52748 228404
rect 51224 228388 51276 228394
rect 51224 228330 51276 228336
rect 51132 228320 51184 228326
rect 51038 228288 51094 228297
rect 51132 228262 51184 228268
rect 51038 228223 51094 228232
rect 50762 227744 50818 227753
rect 50762 227679 50818 227688
rect 50776 226898 50804 227679
rect 51222 227200 51278 227209
rect 51278 227158 51356 227186
rect 51222 227135 51278 227144
rect 50764 226892 50816 226898
rect 50764 226834 50816 226840
rect 51222 226520 51278 226529
rect 51222 226455 51278 226464
rect 51236 225606 51264 226455
rect 51224 225600 51276 225606
rect 51224 225542 51276 225548
rect 51328 225470 51356 227158
rect 52708 226830 52736 228398
rect 55456 228388 55508 228394
rect 55456 228330 55508 228336
rect 55468 227918 55496 228330
rect 58320 228297 58348 229010
rect 58306 228288 58362 228297
rect 58216 228252 58268 228258
rect 58306 228223 58362 228232
rect 58216 228194 58268 228200
rect 55456 227912 55508 227918
rect 55456 227854 55508 227860
rect 58228 227753 58256 228194
rect 58308 227912 58360 227918
rect 58308 227854 58360 227860
rect 58214 227744 58270 227753
rect 58214 227679 58270 227688
rect 58320 227209 58348 227854
rect 58306 227200 58362 227209
rect 58306 227135 58362 227144
rect 55916 226892 55968 226898
rect 55916 226834 55968 226840
rect 52696 226824 52748 226830
rect 52696 226766 52748 226772
rect 55928 226422 55956 226834
rect 58216 226824 58268 226830
rect 58216 226766 58268 226772
rect 58228 226529 58256 226766
rect 58214 226520 58270 226529
rect 58214 226455 58270 226464
rect 55916 226416 55968 226422
rect 55916 226358 55968 226364
rect 58216 226416 58268 226422
rect 58216 226358 58268 226364
rect 58228 225985 58256 226358
rect 58214 225976 58270 225985
rect 58214 225911 58270 225920
rect 58308 225600 58360 225606
rect 58308 225542 58360 225548
rect 51316 225464 51368 225470
rect 51130 225432 51186 225441
rect 51316 225406 51368 225412
rect 58216 225464 58268 225470
rect 58216 225406 58268 225412
rect 51130 225367 51186 225376
rect 51144 224450 51172 225367
rect 58228 225305 58256 225406
rect 58214 225296 58270 225305
rect 58214 225231 58270 225240
rect 51222 224888 51278 224897
rect 51222 224823 51278 224832
rect 51132 224444 51184 224450
rect 51132 224386 51184 224392
rect 51130 224344 51186 224353
rect 51130 224279 51132 224288
rect 51184 224279 51186 224288
rect 51132 224250 51184 224256
rect 51236 224178 51264 224823
rect 58320 224761 58348 225542
rect 58400 225532 58452 225538
rect 58400 225474 58452 225480
rect 58306 224752 58362 224761
rect 58306 224687 58362 224696
rect 56744 224444 56796 224450
rect 56744 224386 56796 224392
rect 52696 224308 52748 224314
rect 52696 224250 52748 224256
rect 51224 224172 51276 224178
rect 51224 224114 51276 224120
rect 51222 223664 51278 223673
rect 51222 223599 51278 223608
rect 51130 223120 51186 223129
rect 51130 223055 51132 223064
rect 51184 223055 51186 223064
rect 51132 223026 51184 223032
rect 51236 222954 51264 223599
rect 51224 222948 51276 222954
rect 51224 222890 51276 222896
rect 52708 222750 52736 224250
rect 56756 224042 56784 224386
rect 58412 224217 58440 225474
rect 58398 224208 58454 224217
rect 58398 224143 58454 224152
rect 58216 224104 58268 224110
rect 58216 224046 58268 224052
rect 56744 224036 56796 224042
rect 56744 223978 56796 223984
rect 52788 223084 52840 223090
rect 52788 223026 52840 223032
rect 52696 222744 52748 222750
rect 52696 222686 52748 222692
rect 51222 222576 51278 222585
rect 51222 222511 51278 222520
rect 51130 222032 51186 222041
rect 51130 221967 51186 221976
rect 51144 221458 51172 221967
rect 51236 221730 51264 222511
rect 51224 221724 51276 221730
rect 51224 221666 51276 221672
rect 51222 221488 51278 221497
rect 51132 221452 51184 221458
rect 51222 221423 51278 221432
rect 51132 221394 51184 221400
rect 51236 221390 51264 221423
rect 51224 221384 51276 221390
rect 51224 221326 51276 221332
rect 52696 221384 52748 221390
rect 52696 221326 52748 221332
rect 51222 220808 51278 220817
rect 51222 220743 51278 220752
rect 51130 220264 51186 220273
rect 51130 220199 51186 220208
rect 51144 220098 51172 220199
rect 51132 220092 51184 220098
rect 51132 220034 51184 220040
rect 51236 220030 51264 220743
rect 51224 220024 51276 220030
rect 51224 219966 51276 219972
rect 52708 219962 52736 221326
rect 52800 221322 52828 223026
rect 58228 222993 58256 224046
rect 58308 224036 58360 224042
rect 58308 223978 58360 223984
rect 58320 223537 58348 223978
rect 58306 223528 58362 223537
rect 58306 223463 58362 223472
rect 58214 222984 58270 222993
rect 55824 222948 55876 222954
rect 58214 222919 58270 222928
rect 55824 222890 55876 222896
rect 55836 222342 55864 222890
rect 58216 222744 58268 222750
rect 58216 222686 58268 222692
rect 55824 222336 55876 222342
rect 58228 222313 58256 222686
rect 58308 222336 58360 222342
rect 55824 222278 55876 222284
rect 58214 222304 58270 222313
rect 58308 222278 58360 222284
rect 58214 222239 58270 222248
rect 58320 221769 58348 222278
rect 58306 221760 58362 221769
rect 56008 221724 56060 221730
rect 58306 221695 58362 221704
rect 56008 221666 56060 221672
rect 52788 221316 52840 221322
rect 52788 221258 52840 221264
rect 56020 221118 56048 221666
rect 56468 221452 56520 221458
rect 56468 221394 56520 221400
rect 56008 221112 56060 221118
rect 56008 221054 56060 221060
rect 56480 220710 56508 221394
rect 58216 221316 58268 221322
rect 58216 221258 58268 221264
rect 58228 221225 58256 221258
rect 58214 221216 58270 221225
rect 58214 221151 58270 221160
rect 58216 221112 58268 221118
rect 58216 221054 58268 221060
rect 56468 220704 56520 220710
rect 56468 220646 56520 220652
rect 58228 220545 58256 221054
rect 58308 220704 58360 220710
rect 58308 220646 58360 220652
rect 58214 220536 58270 220545
rect 58214 220471 58270 220480
rect 52788 220092 52840 220098
rect 52788 220034 52840 220040
rect 52696 219956 52748 219962
rect 52696 219898 52748 219904
rect 50854 219720 50910 219729
rect 50854 219655 50910 219664
rect 50868 218670 50896 219655
rect 52800 219434 52828 220034
rect 55824 220024 55876 220030
rect 58320 220001 58348 220646
rect 55824 219966 55876 219972
rect 58306 219992 58362 220001
rect 52708 219406 52828 219434
rect 51222 219176 51278 219185
rect 51222 219111 51278 219120
rect 51236 218874 51264 219111
rect 51224 218868 51276 218874
rect 51224 218810 51276 218816
rect 51224 218732 51276 218738
rect 51224 218674 51276 218680
rect 50856 218664 50908 218670
rect 51236 218641 51264 218674
rect 50856 218606 50908 218612
rect 51222 218632 51278 218641
rect 52708 218602 52736 219406
rect 55836 219350 55864 219966
rect 58216 219956 58268 219962
rect 58306 219927 58362 219936
rect 58216 219898 58268 219904
rect 55824 219344 55876 219350
rect 58228 219321 58256 219898
rect 58308 219344 58360 219350
rect 55824 219286 55876 219292
rect 58214 219312 58270 219321
rect 58308 219286 58360 219292
rect 58214 219247 58270 219256
rect 53340 218868 53392 218874
rect 53340 218810 53392 218816
rect 52788 218732 52840 218738
rect 52788 218674 52840 218680
rect 51222 218567 51278 218576
rect 52696 218596 52748 218602
rect 52696 218538 52748 218544
rect 50762 217952 50818 217961
rect 50762 217887 50818 217896
rect 50776 217242 50804 217887
rect 51222 217408 51278 217417
rect 51222 217343 51224 217352
rect 51276 217343 51278 217352
rect 51224 217314 51276 217320
rect 50764 217236 50816 217242
rect 50764 217178 50816 217184
rect 52696 217236 52748 217242
rect 52696 217178 52748 217184
rect 51130 216864 51186 216873
rect 51130 216799 51186 216808
rect 51144 215882 51172 216799
rect 51222 216320 51278 216329
rect 51278 216278 51356 216306
rect 51222 216255 51278 216264
rect 51132 215876 51184 215882
rect 51132 215818 51184 215824
rect 51222 215776 51278 215785
rect 51222 215711 51278 215720
rect 51132 214584 51184 214590
rect 51130 214552 51132 214561
rect 51184 214552 51186 214561
rect 51236 214522 51264 215711
rect 51130 214487 51186 214496
rect 51224 214516 51276 214522
rect 51224 214458 51276 214464
rect 51328 214454 51356 216278
rect 52708 215814 52736 217178
rect 52800 217106 52828 218674
rect 52880 217372 52932 217378
rect 52880 217314 52932 217320
rect 52788 217100 52840 217106
rect 52788 217042 52840 217048
rect 52696 215808 52748 215814
rect 52696 215750 52748 215756
rect 52892 215746 52920 217314
rect 53352 217174 53380 218810
rect 58320 218777 58348 219286
rect 58306 218768 58362 218777
rect 58306 218703 58362 218712
rect 55456 218664 55508 218670
rect 55456 218606 55508 218612
rect 55468 218058 55496 218606
rect 58216 218596 58268 218602
rect 58216 218538 58268 218544
rect 58228 218233 58256 218538
rect 58214 218224 58270 218233
rect 58214 218159 58270 218168
rect 55456 218052 55508 218058
rect 55456 217994 55508 218000
rect 58216 218052 58268 218058
rect 58216 217994 58268 218000
rect 58228 217553 58256 217994
rect 58214 217544 58270 217553
rect 58214 217479 58270 217488
rect 53340 217168 53392 217174
rect 53340 217110 53392 217116
rect 58216 217168 58268 217174
rect 58216 217110 58268 217116
rect 58228 217009 58256 217110
rect 58308 217100 58360 217106
rect 58308 217042 58360 217048
rect 58214 217000 58270 217009
rect 58214 216935 58270 216944
rect 58320 216329 58348 217042
rect 58306 216320 58362 216329
rect 58306 216255 58362 216264
rect 56468 215876 56520 215882
rect 56468 215818 56520 215824
rect 52880 215740 52932 215746
rect 52880 215682 52932 215688
rect 56480 215202 56508 215818
rect 58216 215808 58268 215814
rect 58214 215776 58216 215785
rect 58268 215776 58270 215785
rect 58214 215711 58270 215720
rect 58308 215740 58360 215746
rect 58308 215682 58360 215688
rect 58320 215241 58348 215682
rect 58306 215232 58362 215241
rect 56468 215196 56520 215202
rect 56468 215138 56520 215144
rect 58216 215196 58268 215202
rect 58306 215167 58362 215176
rect 58216 215138 58268 215144
rect 52788 214924 52840 214930
rect 52788 214866 52840 214872
rect 52696 214584 52748 214590
rect 52696 214526 52748 214532
rect 51316 214448 51368 214454
rect 51316 214390 51368 214396
rect 51222 213464 51278 213473
rect 51222 213399 51224 213408
rect 51276 213399 51278 213408
rect 51224 213370 51276 213376
rect 52708 213026 52736 214526
rect 52800 213094 52828 214866
rect 58228 214561 58256 215138
rect 58214 214552 58270 214561
rect 58214 214487 58270 214496
rect 58308 214516 58360 214522
rect 58308 214458 58360 214464
rect 58216 214448 58268 214454
rect 58216 214390 58268 214396
rect 58228 214017 58256 214390
rect 58214 214008 58270 214017
rect 58214 213943 58270 213952
rect 52880 213428 52932 213434
rect 52880 213370 52932 213376
rect 52788 213088 52840 213094
rect 52788 213030 52840 213036
rect 52696 213020 52748 213026
rect 52696 212962 52748 212968
rect 51222 212920 51278 212929
rect 51222 212855 51278 212864
rect 51130 212240 51186 212249
rect 51130 212175 51186 212184
rect 51144 212074 51172 212175
rect 51132 212068 51184 212074
rect 51132 212010 51184 212016
rect 51236 211802 51264 212855
rect 52696 212068 52748 212074
rect 52696 212010 52748 212016
rect 51224 211796 51276 211802
rect 51224 211738 51276 211744
rect 51222 211696 51278 211705
rect 51222 211631 51278 211640
rect 50854 211152 50910 211161
rect 50854 211087 50910 211096
rect 50670 210608 50726 210617
rect 50670 210543 50726 210552
rect 50580 207512 50632 207518
rect 50580 207454 50632 207460
rect 50488 196496 50540 196502
rect 50488 196438 50540 196444
rect 50684 195890 50712 210543
rect 50762 210064 50818 210073
rect 50762 209999 50818 210008
rect 50776 195958 50804 209999
rect 50764 195952 50816 195958
rect 50764 195894 50816 195900
rect 50672 195884 50724 195890
rect 50672 195826 50724 195832
rect 50868 195822 50896 211087
rect 51236 210578 51264 211631
rect 51224 210572 51276 210578
rect 51224 210514 51276 210520
rect 52708 210306 52736 212010
rect 52892 211598 52920 213370
rect 58320 213337 58348 214458
rect 58306 213328 58362 213337
rect 58306 213263 58362 213272
rect 52972 213156 53024 213162
rect 52972 213098 53024 213104
rect 52984 211666 53012 213098
rect 58216 213088 58268 213094
rect 58216 213030 58268 213036
rect 58228 212793 58256 213030
rect 58308 213020 58360 213026
rect 58308 212962 58360 212968
rect 58214 212784 58270 212793
rect 58214 212719 58270 212728
rect 58320 212249 58348 212962
rect 58306 212240 58362 212249
rect 58306 212175 58362 212184
rect 56284 211796 56336 211802
rect 56284 211738 56336 211744
rect 52972 211660 53024 211666
rect 52972 211602 53024 211608
rect 52880 211592 52932 211598
rect 52880 211534 52932 211540
rect 56296 211054 56324 211738
rect 58216 211660 58268 211666
rect 58216 211602 58268 211608
rect 58228 211569 58256 211602
rect 58308 211592 58360 211598
rect 58214 211560 58270 211569
rect 58308 211534 58360 211540
rect 58214 211495 58270 211504
rect 56284 211048 56336 211054
rect 58320 211025 58348 211534
rect 58400 211048 58452 211054
rect 56284 210990 56336 210996
rect 58306 211016 58362 211025
rect 58400 210990 58452 210996
rect 58306 210951 58362 210960
rect 56100 210572 56152 210578
rect 56100 210514 56152 210520
rect 52696 210300 52748 210306
rect 52696 210242 52748 210248
rect 56112 209898 56140 210514
rect 58412 210345 58440 210990
rect 58398 210336 58454 210345
rect 58216 210300 58268 210306
rect 58398 210271 58454 210280
rect 58216 210242 58268 210248
rect 56100 209892 56152 209898
rect 56100 209834 56152 209840
rect 58228 209801 58256 210242
rect 58308 209892 58360 209898
rect 58308 209834 58360 209840
rect 58214 209792 58270 209801
rect 58214 209727 58270 209736
rect 50946 209384 51002 209393
rect 50946 209319 51002 209328
rect 50960 196026 50988 209319
rect 58320 209257 58348 209834
rect 58306 209248 58362 209257
rect 90244 209234 90272 233838
rect 92716 233080 92768 233086
rect 92716 233022 92768 233028
rect 92728 232513 92756 233022
rect 92714 232504 92770 232513
rect 92714 232439 92770 232448
rect 94004 232400 94056 232406
rect 94004 232342 94056 232348
rect 94016 231969 94044 232342
rect 94002 231960 94058 231969
rect 94002 231895 94058 231904
rect 92716 231720 92768 231726
rect 92716 231662 92768 231668
rect 92728 231289 92756 231662
rect 92714 231280 92770 231289
rect 92714 231215 92770 231224
rect 92716 230972 92768 230978
rect 92716 230914 92768 230920
rect 92728 230201 92756 230914
rect 93728 230904 93780 230910
rect 93728 230846 93780 230852
rect 93740 230745 93768 230846
rect 93726 230736 93782 230745
rect 93726 230671 93782 230680
rect 92714 230192 92770 230201
rect 92714 230127 92770 230136
rect 92716 229612 92768 229618
rect 92716 229554 92768 229560
rect 92728 229521 92756 229554
rect 92808 229544 92860 229550
rect 92714 229512 92770 229521
rect 92808 229486 92860 229492
rect 92714 229447 92770 229456
rect 92820 228977 92848 229486
rect 92806 228968 92862 228977
rect 92716 228932 92768 228938
rect 92806 228903 92862 228912
rect 92716 228874 92768 228880
rect 92728 228297 92756 228874
rect 92714 228288 92770 228297
rect 92714 228223 92770 228232
rect 93176 228252 93228 228258
rect 93176 228194 93228 228200
rect 92716 228184 92768 228190
rect 92716 228126 92768 228132
rect 92728 227209 92756 228126
rect 93188 227753 93216 228194
rect 93174 227744 93230 227753
rect 93174 227679 93230 227688
rect 92714 227200 92770 227209
rect 92714 227135 92770 227144
rect 92716 226824 92768 226830
rect 92716 226766 92768 226772
rect 92728 226529 92756 226766
rect 92808 226756 92860 226762
rect 92808 226698 92860 226704
rect 92714 226520 92770 226529
rect 92714 226455 92770 226464
rect 92820 225985 92848 226698
rect 92806 225976 92862 225985
rect 92806 225911 92862 225920
rect 93728 225464 93780 225470
rect 93728 225406 93780 225412
rect 92808 225396 92860 225402
rect 92808 225338 92860 225344
rect 92716 225328 92768 225334
rect 92714 225296 92716 225305
rect 92768 225296 92770 225305
rect 92714 225231 92770 225240
rect 92820 224761 92848 225338
rect 92806 224752 92862 224761
rect 92806 224687 92862 224696
rect 93740 224217 93768 225406
rect 93726 224208 93782 224217
rect 93726 224143 93782 224152
rect 93912 224104 93964 224110
rect 93912 224046 93964 224052
rect 93728 224036 93780 224042
rect 93728 223978 93780 223984
rect 93740 223537 93768 223978
rect 93726 223528 93782 223537
rect 93726 223463 93782 223472
rect 93924 222993 93952 224046
rect 93910 222984 93966 222993
rect 93910 222919 93966 222928
rect 92716 222744 92768 222750
rect 92716 222686 92768 222692
rect 92728 222313 92756 222686
rect 92992 222676 93044 222682
rect 92992 222618 93044 222624
rect 92714 222304 92770 222313
rect 92714 222239 92770 222248
rect 93004 221769 93032 222618
rect 92990 221760 93046 221769
rect 92990 221695 93046 221704
rect 92808 221316 92860 221322
rect 92808 221258 92860 221264
rect 92714 221216 92770 221225
rect 92714 221151 92716 221160
rect 92768 221151 92770 221160
rect 92716 221122 92768 221128
rect 92820 220001 92848 221258
rect 93728 221248 93780 221254
rect 93728 221190 93780 221196
rect 93740 220545 93768 221190
rect 93726 220536 93782 220545
rect 93726 220471 93782 220480
rect 92806 219992 92862 220001
rect 92806 219927 92862 219936
rect 93728 219956 93780 219962
rect 93728 219898 93780 219904
rect 93740 219321 93768 219898
rect 93912 219888 93964 219894
rect 93912 219830 93964 219836
rect 93726 219312 93782 219321
rect 93726 219247 93782 219256
rect 93924 218777 93952 219830
rect 93910 218768 93966 218777
rect 93910 218703 93966 218712
rect 93544 218664 93596 218670
rect 93544 218606 93596 218612
rect 93176 218528 93228 218534
rect 93176 218470 93228 218476
rect 93188 218233 93216 218470
rect 93174 218224 93230 218233
rect 93174 218159 93230 218168
rect 92716 217168 92768 217174
rect 92716 217110 92768 217116
rect 92728 216329 92756 217110
rect 93556 217009 93584 218606
rect 93728 218596 93780 218602
rect 93728 218538 93780 218544
rect 93740 217553 93768 218538
rect 93726 217544 93782 217553
rect 93726 217479 93782 217488
rect 93542 217000 93598 217009
rect 93542 216935 93598 216944
rect 92714 216320 92770 216329
rect 92714 216255 92770 216264
rect 93544 215808 93596 215814
rect 92714 215776 92770 215785
rect 93544 215750 93596 215756
rect 92714 215711 92716 215720
rect 92768 215711 92770 215720
rect 92716 215682 92768 215688
rect 92808 215672 92860 215678
rect 92808 215614 92860 215620
rect 92820 215241 92848 215614
rect 92806 215232 92862 215241
rect 92806 215167 92862 215176
rect 93556 214561 93584 215750
rect 93542 214552 93598 214561
rect 93542 214487 93598 214496
rect 93360 214448 93412 214454
rect 93360 214390 93412 214396
rect 92716 214380 92768 214386
rect 92716 214322 92768 214328
rect 92728 214017 92756 214322
rect 92714 214008 92770 214017
rect 92714 213943 92770 213952
rect 93372 213337 93400 214390
rect 93358 213328 93414 213337
rect 93358 213263 93414 213272
rect 93360 213088 93412 213094
rect 93360 213030 93412 213036
rect 92716 213020 92768 213026
rect 92716 212962 92768 212968
rect 92728 212793 92756 212962
rect 92714 212784 92770 212793
rect 92714 212719 92770 212728
rect 93372 212249 93400 213030
rect 93358 212240 93414 212249
rect 93358 212175 93414 212184
rect 92808 211660 92860 211666
rect 92808 211602 92860 211608
rect 92716 211592 92768 211598
rect 92714 211560 92716 211569
rect 92768 211560 92770 211569
rect 92714 211495 92770 211504
rect 92820 211025 92848 211602
rect 92900 211524 92952 211530
rect 92900 211466 92952 211472
rect 92806 211016 92862 211025
rect 92806 210951 92862 210960
rect 92624 210368 92676 210374
rect 92912 210345 92940 211466
rect 94004 210436 94056 210442
rect 94004 210378 94056 210384
rect 92624 210310 92676 210316
rect 92898 210336 92954 210345
rect 90120 209206 90272 209234
rect 58306 209183 58362 209192
rect 83056 209008 83108 209014
rect 61264 208934 61600 208962
rect 64452 208934 65064 208962
rect 51038 208840 51094 208849
rect 51038 208775 51094 208784
rect 51052 196162 51080 208775
rect 51222 208296 51278 208305
rect 51222 208231 51278 208240
rect 51130 207208 51186 207217
rect 51130 207143 51186 207152
rect 51040 196156 51092 196162
rect 51040 196098 51092 196104
rect 50948 196020 51000 196026
rect 50948 195962 51000 195968
rect 50856 195816 50908 195822
rect 50856 195758 50908 195764
rect 51144 195482 51172 207143
rect 51236 196094 51264 208231
rect 61264 207518 61292 208934
rect 61252 207512 61304 207518
rect 61252 207454 61304 207460
rect 57572 196496 57624 196502
rect 57572 196438 57624 196444
rect 51224 196088 51276 196094
rect 51224 196030 51276 196036
rect 51132 195476 51184 195482
rect 51132 195418 51184 195424
rect 56468 195476 56520 195482
rect 56468 195418 56520 195424
rect 56480 193716 56508 195418
rect 57584 193716 57612 196438
rect 59780 196156 59832 196162
rect 59780 196098 59832 196104
rect 58676 196088 58728 196094
rect 58676 196030 58728 196036
rect 58688 193716 58716 196030
rect 59792 193716 59820 196098
rect 60884 196020 60936 196026
rect 60884 195962 60936 195968
rect 60896 193716 60924 195962
rect 61988 195952 62040 195958
rect 61988 195894 62040 195900
rect 62000 193716 62028 195894
rect 63092 195884 63144 195890
rect 63092 195826 63144 195832
rect 63104 193716 63132 195826
rect 65036 195822 65064 208934
rect 65128 208934 65832 208962
rect 66508 208934 67304 208962
rect 67888 208934 68684 208962
rect 69268 208934 70156 208962
rect 70648 208934 71536 208962
rect 72212 208934 73008 208962
rect 74052 208934 74388 208962
rect 75524 208934 75860 208962
rect 76904 208934 77240 208962
rect 78376 208934 78712 208962
rect 79756 208934 80092 208962
rect 81228 208934 81564 208962
rect 81688 208934 82944 208962
rect 83056 208950 83108 208956
rect 84252 209008 84304 209014
rect 91244 209008 91296 209014
rect 88758 208976 88814 208985
rect 84304 208956 84416 208962
rect 84252 208950 84416 208956
rect 64196 195816 64248 195822
rect 64196 195758 64248 195764
rect 65024 195816 65076 195822
rect 65024 195758 65076 195764
rect 64208 193716 64236 195758
rect 65128 193730 65156 208934
rect 66508 196314 66536 208934
rect 66416 196286 66536 196314
rect 65128 193702 65326 193730
rect 66416 193716 66444 196286
rect 67888 195226 67916 208934
rect 69268 195226 69296 208934
rect 70648 196366 70676 208934
rect 72016 196428 72068 196434
rect 72016 196370 72068 196376
rect 69808 196360 69860 196366
rect 69808 196302 69860 196308
rect 70636 196360 70688 196366
rect 70636 196302 70688 196308
rect 70912 196360 70964 196366
rect 70912 196302 70964 196308
rect 67796 195198 67916 195226
rect 68992 195198 69296 195226
rect 67796 193730 67824 195198
rect 68992 193730 69020 195198
rect 67534 193702 67824 193730
rect 68638 193702 69020 193730
rect 69820 193716 69848 196302
rect 70924 193716 70952 196302
rect 72028 193716 72056 196370
rect 72212 196366 72240 208934
rect 73212 206288 73264 206294
rect 73212 206230 73264 206236
rect 72200 196360 72252 196366
rect 72200 196302 72252 196308
rect 73224 193730 73252 206230
rect 74052 206226 74080 208934
rect 75524 206294 75552 208934
rect 76800 206356 76852 206362
rect 76800 206298 76852 206304
rect 75512 206288 75564 206294
rect 75512 206230 75564 206236
rect 73304 206220 73356 206226
rect 73304 206162 73356 206168
rect 74040 206220 74092 206226
rect 74040 206162 74092 206168
rect 74684 206220 74736 206226
rect 74684 206162 74736 206168
rect 73316 196434 73344 206162
rect 73304 196428 73356 196434
rect 73304 196370 73356 196376
rect 74696 193730 74724 206162
rect 76812 196366 76840 206298
rect 76904 206226 76932 208934
rect 78376 206362 78404 208934
rect 78364 206356 78416 206362
rect 78364 206298 78416 206304
rect 79756 206294 79784 208934
rect 78180 206288 78232 206294
rect 78180 206230 78232 206236
rect 79744 206288 79796 206294
rect 79744 206230 79796 206236
rect 76892 206220 76944 206226
rect 76892 206162 76944 206168
rect 75328 196360 75380 196366
rect 75328 196302 75380 196308
rect 76800 196360 76852 196366
rect 76800 196302 76852 196308
rect 73146 193702 73252 193730
rect 74250 193702 74724 193730
rect 75340 193716 75368 196302
rect 77536 195544 77588 195550
rect 77536 195486 77588 195492
rect 76432 195476 76484 195482
rect 76432 195418 76484 195424
rect 76444 193716 76472 195418
rect 77548 193716 77576 195486
rect 78192 195482 78220 206230
rect 81228 206226 81256 208934
rect 79560 206220 79612 206226
rect 79560 206162 79612 206168
rect 81216 206220 81268 206226
rect 81216 206162 81268 206168
rect 78640 196360 78692 196366
rect 78640 196302 78692 196308
rect 78180 195476 78232 195482
rect 78180 195418 78232 195424
rect 78652 193716 78680 196302
rect 79572 195550 79600 206162
rect 81688 196366 81716 208934
rect 81676 196360 81728 196366
rect 81676 196302 81728 196308
rect 80848 196292 80900 196298
rect 80848 196234 80900 196240
rect 79744 195748 79796 195754
rect 79744 195690 79796 195696
rect 79560 195544 79612 195550
rect 79560 195486 79612 195492
rect 79756 193716 79784 195690
rect 80860 193716 80888 196234
rect 81952 195952 82004 195958
rect 81952 195894 82004 195900
rect 81964 193716 81992 195894
rect 83068 195754 83096 208950
rect 84264 208934 84416 208950
rect 84540 208934 85796 208962
rect 87208 208934 87268 208962
rect 88648 208934 88758 208962
rect 84540 196298 84568 208934
rect 85724 206220 85776 206226
rect 85724 206162 85776 206168
rect 84528 196292 84580 196298
rect 84528 196234 84580 196240
rect 83056 195748 83108 195754
rect 83056 195690 83108 195696
rect 85736 193730 85764 206162
rect 87208 195958 87236 208934
rect 91244 208950 91296 208956
rect 88758 208911 88814 208920
rect 89772 196088 89824 196094
rect 89772 196030 89824 196036
rect 88668 196020 88720 196026
rect 88668 195962 88720 195968
rect 87196 195952 87248 195958
rect 87196 195894 87248 195900
rect 87564 195952 87616 195958
rect 87564 195894 87616 195900
rect 86460 195884 86512 195890
rect 86460 195826 86512 195832
rect 85382 193702 85764 193730
rect 86472 193716 86500 195826
rect 87576 193716 87604 195894
rect 88680 193716 88708 195962
rect 89784 193716 89812 196030
rect 91256 193730 91284 208950
rect 92636 195754 92664 210310
rect 92898 210271 92954 210280
rect 93176 210300 93228 210306
rect 93176 210242 93228 210248
rect 92716 210232 92768 210238
rect 92716 210174 92768 210180
rect 92728 209257 92756 210174
rect 93188 209801 93216 210242
rect 93174 209792 93230 209801
rect 93174 209727 93230 209736
rect 92714 209248 92770 209257
rect 92714 209183 92770 209192
rect 94016 196366 94044 210378
rect 93084 196360 93136 196366
rect 93084 196302 93136 196308
rect 94004 196360 94056 196366
rect 94004 196302 94056 196308
rect 91980 195748 92032 195754
rect 91980 195690 92032 195696
rect 92624 195748 92676 195754
rect 92624 195690 92676 195696
rect 90902 193702 91284 193730
rect 91992 193716 92020 195690
rect 93096 193716 93124 196302
rect 94188 195816 94240 195822
rect 94188 195758 94240 195764
rect 94200 193716 94228 195758
rect 53338 173888 53394 173897
rect 53338 173823 53394 173832
rect 44416 168888 44468 168894
rect 44416 168830 44468 168836
rect 49844 168888 49896 168894
rect 49844 168830 49896 168836
rect 44428 168729 44456 168830
rect 44414 168720 44470 168729
rect 44414 168655 44470 168664
rect 49856 167602 49884 168830
rect 49844 167596 49896 167602
rect 49844 167538 49896 167544
rect 53352 163833 53380 173823
rect 53432 167596 53484 167602
rect 53432 167538 53484 167544
rect 53338 163824 53394 163833
rect 53338 163759 53394 163768
rect 53444 160569 53472 167538
rect 53430 160560 53486 160569
rect 53430 160495 53486 160504
rect 44506 158792 44562 158801
rect 44506 158727 44562 158736
rect 25108 153854 26134 153882
rect 25004 151412 25056 151418
rect 25004 151354 25056 151360
rect 24912 151344 24964 151350
rect 24912 151286 24964 151292
rect 23256 143864 23308 143870
rect 23256 143806 23308 143812
rect 22152 143796 22204 143802
rect 22152 143738 22204 143744
rect 20772 143660 20824 143666
rect 20772 143602 20824 143608
rect 20496 143388 20548 143394
rect 20496 143330 20548 143336
rect 20508 140690 20536 143330
rect 20784 140826 20812 143602
rect 21784 142844 21836 142850
rect 21784 142786 21836 142792
rect 20784 140798 20890 140826
rect 21796 140690 21824 142786
rect 22164 140826 22192 143738
rect 22164 140798 22270 140826
rect 23268 140690 23296 143806
rect 24924 143734 24952 151286
rect 24452 143728 24504 143734
rect 24452 143670 24504 143676
rect 24912 143728 24964 143734
rect 24912 143670 24964 143676
rect 23532 143592 23584 143598
rect 23532 143534 23584 143540
rect 23544 140826 23572 143534
rect 23544 140798 23650 140826
rect 24464 140690 24492 143670
rect 25016 140690 25044 151354
rect 25108 143666 25136 153854
rect 26292 151752 26344 151758
rect 26292 151694 26344 151700
rect 25740 151208 25792 151214
rect 25740 151150 25792 151156
rect 25096 143660 25148 143666
rect 25096 143602 25148 143608
rect 25752 143598 25780 151150
rect 26016 151140 26068 151146
rect 26016 151082 26068 151088
rect 25924 151072 25976 151078
rect 25924 151014 25976 151020
rect 25832 151004 25884 151010
rect 25832 150946 25884 150952
rect 25740 143592 25792 143598
rect 25740 143534 25792 143540
rect 25844 142850 25872 150946
rect 25936 143802 25964 151014
rect 26028 143870 26056 151082
rect 26016 143864 26068 143870
rect 26016 143806 26068 143812
rect 25924 143796 25976 143802
rect 25924 143738 25976 143744
rect 26016 143660 26068 143666
rect 26016 143602 26068 143608
rect 25832 142844 25884 142850
rect 25832 142786 25884 142792
rect 26028 140690 26056 143602
rect 26304 140962 26332 151694
rect 26384 151276 26436 151282
rect 26384 151218 26436 151224
rect 26396 143666 26424 151218
rect 26488 151010 26516 153868
rect 26856 151078 26884 153868
rect 27316 151146 27344 153868
rect 27684 151214 27712 153868
rect 27764 152364 27816 152370
rect 27764 152306 27816 152312
rect 27672 151208 27724 151214
rect 27672 151150 27724 151156
rect 27304 151140 27356 151146
rect 27304 151082 27356 151088
rect 26844 151072 26896 151078
rect 26844 151014 26896 151020
rect 27672 151072 27724 151078
rect 27672 151014 27724 151020
rect 26476 151004 26528 151010
rect 26476 150946 26528 150952
rect 26384 143660 26436 143666
rect 26384 143602 26436 143608
rect 27304 143660 27356 143666
rect 27304 143602 27356 143608
rect 26304 140934 26424 140962
rect 26396 140690 26424 140934
rect 27316 140690 27344 143602
rect 27684 140962 27712 151014
rect 27776 143666 27804 152306
rect 28052 151350 28080 153868
rect 28512 151418 28540 153868
rect 28500 151412 28552 151418
rect 28500 151354 28552 151360
rect 28040 151344 28092 151350
rect 28040 151286 28092 151292
rect 28880 151282 28908 153868
rect 29144 152228 29196 152234
rect 29144 152170 29196 152176
rect 29052 151412 29104 151418
rect 29052 151354 29104 151360
rect 28868 151276 28920 151282
rect 28868 151218 28920 151224
rect 29064 143666 29092 151354
rect 27764 143660 27816 143666
rect 27764 143602 27816 143608
rect 28592 143660 28644 143666
rect 28592 143602 28644 143608
rect 29052 143660 29104 143666
rect 29052 143602 29104 143608
rect 27684 140934 27804 140962
rect 27776 140690 27804 140934
rect 28604 140690 28632 143602
rect 29156 140690 29184 152170
rect 29248 151758 29276 153868
rect 29708 152370 29736 153868
rect 29696 152364 29748 152370
rect 29696 152306 29748 152312
rect 29236 151752 29288 151758
rect 29236 151694 29288 151700
rect 30076 151078 30104 153868
rect 30168 153854 30458 153882
rect 30168 151418 30196 153854
rect 30524 152364 30576 152370
rect 30524 152306 30576 152312
rect 30432 152296 30484 152302
rect 30432 152238 30484 152244
rect 30156 151412 30208 151418
rect 30156 151354 30208 151360
rect 30064 151072 30116 151078
rect 30064 151014 30116 151020
rect 30064 143660 30116 143666
rect 30064 143602 30116 143608
rect 30076 140690 30104 143602
rect 30444 140962 30472 152238
rect 30536 143666 30564 152306
rect 30904 152234 30932 153868
rect 31272 152370 31300 153868
rect 31260 152364 31312 152370
rect 31260 152306 31312 152312
rect 31640 152302 31668 153868
rect 32008 153854 32114 153882
rect 31628 152296 31680 152302
rect 32008 152250 32036 153854
rect 32088 152364 32140 152370
rect 32088 152306 32140 152312
rect 31628 152238 31680 152244
rect 30892 152228 30944 152234
rect 30892 152170 30944 152176
rect 31916 152222 32036 152250
rect 31812 151888 31864 151894
rect 31812 151830 31864 151836
rect 30524 143660 30576 143666
rect 30524 143602 30576 143608
rect 31352 142844 31404 142850
rect 31352 142786 31404 142792
rect 30444 140934 30564 140962
rect 30536 140690 30564 140934
rect 31364 140690 31392 142786
rect 31824 140962 31852 151830
rect 31916 142850 31944 152222
rect 31996 151276 32048 151282
rect 31996 151218 32048 151224
rect 32008 143666 32036 151218
rect 31996 143660 32048 143666
rect 31996 143602 32048 143608
rect 31904 142844 31956 142850
rect 31904 142786 31956 142792
rect 31824 140934 31944 140962
rect 31916 140690 31944 140934
rect 32100 140826 32128 152306
rect 32468 151894 32496 153868
rect 32836 152370 32864 153868
rect 32824 152364 32876 152370
rect 32824 152306 32876 152312
rect 32456 151888 32508 151894
rect 32456 151830 32508 151836
rect 33296 151282 33324 153868
rect 33388 153854 33678 153882
rect 33284 151276 33336 151282
rect 33284 151218 33336 151224
rect 32732 143660 32784 143666
rect 32732 143602 32784 143608
rect 32744 140826 32772 143602
rect 33388 140826 33416 153854
rect 34124 151010 34152 153868
rect 33468 151004 33520 151010
rect 33468 150946 33520 150952
rect 34112 151004 34164 151010
rect 34112 150946 34164 150952
rect 33480 140962 33508 150946
rect 34492 143666 34520 153868
rect 34480 143660 34532 143666
rect 34480 143602 34532 143608
rect 34860 143598 34888 153868
rect 35320 151146 35348 153868
rect 35308 151140 35360 151146
rect 35308 151082 35360 151088
rect 34940 143660 34992 143666
rect 34940 143602 34992 143608
rect 34848 143592 34900 143598
rect 34848 143534 34900 143540
rect 33480 140934 33968 140962
rect 32100 140798 32482 140826
rect 32744 140798 33126 140826
rect 33388 140798 33862 140826
rect 20246 140662 20536 140690
rect 21534 140662 21824 140690
rect 22914 140662 23296 140690
rect 24294 140662 24492 140690
rect 24938 140662 25044 140690
rect 25674 140662 26056 140690
rect 26318 140662 26424 140690
rect 27054 140662 27344 140690
rect 27698 140662 27804 140690
rect 28342 140662 28632 140690
rect 29078 140662 29184 140690
rect 29722 140662 30104 140690
rect 30458 140662 30564 140690
rect 31102 140662 31392 140690
rect 31838 140662 31944 140690
rect 33940 140690 33968 140934
rect 34952 140826 34980 143602
rect 35492 143592 35544 143598
rect 35492 143534 35544 143540
rect 35504 140826 35532 143534
rect 35688 143530 35716 153868
rect 36056 151486 36084 153868
rect 36044 151480 36096 151486
rect 36044 151422 36096 151428
rect 36516 151214 36544 153868
rect 36884 152166 36912 153868
rect 37252 152370 37280 153868
rect 37240 152364 37292 152370
rect 37240 152306 37292 152312
rect 36872 152160 36924 152166
rect 36872 152102 36924 152108
rect 37712 151622 37740 153868
rect 38080 151758 38108 153868
rect 38448 152234 38476 153868
rect 38908 152302 38936 153868
rect 39276 152370 39304 153868
rect 38988 152364 39040 152370
rect 38988 152306 39040 152312
rect 39264 152364 39316 152370
rect 39264 152306 39316 152312
rect 38896 152296 38948 152302
rect 38896 152238 38948 152244
rect 38436 152228 38488 152234
rect 38436 152170 38488 152176
rect 38896 152160 38948 152166
rect 38896 152102 38948 152108
rect 38068 151752 38120 151758
rect 38068 151694 38120 151700
rect 37700 151616 37752 151622
rect 37700 151558 37752 151564
rect 37608 151480 37660 151486
rect 37608 151422 37660 151428
rect 36504 151208 36556 151214
rect 36504 151150 36556 151156
rect 37424 151208 37476 151214
rect 37424 151150 37476 151156
rect 36044 151140 36096 151146
rect 36044 151082 36096 151088
rect 35676 143524 35728 143530
rect 35676 143466 35728 143472
rect 36056 142730 36084 151082
rect 36964 143524 37016 143530
rect 36964 143466 37016 143472
rect 36056 142702 36176 142730
rect 36148 140826 36176 142702
rect 36976 140826 37004 143466
rect 37436 142850 37464 151150
rect 37424 142844 37476 142850
rect 37424 142786 37476 142792
rect 37620 140826 37648 151422
rect 38252 142844 38304 142850
rect 38252 142786 38304 142792
rect 38264 140826 38292 142786
rect 38908 140826 38936 152102
rect 39000 142594 39028 152306
rect 39644 143870 39672 153868
rect 39908 152296 39960 152302
rect 39908 152238 39960 152244
rect 39920 144006 39948 152238
rect 39908 144000 39960 144006
rect 39908 143942 39960 143948
rect 40104 143938 40132 153868
rect 40184 152364 40236 152370
rect 40184 152306 40236 152312
rect 40196 144074 40224 152306
rect 40472 151894 40500 153868
rect 40460 151888 40512 151894
rect 40460 151830 40512 151836
rect 40276 151616 40328 151622
rect 40276 151558 40328 151564
rect 40184 144068 40236 144074
rect 40184 144010 40236 144016
rect 40092 143932 40144 143938
rect 40092 143874 40144 143880
rect 39632 143864 39684 143870
rect 39632 143806 39684 143812
rect 39000 142566 39672 142594
rect 39644 140826 39672 142566
rect 40288 140826 40316 151558
rect 40840 151078 40868 153868
rect 40920 151752 40972 151758
rect 40920 151694 40972 151700
rect 40828 151072 40880 151078
rect 40828 151014 40880 151020
rect 40932 140826 40960 151694
rect 41300 151690 41328 153868
rect 41668 152370 41696 153868
rect 41656 152364 41708 152370
rect 41656 152306 41708 152312
rect 43680 152364 43732 152370
rect 43680 152306 43732 152312
rect 41840 152228 41892 152234
rect 41840 152170 41892 152176
rect 41288 151684 41340 151690
rect 41288 151626 41340 151632
rect 41852 140826 41880 152170
rect 43036 144068 43088 144074
rect 43036 144010 43088 144016
rect 42300 144000 42352 144006
rect 42300 143942 42352 143948
rect 42312 140826 42340 143942
rect 43048 140826 43076 144010
rect 43692 143666 43720 152306
rect 44416 143932 44468 143938
rect 44416 143874 44468 143880
rect 43772 143864 43824 143870
rect 43772 143806 43824 143812
rect 43680 143660 43732 143666
rect 43680 143602 43732 143608
rect 43784 140826 43812 143806
rect 44428 140826 44456 143874
rect 44520 143394 44548 158727
rect 44968 151888 45020 151894
rect 44968 151830 45020 151836
rect 44508 143388 44560 143394
rect 44508 143330 44560 143336
rect 44980 140826 45008 151830
rect 45152 151684 45204 151690
rect 45152 151626 45204 151632
rect 45060 151072 45112 151078
rect 45060 151014 45112 151020
rect 45072 142986 45100 151014
rect 45164 143258 45192 151626
rect 59240 146862 59268 153868
rect 69164 151752 69216 151758
rect 69164 151694 69216 151700
rect 59228 146856 59280 146862
rect 59228 146798 59280 146804
rect 59412 146788 59464 146794
rect 59412 146730 59464 146736
rect 59424 144074 59452 146730
rect 59412 144068 59464 144074
rect 59412 144010 59464 144016
rect 47176 143660 47228 143666
rect 47176 143602 47228 143608
rect 45152 143252 45204 143258
rect 45152 143194 45204 143200
rect 46532 143252 46584 143258
rect 46532 143194 46584 143200
rect 45060 142980 45112 142986
rect 45060 142922 45112 142928
rect 45796 142980 45848 142986
rect 45796 142922 45848 142928
rect 45808 140826 45836 142922
rect 46544 140826 46572 143194
rect 47188 140826 47216 143602
rect 69176 142714 69204 151694
rect 72580 151622 72608 153868
rect 79204 151826 79232 153868
rect 79192 151820 79244 151826
rect 79192 151762 79244 151768
rect 92544 151758 92572 153868
rect 92532 151752 92584 151758
rect 92532 151694 92584 151700
rect 95384 151752 95436 151758
rect 95384 151694 95436 151700
rect 72568 151616 72620 151622
rect 72568 151558 72620 151564
rect 68704 142708 68756 142714
rect 68704 142650 68756 142656
rect 69164 142708 69216 142714
rect 69164 142650 69216 142656
rect 34952 140798 35242 140826
rect 35504 140798 35886 140826
rect 36148 140798 36530 140826
rect 36976 140798 37266 140826
rect 37620 140798 37910 140826
rect 38264 140798 38646 140826
rect 38908 140798 39290 140826
rect 39644 140798 40026 140826
rect 40288 140798 40670 140826
rect 40932 140798 41314 140826
rect 41852 140798 42050 140826
rect 42312 140798 42694 140826
rect 43048 140798 43430 140826
rect 43784 140798 44074 140826
rect 44428 140798 44718 140826
rect 44980 140798 45454 140826
rect 45808 140798 46098 140826
rect 46544 140798 46834 140826
rect 47188 140798 47478 140826
rect 33940 140662 34506 140690
rect 51406 140432 51462 140441
rect 51406 140367 51462 140376
rect 49934 140160 49990 140169
rect 49934 140095 49990 140104
rect 49948 139994 49976 140095
rect 49936 139988 49988 139994
rect 49936 139930 49988 139936
rect 50026 139072 50082 139081
rect 50026 139007 50082 139016
rect 49936 138696 49988 138702
rect 49934 138664 49936 138673
rect 49988 138664 49990 138673
rect 50040 138634 50068 139007
rect 49934 138599 49990 138608
rect 50028 138628 50080 138634
rect 50028 138570 50080 138576
rect 51420 138566 51448 140367
rect 56192 139988 56244 139994
rect 56192 139930 56244 139936
rect 51408 138560 51460 138566
rect 51408 138502 51460 138508
rect 56204 138498 56232 139930
rect 68716 138786 68744 142650
rect 68408 138758 68744 138786
rect 58492 138696 58544 138702
rect 58492 138638 58544 138644
rect 58400 138628 58452 138634
rect 58400 138570 58452 138576
rect 56192 138492 56244 138498
rect 56192 138434 56244 138440
rect 50026 137848 50082 137857
rect 50026 137783 50082 137792
rect 49934 137440 49990 137449
rect 49934 137375 49990 137384
rect 49948 137274 49976 137375
rect 49936 137268 49988 137274
rect 49936 137210 49988 137216
rect 50040 137206 50068 137783
rect 58308 137268 58360 137274
rect 58308 137210 58360 137216
rect 50028 137200 50080 137206
rect 50028 137142 50080 137148
rect 58216 137132 58268 137138
rect 58216 137074 58268 137080
rect 50394 136624 50450 136633
rect 50394 136559 50450 136568
rect 18102 135944 18158 135953
rect 18102 135879 18158 135888
rect 18010 126288 18066 126297
rect 18010 126223 18066 126232
rect 18024 117706 18052 126223
rect 17840 117678 18052 117706
rect 17840 113338 17868 117678
rect 18010 117040 18066 117049
rect 18010 116975 18066 116984
rect 17828 113332 17880 113338
rect 17828 113274 17880 113280
rect 18024 112998 18052 116975
rect 18012 112992 18064 112998
rect 18012 112934 18064 112940
rect 18116 63630 18144 135879
rect 50408 135846 50436 136559
rect 51222 136216 51278 136225
rect 51222 136151 51224 136160
rect 51276 136151 51278 136160
rect 52788 136180 52840 136186
rect 51224 136122 51276 136128
rect 52788 136122 52840 136128
rect 51222 136080 51278 136089
rect 51222 136015 51224 136024
rect 51276 136015 51278 136024
rect 52696 136044 52748 136050
rect 51224 135986 51276 135992
rect 52696 135986 52748 135992
rect 50396 135840 50448 135846
rect 50396 135782 50448 135788
rect 51222 134992 51278 135001
rect 51222 134927 51278 134936
rect 51236 134622 51264 134927
rect 51224 134616 51276 134622
rect 51130 134584 51186 134593
rect 51224 134558 51276 134564
rect 51130 134519 51132 134528
rect 51184 134519 51186 134528
rect 51132 134490 51184 134496
rect 52708 134350 52736 135986
rect 52800 134418 52828 136122
rect 58228 136089 58256 137074
rect 58214 136080 58270 136089
rect 58214 136015 58270 136024
rect 58216 135772 58268 135778
rect 58216 135714 58268 135720
rect 58228 134865 58256 135714
rect 58320 135409 58348 137210
rect 58412 137177 58440 138570
rect 58398 137168 58454 137177
rect 58398 137103 58454 137112
rect 58504 136633 58532 138638
rect 59228 138560 59280 138566
rect 59226 138528 59228 138537
rect 92716 138560 92768 138566
rect 59280 138528 59282 138537
rect 58676 138492 58728 138498
rect 59226 138463 59282 138472
rect 92714 138528 92716 138537
rect 92768 138528 92770 138537
rect 92714 138463 92770 138472
rect 92808 138492 92860 138498
rect 58676 138434 58728 138440
rect 92808 138434 92860 138440
rect 58688 138265 58716 138434
rect 58674 138256 58730 138265
rect 58674 138191 58730 138200
rect 92820 138129 92848 138434
rect 92806 138120 92862 138129
rect 92806 138055 92862 138064
rect 92714 137168 92770 137177
rect 92714 137103 92716 137112
rect 92768 137103 92770 137112
rect 92716 137074 92768 137080
rect 92808 137064 92860 137070
rect 92808 137006 92860 137012
rect 92716 136996 92768 137002
rect 92716 136938 92768 136944
rect 58490 136624 58546 136633
rect 58490 136559 58546 136568
rect 92728 136497 92756 136938
rect 92820 136905 92848 137006
rect 92806 136896 92862 136905
rect 92806 136831 92862 136840
rect 92714 136488 92770 136497
rect 92714 136423 92770 136432
rect 92808 135772 92860 135778
rect 92808 135714 92860 135720
rect 92716 135704 92768 135710
rect 92716 135646 92768 135652
rect 92728 135545 92756 135646
rect 92714 135536 92770 135545
rect 92714 135471 92770 135480
rect 58306 135400 58362 135409
rect 58306 135335 58362 135344
rect 92820 135273 92848 135714
rect 92806 135264 92862 135273
rect 92806 135199 92862 135208
rect 58214 134856 58270 134865
rect 58214 134791 58270 134800
rect 56744 134616 56796 134622
rect 56744 134558 56796 134564
rect 52880 134548 52932 134554
rect 52880 134490 52932 134496
rect 52788 134412 52840 134418
rect 52788 134354 52840 134360
rect 52696 134344 52748 134350
rect 52696 134286 52748 134292
rect 50210 133768 50266 133777
rect 50210 133703 50266 133712
rect 50224 133058 50252 133703
rect 50946 133224 51002 133233
rect 50946 133159 51002 133168
rect 50960 133126 50988 133159
rect 50948 133120 51000 133126
rect 50948 133062 51000 133068
rect 52696 133120 52748 133126
rect 52696 133062 52748 133068
rect 50212 133052 50264 133058
rect 50212 132994 50264 133000
rect 51222 132544 51278 132553
rect 51222 132479 51278 132488
rect 50394 132136 50450 132145
rect 50394 132071 50450 132080
rect 50408 132038 50436 132071
rect 50396 132032 50448 132038
rect 50396 131974 50448 131980
rect 51236 131970 51264 132479
rect 51224 131964 51276 131970
rect 51224 131906 51276 131912
rect 51222 131728 51278 131737
rect 51222 131663 51224 131672
rect 51276 131663 51278 131672
rect 51224 131634 51276 131640
rect 52708 131630 52736 133062
rect 52892 132990 52920 134490
rect 56756 133874 56784 134558
rect 59412 134548 59464 134554
rect 59412 134490 59464 134496
rect 58216 134412 58268 134418
rect 58216 134354 58268 134360
rect 58228 134185 58256 134354
rect 58308 134344 58360 134350
rect 58308 134286 58360 134292
rect 58214 134176 58270 134185
rect 58214 134111 58270 134120
rect 56744 133868 56796 133874
rect 56744 133810 56796 133816
rect 58216 133868 58268 133874
rect 58216 133810 58268 133816
rect 58228 133097 58256 133810
rect 58320 133641 58348 134286
rect 58306 133632 58362 133641
rect 58306 133567 58362 133576
rect 58214 133088 58270 133097
rect 56100 133052 56152 133058
rect 58214 133023 58270 133032
rect 56100 132994 56152 133000
rect 52880 132984 52932 132990
rect 52880 132926 52932 132932
rect 56112 132446 56140 132994
rect 59424 132990 59452 134490
rect 92900 134412 92952 134418
rect 92900 134354 92952 134360
rect 92716 134344 92768 134350
rect 92714 134312 92716 134321
rect 92768 134312 92770 134321
rect 92714 134247 92770 134256
rect 92808 134276 92860 134282
rect 92808 134218 92860 134224
rect 92820 133913 92848 134218
rect 92806 133904 92862 133913
rect 92806 133839 92862 133848
rect 92912 133505 92940 134354
rect 92898 133496 92954 133505
rect 92898 133431 92954 133440
rect 58216 132984 58268 132990
rect 58216 132926 58268 132932
rect 59412 132984 59464 132990
rect 59412 132926 59464 132932
rect 92808 132984 92860 132990
rect 92808 132926 92860 132932
rect 56100 132440 56152 132446
rect 58228 132417 58256 132926
rect 92716 132916 92768 132922
rect 92716 132858 92768 132864
rect 92728 132689 92756 132858
rect 92714 132680 92770 132689
rect 92714 132615 92770 132624
rect 58308 132440 58360 132446
rect 56100 132382 56152 132388
rect 58214 132408 58270 132417
rect 58308 132382 58360 132388
rect 58214 132343 58270 132352
rect 53432 132032 53484 132038
rect 53432 131974 53484 131980
rect 52788 131692 52840 131698
rect 52788 131634 52840 131640
rect 52696 131624 52748 131630
rect 52696 131566 52748 131572
rect 51222 130776 51278 130785
rect 51222 130711 51224 130720
rect 51276 130711 51278 130720
rect 51224 130682 51276 130688
rect 51222 130368 51278 130377
rect 51222 130303 51224 130312
rect 51276 130303 51278 130312
rect 52696 130332 52748 130338
rect 51224 130274 51276 130280
rect 52696 130274 52748 130280
rect 50394 129688 50450 129697
rect 50394 129623 50450 129632
rect 50408 129114 50436 129623
rect 50396 129108 50448 129114
rect 50396 129050 50448 129056
rect 51222 129008 51278 129017
rect 51222 128943 51224 128952
rect 51276 128943 51278 128952
rect 51224 128914 51276 128920
rect 52708 128910 52736 130274
rect 52800 130202 52828 131634
rect 52972 130740 53024 130746
rect 52972 130682 53024 130688
rect 52788 130196 52840 130202
rect 52788 130138 52840 130144
rect 52880 128972 52932 128978
rect 52880 128914 52932 128920
rect 52696 128904 52748 128910
rect 52696 128846 52748 128852
rect 50946 128464 51002 128473
rect 50946 128399 51002 128408
rect 50960 127890 50988 128399
rect 51222 127920 51278 127929
rect 50948 127884 51000 127890
rect 51222 127855 51278 127864
rect 50948 127826 51000 127832
rect 51236 127822 51264 127855
rect 51224 127816 51276 127822
rect 51224 127758 51276 127764
rect 52788 127816 52840 127822
rect 52788 127758 52840 127764
rect 51222 127648 51278 127657
rect 51222 127583 51224 127592
rect 51276 127583 51278 127592
rect 52696 127612 52748 127618
rect 51224 127554 51276 127560
rect 52696 127554 52748 127560
rect 51222 126696 51278 126705
rect 51278 126654 51448 126682
rect 51222 126631 51278 126640
rect 51222 126152 51278 126161
rect 51278 126110 51356 126138
rect 51222 126087 51278 126096
rect 50210 125608 50266 125617
rect 50210 125543 50266 125552
rect 50224 124830 50252 125543
rect 51222 125064 51278 125073
rect 51222 124999 51224 125008
rect 51276 124999 51278 125008
rect 51224 124970 51276 124976
rect 51222 124928 51278 124937
rect 51222 124863 51224 124872
rect 51276 124863 51278 124872
rect 51224 124834 51276 124840
rect 50212 124824 50264 124830
rect 50212 124766 50264 124772
rect 51328 124762 51356 126110
rect 51316 124756 51368 124762
rect 51316 124698 51368 124704
rect 51420 124694 51448 126654
rect 52708 126122 52736 127554
rect 52696 126116 52748 126122
rect 52696 126058 52748 126064
rect 52800 126054 52828 127758
rect 52892 127482 52920 128914
rect 52984 128842 53012 130682
rect 53444 130270 53472 131974
rect 55456 131964 55508 131970
rect 55456 131906 55508 131912
rect 55468 131358 55496 131906
rect 58320 131873 58348 132382
rect 92820 132281 92848 132926
rect 92806 132272 92862 132281
rect 92806 132207 92862 132216
rect 58306 131864 58362 131873
rect 58306 131799 58362 131808
rect 58216 131624 58268 131630
rect 58216 131566 58268 131572
rect 92716 131624 92768 131630
rect 92716 131566 92768 131572
rect 55456 131352 55508 131358
rect 55456 131294 55508 131300
rect 58228 131193 58256 131566
rect 92728 131465 92756 131566
rect 92808 131556 92860 131562
rect 92808 131498 92860 131504
rect 92714 131456 92770 131465
rect 92714 131391 92770 131400
rect 58308 131352 58360 131358
rect 58308 131294 58360 131300
rect 58214 131184 58270 131193
rect 58214 131119 58270 131128
rect 58320 130649 58348 131294
rect 92820 131057 92848 131498
rect 92806 131048 92862 131057
rect 92806 130983 92862 130992
rect 58306 130640 58362 130649
rect 58306 130575 58362 130584
rect 53432 130264 53484 130270
rect 53432 130206 53484 130212
rect 58216 130264 58268 130270
rect 92716 130264 92768 130270
rect 58216 130206 58268 130212
rect 92714 130232 92716 130241
rect 92768 130232 92770 130241
rect 58228 130105 58256 130206
rect 58308 130196 58360 130202
rect 92714 130167 92770 130176
rect 92808 130196 92860 130202
rect 58308 130138 58360 130144
rect 92808 130138 92860 130144
rect 58214 130096 58270 130105
rect 58214 130031 58270 130040
rect 58320 129425 58348 130138
rect 92820 129833 92848 130138
rect 92806 129824 92862 129833
rect 92806 129759 92862 129768
rect 58306 129416 58362 129425
rect 58306 129351 58362 129360
rect 56468 129108 56520 129114
rect 56468 129050 56520 129056
rect 52972 128836 53024 128842
rect 52972 128778 53024 128784
rect 56480 128366 56508 129050
rect 58308 128904 58360 128910
rect 58214 128872 58270 128881
rect 92716 128904 92768 128910
rect 58308 128846 58360 128852
rect 92714 128872 92716 128881
rect 92768 128872 92770 128881
rect 58214 128807 58216 128816
rect 58268 128807 58270 128816
rect 58216 128778 58268 128784
rect 56468 128360 56520 128366
rect 56468 128302 56520 128308
rect 58216 128360 58268 128366
rect 58216 128302 58268 128308
rect 56744 127884 56796 127890
rect 56744 127826 56796 127832
rect 52880 127476 52932 127482
rect 52880 127418 52932 127424
rect 56756 127210 56784 127826
rect 58228 127657 58256 128302
rect 58320 128201 58348 128846
rect 92714 128807 92770 128816
rect 92808 128836 92860 128842
rect 92808 128778 92860 128784
rect 92716 128768 92768 128774
rect 92716 128710 92768 128716
rect 58306 128192 58362 128201
rect 58306 128127 58362 128136
rect 92728 128065 92756 128710
rect 92820 128473 92848 128778
rect 92806 128464 92862 128473
rect 92806 128399 92862 128408
rect 92714 128056 92770 128065
rect 92714 127991 92770 128000
rect 58214 127648 58270 127657
rect 58214 127583 58270 127592
rect 58216 127476 58268 127482
rect 58216 127418 58268 127424
rect 92808 127476 92860 127482
rect 92808 127418 92860 127424
rect 56744 127204 56796 127210
rect 56744 127146 56796 127152
rect 58228 127113 58256 127418
rect 92716 127408 92768 127414
rect 92716 127350 92768 127356
rect 92728 127249 92756 127350
rect 92714 127240 92770 127249
rect 58308 127204 58360 127210
rect 92714 127175 92770 127184
rect 58308 127146 58360 127152
rect 58214 127104 58270 127113
rect 58214 127039 58270 127048
rect 58320 126433 58348 127146
rect 92820 126977 92848 127418
rect 92806 126968 92862 126977
rect 92806 126903 92862 126912
rect 58306 126424 58362 126433
rect 58306 126359 58362 126368
rect 58308 126116 58360 126122
rect 58308 126058 58360 126064
rect 92808 126116 92860 126122
rect 92808 126058 92860 126064
rect 52788 126048 52840 126054
rect 52788 125990 52840 125996
rect 58216 126048 58268 126054
rect 58216 125990 58268 125996
rect 58228 125889 58256 125990
rect 58214 125880 58270 125889
rect 58214 125815 58270 125824
rect 58320 125209 58348 126058
rect 92716 126048 92768 126054
rect 92714 126016 92716 126025
rect 92768 126016 92770 126025
rect 92714 125951 92770 125960
rect 92820 125617 92848 126058
rect 92806 125608 92862 125617
rect 92806 125543 92862 125552
rect 58306 125200 58362 125209
rect 58306 125135 58362 125144
rect 52972 125028 53024 125034
rect 52972 124970 53024 124976
rect 52880 124892 52932 124898
rect 52880 124834 52932 124840
rect 51408 124688 51460 124694
rect 51408 124630 51460 124636
rect 50578 123840 50634 123849
rect 50578 123775 50634 123784
rect 50592 123470 50620 123775
rect 50580 123464 50632 123470
rect 52696 123464 52748 123470
rect 50580 123406 50632 123412
rect 51130 123432 51186 123441
rect 52696 123406 52748 123412
rect 51130 123367 51132 123376
rect 51184 123367 51186 123376
rect 51132 123338 51184 123344
rect 50854 122616 50910 122625
rect 50854 122551 50910 122560
rect 50868 122382 50896 122551
rect 50856 122376 50908 122382
rect 50210 122344 50266 122353
rect 50856 122318 50908 122324
rect 50210 122279 50266 122288
rect 50224 122246 50252 122279
rect 50212 122240 50264 122246
rect 50212 122182 50264 122188
rect 52708 121906 52736 123406
rect 52788 123396 52840 123402
rect 52788 123338 52840 123344
rect 52800 121974 52828 123338
rect 52892 123266 52920 124834
rect 52984 123334 53012 124970
rect 58400 124824 58452 124830
rect 58400 124766 58452 124772
rect 58308 124756 58360 124762
rect 58308 124698 58360 124704
rect 58216 124688 58268 124694
rect 58214 124656 58216 124665
rect 58268 124656 58270 124665
rect 58214 124591 58270 124600
rect 58320 124121 58348 124698
rect 58306 124112 58362 124121
rect 58306 124047 58362 124056
rect 58412 123441 58440 124766
rect 92900 124756 92952 124762
rect 92900 124698 92952 124704
rect 92716 124688 92768 124694
rect 92714 124656 92716 124665
rect 92768 124656 92770 124665
rect 92714 124591 92770 124600
rect 92808 124620 92860 124626
rect 92808 124562 92860 124568
rect 92820 124393 92848 124562
rect 92806 124384 92862 124393
rect 92806 124319 92862 124328
rect 92912 123985 92940 124698
rect 92898 123976 92954 123985
rect 92898 123911 92954 123920
rect 58398 123432 58454 123441
rect 58398 123367 58454 123376
rect 52972 123328 53024 123334
rect 52972 123270 53024 123276
rect 58216 123328 58268 123334
rect 58216 123270 58268 123276
rect 92716 123328 92768 123334
rect 92716 123270 92768 123276
rect 52880 123260 52932 123266
rect 52880 123202 52932 123208
rect 58228 122897 58256 123270
rect 58308 123260 58360 123266
rect 58308 123202 58360 123208
rect 58214 122888 58270 122897
rect 58214 122823 58270 122832
rect 52972 122376 53024 122382
rect 52972 122318 53024 122324
rect 52880 122240 52932 122246
rect 52880 122182 52932 122188
rect 52788 121968 52840 121974
rect 52788 121910 52840 121916
rect 52696 121900 52748 121906
rect 52696 121842 52748 121848
rect 50210 121528 50266 121537
rect 50210 121463 50266 121472
rect 50224 120682 50252 121463
rect 51222 120984 51278 120993
rect 51222 120919 51224 120928
rect 51276 120919 51278 120928
rect 51224 120890 51276 120896
rect 51222 120848 51278 120857
rect 51222 120783 51278 120792
rect 51236 120750 51264 120783
rect 51224 120744 51276 120750
rect 51224 120686 51276 120692
rect 52696 120744 52748 120750
rect 52696 120686 52748 120692
rect 50212 120676 50264 120682
rect 50212 120618 50264 120624
rect 51222 119760 51278 119769
rect 51222 119695 51278 119704
rect 51236 119594 51264 119695
rect 51224 119588 51276 119594
rect 51224 119530 51276 119536
rect 51222 119352 51278 119361
rect 51222 119287 51224 119296
rect 51276 119287 51278 119296
rect 51224 119258 51276 119264
rect 52708 119254 52736 120686
rect 52892 120546 52920 122182
rect 52984 120614 53012 122318
rect 58320 122217 58348 123202
rect 92728 123169 92756 123270
rect 92808 123260 92860 123266
rect 92808 123202 92860 123208
rect 92714 123160 92770 123169
rect 92714 123095 92770 123104
rect 92820 122761 92848 123202
rect 92806 122752 92862 122761
rect 92806 122687 92862 122696
rect 58306 122208 58362 122217
rect 58306 122143 58362 122152
rect 58308 121968 58360 121974
rect 58308 121910 58360 121916
rect 92808 121968 92860 121974
rect 92808 121910 92860 121916
rect 58216 121900 58268 121906
rect 58216 121842 58268 121848
rect 58228 121673 58256 121842
rect 58214 121664 58270 121673
rect 58214 121599 58270 121608
rect 58320 121129 58348 121910
rect 92716 121900 92768 121906
rect 92716 121842 92768 121848
rect 92728 121809 92756 121842
rect 92714 121800 92770 121809
rect 92714 121735 92770 121744
rect 92820 121537 92848 121910
rect 92806 121528 92862 121537
rect 92806 121463 92862 121472
rect 58306 121120 58362 121129
rect 58306 121055 58362 121064
rect 53064 120948 53116 120954
rect 53064 120890 53116 120896
rect 52972 120608 53024 120614
rect 52972 120550 53024 120556
rect 52880 120540 52932 120546
rect 52880 120482 52932 120488
rect 52880 119588 52932 119594
rect 52880 119530 52932 119536
rect 52788 119316 52840 119322
rect 52788 119258 52840 119264
rect 52696 119248 52748 119254
rect 52696 119190 52748 119196
rect 51222 118536 51278 118545
rect 51222 118471 51278 118480
rect 51236 118234 51264 118471
rect 51224 118228 51276 118234
rect 51224 118170 51276 118176
rect 51222 117992 51278 118001
rect 51222 117927 51224 117936
rect 51276 117927 51278 117936
rect 52696 117956 52748 117962
rect 51224 117898 51276 117904
rect 52696 117898 52748 117904
rect 51222 117448 51278 117457
rect 51222 117383 51278 117392
rect 50578 116768 50634 116777
rect 51236 116738 51264 117383
rect 50578 116703 50634 116712
rect 51224 116732 51276 116738
rect 29722 113054 30288 113082
rect 20232 110278 20260 112932
rect 20220 110272 20272 110278
rect 20220 110214 20272 110220
rect 20876 109598 20904 112932
rect 21520 109734 21548 112932
rect 21508 109728 21560 109734
rect 21508 109670 21560 109676
rect 22256 109666 22284 112932
rect 22900 109870 22928 112932
rect 22888 109864 22940 109870
rect 22888 109806 22940 109812
rect 23636 109802 23664 112932
rect 23624 109796 23676 109802
rect 23624 109738 23676 109744
rect 22244 109660 22296 109666
rect 22244 109602 22296 109608
rect 24280 109598 24308 112932
rect 24924 109938 24952 112932
rect 25674 112918 25964 112946
rect 26318 112918 26424 112946
rect 25936 110006 25964 112918
rect 25924 110000 25976 110006
rect 25924 109942 25976 109948
rect 26292 110000 26344 110006
rect 26292 109942 26344 109948
rect 24912 109932 24964 109938
rect 24912 109874 24964 109880
rect 20864 109592 20916 109598
rect 20864 109534 20916 109540
rect 22980 109592 23032 109598
rect 22980 109534 23032 109540
rect 24268 109592 24320 109598
rect 24268 109534 24320 109540
rect 22992 102458 23020 109534
rect 22980 102452 23032 102458
rect 22980 102394 23032 102400
rect 26108 102452 26160 102458
rect 26108 102394 26160 102400
rect 26120 99740 26148 102394
rect 26304 102050 26332 109942
rect 26292 102044 26344 102050
rect 26292 101986 26344 101992
rect 26396 101778 26424 112918
rect 26476 109728 26528 109734
rect 26476 109670 26528 109676
rect 26384 101772 26436 101778
rect 26384 101714 26436 101720
rect 26488 99740 26516 109670
rect 27040 109666 27068 112932
rect 27684 109938 27712 112932
rect 27672 109932 27724 109938
rect 27672 109874 27724 109880
rect 27304 109864 27356 109870
rect 27304 109806 27356 109812
rect 26844 109660 26896 109666
rect 26844 109602 26896 109608
rect 27028 109660 27080 109666
rect 27028 109602 27080 109608
rect 26856 99740 26884 109602
rect 27316 99740 27344 109806
rect 27672 109796 27724 109802
rect 27672 109738 27724 109744
rect 27684 99740 27712 109738
rect 28328 109598 28356 112932
rect 29064 110006 29092 112932
rect 29052 110000 29104 110006
rect 29052 109942 29104 109948
rect 30064 109932 30116 109938
rect 30064 109874 30116 109880
rect 28500 109864 28552 109870
rect 28500 109806 28552 109812
rect 28132 109592 28184 109598
rect 28132 109534 28184 109540
rect 28316 109592 28368 109598
rect 28316 109534 28368 109540
rect 28144 99754 28172 109534
rect 28066 99726 28172 99754
rect 28512 99740 28540 109806
rect 29696 109660 29748 109666
rect 29696 109602 29748 109608
rect 29144 109592 29196 109598
rect 29144 109534 29196 109540
rect 29156 102050 29184 109534
rect 28868 102044 28920 102050
rect 28868 101986 28920 101992
rect 29144 102044 29196 102050
rect 29144 101986 29196 101992
rect 28880 99740 28908 101986
rect 29236 101772 29288 101778
rect 29236 101714 29288 101720
rect 29248 99740 29276 101714
rect 29708 99740 29736 109602
rect 30076 99740 30104 109874
rect 30260 102662 30288 113054
rect 35320 113054 35886 113082
rect 30458 112918 30564 112946
rect 30248 102656 30300 102662
rect 30248 102598 30300 102604
rect 30432 102044 30484 102050
rect 30432 101986 30484 101992
rect 30444 99740 30472 101986
rect 30536 101846 30564 112918
rect 31088 110482 31116 112932
rect 31076 110476 31128 110482
rect 31076 110418 31128 110424
rect 30892 110000 30944 110006
rect 30892 109942 30944 109948
rect 30524 101840 30576 101846
rect 30524 101782 30576 101788
rect 30904 99740 30932 109942
rect 31260 102656 31312 102662
rect 31260 102598 31312 102604
rect 31272 99740 31300 102598
rect 31628 101840 31680 101846
rect 31628 101782 31680 101788
rect 31640 99740 31668 101782
rect 31824 101438 31852 112932
rect 32100 112918 32482 112946
rect 32744 112918 33126 112946
rect 33480 112918 33862 112946
rect 34216 112918 34506 112946
rect 34768 112918 35242 112946
rect 31904 110476 31956 110482
rect 31904 110418 31956 110424
rect 31812 101432 31864 101438
rect 31812 101374 31864 101380
rect 31916 101386 31944 110418
rect 32100 102662 32128 112918
rect 32088 102656 32140 102662
rect 32088 102598 32140 102604
rect 32744 102594 32772 112918
rect 32824 102656 32876 102662
rect 32824 102598 32876 102604
rect 32732 102588 32784 102594
rect 32732 102530 32784 102536
rect 32456 101432 32508 101438
rect 31916 101358 32036 101386
rect 32456 101374 32508 101380
rect 32008 99754 32036 101358
rect 32008 99726 32114 99754
rect 32468 99740 32496 101374
rect 32836 99740 32864 102598
rect 33284 102588 33336 102594
rect 33284 102530 33336 102536
rect 33296 99740 33324 102530
rect 33480 99754 33508 112918
rect 34216 99754 34244 112918
rect 34768 101352 34796 112918
rect 35320 112674 35348 113054
rect 34676 101324 34796 101352
rect 34860 112646 35348 112674
rect 36148 112918 36530 112946
rect 36792 112918 37266 112946
rect 37620 112918 37910 112946
rect 38264 112918 38646 112946
rect 34676 99754 34704 101324
rect 33480 99726 33678 99754
rect 34138 99726 34244 99754
rect 34506 99726 34704 99754
rect 34860 99740 34888 112646
rect 36148 102662 36176 112918
rect 35308 102656 35360 102662
rect 35308 102598 35360 102604
rect 36136 102656 36188 102662
rect 36136 102598 36188 102604
rect 35320 99740 35348 102598
rect 36792 102594 36820 112918
rect 37516 109728 37568 109734
rect 37516 109670 37568 109676
rect 36872 102656 36924 102662
rect 36872 102598 36924 102604
rect 35676 102588 35728 102594
rect 35676 102530 35728 102536
rect 36780 102588 36832 102594
rect 36780 102530 36832 102536
rect 35688 99740 35716 102530
rect 36044 102520 36096 102526
rect 36044 102462 36096 102468
rect 36056 99740 36084 102462
rect 36504 102044 36556 102050
rect 36504 101986 36556 101992
rect 36516 99740 36544 101986
rect 36884 99740 36912 102598
rect 37528 102050 37556 109670
rect 37620 102526 37648 112918
rect 38264 109734 38292 112918
rect 38252 109728 38304 109734
rect 38252 109670 38304 109676
rect 38160 109660 38212 109666
rect 38160 109602 38212 109608
rect 37700 102588 37752 102594
rect 37700 102530 37752 102536
rect 37608 102520 37660 102526
rect 37608 102462 37660 102468
rect 37516 102044 37568 102050
rect 37516 101986 37568 101992
rect 37240 101840 37292 101846
rect 37240 101782 37292 101788
rect 37252 99740 37280 101782
rect 37712 99740 37740 102530
rect 38068 102520 38120 102526
rect 38068 102462 38120 102468
rect 38080 99740 38108 102462
rect 38172 101846 38200 109602
rect 39276 109598 39304 112932
rect 40012 109666 40040 112932
rect 40288 112918 40670 112946
rect 40840 112918 41314 112946
rect 41852 112918 42050 112946
rect 42312 112918 42694 112946
rect 43140 112918 43430 112946
rect 43784 112918 44074 112946
rect 44520 112918 44718 112946
rect 45072 112918 45454 112946
rect 40000 109660 40052 109666
rect 40000 109602 40052 109608
rect 38252 109592 38304 109598
rect 38252 109534 38304 109540
rect 39264 109592 39316 109598
rect 39264 109534 39316 109540
rect 38264 102662 38292 109534
rect 38252 102656 38304 102662
rect 38252 102598 38304 102604
rect 40288 102594 40316 112918
rect 40276 102588 40328 102594
rect 40276 102530 40328 102536
rect 40840 102526 40868 112918
rect 41748 110272 41800 110278
rect 41748 110214 41800 110220
rect 41656 107552 41708 107558
rect 41656 107494 41708 107500
rect 40828 102520 40880 102526
rect 40828 102462 40880 102468
rect 40092 101908 40144 101914
rect 40092 101850 40144 101856
rect 38160 101840 38212 101846
rect 38160 101782 38212 101788
rect 39264 101840 39316 101846
rect 39264 101782 39316 101788
rect 38436 101772 38488 101778
rect 38436 101714 38488 101720
rect 38448 99740 38476 101714
rect 38896 101500 38948 101506
rect 38896 101442 38948 101448
rect 38908 99740 38936 101442
rect 39276 99740 39304 101782
rect 39632 101636 39684 101642
rect 39632 101578 39684 101584
rect 39644 99740 39672 101578
rect 40104 99740 40132 101850
rect 40828 101704 40880 101710
rect 40828 101646 40880 101652
rect 40460 101568 40512 101574
rect 40460 101510 40512 101516
rect 40472 99740 40500 101510
rect 40840 99740 40868 101646
rect 41668 101506 41696 107494
rect 41656 101500 41708 101506
rect 41656 101442 41708 101448
rect 41288 101432 41340 101438
rect 41288 101374 41340 101380
rect 41300 99740 41328 101374
rect 41656 101364 41708 101370
rect 41656 101306 41708 101312
rect 41668 99740 41696 101306
rect 22336 97148 22388 97154
rect 22336 97090 22388 97096
rect 22348 96513 22376 97090
rect 22334 96504 22390 96513
rect 22334 96439 22390 96448
rect 41760 95266 41788 110214
rect 41852 101778 41880 112918
rect 42312 107558 42340 112918
rect 42944 109728 42996 109734
rect 42944 109670 42996 109676
rect 42300 107552 42352 107558
rect 42300 107494 42352 107500
rect 41840 101772 41892 101778
rect 41840 101714 41892 101720
rect 42956 101370 42984 109670
rect 43036 107552 43088 107558
rect 43036 107494 43088 107500
rect 43048 101642 43076 107494
rect 43140 101846 43168 112918
rect 43784 107558 43812 112918
rect 44416 109796 44468 109802
rect 44416 109738 44468 109744
rect 43772 107552 43824 107558
rect 43772 107494 43824 107500
rect 43128 101840 43180 101846
rect 43128 101782 43180 101788
rect 43036 101636 43088 101642
rect 43036 101578 43088 101584
rect 44428 101574 44456 109738
rect 44520 101914 44548 112918
rect 45072 109802 45100 112918
rect 45060 109796 45112 109802
rect 45060 109738 45112 109744
rect 45060 109660 45112 109666
rect 45060 109602 45112 109608
rect 44508 101908 44560 101914
rect 44508 101850 44560 101856
rect 44416 101568 44468 101574
rect 44416 101510 44468 101516
rect 45072 101438 45100 109602
rect 46084 109598 46112 112932
rect 46820 109666 46848 112932
rect 47464 109734 47492 112932
rect 47452 109728 47504 109734
rect 47452 109670 47504 109676
rect 46808 109660 46860 109666
rect 46808 109602 46860 109608
rect 45152 109592 45204 109598
rect 45152 109534 45204 109540
rect 46072 109592 46124 109598
rect 46072 109534 46124 109540
rect 45164 101710 45192 109534
rect 50592 102050 50620 116703
rect 51224 116674 51276 116680
rect 50762 116496 50818 116505
rect 50762 116431 50818 116440
rect 50670 115136 50726 115145
rect 50670 115071 50726 115080
rect 50684 102254 50712 115071
rect 50672 102248 50724 102254
rect 50672 102190 50724 102196
rect 50776 102118 50804 116431
rect 52708 116398 52736 117898
rect 52800 117758 52828 119258
rect 52892 117826 52920 119530
rect 53076 119118 53104 120890
rect 53156 120676 53208 120682
rect 53156 120618 53208 120624
rect 53168 119186 53196 120618
rect 58216 120608 58268 120614
rect 92716 120608 92768 120614
rect 58216 120550 58268 120556
rect 92714 120576 92716 120585
rect 92768 120576 92770 120585
rect 58228 120449 58256 120550
rect 58308 120540 58360 120546
rect 92714 120511 92770 120520
rect 92808 120540 92860 120546
rect 58308 120482 58360 120488
rect 92808 120482 92860 120488
rect 58214 120440 58270 120449
rect 58214 120375 58270 120384
rect 58320 119905 58348 120482
rect 92820 120177 92848 120482
rect 92806 120168 92862 120177
rect 92806 120103 92862 120112
rect 58306 119896 58362 119905
rect 58306 119831 58362 119840
rect 58400 119248 58452 119254
rect 58214 119216 58270 119225
rect 53156 119180 53208 119186
rect 92900 119248 92952 119254
rect 58400 119190 58452 119196
rect 92714 119216 92770 119225
rect 58214 119151 58216 119160
rect 53156 119122 53208 119128
rect 58268 119151 58270 119160
rect 58216 119122 58268 119128
rect 53064 119112 53116 119118
rect 53064 119054 53116 119060
rect 58308 119112 58360 119118
rect 58308 119054 58360 119060
rect 58320 118681 58348 119054
rect 58306 118672 58362 118681
rect 58306 118607 58362 118616
rect 52972 118228 53024 118234
rect 52972 118170 53024 118176
rect 52880 117820 52932 117826
rect 52880 117762 52932 117768
rect 52788 117752 52840 117758
rect 52788 117694 52840 117700
rect 52984 116466 53012 118170
rect 58412 118137 58440 119190
rect 92900 119190 92952 119196
rect 92714 119151 92770 119160
rect 92808 119180 92860 119186
rect 92728 119118 92756 119151
rect 92808 119122 92860 119128
rect 92716 119112 92768 119118
rect 92716 119054 92768 119060
rect 92820 118953 92848 119122
rect 92806 118944 92862 118953
rect 92806 118879 92862 118888
rect 92912 118545 92940 119190
rect 92898 118536 92954 118545
rect 92898 118471 92954 118480
rect 58398 118128 58454 118137
rect 58398 118063 58454 118072
rect 58216 117820 58268 117826
rect 58216 117762 58268 117768
rect 92716 117820 92768 117826
rect 92716 117762 92768 117768
rect 58228 117457 58256 117762
rect 58308 117752 58360 117758
rect 58308 117694 58360 117700
rect 58214 117448 58270 117457
rect 58214 117383 58270 117392
rect 58320 116913 58348 117694
rect 92728 117593 92756 117762
rect 92808 117752 92860 117758
rect 92808 117694 92860 117700
rect 92714 117584 92770 117593
rect 92714 117519 92770 117528
rect 92820 117321 92848 117694
rect 92806 117312 92862 117321
rect 92806 117247 92862 117256
rect 58306 116904 58362 116913
rect 58306 116839 58362 116848
rect 56468 116732 56520 116738
rect 56468 116674 56520 116680
rect 52972 116460 53024 116466
rect 52972 116402 53024 116408
rect 52696 116392 52748 116398
rect 52696 116334 52748 116340
rect 56480 116330 56508 116674
rect 94004 116596 94056 116602
rect 94004 116538 94056 116544
rect 92624 116528 92676 116534
rect 92624 116470 92676 116476
rect 58216 116460 58268 116466
rect 58216 116402 58268 116408
rect 56468 116324 56520 116330
rect 56468 116266 56520 116272
rect 58228 116233 58256 116402
rect 58308 116392 58360 116398
rect 58308 116334 58360 116340
rect 58214 116224 58270 116233
rect 58214 116159 58270 116168
rect 58320 115689 58348 116334
rect 58400 116324 58452 116330
rect 58400 116266 58452 116272
rect 50854 115680 50910 115689
rect 50854 115615 50910 115624
rect 58306 115680 58362 115689
rect 58306 115615 58362 115624
rect 50868 102186 50896 115615
rect 58412 115145 58440 116266
rect 91244 115236 91296 115242
rect 91244 115178 91296 115184
rect 59320 115168 59372 115174
rect 58398 115136 58454 115145
rect 59320 115110 59372 115116
rect 90600 115168 90652 115174
rect 90600 115110 90652 115116
rect 58398 115071 58454 115080
rect 50946 114456 51002 114465
rect 50946 114391 51002 114400
rect 50960 102390 50988 114391
rect 51130 114048 51186 114057
rect 51130 113983 51186 113992
rect 51038 112824 51094 112833
rect 51038 112759 51094 112768
rect 50948 102384 51000 102390
rect 50948 102326 51000 102332
rect 50856 102180 50908 102186
rect 50856 102122 50908 102128
rect 50764 102112 50816 102118
rect 50764 102054 50816 102060
rect 50580 102044 50632 102050
rect 50580 101986 50632 101992
rect 51052 101778 51080 112759
rect 51144 101982 51172 113983
rect 51222 113912 51278 113921
rect 51222 113847 51224 113856
rect 51276 113847 51278 113856
rect 57572 113876 57624 113882
rect 51224 113818 51276 113824
rect 57572 113818 57624 113824
rect 52604 112992 52656 112998
rect 52604 112934 52656 112940
rect 52616 112318 52644 112934
rect 52604 112312 52656 112318
rect 52604 112254 52656 112260
rect 51132 101976 51184 101982
rect 51132 101918 51184 101924
rect 51040 101772 51092 101778
rect 51040 101714 51092 101720
rect 45152 101704 45204 101710
rect 45152 101646 45204 101652
rect 45060 101432 45112 101438
rect 45060 101374 45112 101380
rect 42944 101364 42996 101370
rect 42944 101306 42996 101312
rect 41838 95280 41894 95289
rect 41760 95238 41838 95266
rect 41838 95215 41894 95224
rect 22336 90280 22388 90286
rect 22336 90222 22388 90228
rect 22348 89849 22376 90222
rect 22334 89840 22390 89849
rect 22334 89775 22390 89784
rect 44414 84808 44470 84817
rect 44414 84743 44470 84752
rect 22334 83176 22390 83185
rect 22334 83111 22390 83120
rect 22348 82058 22376 83111
rect 22336 82052 22388 82058
rect 22336 81994 22388 82000
rect 44428 76521 44456 84743
rect 44414 76512 44470 76521
rect 44414 76447 44470 76456
rect 52616 75054 52644 112254
rect 56468 101772 56520 101778
rect 56468 101714 56520 101720
rect 56480 99740 56508 101714
rect 57584 99740 57612 113818
rect 59332 108238 59360 115110
rect 61600 114822 61936 114850
rect 62980 114822 63316 114850
rect 61908 112318 61936 114822
rect 61896 112312 61948 112318
rect 61896 112254 61948 112260
rect 61908 111201 61936 112254
rect 61894 111192 61950 111201
rect 61894 111127 61950 111136
rect 63288 110890 63316 114822
rect 64116 114822 64452 114850
rect 65312 114822 65832 114850
rect 66508 114822 67304 114850
rect 67888 114822 68684 114850
rect 69268 114822 70156 114850
rect 70648 114822 71536 114850
rect 72028 114822 73008 114850
rect 73500 114822 74388 114850
rect 75524 114822 75860 114850
rect 76904 114822 77240 114850
rect 77548 114822 78712 114850
rect 79756 114822 80092 114850
rect 81228 114822 81564 114850
rect 82608 114822 82944 114850
rect 84080 114822 84416 114850
rect 85460 114822 85796 114850
rect 87208 114822 87268 114850
rect 90120 114822 90456 114850
rect 64116 113338 64144 114822
rect 64104 113332 64156 113338
rect 64104 113274 64156 113280
rect 63276 110884 63328 110890
rect 63276 110826 63328 110832
rect 59320 108232 59372 108238
rect 59320 108174 59372 108180
rect 59412 108164 59464 108170
rect 59412 108106 59464 108112
rect 59424 101982 59452 108106
rect 59780 102384 59832 102390
rect 59780 102326 59832 102332
rect 58676 101976 58728 101982
rect 58676 101918 58728 101924
rect 59412 101976 59464 101982
rect 59412 101918 59464 101924
rect 58688 99740 58716 101918
rect 59792 99740 59820 102326
rect 60884 102248 60936 102254
rect 60884 102190 60936 102196
rect 60896 99740 60924 102190
rect 61988 102180 62040 102186
rect 61988 102122 62040 102128
rect 62000 99740 62028 102122
rect 63092 102112 63144 102118
rect 63092 102054 63144 102060
rect 63104 99740 63132 102054
rect 64196 102044 64248 102050
rect 64196 101986 64248 101992
rect 64208 99740 64236 101986
rect 65312 99740 65340 114822
rect 66508 101386 66536 114822
rect 67888 101386 67916 114822
rect 66416 101358 66536 101386
rect 67704 101358 67916 101386
rect 69268 101370 69296 114822
rect 70648 101370 70676 114822
rect 72028 101370 72056 114822
rect 73500 101438 73528 114822
rect 75524 111094 75552 114822
rect 74040 111088 74092 111094
rect 74040 111030 74092 111036
rect 75512 111088 75564 111094
rect 75512 111030 75564 111036
rect 72384 101432 72436 101438
rect 72384 101374 72436 101380
rect 73488 101432 73540 101438
rect 73488 101374 73540 101380
rect 68612 101364 68664 101370
rect 66416 99740 66444 101358
rect 67704 99754 67732 101358
rect 68612 101306 68664 101312
rect 69256 101364 69308 101370
rect 69256 101306 69308 101312
rect 69808 101364 69860 101370
rect 69808 101306 69860 101312
rect 70636 101364 70688 101370
rect 70636 101306 70688 101312
rect 70912 101364 70964 101370
rect 70912 101306 70964 101312
rect 72016 101364 72068 101370
rect 72016 101306 72068 101312
rect 67534 99726 67732 99754
rect 68624 99740 68652 101306
rect 69820 99740 69848 101306
rect 70924 99740 70952 101306
rect 72396 99754 72424 101374
rect 74052 101370 74080 111030
rect 76904 111026 76932 114822
rect 77444 111088 77496 111094
rect 77444 111030 77496 111036
rect 74684 111020 74736 111026
rect 74684 110962 74736 110968
rect 76892 111020 76944 111026
rect 76892 110962 76944 110968
rect 73120 101364 73172 101370
rect 73120 101306 73172 101312
rect 74040 101364 74092 101370
rect 74040 101306 74092 101312
rect 72042 99726 72424 99754
rect 73132 99740 73160 101306
rect 74696 99754 74724 110962
rect 75328 101568 75380 101574
rect 75328 101510 75380 101516
rect 74250 99726 74724 99754
rect 75340 99740 75368 101510
rect 77456 101370 77484 111030
rect 77548 101574 77576 114822
rect 79652 111156 79704 111162
rect 79652 111098 79704 111104
rect 79560 111020 79612 111026
rect 79560 110962 79612 110968
rect 77536 101568 77588 101574
rect 77536 101510 77588 101516
rect 79572 101438 79600 110962
rect 77536 101432 77588 101438
rect 77536 101374 77588 101380
rect 79560 101432 79612 101438
rect 79560 101374 79612 101380
rect 76432 101364 76484 101370
rect 76432 101306 76484 101312
rect 77444 101364 77496 101370
rect 77444 101306 77496 101312
rect 76444 99740 76472 101306
rect 77548 99740 77576 101374
rect 79664 101370 79692 111098
rect 79756 111094 79784 114822
rect 80940 111496 80992 111502
rect 80940 111438 80992 111444
rect 79744 111088 79796 111094
rect 79744 111030 79796 111036
rect 80848 101432 80900 101438
rect 80848 101374 80900 101380
rect 78640 101364 78692 101370
rect 78640 101306 78692 101312
rect 79652 101364 79704 101370
rect 79652 101306 79704 101312
rect 79744 101364 79796 101370
rect 79744 101306 79796 101312
rect 78652 99740 78680 101306
rect 79756 99740 79784 101306
rect 80860 99740 80888 101374
rect 80952 101370 80980 111438
rect 81228 111026 81256 114822
rect 82320 111632 82372 111638
rect 82320 111574 82372 111580
rect 81216 111020 81268 111026
rect 81216 110962 81268 110968
rect 82332 101438 82360 111574
rect 82608 111162 82636 114822
rect 83700 111564 83752 111570
rect 83700 111506 83752 111512
rect 82596 111156 82648 111162
rect 82596 111098 82648 111104
rect 83148 101976 83200 101982
rect 83148 101918 83200 101924
rect 82320 101432 82372 101438
rect 82320 101374 82372 101380
rect 80940 101364 80992 101370
rect 80940 101306 80992 101312
rect 81952 101364 82004 101370
rect 81952 101306 82004 101312
rect 81964 99740 81992 101306
rect 83160 99740 83188 101918
rect 83712 101370 83740 111506
rect 84080 111502 84108 114822
rect 85460 111638 85488 114822
rect 85724 112380 85776 112386
rect 85724 112322 85776 112328
rect 85448 111632 85500 111638
rect 85448 111574 85500 111580
rect 84068 111496 84120 111502
rect 84068 111438 84120 111444
rect 83700 101364 83752 101370
rect 83700 101306 83752 101312
rect 85736 99754 85764 112322
rect 87208 111570 87236 114822
rect 90428 112250 90456 114822
rect 90416 112244 90468 112250
rect 90416 112186 90468 112192
rect 87196 111564 87248 111570
rect 87196 111506 87248 111512
rect 88668 102112 88720 102118
rect 88668 102054 88720 102060
rect 87564 102044 87616 102050
rect 87564 101986 87616 101992
rect 86460 101976 86512 101982
rect 86460 101918 86512 101924
rect 85382 99726 85764 99754
rect 86472 99740 86500 101918
rect 87576 99740 87604 101986
rect 88680 99740 88708 102054
rect 90612 101370 90640 115110
rect 89772 101364 89824 101370
rect 89772 101306 89824 101312
rect 90600 101364 90652 101370
rect 90600 101306 90652 101312
rect 89784 99740 89812 101306
rect 91256 99754 91284 115178
rect 92636 101370 92664 116470
rect 92900 116460 92952 116466
rect 92900 116402 92952 116408
rect 92716 116392 92768 116398
rect 92714 116360 92716 116369
rect 92768 116360 92770 116369
rect 92714 116295 92770 116304
rect 92808 116324 92860 116330
rect 92808 116266 92860 116272
rect 92820 115961 92848 116266
rect 92806 115952 92862 115961
rect 92806 115887 92862 115896
rect 92912 115553 92940 116402
rect 92898 115544 92954 115553
rect 92898 115479 92954 115488
rect 93360 112244 93412 112250
rect 93360 112186 93412 112192
rect 93372 102458 93400 112186
rect 93360 102452 93412 102458
rect 93360 102394 93412 102400
rect 94016 101370 94044 116538
rect 94188 102452 94240 102458
rect 94188 102394 94240 102400
rect 91980 101364 92032 101370
rect 91980 101306 92032 101312
rect 92624 101364 92676 101370
rect 92624 101306 92676 101312
rect 93084 101364 93136 101370
rect 93084 101306 93136 101312
rect 94004 101364 94056 101370
rect 94004 101306 94056 101312
rect 90902 99726 91284 99754
rect 91992 99740 92020 101306
rect 93096 99740 93124 101306
rect 94200 99740 94228 102394
rect 53338 79912 53394 79921
rect 53338 79847 53394 79856
rect 44416 75048 44468 75054
rect 44416 74990 44468 74996
rect 52604 75048 52656 75054
rect 52604 74990 52656 74996
rect 44428 74753 44456 74990
rect 44414 74744 44470 74753
rect 52616 74714 52644 74990
rect 44414 74679 44470 74688
rect 52604 74708 52656 74714
rect 52604 74650 52656 74656
rect 53352 69857 53380 79847
rect 53432 74708 53484 74714
rect 53432 74650 53484 74656
rect 53338 69848 53394 69857
rect 53338 69783 53394 69792
rect 53444 66593 53472 74650
rect 53430 66584 53486 66593
rect 53430 66519 53486 66528
rect 53982 66584 54038 66593
rect 53982 66519 54038 66528
rect 44506 64816 44562 64825
rect 44506 64751 44562 64760
rect 18104 63624 18156 63630
rect 18104 63566 18156 63572
rect 22336 63624 22388 63630
rect 22336 63566 22388 63572
rect 22348 63193 22376 63566
rect 22334 63184 22390 63193
rect 22334 63119 22390 63128
rect 25108 59878 26134 59906
rect 26502 59878 26608 59906
rect 22888 50228 22940 50234
rect 22888 50170 22940 50176
rect 22244 50024 22296 50030
rect 22244 49966 22296 49972
rect 20220 49548 20272 49554
rect 20220 49490 20272 49496
rect 20232 46428 20260 49490
rect 21508 49480 21560 49486
rect 21508 49422 21560 49428
rect 20864 49072 20916 49078
rect 20864 49014 20916 49020
rect 20876 46428 20904 49014
rect 21520 46428 21548 49422
rect 22256 46428 22284 49966
rect 22900 46428 22928 50170
rect 24912 50160 24964 50166
rect 24912 50102 24964 50108
rect 24268 50092 24320 50098
rect 24268 50034 24320 50040
rect 23624 49956 23676 49962
rect 23624 49898 23676 49904
rect 23636 46428 23664 49898
rect 24280 46428 24308 50034
rect 24924 46428 24952 50102
rect 25108 49078 25136 59878
rect 26476 57164 26528 57170
rect 26476 57106 26528 57112
rect 26488 49962 26516 57106
rect 26476 49956 26528 49962
rect 26476 49898 26528 49904
rect 26292 49684 26344 49690
rect 26292 49626 26344 49632
rect 25648 49140 25700 49146
rect 25648 49082 25700 49088
rect 25096 49072 25148 49078
rect 25096 49014 25148 49020
rect 25660 46428 25688 49082
rect 26304 46428 26332 49626
rect 26580 49486 26608 59878
rect 26672 59878 26870 59906
rect 26948 59878 27330 59906
rect 27408 59878 27698 59906
rect 27868 59878 28066 59906
rect 28144 59878 28526 59906
rect 28604 59878 28894 59906
rect 29262 59878 29368 59906
rect 26672 54450 26700 59878
rect 26948 57050 26976 59878
rect 27408 57170 27436 59878
rect 27396 57164 27448 57170
rect 27396 57106 27448 57112
rect 26764 57022 26976 57050
rect 26660 54444 26712 54450
rect 26660 54386 26712 54392
rect 26764 50234 26792 57022
rect 26844 54444 26896 54450
rect 26844 54386 26896 54392
rect 26752 50228 26804 50234
rect 26752 50170 26804 50176
rect 26856 50030 26884 54386
rect 27868 50098 27896 59878
rect 28144 57186 28172 59878
rect 27960 57158 28172 57186
rect 27960 50166 27988 57158
rect 28604 57050 28632 59878
rect 29144 57368 29196 57374
rect 29144 57310 29196 57316
rect 28052 57022 28632 57050
rect 27948 50160 28000 50166
rect 27948 50102 28000 50108
rect 27856 50092 27908 50098
rect 27856 50034 27908 50040
rect 26844 50024 26896 50030
rect 26844 49966 26896 49972
rect 27672 50024 27724 50030
rect 27672 49966 27724 49972
rect 26568 49480 26620 49486
rect 26568 49422 26620 49428
rect 27028 49140 27080 49146
rect 27028 49082 27080 49088
rect 27040 46428 27068 49082
rect 27684 46428 27712 49966
rect 28052 49214 28080 57022
rect 29156 50234 29184 57310
rect 28316 50228 28368 50234
rect 28316 50170 28368 50176
rect 29144 50228 29196 50234
rect 29144 50170 29196 50176
rect 28040 49208 28092 49214
rect 28040 49150 28092 49156
rect 28328 46428 28356 50170
rect 29052 50092 29104 50098
rect 29052 50034 29104 50040
rect 29064 46428 29092 50034
rect 29340 49690 29368 59878
rect 29524 59878 29722 59906
rect 29800 59878 30090 59906
rect 29420 57164 29472 57170
rect 29420 57106 29472 57112
rect 29432 50030 29460 57106
rect 29420 50024 29472 50030
rect 29420 49966 29472 49972
rect 29328 49684 29380 49690
rect 29328 49626 29380 49632
rect 29524 49146 29552 59878
rect 29800 57170 29828 59878
rect 30444 57374 30472 59892
rect 30720 59878 30918 59906
rect 30432 57368 30484 57374
rect 30432 57310 30484 57316
rect 30432 57232 30484 57238
rect 30432 57174 30484 57180
rect 29788 57164 29840 57170
rect 29788 57106 29840 57112
rect 30444 50234 30472 57174
rect 30524 57164 30576 57170
rect 30524 57106 30576 57112
rect 29696 50228 29748 50234
rect 29696 50170 29748 50176
rect 30432 50228 30484 50234
rect 30432 50170 30484 50176
rect 29512 49140 29564 49146
rect 29512 49082 29564 49088
rect 29708 46428 29736 50170
rect 30536 46442 30564 57106
rect 30720 50098 30748 59878
rect 31272 57238 31300 59892
rect 31260 57232 31312 57238
rect 31260 57174 31312 57180
rect 31640 57170 31668 59892
rect 32008 59878 32114 59906
rect 32008 57186 32036 59878
rect 32468 57238 32496 59892
rect 31628 57164 31680 57170
rect 31628 57106 31680 57112
rect 31824 57158 32036 57186
rect 32456 57232 32508 57238
rect 32456 57174 32508 57180
rect 32836 57170 32864 59892
rect 33296 57170 33324 59892
rect 33480 59878 33678 59906
rect 32088 57164 32140 57170
rect 31824 50234 31852 57158
rect 32088 57106 32140 57112
rect 32824 57164 32876 57170
rect 32824 57106 32876 57112
rect 33284 57164 33336 57170
rect 33284 57106 33336 57112
rect 33376 57164 33428 57170
rect 33376 57106 33428 57112
rect 31904 57096 31956 57102
rect 31904 57038 31956 57044
rect 31996 57096 32048 57102
rect 31996 57038 32048 57044
rect 31076 50228 31128 50234
rect 31076 50170 31128 50176
rect 31812 50228 31864 50234
rect 31812 50170 31864 50176
rect 30708 50092 30760 50098
rect 30708 50034 30760 50040
rect 30458 46414 30564 46442
rect 31088 46428 31116 50170
rect 31916 46442 31944 57038
rect 32008 50302 32036 57038
rect 31996 50296 32048 50302
rect 31996 50238 32048 50244
rect 31838 46414 31944 46442
rect 32100 46442 32128 57106
rect 33388 50302 33416 57106
rect 32732 50296 32784 50302
rect 32732 50238 32784 50244
rect 33376 50296 33428 50302
rect 33376 50238 33428 50244
rect 32744 46442 32772 50238
rect 33480 46442 33508 59878
rect 34124 57170 34152 59892
rect 34506 59878 34704 59906
rect 34112 57164 34164 57170
rect 34112 57106 34164 57112
rect 34204 50296 34256 50302
rect 34204 50238 34256 50244
rect 34216 46442 34244 50238
rect 34676 48890 34704 59878
rect 34860 49026 34888 59892
rect 35320 57170 35348 59892
rect 35702 59878 35992 59906
rect 35308 57164 35360 57170
rect 35308 57106 35360 57112
rect 35964 50114 35992 59878
rect 36056 58682 36084 59892
rect 36056 58654 36176 58682
rect 36148 58530 36176 58654
rect 36136 58524 36188 58530
rect 36136 58466 36188 58472
rect 36516 57170 36544 59892
rect 36884 57306 36912 59892
rect 36872 57300 36924 57306
rect 36872 57242 36924 57248
rect 37252 57238 37280 59892
rect 37516 58524 37568 58530
rect 37516 58466 37568 58472
rect 37240 57232 37292 57238
rect 37240 57174 37292 57180
rect 36044 57164 36096 57170
rect 36044 57106 36096 57112
rect 36504 57164 36556 57170
rect 36504 57106 36556 57112
rect 36056 50250 36084 57106
rect 36056 50222 36268 50250
rect 35964 50086 36176 50114
rect 34860 48998 35624 49026
rect 34676 48862 34888 48890
rect 34860 46442 34888 48862
rect 35596 46442 35624 48998
rect 36148 48942 36176 50086
rect 36136 48936 36188 48942
rect 36136 48878 36188 48884
rect 36240 46442 36268 50222
rect 37240 48936 37292 48942
rect 37240 48878 37292 48884
rect 32100 46414 32482 46442
rect 32744 46414 33126 46442
rect 33480 46414 33862 46442
rect 34216 46414 34506 46442
rect 34860 46414 35242 46442
rect 35596 46414 35886 46442
rect 36240 46414 36530 46442
rect 37252 46428 37280 48878
rect 37528 46442 37556 58466
rect 37712 57374 37740 59892
rect 37700 57368 37752 57374
rect 37700 57310 37752 57316
rect 38080 57170 38108 59892
rect 38160 57300 38212 57306
rect 38160 57242 38212 57248
rect 37608 57164 37660 57170
rect 37608 57106 37660 57112
rect 38068 57164 38120 57170
rect 38068 57106 38120 57112
rect 37620 46714 37648 57106
rect 38172 49146 38200 57242
rect 38448 57238 38476 59892
rect 38908 57442 38936 59892
rect 39276 57646 39304 59892
rect 39264 57640 39316 57646
rect 39264 57582 39316 57588
rect 39644 57510 39672 59892
rect 40104 57578 40132 59892
rect 40092 57572 40144 57578
rect 40092 57514 40144 57520
rect 39632 57504 39684 57510
rect 39632 57446 39684 57452
rect 38896 57436 38948 57442
rect 38896 57378 38948 57384
rect 40276 57368 40328 57374
rect 40276 57310 40328 57316
rect 38252 57232 38304 57238
rect 38252 57174 38304 57180
rect 38436 57232 38488 57238
rect 38436 57174 38488 57180
rect 38160 49140 38212 49146
rect 38160 49082 38212 49088
rect 38264 49078 38292 57174
rect 39264 49140 39316 49146
rect 39264 49082 39316 49088
rect 38252 49072 38304 49078
rect 38252 49014 38304 49020
rect 37620 46686 38200 46714
rect 38172 46442 38200 46686
rect 37528 46414 37910 46442
rect 38172 46414 38646 46442
rect 39276 46428 39304 49082
rect 40000 49072 40052 49078
rect 40000 49014 40052 49020
rect 40012 46428 40040 49014
rect 40288 46442 40316 57310
rect 40472 57306 40500 59892
rect 40840 57374 40868 59892
rect 40828 57368 40880 57374
rect 40828 57310 40880 57316
rect 40460 57300 40512 57306
rect 40460 57242 40512 57248
rect 40920 57232 40972 57238
rect 40920 57174 40972 57180
rect 40368 57164 40420 57170
rect 40368 57106 40420 57112
rect 40380 46714 40408 57106
rect 40932 50234 40960 57174
rect 41300 57170 41328 59892
rect 41668 58258 41696 59892
rect 41656 58252 41708 58258
rect 41656 58194 41708 58200
rect 43036 57640 43088 57646
rect 43036 57582 43088 57588
rect 41840 57436 41892 57442
rect 41840 57378 41892 57384
rect 41288 57164 41340 57170
rect 41288 57106 41340 57112
rect 41852 50302 41880 57378
rect 41840 50296 41892 50302
rect 41840 50238 41892 50244
rect 42300 50296 42352 50302
rect 42300 50238 42352 50244
rect 40920 50228 40972 50234
rect 40920 50170 40972 50176
rect 42024 50228 42076 50234
rect 42024 50170 42076 50176
rect 40380 46686 40960 46714
rect 40932 46442 40960 46686
rect 40288 46414 40670 46442
rect 40932 46414 41314 46442
rect 42036 46428 42064 50170
rect 42312 46442 42340 50238
rect 43048 46442 43076 57582
rect 43680 57572 43732 57578
rect 43680 57514 43732 57520
rect 43128 57504 43180 57510
rect 43128 57446 43180 57452
rect 43140 46714 43168 57446
rect 43692 48942 43720 57514
rect 44520 49554 44548 64751
rect 46440 58252 46492 58258
rect 46440 58194 46492 58200
rect 45152 57368 45204 57374
rect 45152 57310 45204 57316
rect 44600 57300 44652 57306
rect 44600 57242 44652 57248
rect 44612 50386 44640 57242
rect 45060 57164 45112 57170
rect 45060 57106 45112 57112
rect 44612 50358 45008 50386
rect 44508 49548 44560 49554
rect 44508 49490 44560 49496
rect 43680 48936 43732 48942
rect 43680 48878 43732 48884
rect 44692 48936 44744 48942
rect 44692 48878 44744 48884
rect 43140 46686 43720 46714
rect 43692 46442 43720 46686
rect 42312 46414 42694 46442
rect 43048 46414 43430 46442
rect 43692 46414 44074 46442
rect 44704 46428 44732 48878
rect 44980 46442 45008 50358
rect 45072 49010 45100 57106
rect 45060 49004 45112 49010
rect 45060 48946 45112 48952
rect 45164 48942 45192 57310
rect 46452 48942 46480 58194
rect 46808 49004 46860 49010
rect 46808 48946 46860 48952
rect 45152 48936 45204 48942
rect 45152 48878 45204 48884
rect 46072 48936 46124 48942
rect 46072 48878 46124 48884
rect 46440 48936 46492 48942
rect 46440 48878 46492 48884
rect 44980 46414 45454 46442
rect 46084 46428 46112 48878
rect 46820 46428 46848 48946
rect 47452 48936 47504 48942
rect 47452 48878 47504 48884
rect 47464 46428 47492 48878
rect 50764 46556 50816 46562
rect 50764 46498 50816 46504
rect 49936 46488 49988 46494
rect 49936 46430 49988 46436
rect 49948 46329 49976 46430
rect 50580 46420 50632 46426
rect 50580 46362 50632 46368
rect 49934 46320 49990 46329
rect 49934 46255 49990 46264
rect 50026 44008 50082 44017
rect 50026 43943 50082 43952
rect 49934 43600 49990 43609
rect 50040 43570 50068 43943
rect 49934 43535 49990 43544
rect 50028 43564 50080 43570
rect 49948 43366 49976 43535
rect 50028 43506 50080 43512
rect 49936 43360 49988 43366
rect 49936 43302 49988 43308
rect 50026 42784 50082 42793
rect 50026 42719 50082 42728
rect 49934 42512 49990 42521
rect 49934 42447 49936 42456
rect 49988 42447 49990 42456
rect 49936 42418 49988 42424
rect 50040 42346 50068 42719
rect 50028 42340 50080 42346
rect 50028 42282 50080 42288
rect 49934 42104 49990 42113
rect 49934 42039 49990 42048
rect 49948 42006 49976 42039
rect 49936 42000 49988 42006
rect 18102 41968 18158 41977
rect 14700 41932 14752 41938
rect 49936 41942 49988 41948
rect 18102 41903 18104 41912
rect 14700 41874 14752 41880
rect 18156 41903 18158 41912
rect 18104 41874 18156 41880
rect 50026 41016 50082 41025
rect 50026 40951 50082 40960
rect 49934 40744 49990 40753
rect 49934 40679 49936 40688
rect 49988 40679 49990 40688
rect 49936 40650 49988 40656
rect 50040 40646 50068 40951
rect 50028 40640 50080 40646
rect 50028 40582 50080 40588
rect 50210 37344 50266 37353
rect 50210 37279 50266 37288
rect 50224 36498 50252 37279
rect 50212 36492 50264 36498
rect 50212 36434 50264 36440
rect 50026 33128 50082 33137
rect 50026 33063 50082 33072
rect 50040 32554 50068 33063
rect 50028 32548 50080 32554
rect 50028 32490 50080 32496
rect 18102 32448 18158 32457
rect 18102 32383 18158 32392
rect 13318 20616 13374 20625
rect 13318 20551 13374 20560
rect 18116 18478 18144 32383
rect 50026 31904 50082 31913
rect 50026 31839 50082 31848
rect 50040 31330 50068 31839
rect 50028 31324 50080 31330
rect 50028 31266 50080 31272
rect 50026 27552 50082 27561
rect 50026 27487 50082 27496
rect 50040 26842 50068 27487
rect 50028 26836 50080 26842
rect 50028 26778 50080 26784
rect 50304 25408 50356 25414
rect 50304 25350 50356 25356
rect 50316 21169 50344 25350
rect 50394 23336 50450 23345
rect 50394 23271 50450 23280
rect 50408 22694 50436 23271
rect 50396 22688 50448 22694
rect 50396 22630 50448 22636
rect 50592 22234 50620 46362
rect 50672 46216 50724 46222
rect 50672 46158 50724 46164
rect 50684 25414 50712 46158
rect 50672 25408 50724 25414
rect 50672 25350 50724 25356
rect 50500 22206 50620 22234
rect 50302 21160 50358 21169
rect 50302 21095 50358 21104
rect 50500 19809 50528 22206
rect 50578 22112 50634 22121
rect 50578 22047 50634 22056
rect 50592 21334 50620 22047
rect 50580 21328 50632 21334
rect 50580 21270 50632 21276
rect 50486 19800 50542 19809
rect 50486 19735 50542 19744
rect 50776 19265 50804 46498
rect 51040 46352 51092 46358
rect 51040 46294 51092 46300
rect 50856 46284 50908 46290
rect 50856 46226 50908 46232
rect 50868 21033 50896 46226
rect 50948 46148 51000 46154
rect 50948 46090 51000 46096
rect 50960 21985 50988 46090
rect 50946 21976 51002 21985
rect 50946 21911 51002 21920
rect 50854 21024 50910 21033
rect 50854 20959 50910 20968
rect 51052 20489 51080 46294
rect 53338 45232 53394 45241
rect 53338 45167 53394 45176
rect 53246 44960 53302 44969
rect 53246 44895 53302 44904
rect 53260 44794 53288 44895
rect 53248 44788 53300 44794
rect 53248 44730 53300 44736
rect 53352 44726 53380 45167
rect 53340 44720 53392 44726
rect 53340 44662 53392 44668
rect 51130 39792 51186 39801
rect 51130 39727 51186 39736
rect 51144 39218 51172 39727
rect 51222 39384 51278 39393
rect 51222 39319 51278 39328
rect 51236 39286 51264 39319
rect 51224 39280 51276 39286
rect 51224 39222 51276 39228
rect 51132 39212 51184 39218
rect 51132 39154 51184 39160
rect 51130 38568 51186 38577
rect 51130 38503 51186 38512
rect 51144 37858 51172 38503
rect 51222 38160 51278 38169
rect 51222 38095 51278 38104
rect 51236 37926 51264 38095
rect 51224 37920 51276 37926
rect 51224 37862 51276 37868
rect 51132 37852 51184 37858
rect 51132 37794 51184 37800
rect 51222 36800 51278 36809
rect 51222 36735 51278 36744
rect 51132 36628 51184 36634
rect 51132 36570 51184 36576
rect 51144 36537 51172 36570
rect 51236 36566 51264 36735
rect 51224 36560 51276 36566
rect 51130 36528 51186 36537
rect 51224 36502 51276 36508
rect 51130 36463 51186 36472
rect 51222 35712 51278 35721
rect 51222 35647 51278 35656
rect 51236 35410 51264 35647
rect 51224 35404 51276 35410
rect 51224 35346 51276 35352
rect 51222 35168 51278 35177
rect 51222 35103 51224 35112
rect 51276 35103 51278 35112
rect 51224 35074 51276 35080
rect 51130 34216 51186 34225
rect 51130 34151 51186 34160
rect 51144 33710 51172 34151
rect 51222 33944 51278 33953
rect 51222 33879 51278 33888
rect 51236 33778 51264 33879
rect 51224 33772 51276 33778
rect 51224 33714 51276 33720
rect 51132 33704 51184 33710
rect 51132 33646 51184 33652
rect 51222 32584 51278 32593
rect 51222 32519 51278 32528
rect 51236 32350 51264 32519
rect 51224 32344 51276 32350
rect 51224 32286 51276 32292
rect 51222 31496 51278 31505
rect 51222 31431 51278 31440
rect 51236 31194 51264 31431
rect 51224 31188 51276 31194
rect 51224 31130 51276 31136
rect 51224 30984 51276 30990
rect 51222 30952 51224 30961
rect 51276 30952 51278 30961
rect 51222 30887 51278 30896
rect 51130 30000 51186 30009
rect 51130 29935 51186 29944
rect 51144 29562 51172 29935
rect 51222 29728 51278 29737
rect 51222 29663 51224 29672
rect 51276 29663 51278 29672
rect 51224 29634 51276 29640
rect 51132 29556 51184 29562
rect 51132 29498 51184 29504
rect 51130 28776 51186 28785
rect 51130 28711 51186 28720
rect 51144 28338 51172 28711
rect 51222 28368 51278 28377
rect 51132 28332 51184 28338
rect 51222 28303 51278 28312
rect 51132 28274 51184 28280
rect 51236 28202 51264 28303
rect 51224 28196 51276 28202
rect 51224 28138 51276 28144
rect 51222 27144 51278 27153
rect 51222 27079 51278 27088
rect 51132 26972 51184 26978
rect 51132 26914 51184 26920
rect 51144 26881 51172 26914
rect 51236 26910 51264 27079
rect 51224 26904 51276 26910
rect 51130 26872 51186 26881
rect 51224 26846 51276 26852
rect 51130 26807 51186 26816
rect 51130 25784 51186 25793
rect 51130 25719 51186 25728
rect 51144 25482 51172 25719
rect 51224 25544 51276 25550
rect 51222 25512 51224 25521
rect 51276 25512 51278 25521
rect 51132 25476 51184 25482
rect 51222 25447 51278 25456
rect 51132 25418 51184 25424
rect 51130 24560 51186 24569
rect 51130 24495 51186 24504
rect 51144 24054 51172 24495
rect 51222 24288 51278 24297
rect 51222 24223 51278 24232
rect 51236 24122 51264 24223
rect 51224 24116 51276 24122
rect 51224 24058 51276 24064
rect 51132 24048 51184 24054
rect 51132 23990 51184 23996
rect 51222 22928 51278 22937
rect 51222 22863 51278 22872
rect 51236 22762 51264 22863
rect 53996 22801 54024 66519
rect 59240 58433 59268 59892
rect 59226 58424 59282 58433
rect 72580 58394 72608 59892
rect 79204 58394 79232 59892
rect 59226 58359 59282 58368
rect 72568 58388 72620 58394
rect 72568 58330 72620 58336
rect 79192 58388 79244 58394
rect 79192 58330 79244 58336
rect 70544 57980 70596 57986
rect 70544 57922 70596 57928
rect 61344 46556 61396 46562
rect 61344 46498 61396 46504
rect 58952 46488 59004 46494
rect 58952 46430 59004 46436
rect 58216 44720 58268 44726
rect 58216 44662 58268 44668
rect 58228 43881 58256 44662
rect 58964 44425 58992 46430
rect 61356 44810 61384 46498
rect 62816 46420 62868 46426
rect 62816 46362 62868 46368
rect 62828 44810 62856 46362
rect 64288 46352 64340 46358
rect 64288 46294 64340 46300
rect 64300 44810 64328 46294
rect 65760 46284 65812 46290
rect 65760 46226 65812 46232
rect 65772 44810 65800 46226
rect 67324 46216 67376 46222
rect 67324 46158 67376 46164
rect 67336 44810 67364 46158
rect 68796 46148 68848 46154
rect 68796 46090 68848 46096
rect 68808 44810 68836 46090
rect 70556 44810 70584 57922
rect 72580 57918 72608 58330
rect 72568 57912 72620 57918
rect 72568 57854 72620 57860
rect 79204 57850 79232 58330
rect 92544 57986 92572 59892
rect 95396 58326 95424 151694
rect 95384 58320 95436 58326
rect 95384 58262 95436 58268
rect 92532 57980 92584 57986
rect 92532 57922 92584 57928
rect 79192 57844 79244 57850
rect 79192 57786 79244 57792
rect 96132 48874 96160 236558
rect 99628 235942 99656 244242
rect 121420 236684 121472 236690
rect 121420 236626 121472 236632
rect 99616 235936 99668 235942
rect 99616 235878 99668 235884
rect 107436 235392 107488 235398
rect 107436 235334 107488 235340
rect 107448 235058 107476 235334
rect 114428 235256 114480 235262
rect 114428 235198 114480 235204
rect 107436 235052 107488 235058
rect 107436 234994 107488 235000
rect 107448 234788 107476 234994
rect 114440 234788 114468 235198
rect 121432 234788 121460 236626
rect 135876 235942 135904 244344
rect 171848 241382 171876 244344
rect 207820 241382 207848 244344
rect 171836 241376 171888 241382
rect 171836 241318 171888 241324
rect 174044 241376 174096 241382
rect 174044 241318 174096 241324
rect 207808 241376 207860 241382
rect 207808 241318 207860 241324
rect 135864 235936 135916 235942
rect 135864 235878 135916 235884
rect 169536 235936 169588 235942
rect 169536 235878 169588 235884
rect 166224 235868 166276 235874
rect 166224 235810 166276 235816
rect 139452 235392 139504 235398
rect 139452 235334 139504 235340
rect 139464 235233 139492 235334
rect 159508 235256 159560 235262
rect 139450 235224 139506 235233
rect 159508 235198 159560 235204
rect 163554 235224 163610 235233
rect 139450 235159 139506 235168
rect 146536 235188 146588 235194
rect 146536 235130 146588 235136
rect 156840 235188 156892 235194
rect 156840 235130 156892 235136
rect 134758 234544 134814 234553
rect 134758 234479 134760 234488
rect 134812 234479 134814 234488
rect 134760 234450 134812 234456
rect 101178 234000 101234 234009
rect 101178 233935 101234 233944
rect 134758 234000 134814 234009
rect 134758 233935 134814 233944
rect 101192 233902 101220 233935
rect 134772 233902 134800 233935
rect 101180 233896 101232 233902
rect 101180 233838 101232 233844
rect 134760 233896 134812 233902
rect 134760 233838 134812 233844
rect 142304 233896 142356 233902
rect 142304 233838 142356 233844
rect 134850 233456 134906 233465
rect 134850 233391 134906 233400
rect 101362 233184 101418 233193
rect 101362 233119 101418 233128
rect 101376 233086 101404 233119
rect 101364 233080 101416 233086
rect 101364 233022 101416 233028
rect 101730 232912 101786 232921
rect 101730 232847 101786 232856
rect 134758 232912 134814 232921
rect 134758 232847 134814 232856
rect 101744 232474 101772 232847
rect 134772 232746 134800 232847
rect 134760 232740 134812 232746
rect 134760 232682 134812 232688
rect 134864 232678 134892 233391
rect 142316 233057 142344 233838
rect 142302 233048 142358 233057
rect 142302 232983 142358 232992
rect 146548 232762 146576 235130
rect 156852 232762 156880 235130
rect 142212 232740 142264 232746
rect 146548 232734 146608 232762
rect 156544 232734 156880 232762
rect 159520 232762 159548 235198
rect 163554 235159 163610 235168
rect 163568 232762 163596 235159
rect 159520 232734 159856 232762
rect 163260 232734 163596 232762
rect 166236 232762 166264 235810
rect 169548 232762 169576 235878
rect 174056 235262 174084 241318
rect 173492 235256 173544 235262
rect 173492 235198 173544 235204
rect 174044 235256 174096 235262
rect 174044 235198 174096 235204
rect 173504 232762 173532 235198
rect 215628 235188 215680 235194
rect 215628 235130 215680 235136
rect 185266 234544 185322 234553
rect 185266 234479 185322 234488
rect 185174 234000 185230 234009
rect 185174 233935 185230 233944
rect 185188 233902 185216 233935
rect 180300 233896 180352 233902
rect 180300 233838 180352 233844
rect 185176 233896 185228 233902
rect 185176 233838 185228 233844
rect 177724 233080 177776 233086
rect 177724 233022 177776 233028
rect 177736 232785 177764 233022
rect 166236 232734 166572 232762
rect 169548 232734 169884 232762
rect 173196 232734 173532 232762
rect 177722 232776 177778 232785
rect 177722 232711 177778 232720
rect 142212 232682 142264 232688
rect 134852 232672 134904 232678
rect 134852 232614 134904 232620
rect 101732 232468 101784 232474
rect 101732 232410 101784 232416
rect 134850 232232 134906 232241
rect 134850 232167 134906 232176
rect 101270 231960 101326 231969
rect 101270 231895 101326 231904
rect 101284 231726 101312 231895
rect 101272 231720 101324 231726
rect 101272 231662 101324 231668
rect 134758 231688 134814 231697
rect 134758 231623 134814 231632
rect 101454 231552 101510 231561
rect 134772 231522 134800 231623
rect 101454 231487 101510 231496
rect 134760 231516 134812 231522
rect 101468 231114 101496 231487
rect 134760 231458 134812 231464
rect 101730 231280 101786 231289
rect 101730 231215 101786 231224
rect 98880 231108 98932 231114
rect 98880 231050 98932 231056
rect 101456 231108 101508 231114
rect 101456 231050 101508 231056
rect 98892 230910 98920 231050
rect 101744 231046 101772 231215
rect 134758 231144 134814 231153
rect 134758 231079 134760 231088
rect 134812 231079 134814 231088
rect 134760 231050 134812 231056
rect 134864 231046 134892 232167
rect 139636 231516 139688 231522
rect 139636 231458 139688 231464
rect 136876 231108 136928 231114
rect 136876 231050 136928 231056
rect 101732 231040 101784 231046
rect 101732 230982 101784 230988
rect 134852 231040 134904 231046
rect 134852 230982 134904 230988
rect 98880 230904 98932 230910
rect 98880 230846 98932 230852
rect 134390 230600 134446 230609
rect 134390 230535 134446 230544
rect 101730 230192 101786 230201
rect 101730 230127 101786 230136
rect 101546 229784 101602 229793
rect 101546 229719 101602 229728
rect 101560 229550 101588 229719
rect 101744 229618 101772 230127
rect 134298 230056 134354 230065
rect 134298 229991 134300 230000
rect 134352 229991 134354 230000
rect 134300 229962 134352 229968
rect 134404 229686 134432 230535
rect 134392 229680 134444 229686
rect 134392 229622 134444 229628
rect 101732 229612 101784 229618
rect 101732 229554 101784 229560
rect 136888 229550 136916 231050
rect 139648 230638 139676 231458
rect 142224 231289 142252 232682
rect 142304 232672 142356 232678
rect 142304 232614 142356 232620
rect 142316 231969 142344 232614
rect 177724 232400 177776 232406
rect 177724 232342 177776 232348
rect 177736 232241 177764 232342
rect 177722 232232 177778 232241
rect 177722 232167 177778 232176
rect 142302 231960 142358 231969
rect 142302 231895 142358 231904
rect 177724 231720 177776 231726
rect 177724 231662 177776 231668
rect 177736 231561 177764 231662
rect 177722 231552 177778 231561
rect 177722 231487 177778 231496
rect 142210 231280 142266 231289
rect 142210 231215 142266 231224
rect 143684 230904 143736 230910
rect 177724 230904 177776 230910
rect 143684 230846 143736 230852
rect 177722 230872 177724 230881
rect 177776 230872 177778 230881
rect 143696 230745 143724 230846
rect 177722 230807 177778 230816
rect 143682 230736 143738 230745
rect 143682 230671 143738 230680
rect 139636 230632 139688 230638
rect 139636 230574 139688 230580
rect 142948 230632 143000 230638
rect 142948 230574 143000 230580
rect 177724 230632 177776 230638
rect 177724 230574 177776 230580
rect 142960 230201 142988 230574
rect 177736 230473 177764 230574
rect 177722 230464 177778 230473
rect 177722 230399 177778 230408
rect 142946 230192 143002 230201
rect 142946 230127 143002 230136
rect 139636 230020 139688 230026
rect 139636 229962 139688 229968
rect 101548 229544 101600 229550
rect 101548 229486 101600 229492
rect 136876 229544 136928 229550
rect 136876 229486 136928 229492
rect 139648 229482 139676 229962
rect 177722 229648 177778 229657
rect 143592 229612 143644 229618
rect 143592 229554 143644 229560
rect 177632 229612 177684 229618
rect 177722 229583 177778 229592
rect 177632 229554 177684 229560
rect 139636 229476 139688 229482
rect 139636 229418 139688 229424
rect 143500 229476 143552 229482
rect 143500 229418 143552 229424
rect 134390 229376 134446 229385
rect 134390 229311 134446 229320
rect 101730 229240 101786 229249
rect 101730 229175 101786 229184
rect 101744 228938 101772 229175
rect 101732 228932 101784 228938
rect 101732 228874 101784 228880
rect 101454 228696 101510 228705
rect 101454 228631 101510 228640
rect 101468 228394 101496 228631
rect 134404 228462 134432 229311
rect 134758 228832 134814 228841
rect 134758 228767 134814 228776
rect 134392 228456 134444 228462
rect 101730 228424 101786 228433
rect 101456 228388 101508 228394
rect 134392 228398 134444 228404
rect 134772 228394 134800 228767
rect 101730 228359 101786 228368
rect 134760 228388 134812 228394
rect 101456 228330 101508 228336
rect 101744 228326 101772 228359
rect 134760 228330 134812 228336
rect 101732 228320 101784 228326
rect 134852 228320 134904 228326
rect 101732 228262 101784 228268
rect 134850 228288 134852 228297
rect 136876 228320 136928 228326
rect 134904 228288 134906 228297
rect 143512 228297 143540 229418
rect 143604 228977 143632 229554
rect 143684 229544 143736 229550
rect 143682 229512 143684 229521
rect 143736 229512 143738 229521
rect 143682 229447 143738 229456
rect 177644 229249 177672 229554
rect 177736 229550 177764 229583
rect 177724 229544 177776 229550
rect 177724 229486 177776 229492
rect 177630 229240 177686 229249
rect 177630 229175 177686 229184
rect 143590 228968 143646 228977
rect 143590 228903 143646 228912
rect 176988 228932 177040 228938
rect 176988 228874 177040 228880
rect 177000 228569 177028 228874
rect 176986 228560 177042 228569
rect 176986 228495 177042 228504
rect 136876 228262 136928 228268
rect 143498 228288 143554 228297
rect 134850 228223 134906 228232
rect 134758 227744 134814 227753
rect 134758 227679 134814 227688
rect 101362 227472 101418 227481
rect 101362 227407 101418 227416
rect 101376 226830 101404 227407
rect 101454 227064 101510 227073
rect 101454 226999 101510 227008
rect 101364 226824 101416 226830
rect 101364 226766 101416 226772
rect 101468 226762 101496 226999
rect 134772 226898 134800 227679
rect 135402 227200 135458 227209
rect 135458 227158 135536 227186
rect 135402 227135 135458 227144
rect 134760 226892 134812 226898
rect 134760 226834 134812 226840
rect 101456 226756 101508 226762
rect 101456 226698 101508 226704
rect 134390 226520 134446 226529
rect 134390 226455 134446 226464
rect 101638 226384 101694 226393
rect 101638 226319 101694 226328
rect 101546 225568 101602 225577
rect 101546 225503 101602 225512
rect 101560 225470 101588 225503
rect 101548 225464 101600 225470
rect 101548 225406 101600 225412
rect 101652 225334 101680 226319
rect 101822 225704 101878 225713
rect 101822 225639 101878 225648
rect 101836 225402 101864 225639
rect 134404 225606 134432 226455
rect 134758 225976 134814 225985
rect 134758 225911 134814 225920
rect 134392 225600 134444 225606
rect 134392 225542 134444 225548
rect 134772 225538 134800 225911
rect 134760 225532 134812 225538
rect 134760 225474 134812 225480
rect 135508 225470 135536 227158
rect 136888 226762 136916 228262
rect 143498 228223 143554 228232
rect 143684 228252 143736 228258
rect 143684 228194 143736 228200
rect 177724 228252 177776 228258
rect 177724 228194 177776 228200
rect 143316 228184 143368 228190
rect 143316 228126 143368 228132
rect 143328 227209 143356 228126
rect 143696 227753 143724 228194
rect 177632 228184 177684 228190
rect 177632 228126 177684 228132
rect 143682 227744 143738 227753
rect 143682 227679 143738 227688
rect 177644 227481 177672 228126
rect 177736 228025 177764 228194
rect 177722 228016 177778 228025
rect 177722 227951 177778 227960
rect 177630 227472 177686 227481
rect 177630 227407 177686 227416
rect 143314 227200 143370 227209
rect 143314 227135 143370 227144
rect 143316 226824 143368 226830
rect 143316 226766 143368 226772
rect 177172 226824 177224 226830
rect 177172 226766 177224 226772
rect 136876 226756 136928 226762
rect 136876 226698 136928 226704
rect 143328 225985 143356 226766
rect 143684 226756 143736 226762
rect 143684 226698 143736 226704
rect 143696 226529 143724 226698
rect 177184 226665 177212 226766
rect 177724 226756 177776 226762
rect 177724 226698 177776 226704
rect 177170 226656 177226 226665
rect 177170 226591 177226 226600
rect 143682 226520 143738 226529
rect 143682 226455 143738 226464
rect 177736 226257 177764 226698
rect 177722 226248 177778 226257
rect 177722 226183 177778 226192
rect 143314 225976 143370 225985
rect 143314 225911 143370 225920
rect 143316 225600 143368 225606
rect 143316 225542 143368 225548
rect 142580 225532 142632 225538
rect 142580 225474 142632 225480
rect 135496 225464 135548 225470
rect 134666 225432 134722 225441
rect 101824 225396 101876 225402
rect 135496 225406 135548 225412
rect 134666 225367 134722 225376
rect 101824 225338 101876 225344
rect 101640 225328 101692 225334
rect 101640 225270 101692 225276
rect 134298 224888 134354 224897
rect 134298 224823 134354 224832
rect 101086 224616 101142 224625
rect 101086 224551 101142 224560
rect 100994 224480 101050 224489
rect 100994 224415 101050 224424
rect 101008 224110 101036 224415
rect 100996 224104 101048 224110
rect 100996 224046 101048 224052
rect 101100 224042 101128 224551
rect 134312 224178 134340 224823
rect 134680 224314 134708 225367
rect 135402 224344 135458 224353
rect 134668 224308 134720 224314
rect 135402 224279 135458 224288
rect 134668 224250 134720 224256
rect 135416 224246 135444 224279
rect 135404 224240 135456 224246
rect 135404 224182 135456 224188
rect 136876 224240 136928 224246
rect 142592 224217 142620 225474
rect 143328 224761 143356 225542
rect 143684 225464 143736 225470
rect 177724 225464 177776 225470
rect 143684 225406 143736 225412
rect 177722 225432 177724 225441
rect 177776 225432 177778 225441
rect 143696 225305 143724 225406
rect 177172 225396 177224 225402
rect 177722 225367 177778 225376
rect 177172 225338 177224 225344
rect 143682 225296 143738 225305
rect 143682 225231 143738 225240
rect 143314 224752 143370 224761
rect 143314 224687 143370 224696
rect 177184 224489 177212 225338
rect 177724 225328 177776 225334
rect 177724 225270 177776 225276
rect 177736 225033 177764 225270
rect 177722 225024 177778 225033
rect 177722 224959 177778 224968
rect 177170 224480 177226 224489
rect 177170 224415 177226 224424
rect 136876 224182 136928 224188
rect 142578 224208 142634 224217
rect 134300 224172 134352 224178
rect 134300 224114 134352 224120
rect 101088 224036 101140 224042
rect 101088 223978 101140 223984
rect 134760 224036 134812 224042
rect 134760 223978 134812 223984
rect 101454 223528 101510 223537
rect 101454 223463 101510 223472
rect 101362 222984 101418 222993
rect 101362 222919 101418 222928
rect 100902 222848 100958 222857
rect 100902 222783 100958 222792
rect 100916 221186 100944 222783
rect 101376 222682 101404 222919
rect 101468 222750 101496 223463
rect 134482 223120 134538 223129
rect 134482 223055 134484 223064
rect 134536 223055 134538 223064
rect 134484 223026 134536 223032
rect 101456 222744 101508 222750
rect 101456 222686 101508 222692
rect 101364 222676 101416 222682
rect 101364 222618 101416 222624
rect 134666 222032 134722 222041
rect 134666 221967 134722 221976
rect 101638 221896 101694 221905
rect 101638 221831 101694 221840
rect 101546 221488 101602 221497
rect 101546 221423 101602 221432
rect 101560 221322 101588 221423
rect 101548 221316 101600 221322
rect 101548 221258 101600 221264
rect 101652 221254 101680 221831
rect 134680 221458 134708 221967
rect 134668 221452 134720 221458
rect 134668 221394 134720 221400
rect 101640 221248 101692 221254
rect 101640 221190 101692 221196
rect 100904 221180 100956 221186
rect 100904 221122 100956 221128
rect 101822 220672 101878 220681
rect 101822 220607 101878 220616
rect 101270 220128 101326 220137
rect 101270 220063 101326 220072
rect 100902 219992 100958 220001
rect 100902 219927 100958 219936
rect 100916 218534 100944 219927
rect 101284 219894 101312 220063
rect 101836 219962 101864 220607
rect 101824 219956 101876 219962
rect 101824 219898 101876 219904
rect 101272 219888 101324 219894
rect 101272 219830 101324 219836
rect 101362 219040 101418 219049
rect 101362 218975 101418 218984
rect 101376 218602 101404 218975
rect 101730 218904 101786 218913
rect 101730 218839 101786 218848
rect 101744 218670 101772 218839
rect 101732 218664 101784 218670
rect 101732 218606 101784 218612
rect 101364 218596 101416 218602
rect 101364 218538 101416 218544
rect 100904 218528 100956 218534
rect 100904 218470 100956 218476
rect 101178 217952 101234 217961
rect 101178 217887 101234 217896
rect 100810 217408 100866 217417
rect 100810 217343 100866 217352
rect 100718 216048 100774 216057
rect 100718 215983 100774 215992
rect 100732 214386 100760 215983
rect 100824 215746 100852 217343
rect 100902 217272 100958 217281
rect 101192 217242 101220 217887
rect 134482 217408 134538 217417
rect 134482 217343 134484 217352
rect 134536 217343 134538 217352
rect 134484 217314 134536 217320
rect 100902 217207 100958 217216
rect 101180 217236 101232 217242
rect 100812 215740 100864 215746
rect 100812 215682 100864 215688
rect 100916 215678 100944 217207
rect 101180 217178 101232 217184
rect 101362 216184 101418 216193
rect 101362 216119 101418 216128
rect 101376 215814 101404 216119
rect 101364 215808 101416 215814
rect 101364 215750 101416 215756
rect 100904 215672 100956 215678
rect 100904 215614 100956 215620
rect 100994 215096 101050 215105
rect 100994 215031 101050 215040
rect 100810 214688 100866 214697
rect 100810 214623 100866 214632
rect 100720 214380 100772 214386
rect 100720 214322 100772 214328
rect 100718 213464 100774 213473
rect 100718 213399 100774 213408
rect 97500 212000 97552 212006
rect 97500 211942 97552 211948
rect 97512 211530 97540 211942
rect 100732 211598 100760 213399
rect 100824 213026 100852 214623
rect 101008 214454 101036 215031
rect 134772 214454 134800 223978
rect 135402 223664 135458 223673
rect 135402 223599 135458 223608
rect 135416 222818 135444 223599
rect 135404 222812 135456 222818
rect 135404 222754 135456 222760
rect 136888 222682 136916 224182
rect 142578 224143 142634 224152
rect 143684 224104 143736 224110
rect 143684 224046 143736 224052
rect 177724 224104 177776 224110
rect 177724 224046 177776 224052
rect 143316 224036 143368 224042
rect 143316 223978 143368 223984
rect 136968 223084 137020 223090
rect 136968 223026 137020 223032
rect 136876 222676 136928 222682
rect 136876 222618 136928 222624
rect 134850 222576 134906 222585
rect 134850 222511 134906 222520
rect 134864 221730 134892 222511
rect 134852 221724 134904 221730
rect 134852 221666 134904 221672
rect 135402 221488 135458 221497
rect 135402 221423 135458 221432
rect 135416 221390 135444 221423
rect 135404 221384 135456 221390
rect 135404 221326 135456 221332
rect 136876 221384 136928 221390
rect 136876 221326 136928 221332
rect 135402 220808 135458 220817
rect 135402 220743 135458 220752
rect 135310 220264 135366 220273
rect 135310 220199 135366 220208
rect 135324 220166 135352 220199
rect 135312 220160 135364 220166
rect 135312 220102 135364 220108
rect 135416 220030 135444 220743
rect 135404 220024 135456 220030
rect 135404 219966 135456 219972
rect 136888 219894 136916 221326
rect 136980 221322 137008 223026
rect 143328 222993 143356 223978
rect 143696 223537 143724 224046
rect 177632 224036 177684 224042
rect 177632 223978 177684 223984
rect 143682 223528 143738 223537
rect 143682 223463 143738 223472
rect 177644 223265 177672 223978
rect 177736 223809 177764 224046
rect 177722 223800 177778 223809
rect 177722 223735 177778 223744
rect 177630 223256 177686 223265
rect 177630 223191 177686 223200
rect 143314 222984 143370 222993
rect 143314 222919 143370 222928
rect 143316 222744 143368 222750
rect 143316 222686 143368 222692
rect 177632 222744 177684 222750
rect 177632 222686 177684 222692
rect 143328 221769 143356 222686
rect 143684 222676 143736 222682
rect 143684 222618 143736 222624
rect 143696 222313 143724 222618
rect 143682 222304 143738 222313
rect 143682 222239 143738 222248
rect 177644 222041 177672 222686
rect 177724 222676 177776 222682
rect 177724 222618 177776 222624
rect 177736 222449 177764 222618
rect 177722 222440 177778 222449
rect 177722 222375 177778 222384
rect 177630 222032 177686 222041
rect 177630 221967 177686 221976
rect 143314 221760 143370 221769
rect 139636 221724 139688 221730
rect 143314 221695 143370 221704
rect 139636 221666 139688 221672
rect 136968 221316 137020 221322
rect 136968 221258 137020 221264
rect 139648 220982 139676 221666
rect 139728 221452 139780 221458
rect 139728 221394 139780 221400
rect 139636 220976 139688 220982
rect 139636 220918 139688 220924
rect 139740 220642 139768 221394
rect 143684 221316 143736 221322
rect 143684 221258 143736 221264
rect 177172 221316 177224 221322
rect 177172 221258 177224 221264
rect 143696 221225 143724 221258
rect 143682 221216 143738 221225
rect 143682 221151 143738 221160
rect 143316 220976 143368 220982
rect 143316 220918 143368 220924
rect 139728 220636 139780 220642
rect 139728 220578 139780 220584
rect 143328 220545 143356 220918
rect 143684 220636 143736 220642
rect 143684 220578 143736 220584
rect 143314 220536 143370 220545
rect 143314 220471 143370 220480
rect 138164 220160 138216 220166
rect 138164 220102 138216 220108
rect 136876 219888 136928 219894
rect 136876 219830 136928 219836
rect 135402 219720 135458 219729
rect 135402 219655 135458 219664
rect 135034 219176 135090 219185
rect 135034 219111 135090 219120
rect 135048 218874 135076 219111
rect 135036 218868 135088 218874
rect 135036 218810 135088 218816
rect 135416 218738 135444 219655
rect 137520 218868 137572 218874
rect 137520 218810 137572 218816
rect 135404 218732 135456 218738
rect 135404 218674 135456 218680
rect 135312 218664 135364 218670
rect 135310 218632 135312 218641
rect 135364 218632 135366 218641
rect 135310 218567 135366 218576
rect 135402 217952 135458 217961
rect 135402 217887 135458 217896
rect 135416 217310 135444 217887
rect 135404 217304 135456 217310
rect 135404 217246 135456 217252
rect 137532 217174 137560 218810
rect 137980 218664 138032 218670
rect 137980 218606 138032 218612
rect 137612 217372 137664 217378
rect 137612 217314 137664 217320
rect 137520 217168 137572 217174
rect 137520 217110 137572 217116
rect 135402 216864 135458 216873
rect 135402 216799 135458 216808
rect 135416 215882 135444 216799
rect 135494 216320 135550 216329
rect 135494 216255 135550 216264
rect 135404 215876 135456 215882
rect 135404 215818 135456 215824
rect 135402 215776 135458 215785
rect 135402 215711 135458 215720
rect 134850 215096 134906 215105
rect 134850 215031 134906 215040
rect 134864 214930 134892 215031
rect 134852 214924 134904 214930
rect 134852 214866 134904 214872
rect 135312 214584 135364 214590
rect 135310 214552 135312 214561
rect 135364 214552 135366 214561
rect 135416 214522 135444 215711
rect 135310 214487 135366 214496
rect 135404 214516 135456 214522
rect 135404 214458 135456 214464
rect 135508 214454 135536 216255
rect 137624 215678 137652 217314
rect 137704 217304 137756 217310
rect 137704 217246 137756 217252
rect 137716 215746 137744 217246
rect 137992 217106 138020 218606
rect 138176 218534 138204 220102
rect 143696 220001 143724 220578
rect 177184 220273 177212 221258
rect 177632 221248 177684 221254
rect 177632 221190 177684 221196
rect 177644 220953 177672 221190
rect 177724 221180 177776 221186
rect 177724 221122 177776 221128
rect 177736 221089 177764 221122
rect 177722 221080 177778 221089
rect 177722 221015 177778 221024
rect 177630 220944 177686 220953
rect 177630 220879 177686 220888
rect 177170 220264 177226 220273
rect 177170 220199 177226 220208
rect 143682 219992 143738 220001
rect 143132 219956 143184 219962
rect 143682 219927 143738 219936
rect 177172 219956 177224 219962
rect 143132 219898 143184 219904
rect 177172 219898 177224 219904
rect 143144 218777 143172 219898
rect 143684 219888 143736 219894
rect 143684 219830 143736 219836
rect 143696 219321 143724 219830
rect 143682 219312 143738 219321
rect 143682 219247 143738 219256
rect 177184 219049 177212 219898
rect 177724 219888 177776 219894
rect 177724 219830 177776 219836
rect 177736 219593 177764 219830
rect 177722 219584 177778 219593
rect 177722 219519 177778 219528
rect 177170 219040 177226 219049
rect 177170 218975 177226 218984
rect 143130 218768 143186 218777
rect 143130 218703 143186 218712
rect 178000 218664 178052 218670
rect 178000 218606 178052 218612
rect 143500 218596 143552 218602
rect 143500 218538 143552 218544
rect 177172 218596 177224 218602
rect 177172 218538 177224 218544
rect 138164 218528 138216 218534
rect 138164 218470 138216 218476
rect 143512 217553 143540 218538
rect 143684 218528 143736 218534
rect 143684 218470 143736 218476
rect 143696 218233 143724 218470
rect 143682 218224 143738 218233
rect 143682 218159 143738 218168
rect 177184 217961 177212 218538
rect 177724 218528 177776 218534
rect 177724 218470 177776 218476
rect 177736 218369 177764 218470
rect 177722 218360 177778 218369
rect 177722 218295 177778 218304
rect 177170 217952 177226 217961
rect 177170 217887 177226 217896
rect 143498 217544 143554 217553
rect 143498 217479 143554 217488
rect 143684 217168 143736 217174
rect 143684 217110 143736 217116
rect 177724 217168 177776 217174
rect 178012 217145 178040 218606
rect 177724 217110 177776 217116
rect 177998 217136 178054 217145
rect 137980 217100 138032 217106
rect 137980 217042 138032 217048
rect 143132 217100 143184 217106
rect 143132 217042 143184 217048
rect 143144 216329 143172 217042
rect 143696 217009 143724 217110
rect 143682 217000 143738 217009
rect 143682 216935 143738 216944
rect 177736 216737 177764 217110
rect 177998 217071 178054 217080
rect 177722 216728 177778 216737
rect 177722 216663 177778 216672
rect 143130 216320 143186 216329
rect 143130 216255 143186 216264
rect 143500 215808 143552 215814
rect 143130 215776 143186 215785
rect 137704 215740 137756 215746
rect 143500 215750 143552 215756
rect 177172 215808 177224 215814
rect 177172 215750 177224 215756
rect 143130 215711 143132 215720
rect 137704 215682 137756 215688
rect 143184 215711 143186 215720
rect 143132 215682 143184 215688
rect 137612 215672 137664 215678
rect 137612 215614 137664 215620
rect 142948 215672 143000 215678
rect 142948 215614 143000 215620
rect 142960 215241 142988 215614
rect 142946 215232 143002 215241
rect 142946 215167 143002 215176
rect 137612 214924 137664 214930
rect 137612 214866 137664 214872
rect 136876 214584 136928 214590
rect 136876 214526 136928 214532
rect 100996 214448 101048 214454
rect 100996 214390 101048 214396
rect 134760 214448 134812 214454
rect 134760 214390 134812 214396
rect 135312 214448 135364 214454
rect 135312 214390 135364 214396
rect 135496 214448 135548 214454
rect 135496 214390 135548 214396
rect 100994 214008 101050 214017
rect 100994 213943 101050 213952
rect 134482 214008 134538 214017
rect 134482 213943 134538 213952
rect 100902 213192 100958 213201
rect 100902 213127 100958 213136
rect 100812 213020 100864 213026
rect 100812 212962 100864 212968
rect 100916 211666 100944 213127
rect 101008 213094 101036 213943
rect 134496 213570 134524 213943
rect 134484 213564 134536 213570
rect 134484 213506 134536 213512
rect 134482 213464 134538 213473
rect 134482 213399 134538 213408
rect 134496 213162 134524 213399
rect 134484 213156 134536 213162
rect 134484 213098 134536 213104
rect 100996 213088 101048 213094
rect 100996 213030 101048 213036
rect 134482 212920 134538 212929
rect 134482 212855 134538 212864
rect 100994 212376 101050 212385
rect 100994 212311 101050 212320
rect 101008 212006 101036 212311
rect 100996 212000 101048 212006
rect 100996 211942 101048 211948
rect 101270 211968 101326 211977
rect 134496 211938 134524 212855
rect 134666 212240 134722 212249
rect 134666 212175 134722 212184
rect 101270 211903 101326 211912
rect 134484 211932 134536 211938
rect 100904 211660 100956 211666
rect 100904 211602 100956 211608
rect 100720 211592 100772 211598
rect 100720 211534 100772 211540
rect 97500 211524 97552 211530
rect 97500 211466 97552 211472
rect 101178 211152 101234 211161
rect 101178 211087 101234 211096
rect 101086 210744 101142 210753
rect 101086 210679 101142 210688
rect 100994 210472 101050 210481
rect 101100 210442 101128 210679
rect 100994 210407 101050 210416
rect 101088 210436 101140 210442
rect 101008 210374 101036 210407
rect 101088 210378 101140 210384
rect 100996 210368 101048 210374
rect 100996 210310 101048 210316
rect 101192 210238 101220 211087
rect 101284 210306 101312 211903
rect 134484 211874 134536 211880
rect 134680 211802 134708 212175
rect 134668 211796 134720 211802
rect 134668 211738 134720 211744
rect 134574 211696 134630 211705
rect 134574 211631 134630 211640
rect 134588 210374 134616 211631
rect 135034 211152 135090 211161
rect 135034 211087 135090 211096
rect 134850 210608 134906 210617
rect 134850 210543 134906 210552
rect 134576 210368 134628 210374
rect 134576 210310 134628 210316
rect 101272 210300 101324 210306
rect 101272 210242 101324 210248
rect 101180 210232 101232 210238
rect 101180 210174 101232 210180
rect 100994 209520 101050 209529
rect 100994 209455 101050 209464
rect 101008 209014 101036 209455
rect 100996 209008 101048 209014
rect 100996 208950 101048 208956
rect 101638 208976 101694 208985
rect 101638 208911 101694 208920
rect 100994 206528 101050 206537
rect 100994 206463 101050 206472
rect 101008 206226 101036 206463
rect 100996 206220 101048 206226
rect 100996 206162 101048 206168
rect 98972 204452 99024 204458
rect 98972 204394 99024 204400
rect 98880 203500 98932 203506
rect 98880 203442 98932 203448
rect 98892 185321 98920 203442
rect 98984 186545 99012 204394
rect 99432 204316 99484 204322
rect 99432 204258 99484 204264
rect 99248 204180 99300 204186
rect 99248 204122 99300 204128
rect 99156 203840 99208 203846
rect 99156 203782 99208 203788
rect 99064 203568 99116 203574
rect 99064 203510 99116 203516
rect 99076 187769 99104 203510
rect 99168 189537 99196 203782
rect 99260 190761 99288 204122
rect 99340 203636 99392 203642
rect 99340 203578 99392 203584
rect 99246 190752 99302 190761
rect 99246 190687 99302 190696
rect 99154 189528 99210 189537
rect 99154 189463 99210 189472
rect 99352 188993 99380 203578
rect 99444 192393 99472 204258
rect 99524 204112 99576 204118
rect 99524 204054 99576 204060
rect 99536 193753 99564 204054
rect 101652 196094 101680 208911
rect 101730 208432 101786 208441
rect 101730 208367 101786 208376
rect 101640 196088 101692 196094
rect 101640 196030 101692 196036
rect 101744 196026 101772 208367
rect 102098 207888 102154 207897
rect 102098 207823 102154 207832
rect 101914 207616 101970 207625
rect 101914 207551 101970 207560
rect 101732 196020 101784 196026
rect 101732 195962 101784 195968
rect 101928 195890 101956 207551
rect 102112 195958 102140 207823
rect 134206 207752 134262 207761
rect 134206 207687 134208 207696
rect 134260 207687 134262 207696
rect 134208 207658 134260 207664
rect 104228 203506 104256 206908
rect 104780 204458 104808 206908
rect 104768 204452 104820 204458
rect 104768 204394 104820 204400
rect 105332 203574 105360 206908
rect 105884 203642 105912 206908
rect 106436 203846 106464 206908
rect 106988 204186 107016 206908
rect 107540 204322 107568 206908
rect 107528 204316 107580 204322
rect 107528 204258 107580 204264
rect 106976 204180 107028 204186
rect 106976 204122 107028 204128
rect 108092 204118 108120 206908
rect 108080 204112 108132 204118
rect 108080 204054 108132 204060
rect 106424 203840 106476 203846
rect 106424 203782 106476 203788
rect 105872 203636 105924 203642
rect 105872 203578 105924 203584
rect 105320 203568 105372 203574
rect 105320 203510 105372 203516
rect 104216 203500 104268 203506
rect 104216 203442 104268 203448
rect 108644 203438 108672 206908
rect 109196 203522 109224 206908
rect 109276 203568 109328 203574
rect 109196 203516 109276 203522
rect 109196 203510 109328 203516
rect 109196 203494 109316 203510
rect 109748 203438 109776 206908
rect 110300 203710 110328 206908
rect 110288 203704 110340 203710
rect 110288 203646 110340 203652
rect 110288 203568 110340 203574
rect 110288 203510 110340 203516
rect 108632 203432 108684 203438
rect 108632 203374 108684 203380
rect 109276 203432 109328 203438
rect 109276 203374 109328 203380
rect 109736 203432 109788 203438
rect 109736 203374 109788 203380
rect 102100 195952 102152 195958
rect 102100 195894 102152 195900
rect 101916 195884 101968 195890
rect 101916 195826 101968 195832
rect 109288 193866 109316 203374
rect 109288 193838 109868 193866
rect 99522 193744 99578 193753
rect 109840 193730 109868 193838
rect 110300 193730 110328 203510
rect 110748 203432 110800 203438
rect 110748 203374 110800 203380
rect 110760 196314 110788 203374
rect 110852 196502 110880 206908
rect 111024 203704 111076 203710
rect 111024 203646 111076 203652
rect 110840 196496 110892 196502
rect 110840 196438 110892 196444
rect 110760 196286 110880 196314
rect 109840 193702 110130 193730
rect 110300 193702 110498 193730
rect 110852 193716 110880 196286
rect 111036 193730 111064 203646
rect 111496 203438 111524 206908
rect 111484 203432 111536 203438
rect 111484 203374 111536 203380
rect 112048 196502 112076 206908
rect 112312 203432 112364 203438
rect 112312 203374 112364 203380
rect 111668 196496 111720 196502
rect 111668 196438 111720 196444
rect 112036 196496 112088 196502
rect 112036 196438 112088 196444
rect 111036 193702 111326 193730
rect 111680 193716 111708 196438
rect 112324 193730 112352 203374
rect 112496 196496 112548 196502
rect 112496 196438 112548 196444
rect 112062 193702 112352 193730
rect 112508 193716 112536 196438
rect 112600 193730 112628 206908
rect 113152 193730 113180 206908
rect 112600 193702 112890 193730
rect 113152 193702 113258 193730
rect 113704 193716 113732 206908
rect 114256 193730 114284 206908
rect 114808 203438 114836 206908
rect 114612 203432 114664 203438
rect 114612 203374 114664 203380
rect 114796 203432 114848 203438
rect 114796 203374 114848 203380
rect 114624 193730 114652 203374
rect 115360 196502 115388 206908
rect 114888 196496 114940 196502
rect 114888 196438 114940 196444
rect 115348 196496 115400 196502
rect 115348 196438 115400 196444
rect 114086 193702 114284 193730
rect 114454 193702 114652 193730
rect 114900 193716 114928 196438
rect 115912 196434 115940 206908
rect 116360 203568 116412 203574
rect 116360 203510 116412 203516
rect 116084 203500 116136 203506
rect 116084 203442 116136 203448
rect 115992 203432 116044 203438
rect 115992 203374 116044 203380
rect 115256 196428 115308 196434
rect 115256 196370 115308 196376
rect 115900 196428 115952 196434
rect 115900 196370 115952 196376
rect 115268 193716 115296 196370
rect 116004 193730 116032 203374
rect 115650 193702 116032 193730
rect 116096 193716 116124 203442
rect 116372 199986 116400 203510
rect 116464 203438 116492 206908
rect 117016 203506 117044 206908
rect 117464 203840 117516 203846
rect 117464 203782 117516 203788
rect 117004 203500 117056 203506
rect 117004 203442 117056 203448
rect 116452 203432 116504 203438
rect 116452 203374 116504 203380
rect 117372 203432 117424 203438
rect 117372 203374 117424 203380
rect 116372 199958 116492 199986
rect 116464 193716 116492 199958
rect 117384 194002 117412 203374
rect 117016 193974 117412 194002
rect 117016 193730 117044 193974
rect 117476 193730 117504 203782
rect 117568 203574 117596 206908
rect 117556 203568 117608 203574
rect 117556 203510 117608 203516
rect 117648 203500 117700 203506
rect 117648 203442 117700 203448
rect 116846 193702 117044 193730
rect 117306 193702 117504 193730
rect 117660 193716 117688 203442
rect 118212 203438 118240 206908
rect 118764 203846 118792 206908
rect 118752 203840 118804 203846
rect 118752 203782 118804 203788
rect 118752 203704 118804 203710
rect 118752 203646 118804 203652
rect 118660 203500 118712 203506
rect 118660 203442 118712 203448
rect 118200 203432 118252 203438
rect 118200 203374 118252 203380
rect 118672 194274 118700 203442
rect 118304 194246 118700 194274
rect 118304 193730 118332 194246
rect 118660 194184 118712 194190
rect 118660 194126 118712 194132
rect 118672 193730 118700 194126
rect 118134 193702 118332 193730
rect 118502 193702 118700 193730
rect 118764 193730 118792 203646
rect 118844 203568 118896 203574
rect 118844 203510 118896 203516
rect 118856 194190 118884 203510
rect 119316 203438 119344 206908
rect 119868 203506 119896 206908
rect 120132 204384 120184 204390
rect 120132 204326 120184 204332
rect 119856 203500 119908 203506
rect 119856 203442 119908 203448
rect 120040 203500 120092 203506
rect 120040 203442 120092 203448
rect 119304 203432 119356 203438
rect 119304 203374 119356 203380
rect 120052 196366 120080 203442
rect 119672 196360 119724 196366
rect 119672 196302 119724 196308
rect 120040 196360 120092 196366
rect 120040 196302 120092 196308
rect 119304 195476 119356 195482
rect 119304 195418 119356 195424
rect 118844 194184 118896 194190
rect 118844 194126 118896 194132
rect 118764 193702 118870 193730
rect 119316 193716 119344 195418
rect 119684 193716 119712 196302
rect 120144 195482 120172 204326
rect 120420 203574 120448 206908
rect 120972 203710 121000 206908
rect 121420 204588 121472 204594
rect 121420 204530 121472 204536
rect 120960 203704 121012 203710
rect 120960 203646 121012 203652
rect 120408 203568 120460 203574
rect 120408 203510 120460 203516
rect 120224 203432 120276 203438
rect 120224 203374 120276 203380
rect 120132 195476 120184 195482
rect 120132 195418 120184 195424
rect 120236 193730 120264 203374
rect 120868 196428 120920 196434
rect 120868 196370 120920 196376
rect 120500 196360 120552 196366
rect 120500 196302 120552 196308
rect 120066 193702 120264 193730
rect 120512 193716 120540 196302
rect 120880 193716 120908 196370
rect 121432 196366 121460 204530
rect 121524 204390 121552 206908
rect 121604 204452 121656 204458
rect 121604 204394 121656 204400
rect 121512 204384 121564 204390
rect 121512 204326 121564 204332
rect 121512 204248 121564 204254
rect 121512 204190 121564 204196
rect 121420 196360 121472 196366
rect 121420 196302 121472 196308
rect 121524 193730 121552 204190
rect 121616 196434 121644 204394
rect 122076 203506 122104 206908
rect 122064 203500 122116 203506
rect 122064 203442 122116 203448
rect 122628 203438 122656 206908
rect 123180 204594 123208 206908
rect 123168 204588 123220 204594
rect 123168 204530 123220 204536
rect 123732 204458 123760 206908
rect 123720 204452 123772 204458
rect 123720 204394 123772 204400
rect 124284 204254 124312 206908
rect 124272 204248 124324 204254
rect 124272 204190 124324 204196
rect 124272 203840 124324 203846
rect 124272 203782 124324 203788
rect 123720 203772 123772 203778
rect 123720 203714 123772 203720
rect 122616 203432 122668 203438
rect 122616 203374 122668 203380
rect 123628 196496 123680 196502
rect 123628 196438 123680 196444
rect 121604 196428 121656 196434
rect 121604 196370 121656 196376
rect 121696 196428 121748 196434
rect 121696 196370 121748 196376
rect 121262 193702 121552 193730
rect 121708 193716 121736 196370
rect 123260 196360 123312 196366
rect 123260 196302 123312 196308
rect 122432 196292 122484 196298
rect 122432 196234 122484 196240
rect 122064 195884 122116 195890
rect 122064 195826 122116 195832
rect 122076 193716 122104 195826
rect 122444 193716 122472 196234
rect 122892 195748 122944 195754
rect 122892 195690 122944 195696
rect 122904 193716 122932 195690
rect 123272 193716 123300 196302
rect 123640 193716 123668 196438
rect 123732 195890 123760 203714
rect 123904 203704 123956 203710
rect 123904 203646 123956 203652
rect 123812 203500 123864 203506
rect 123812 203442 123864 203448
rect 123824 196434 123852 203442
rect 123812 196428 123864 196434
rect 123812 196370 123864 196376
rect 123720 195884 123772 195890
rect 123720 195826 123772 195832
rect 123916 195754 123944 203646
rect 124180 203636 124232 203642
rect 124180 203578 124232 203584
rect 123996 203568 124048 203574
rect 123996 203510 124048 203516
rect 124008 196298 124036 203510
rect 124192 196366 124220 203578
rect 124180 196360 124232 196366
rect 124180 196302 124232 196308
rect 123996 196292 124048 196298
rect 123996 196234 124048 196240
rect 123904 195748 123956 195754
rect 123904 195690 123956 195696
rect 124284 193730 124312 203782
rect 124836 203506 124864 206908
rect 125480 203778 125508 206908
rect 125468 203772 125520 203778
rect 125468 203714 125520 203720
rect 126032 203574 126060 206908
rect 126584 203710 126612 206908
rect 126572 203704 126624 203710
rect 126572 203646 126624 203652
rect 127136 203642 127164 206908
rect 127124 203636 127176 203642
rect 127124 203578 127176 203584
rect 126020 203568 126072 203574
rect 126020 203510 126072 203516
rect 124824 203500 124876 203506
rect 124824 203442 124876 203448
rect 127688 203438 127716 206908
rect 128240 203846 128268 206908
rect 128228 203840 128280 203846
rect 128228 203782 128280 203788
rect 127952 203636 128004 203642
rect 127952 203578 128004 203584
rect 127860 203568 127912 203574
rect 127860 203510 127912 203516
rect 124364 203432 124416 203438
rect 124364 203374 124416 203380
rect 127676 203432 127728 203438
rect 127676 203374 127728 203380
rect 124376 196502 124404 203374
rect 124364 196496 124416 196502
rect 124364 196438 124416 196444
rect 127872 196026 127900 203510
rect 124456 196020 124508 196026
rect 124456 195962 124508 195968
rect 127860 196020 127912 196026
rect 127860 195962 127912 195968
rect 124114 193702 124312 193730
rect 124468 193716 124496 195962
rect 127964 195822 127992 203578
rect 128792 203574 128820 206908
rect 128780 203568 128832 203574
rect 128780 203510 128832 203516
rect 128136 203500 128188 203506
rect 128136 203442 128188 203448
rect 128044 203432 128096 203438
rect 128044 203374 128096 203380
rect 125652 195816 125704 195822
rect 125652 195758 125704 195764
rect 127952 195816 128004 195822
rect 127952 195758 128004 195764
rect 125284 195680 125336 195686
rect 125284 195622 125336 195628
rect 124824 195612 124876 195618
rect 124824 195554 124876 195560
rect 124836 193716 124864 195554
rect 125296 193716 125324 195622
rect 125664 193716 125692 195758
rect 128056 195618 128084 203374
rect 128148 195686 128176 203442
rect 129344 203438 129372 206908
rect 129896 203506 129924 206908
rect 130448 203642 130476 206908
rect 130436 203636 130488 203642
rect 130436 203578 130488 203584
rect 129884 203500 129936 203506
rect 129884 203442 129936 203448
rect 129332 203432 129384 203438
rect 129332 203374 129384 203380
rect 134864 195822 134892 210543
rect 134942 209384 134998 209393
rect 134942 209319 134998 209328
rect 134956 196026 134984 209319
rect 134944 196020 134996 196026
rect 134944 195962 134996 195968
rect 135048 195890 135076 211087
rect 135126 210064 135182 210073
rect 135126 209999 135182 210008
rect 135140 195958 135168 209999
rect 135218 208296 135274 208305
rect 135218 208231 135274 208240
rect 135232 196094 135260 208231
rect 135324 207518 135352 214390
rect 136888 213026 136916 214526
rect 137060 213564 137112 213570
rect 137060 213506 137112 213512
rect 136968 213156 137020 213162
rect 136968 213098 137020 213104
rect 136876 213020 136928 213026
rect 136876 212962 136928 212968
rect 136876 211796 136928 211802
rect 136876 211738 136928 211744
rect 136888 210238 136916 211738
rect 136980 211394 137008 213098
rect 137072 211666 137100 213506
rect 137624 213094 137652 214866
rect 143512 214561 143540 215750
rect 177184 214969 177212 215750
rect 177724 215740 177776 215746
rect 177724 215682 177776 215688
rect 177632 215672 177684 215678
rect 177736 215649 177764 215682
rect 177632 215614 177684 215620
rect 177722 215640 177778 215649
rect 177644 215513 177672 215614
rect 177722 215575 177778 215584
rect 177630 215504 177686 215513
rect 177630 215439 177686 215448
rect 177170 214960 177226 214969
rect 177170 214895 177226 214904
rect 143498 214552 143554 214561
rect 143498 214487 143554 214496
rect 143684 214516 143736 214522
rect 143684 214458 143736 214464
rect 142948 214448 143000 214454
rect 142948 214390 143000 214396
rect 142960 214017 142988 214390
rect 142946 214008 143002 214017
rect 142946 213943 143002 213952
rect 143696 213337 143724 214458
rect 177632 214448 177684 214454
rect 177632 214390 177684 214396
rect 177644 213745 177672 214390
rect 177724 214380 177776 214386
rect 177724 214322 177776 214328
rect 177736 214153 177764 214322
rect 177722 214144 177778 214153
rect 177722 214079 177778 214088
rect 177630 213736 177686 213745
rect 177630 213671 177686 213680
rect 143682 213328 143738 213337
rect 143682 213263 143738 213272
rect 137612 213088 137664 213094
rect 137612 213030 137664 213036
rect 143684 213088 143736 213094
rect 143684 213030 143736 213036
rect 177172 213088 177224 213094
rect 177172 213030 177224 213036
rect 143500 213020 143552 213026
rect 143500 212962 143552 212968
rect 143512 212249 143540 212962
rect 143696 212793 143724 213030
rect 143682 212784 143738 212793
rect 143682 212719 143738 212728
rect 177184 212521 177212 213030
rect 177724 213020 177776 213026
rect 177724 212962 177776 212968
rect 177736 212929 177764 212962
rect 177722 212920 177778 212929
rect 177722 212855 177778 212864
rect 177170 212512 177226 212521
rect 177170 212447 177226 212456
rect 143498 212240 143554 212249
rect 143498 212175 143554 212184
rect 139636 211932 139688 211938
rect 139636 211874 139688 211880
rect 137060 211660 137112 211666
rect 137060 211602 137112 211608
rect 136968 211388 137020 211394
rect 136968 211330 137020 211336
rect 139648 210986 139676 211874
rect 177722 211696 177778 211705
rect 143684 211660 143736 211666
rect 177722 211631 177724 211640
rect 143684 211602 143736 211608
rect 177776 211631 177778 211640
rect 177724 211602 177776 211608
rect 143696 211569 143724 211602
rect 177172 211592 177224 211598
rect 143682 211560 143738 211569
rect 177172 211534 177224 211540
rect 143682 211495 143738 211504
rect 143684 211388 143736 211394
rect 143684 211330 143736 211336
rect 143696 211025 143724 211330
rect 177184 211297 177212 211534
rect 177170 211288 177226 211297
rect 177170 211223 177226 211232
rect 143682 211016 143738 211025
rect 139636 210980 139688 210986
rect 139636 210922 139688 210928
rect 143592 210980 143644 210986
rect 143682 210951 143738 210960
rect 143592 210922 143644 210928
rect 143604 210345 143632 210922
rect 177724 210844 177776 210850
rect 177724 210786 177776 210792
rect 177736 210617 177764 210786
rect 177722 210608 177778 210617
rect 177722 210543 177778 210552
rect 178184 210436 178236 210442
rect 178184 210378 178236 210384
rect 176804 210368 176856 210374
rect 143590 210336 143646 210345
rect 176804 210310 176856 210316
rect 143590 210271 143646 210280
rect 143684 210300 143736 210306
rect 143684 210242 143736 210248
rect 136876 210232 136928 210238
rect 136876 210174 136928 210180
rect 142948 210232 143000 210238
rect 142948 210174 143000 210180
rect 142960 209801 142988 210174
rect 142946 209792 143002 209801
rect 142946 209727 143002 209736
rect 143696 209257 143724 210242
rect 143682 209248 143738 209257
rect 143682 209183 143738 209192
rect 175424 209008 175476 209014
rect 172294 208976 172350 208985
rect 145352 208934 145596 208962
rect 146976 208934 147312 208962
rect 148448 208934 148784 208962
rect 135402 208840 135458 208849
rect 135402 208775 135458 208784
rect 135312 207512 135364 207518
rect 135312 207454 135364 207460
rect 135310 207208 135366 207217
rect 135310 207143 135366 207152
rect 135324 196434 135352 207143
rect 135312 196428 135364 196434
rect 135312 196370 135364 196376
rect 135416 196162 135444 208775
rect 140280 207716 140332 207722
rect 140280 207658 140332 207664
rect 140292 196366 140320 207658
rect 145352 207518 145380 208934
rect 145340 207512 145392 207518
rect 145340 207454 145392 207460
rect 147284 206226 147312 208934
rect 147272 206220 147324 206226
rect 147272 206162 147324 206168
rect 147824 206220 147876 206226
rect 147824 206162 147876 206168
rect 140464 196428 140516 196434
rect 140464 196370 140516 196376
rect 140280 196360 140332 196366
rect 140280 196302 140332 196308
rect 135404 196156 135456 196162
rect 135404 196098 135456 196104
rect 135220 196088 135272 196094
rect 135220 196030 135272 196036
rect 135128 195952 135180 195958
rect 135128 195894 135180 195900
rect 135036 195884 135088 195890
rect 135036 195826 135088 195832
rect 134852 195816 134904 195822
rect 134852 195758 134904 195764
rect 128136 195680 128188 195686
rect 128136 195622 128188 195628
rect 128044 195612 128096 195618
rect 128044 195554 128096 195560
rect 140476 193716 140504 196370
rect 141568 196360 141620 196366
rect 141568 196302 141620 196308
rect 141580 193716 141608 196302
rect 143776 196156 143828 196162
rect 143776 196098 143828 196104
rect 142672 196088 142724 196094
rect 142672 196030 142724 196036
rect 142684 193716 142712 196030
rect 143788 193716 143816 196098
rect 144880 196020 144932 196026
rect 144880 195962 144932 195968
rect 144892 193716 144920 195962
rect 145984 195952 146036 195958
rect 145984 195894 146036 195900
rect 145996 193716 146024 195894
rect 147836 195822 147864 206162
rect 148756 204798 148784 208934
rect 149308 208934 149828 208962
rect 150688 208934 151300 208962
rect 152068 208934 152680 208962
rect 153448 208934 154152 208962
rect 154828 208934 155532 208962
rect 156208 208934 157004 208962
rect 158048 208934 158384 208962
rect 159520 208934 159856 208962
rect 160900 208934 161236 208962
rect 162464 208934 162708 208962
rect 163752 208934 164088 208962
rect 164488 208934 165560 208962
rect 165868 208934 166940 208962
rect 167248 208934 168412 208962
rect 168628 208934 169792 208962
rect 170008 208934 171264 208962
rect 148744 204792 148796 204798
rect 148744 204734 148796 204740
rect 148192 195884 148244 195890
rect 148192 195826 148244 195832
rect 147088 195816 147140 195822
rect 147088 195758 147140 195764
rect 147824 195816 147876 195822
rect 147824 195758 147876 195764
rect 147100 193716 147128 195758
rect 148204 193716 148232 195826
rect 149308 193716 149336 208934
rect 150688 195226 150716 208934
rect 152068 195226 152096 208934
rect 153448 196366 153476 208934
rect 154828 196366 154856 208934
rect 152608 196360 152660 196366
rect 152608 196302 152660 196308
rect 153436 196360 153488 196366
rect 153436 196302 153488 196308
rect 153804 196360 153856 196366
rect 153804 196302 153856 196308
rect 154816 196360 154868 196366
rect 154816 196302 154868 196308
rect 156012 196360 156064 196366
rect 156012 196302 156064 196308
rect 150596 195198 150716 195226
rect 151976 195198 152096 195226
rect 150596 193730 150624 195198
rect 151976 193730 152004 195198
rect 150426 193702 150624 193730
rect 151530 193702 152004 193730
rect 152620 193716 152648 196302
rect 153816 193716 153844 196302
rect 154908 196156 154960 196162
rect 154908 196098 154960 196104
rect 154920 193716 154948 196098
rect 156024 193716 156052 196302
rect 156208 196162 156236 208934
rect 157484 206288 157536 206294
rect 157484 206230 157536 206236
rect 156840 206220 156892 206226
rect 156840 206162 156892 206168
rect 156852 196366 156880 206162
rect 156840 196360 156892 196366
rect 156840 196302 156892 196308
rect 156196 196156 156248 196162
rect 156196 196098 156248 196104
rect 157496 193730 157524 206230
rect 158048 206226 158076 208934
rect 159520 206294 159548 208934
rect 159508 206288 159560 206294
rect 159508 206230 159560 206236
rect 160900 206226 160928 208934
rect 162464 206294 162492 208934
rect 160980 206288 161032 206294
rect 160980 206230 161032 206236
rect 162452 206288 162504 206294
rect 162452 206230 162504 206236
rect 158036 206220 158088 206226
rect 158036 206162 158088 206168
rect 158864 206220 158916 206226
rect 158864 206162 158916 206168
rect 160888 206220 160940 206226
rect 160888 206162 160940 206168
rect 158876 193866 158904 206162
rect 160428 196156 160480 196162
rect 160428 196098 160480 196104
rect 159324 195340 159376 195346
rect 159324 195282 159376 195288
rect 158508 193838 158904 193866
rect 158508 193730 158536 193838
rect 157142 193702 157524 193730
rect 158246 193702 158536 193730
rect 159336 193716 159364 195282
rect 160440 193716 160468 196098
rect 160992 195346 161020 206230
rect 163752 206226 163780 208934
rect 162360 206220 162412 206226
rect 162360 206162 162412 206168
rect 163740 206220 163792 206226
rect 163740 206162 163792 206168
rect 162372 196162 162400 206162
rect 162636 196360 162688 196366
rect 162636 196302 162688 196308
rect 162360 196156 162412 196162
rect 162360 196098 162412 196104
rect 161532 196020 161584 196026
rect 161532 195962 161584 195968
rect 160980 195340 161032 195346
rect 160980 195282 161032 195288
rect 161544 193716 161572 195962
rect 162648 193716 162676 196302
rect 164488 196026 164516 208934
rect 165868 196366 165896 208934
rect 165856 196360 165908 196366
rect 165856 196302 165908 196308
rect 165948 196360 166000 196366
rect 165948 196302 166000 196308
rect 164476 196020 164528 196026
rect 164476 195962 164528 195968
rect 164844 196020 164896 196026
rect 164844 195962 164896 195968
rect 163740 195884 163792 195890
rect 163740 195826 163792 195832
rect 163752 193716 163780 195826
rect 164856 193716 164884 195962
rect 165960 193716 165988 196302
rect 167248 195890 167276 208934
rect 168628 196026 168656 208934
rect 169904 206220 169956 206226
rect 169904 206162 169956 206168
rect 168616 196020 168668 196026
rect 168616 195962 168668 195968
rect 167236 195884 167288 195890
rect 167236 195826 167288 195832
rect 167142 195240 167198 195249
rect 167142 195175 167198 195184
rect 167156 193716 167184 195175
rect 169916 193866 169944 206162
rect 170008 196366 170036 208934
rect 172350 208934 172644 208962
rect 174056 208934 174116 208962
rect 175424 208950 175476 208956
rect 172294 208911 172350 208920
rect 174056 207518 174084 208934
rect 174044 207512 174096 207518
rect 174044 207454 174096 207460
rect 169996 196360 170048 196366
rect 169996 196302 170048 196308
rect 173768 196088 173820 196094
rect 173768 196030 173820 196036
rect 172664 196020 172716 196026
rect 172664 195962 172716 195968
rect 171560 195952 171612 195958
rect 171560 195894 171612 195900
rect 170456 195884 170508 195890
rect 170456 195826 170508 195832
rect 169732 193838 169944 193866
rect 169732 193730 169760 193838
rect 169378 193702 169760 193730
rect 170468 193716 170496 195826
rect 171572 193716 171600 195894
rect 172676 193716 172704 195962
rect 173780 193716 173808 196030
rect 175436 193866 175464 208950
rect 176816 196366 176844 210310
rect 177172 210300 177224 210306
rect 177172 210242 177224 210248
rect 177184 210073 177212 210242
rect 177724 210232 177776 210238
rect 177724 210174 177776 210180
rect 177170 210064 177226 210073
rect 177170 209999 177226 210008
rect 177736 209529 177764 210174
rect 177722 209520 177778 209529
rect 177722 209455 177778 209464
rect 178196 196366 178224 210378
rect 180312 207518 180340 233838
rect 185280 233834 185308 234479
rect 185268 233828 185320 233834
rect 185268 233770 185320 233776
rect 185174 233456 185230 233465
rect 185174 233391 185230 233400
rect 185188 233086 185216 233391
rect 185176 233080 185228 233086
rect 185176 233022 185228 233028
rect 185174 232912 185230 232921
rect 185174 232847 185230 232856
rect 185188 232474 185216 232847
rect 185176 232468 185228 232474
rect 185176 232410 185228 232416
rect 185174 232368 185230 232377
rect 185174 232303 185230 232312
rect 185188 231726 185216 232303
rect 185266 231824 185322 231833
rect 185266 231759 185322 231768
rect 185176 231720 185228 231726
rect 185176 231662 185228 231668
rect 185174 231280 185230 231289
rect 185174 231215 185230 231224
rect 185188 231046 185216 231215
rect 185280 231114 185308 231759
rect 185268 231108 185320 231114
rect 185268 231050 185320 231056
rect 183704 231040 183756 231046
rect 183704 230982 183756 230988
rect 185176 231040 185228 231046
rect 185176 230982 185228 230988
rect 183716 230638 183744 230982
rect 185266 230736 185322 230745
rect 185266 230671 185322 230680
rect 183704 230632 183756 230638
rect 183704 230574 183756 230580
rect 185174 230056 185230 230065
rect 185174 229991 185230 230000
rect 185188 229618 185216 229991
rect 185176 229612 185228 229618
rect 185176 229554 185228 229560
rect 185280 229550 185308 230671
rect 185268 229544 185320 229550
rect 185174 229512 185230 229521
rect 185268 229486 185320 229492
rect 185174 229447 185230 229456
rect 185188 228938 185216 229447
rect 185266 228968 185322 228977
rect 185176 228932 185228 228938
rect 185266 228903 185322 228912
rect 185176 228874 185228 228880
rect 185174 228424 185230 228433
rect 185280 228394 185308 228903
rect 185174 228359 185230 228368
rect 185268 228388 185320 228394
rect 185188 228326 185216 228359
rect 185268 228330 185320 228336
rect 185176 228320 185228 228326
rect 185176 228262 185228 228268
rect 185174 227880 185230 227889
rect 185174 227815 185230 227824
rect 185188 226830 185216 227815
rect 185266 227336 185322 227345
rect 185266 227271 185322 227280
rect 185176 226824 185228 226830
rect 185176 226766 185228 226772
rect 185280 226762 185308 227271
rect 185358 226792 185414 226801
rect 185268 226756 185320 226762
rect 185358 226727 185414 226736
rect 185268 226698 185320 226704
rect 185266 226248 185322 226257
rect 185266 226183 185322 226192
rect 185174 225568 185230 225577
rect 185174 225503 185230 225512
rect 185188 225402 185216 225503
rect 185176 225396 185228 225402
rect 185176 225338 185228 225344
rect 185280 225334 185308 226183
rect 185372 225470 185400 226727
rect 185360 225464 185412 225470
rect 185360 225406 185412 225412
rect 185268 225328 185320 225334
rect 185268 225270 185320 225276
rect 185266 225024 185322 225033
rect 185266 224959 185322 224968
rect 185174 224480 185230 224489
rect 185174 224415 185230 224424
rect 185188 224042 185216 224415
rect 185280 224110 185308 224959
rect 185268 224104 185320 224110
rect 185268 224046 185320 224052
rect 185176 224036 185228 224042
rect 185176 223978 185228 223984
rect 185266 223936 185322 223945
rect 185266 223871 185322 223880
rect 185174 223392 185230 223401
rect 185174 223327 185230 223336
rect 185082 222848 185138 222857
rect 185082 222783 185138 222792
rect 185096 221186 185124 222783
rect 185188 222750 185216 223327
rect 185176 222744 185228 222750
rect 185176 222686 185228 222692
rect 185280 222682 185308 223871
rect 185268 222676 185320 222682
rect 185268 222618 185320 222624
rect 185266 222304 185322 222313
rect 185266 222239 185322 222248
rect 185174 221760 185230 221769
rect 185174 221695 185230 221704
rect 185188 221322 185216 221695
rect 185176 221316 185228 221322
rect 185176 221258 185228 221264
rect 185280 221254 185308 222239
rect 185268 221248 185320 221254
rect 185268 221190 185320 221196
rect 185358 221216 185414 221225
rect 185084 221180 185136 221186
rect 215640 221202 215668 235130
rect 222342 231688 222398 231697
rect 222342 231623 222398 231632
rect 222356 231114 222384 231623
rect 217560 231108 217612 231114
rect 217560 231050 217612 231056
rect 222344 231108 222396 231114
rect 222344 231050 222396 231056
rect 215718 221216 215774 221225
rect 215640 221174 215718 221202
rect 185358 221151 185414 221160
rect 215718 221151 215774 221160
rect 185084 221122 185136 221128
rect 185174 220536 185230 220545
rect 185174 220471 185230 220480
rect 185082 219992 185138 220001
rect 185188 219962 185216 220471
rect 185082 219927 185138 219936
rect 185176 219956 185228 219962
rect 185096 218534 185124 219927
rect 185176 219898 185228 219904
rect 185372 219894 185400 221151
rect 185360 219888 185412 219894
rect 185360 219830 185412 219836
rect 185818 219448 185874 219457
rect 185818 219383 185874 219392
rect 185174 218904 185230 218913
rect 185174 218839 185230 218848
rect 185188 218670 185216 218839
rect 185176 218664 185228 218670
rect 185176 218606 185228 218612
rect 185832 218602 185860 219383
rect 185820 218596 185872 218602
rect 185820 218538 185872 218544
rect 185084 218528 185136 218534
rect 185084 218470 185136 218476
rect 185174 218360 185230 218369
rect 185174 218295 185230 218304
rect 184990 217816 185046 217825
rect 184990 217751 185046 217760
rect 184806 216048 184862 216057
rect 184806 215983 184862 215992
rect 184820 214386 184848 215983
rect 185004 215746 185032 217751
rect 185082 217272 185138 217281
rect 185188 217242 185216 218295
rect 185082 217207 185138 217216
rect 185176 217236 185228 217242
rect 184992 215740 185044 215746
rect 184992 215682 185044 215688
rect 185096 215678 185124 217207
rect 185176 217178 185228 217184
rect 185174 216728 185230 216737
rect 185174 216663 185230 216672
rect 185188 215814 185216 216663
rect 185176 215808 185228 215814
rect 185176 215750 185228 215756
rect 185084 215672 185136 215678
rect 185084 215614 185136 215620
rect 185174 215504 185230 215513
rect 185174 215439 185230 215448
rect 184898 214960 184954 214969
rect 184898 214895 184954 214904
rect 184808 214380 184860 214386
rect 184808 214322 184860 214328
rect 184912 213026 184940 214895
rect 185188 214454 185216 215439
rect 185176 214448 185228 214454
rect 185176 214390 185228 214396
rect 185266 214416 185322 214425
rect 185266 214351 185322 214360
rect 184990 213872 185046 213881
rect 184990 213807 185046 213816
rect 184900 213020 184952 213026
rect 184900 212962 184952 212968
rect 181772 211728 181824 211734
rect 181772 211670 181824 211676
rect 181784 210850 181812 211670
rect 185004 211666 185032 213807
rect 185082 213328 185138 213337
rect 185082 213263 185138 213272
rect 184992 211660 185044 211666
rect 184992 211602 185044 211608
rect 185096 211598 185124 213263
rect 185280 213094 185308 214351
rect 185268 213088 185320 213094
rect 185268 213030 185320 213036
rect 185174 212784 185230 212793
rect 185174 212719 185230 212728
rect 185188 211734 185216 212719
rect 185450 212240 185506 212249
rect 185450 212175 185506 212184
rect 185176 211728 185228 211734
rect 185176 211670 185228 211676
rect 185084 211592 185136 211598
rect 185084 211534 185136 211540
rect 185358 211560 185414 211569
rect 185358 211495 185414 211504
rect 185266 211016 185322 211025
rect 185266 210951 185322 210960
rect 181772 210844 181824 210850
rect 181772 210786 181824 210792
rect 185174 210472 185230 210481
rect 185280 210442 185308 210951
rect 185174 210407 185230 210416
rect 185268 210436 185320 210442
rect 185188 210374 185216 210407
rect 185268 210378 185320 210384
rect 185176 210368 185228 210374
rect 185176 210310 185228 210316
rect 185372 210238 185400 211495
rect 185464 210306 185492 212175
rect 185452 210300 185504 210306
rect 185452 210242 185504 210248
rect 185360 210232 185412 210238
rect 185360 210174 185412 210180
rect 185174 209928 185230 209937
rect 185174 209863 185230 209872
rect 185188 209014 185216 209863
rect 185726 209384 185782 209393
rect 185726 209319 185782 209328
rect 185176 209008 185228 209014
rect 185176 208950 185228 208956
rect 180300 207512 180352 207518
rect 180300 207454 180352 207460
rect 185174 207208 185230 207217
rect 185174 207143 185230 207152
rect 185188 206226 185216 207143
rect 185176 206220 185228 206226
rect 185176 206162 185228 206168
rect 183612 204248 183664 204254
rect 183612 204190 183664 204196
rect 183428 204112 183480 204118
rect 183428 204054 183480 204060
rect 183336 203704 183388 203710
rect 183336 203646 183388 203652
rect 183244 203636 183296 203642
rect 183244 203578 183296 203584
rect 183152 203568 183204 203574
rect 183152 203510 183204 203516
rect 183060 203500 183112 203506
rect 183060 203442 183112 203448
rect 175976 196360 176028 196366
rect 175976 196302 176028 196308
rect 176804 196360 176856 196366
rect 176804 196302 176856 196308
rect 177080 196360 177132 196366
rect 177080 196302 177132 196308
rect 178184 196360 178236 196366
rect 178184 196302 178236 196308
rect 175252 193838 175464 193866
rect 175252 193730 175280 193838
rect 174898 193702 175280 193730
rect 175988 193716 176016 196302
rect 177092 193716 177120 196302
rect 179288 195816 179340 195822
rect 179288 195758 179340 195764
rect 179300 193716 179328 195758
rect 99522 193679 99578 193688
rect 105778 192520 105834 192529
rect 105778 192455 105834 192464
rect 99430 192384 99486 192393
rect 99430 192319 99486 192328
rect 99338 188984 99394 188993
rect 99338 188919 99394 188928
rect 99062 187760 99118 187769
rect 99062 187695 99118 187704
rect 99432 186908 99484 186914
rect 99432 186850 99484 186856
rect 98970 186536 99026 186545
rect 98970 186471 99026 186480
rect 98878 185312 98934 185321
rect 98878 185247 98934 185256
rect 98604 182692 98656 182698
rect 98604 182634 98656 182640
rect 98616 182465 98644 182634
rect 98602 182456 98658 182465
rect 98602 182391 98658 182400
rect 99444 181105 99472 186850
rect 104400 184120 104452 184126
rect 104400 184062 104452 184068
rect 99524 184052 99576 184058
rect 99524 183994 99576 184000
rect 99536 183689 99564 183994
rect 99522 183680 99578 183689
rect 99522 183615 99578 183624
rect 99430 181096 99486 181105
rect 99430 181031 99486 181040
rect 98420 179904 98472 179910
rect 98420 179846 98472 179852
rect 99522 179872 99578 179881
rect 98432 179337 98460 179846
rect 99522 179807 99578 179816
rect 99536 179570 99564 179807
rect 104412 179570 104440 184062
rect 105792 184058 105820 192455
rect 107158 190208 107214 190217
rect 107158 190143 107214 190152
rect 106790 187896 106846 187905
rect 106790 187831 106846 187840
rect 106804 186914 106832 187831
rect 106792 186908 106844 186914
rect 106792 186850 106844 186856
rect 106790 185448 106846 185457
rect 106790 185383 106846 185392
rect 106804 184126 106832 185383
rect 106792 184120 106844 184126
rect 106792 184062 106844 184068
rect 105780 184052 105832 184058
rect 105780 183994 105832 184000
rect 107172 183258 107200 190143
rect 183072 184641 183100 203442
rect 183164 185865 183192 203510
rect 183256 187089 183284 203578
rect 183348 188313 183376 203646
rect 183440 190761 183468 204054
rect 183520 203432 183572 203438
rect 183520 203374 183572 203380
rect 183426 190752 183482 190761
rect 183426 190687 183482 190696
rect 183532 189537 183560 203374
rect 183624 191985 183652 204190
rect 183704 204180 183756 204186
rect 183704 204122 183756 204128
rect 183716 193209 183744 204122
rect 185740 204100 185768 209319
rect 185910 208840 185966 208849
rect 185910 208775 185966 208784
rect 185740 204072 185860 204100
rect 185832 196094 185860 204072
rect 185820 196088 185872 196094
rect 185820 196030 185872 196036
rect 185924 196026 185952 208775
rect 186278 208296 186334 208305
rect 186278 208231 186334 208240
rect 186094 207752 186150 207761
rect 186094 207687 186150 207696
rect 185912 196020 185964 196026
rect 185912 195962 185964 195968
rect 186108 195890 186136 207687
rect 186292 195958 186320 208231
rect 201104 207030 201578 207058
rect 188224 203506 188252 206908
rect 188776 203574 188804 206908
rect 189328 203642 189356 206908
rect 189880 203710 189908 206908
rect 189868 203704 189920 203710
rect 189868 203646 189920 203652
rect 189316 203636 189368 203642
rect 189316 203578 189368 203584
rect 188764 203568 188816 203574
rect 188764 203510 188816 203516
rect 188212 203500 188264 203506
rect 188212 203442 188264 203448
rect 190432 203438 190460 206908
rect 190984 204118 191012 206908
rect 191536 204254 191564 206908
rect 191524 204248 191576 204254
rect 191524 204190 191576 204196
rect 192088 204186 192116 206908
rect 192076 204180 192128 204186
rect 192076 204122 192128 204128
rect 190972 204112 191024 204118
rect 190972 204054 191024 204060
rect 191984 204112 192036 204118
rect 191984 204054 192036 204060
rect 190420 203432 190472 203438
rect 190420 203374 190472 203380
rect 186280 195952 186332 195958
rect 186280 195894 186332 195900
rect 186096 195884 186148 195890
rect 186096 195826 186148 195832
rect 183702 193200 183758 193209
rect 183702 193135 183758 193144
rect 191996 192801 192024 204054
rect 192640 203438 192668 206908
rect 193206 206894 193312 206922
rect 192628 203432 192680 203438
rect 192628 203374 192680 203380
rect 193284 196026 193312 206894
rect 193744 203438 193772 206908
rect 194310 206894 194692 206922
rect 194862 206894 194968 206922
rect 193364 203432 193416 203438
rect 193364 203374 193416 203380
rect 193732 203432 193784 203438
rect 193732 203374 193784 203380
rect 193272 196020 193324 196026
rect 193272 195962 193324 195968
rect 193376 195226 193404 203374
rect 194468 196020 194520 196026
rect 194468 195962 194520 195968
rect 193376 195198 193680 195226
rect 193652 193730 193680 195198
rect 193652 193702 194126 193730
rect 194480 193716 194508 195962
rect 194664 195278 194692 206894
rect 194744 203432 194796 203438
rect 194744 203374 194796 203380
rect 194756 196314 194784 203374
rect 194756 196286 194876 196314
rect 194652 195272 194704 195278
rect 194652 195214 194704 195220
rect 194848 193716 194876 196286
rect 194940 195754 194968 206894
rect 195124 206894 195506 206922
rect 196058 206894 196164 206922
rect 195124 196366 195152 206894
rect 195112 196360 195164 196366
rect 195112 196302 195164 196308
rect 196032 196360 196084 196366
rect 196032 196302 196084 196308
rect 194928 195748 194980 195754
rect 194928 195690 194980 195696
rect 195664 195748 195716 195754
rect 195664 195690 195716 195696
rect 195296 195272 195348 195278
rect 195296 195214 195348 195220
rect 195308 193716 195336 195214
rect 195676 193716 195704 195690
rect 196044 193716 196072 196302
rect 196136 195226 196164 206894
rect 196320 206894 196610 206922
rect 196872 206894 197162 206922
rect 197516 206894 197714 206922
rect 197792 206894 198266 206922
rect 198344 206894 198818 206922
rect 198988 206894 199370 206922
rect 199540 206894 199922 206922
rect 200368 206894 200474 206922
rect 196216 201460 196268 201466
rect 196216 201402 196268 201408
rect 196228 196366 196256 201402
rect 196320 196434 196348 206894
rect 196872 201466 196900 206894
rect 197516 202894 197544 206894
rect 197792 204474 197820 206894
rect 197608 204446 197820 204474
rect 197504 202888 197556 202894
rect 197504 202830 197556 202836
rect 196860 201460 196912 201466
rect 196860 201402 196912 201408
rect 196308 196428 196360 196434
rect 196308 196370 196360 196376
rect 196860 196428 196912 196434
rect 196860 196370 196912 196376
rect 196216 196360 196268 196366
rect 196216 196302 196268 196308
rect 196136 195198 196256 195226
rect 196228 193730 196256 195198
rect 196228 193702 196518 193730
rect 196872 193716 196900 196370
rect 197228 196360 197280 196366
rect 197228 196302 197280 196308
rect 197240 193716 197268 196302
rect 197608 195414 197636 204446
rect 198344 203114 198372 206894
rect 198988 203420 199016 206894
rect 197976 203086 198372 203114
rect 198896 203392 199016 203420
rect 197780 202888 197832 202894
rect 197780 202830 197832 202836
rect 197596 195408 197648 195414
rect 197596 195350 197648 195356
rect 197792 193730 197820 202830
rect 197976 195498 198004 203086
rect 197976 195470 198188 195498
rect 198056 195408 198108 195414
rect 198056 195350 198108 195356
rect 197714 193702 197820 193730
rect 198068 193716 198096 195350
rect 198160 193730 198188 195470
rect 198160 193702 198450 193730
rect 198896 193716 198924 203392
rect 199540 203114 199568 206894
rect 200368 204474 200396 206894
rect 199172 203086 199568 203114
rect 200184 204446 200396 204474
rect 199172 193730 199200 203086
rect 200184 194002 200212 204446
rect 201012 204390 201040 206908
rect 200264 204384 200316 204390
rect 200264 204326 200316 204332
rect 201000 204384 201052 204390
rect 201000 204326 201052 204332
rect 200000 193974 200212 194002
rect 200000 193730 200028 193974
rect 200276 193730 200304 204326
rect 201104 203114 201132 207030
rect 201748 206894 202222 206922
rect 201460 203636 201512 203642
rect 201460 203578 201512 203584
rect 200552 203086 201132 203114
rect 200552 193730 200580 203086
rect 200816 196428 200868 196434
rect 200816 196370 200868 196376
rect 199172 193702 199278 193730
rect 199646 193702 200028 193730
rect 200106 193702 200304 193730
rect 200474 193702 200580 193730
rect 200828 193716 200856 196370
rect 201472 196298 201500 203578
rect 201748 203522 201776 206894
rect 201656 203494 201776 203522
rect 201552 203432 201604 203438
rect 201552 203374 201604 203380
rect 201460 196292 201512 196298
rect 201460 196234 201512 196240
rect 201564 193730 201592 203374
rect 201656 196434 201684 203494
rect 202760 203438 202788 206908
rect 203312 203642 203340 206908
rect 203300 203636 203352 203642
rect 203300 203578 203352 203584
rect 202932 203568 202984 203574
rect 202932 203510 202984 203516
rect 202748 203432 202800 203438
rect 202748 203374 202800 203380
rect 202840 203432 202892 203438
rect 202840 203374 202892 203380
rect 201644 196428 201696 196434
rect 201644 196370 201696 196376
rect 201644 196292 201696 196298
rect 201644 196234 201696 196240
rect 201302 193702 201592 193730
rect 201656 193716 201684 196234
rect 202852 196026 202880 203374
rect 202104 196020 202156 196026
rect 202104 195962 202156 195968
rect 202840 196020 202892 196026
rect 202840 195962 202892 195968
rect 202116 193716 202144 195962
rect 202944 194002 202972 203510
rect 203024 203500 203076 203506
rect 203024 203442 203076 203448
rect 202760 193974 202972 194002
rect 202760 193730 202788 193974
rect 203036 193730 203064 203442
rect 203864 203438 203892 206908
rect 204312 203704 204364 203710
rect 204312 203646 204364 203652
rect 204220 203636 204272 203642
rect 204220 203578 204272 203584
rect 203852 203432 203904 203438
rect 203852 203374 203904 203380
rect 204232 196434 204260 203578
rect 203668 196428 203720 196434
rect 203668 196370 203720 196376
rect 204220 196428 204272 196434
rect 204220 196370 204272 196376
rect 203300 196360 203352 196366
rect 203300 196302 203352 196308
rect 202498 193702 202788 193730
rect 202866 193702 203064 193730
rect 203312 193716 203340 196302
rect 203680 193716 203708 196370
rect 204324 193730 204352 203646
rect 204416 203574 204444 206908
rect 204404 203568 204456 203574
rect 204404 203510 204456 203516
rect 204968 203506 204996 206908
rect 204956 203500 205008 203506
rect 204956 203442 205008 203448
rect 205416 203500 205468 203506
rect 205416 203442 205468 203448
rect 204404 203432 204456 203438
rect 204404 203374 204456 203380
rect 204416 196366 204444 203374
rect 205428 203114 205456 203442
rect 205520 203438 205548 206908
rect 205692 203772 205744 203778
rect 205692 203714 205744 203720
rect 205508 203432 205560 203438
rect 205508 203374 205560 203380
rect 205600 203432 205652 203438
rect 205600 203374 205652 203380
rect 205428 203086 205548 203114
rect 205520 196434 205548 203086
rect 204496 196428 204548 196434
rect 204496 196370 204548 196376
rect 205508 196428 205560 196434
rect 205508 196370 205560 196376
rect 204404 196360 204456 196366
rect 204404 196302 204456 196308
rect 204062 193702 204352 193730
rect 204508 193716 204536 196370
rect 205612 196366 205640 203374
rect 204864 196360 204916 196366
rect 204864 196302 204916 196308
rect 205600 196360 205652 196366
rect 205600 196302 205652 196308
rect 204876 193716 204904 196302
rect 205232 196292 205284 196298
rect 205232 196234 205284 196240
rect 205244 193716 205272 196234
rect 205704 193716 205732 203714
rect 206072 203642 206100 206908
rect 206624 203710 206652 206908
rect 206612 203704 206664 203710
rect 206612 203646 206664 203652
rect 206060 203636 206112 203642
rect 206060 203578 206112 203584
rect 205784 203568 205836 203574
rect 205784 203510 205836 203516
rect 205796 196298 205824 203510
rect 207176 203506 207204 206908
rect 207164 203500 207216 203506
rect 207164 203442 207216 203448
rect 207728 203438 207756 206908
rect 207900 204452 207952 204458
rect 207900 204394 207952 204400
rect 207716 203432 207768 203438
rect 207716 203374 207768 203380
rect 207624 196360 207676 196366
rect 207624 196302 207676 196308
rect 205784 196292 205836 196298
rect 205784 196234 205836 196240
rect 206428 196156 206480 196162
rect 206428 196098 206480 196104
rect 206060 195748 206112 195754
rect 206060 195690 206112 195696
rect 206072 193716 206100 195690
rect 206440 193716 206468 196098
rect 207256 195680 207308 195686
rect 207256 195622 207308 195628
rect 206888 195612 206940 195618
rect 206888 195554 206940 195560
rect 206900 193716 206928 195554
rect 207268 193716 207296 195622
rect 207636 193716 207664 196302
rect 207912 195618 207940 204394
rect 208084 204316 208136 204322
rect 208084 204258 208136 204264
rect 207992 203432 208044 203438
rect 207992 203374 208044 203380
rect 208004 195754 208032 203374
rect 208096 196162 208124 204258
rect 208280 203574 208308 206908
rect 208544 204588 208596 204594
rect 208544 204530 208596 204536
rect 208452 204248 208504 204254
rect 208452 204190 208504 204196
rect 208360 204180 208412 204186
rect 208360 204122 208412 204128
rect 208268 203568 208320 203574
rect 208268 203510 208320 203516
rect 208084 196156 208136 196162
rect 208084 196098 208136 196104
rect 207992 195748 208044 195754
rect 207992 195690 208044 195696
rect 207900 195612 207952 195618
rect 207900 195554 207952 195560
rect 208372 193730 208400 204122
rect 208464 196366 208492 204190
rect 208452 196360 208504 196366
rect 208452 196302 208504 196308
rect 208452 195816 208504 195822
rect 208452 195758 208504 195764
rect 208110 193702 208400 193730
rect 208464 193716 208492 195758
rect 208556 195686 208584 204530
rect 208832 203778 208860 206908
rect 208820 203772 208872 203778
rect 208820 203714 208872 203720
rect 209476 203438 209504 206908
rect 210028 204322 210056 206908
rect 210580 204458 210608 206908
rect 211132 204594 211160 206908
rect 211120 204588 211172 204594
rect 211120 204530 211172 204536
rect 210568 204452 210620 204458
rect 210568 204394 210620 204400
rect 210016 204316 210068 204322
rect 210016 204258 210068 204264
rect 211684 204254 211712 206908
rect 211672 204248 211724 204254
rect 211672 204190 211724 204196
rect 212236 204186 212264 206908
rect 212802 206894 213000 206922
rect 212224 204180 212276 204186
rect 212224 204122 212276 204128
rect 209464 203432 209516 203438
rect 209464 203374 209516 203380
rect 212868 203092 212920 203098
rect 212868 203034 212920 203040
rect 209280 196020 209332 196026
rect 209280 195962 209332 195968
rect 208820 195952 208872 195958
rect 208820 195894 208872 195900
rect 208544 195680 208596 195686
rect 208544 195622 208596 195628
rect 208832 193716 208860 195894
rect 209292 193716 209320 195962
rect 212880 195958 212908 203034
rect 212868 195952 212920 195958
rect 212868 195894 212920 195900
rect 209648 195884 209700 195890
rect 209648 195826 209700 195832
rect 209660 193716 209688 195826
rect 212972 195822 213000 206894
rect 213064 206894 213354 206922
rect 213432 206894 213906 206922
rect 213064 203098 213092 206894
rect 213432 203658 213460 206894
rect 213156 203630 213460 203658
rect 213052 203092 213104 203098
rect 213052 203034 213104 203040
rect 213156 202978 213184 203630
rect 214444 203438 214472 206908
rect 214996 204118 215024 206908
rect 215548 204798 215576 206908
rect 216180 204860 216232 204866
rect 216180 204802 216232 204808
rect 215536 204792 215588 204798
rect 215536 204734 215588 204740
rect 214984 204112 215036 204118
rect 214984 204054 215036 204060
rect 213420 203432 213472 203438
rect 213420 203374 213472 203380
rect 214432 203432 214484 203438
rect 214432 203374 214484 203380
rect 213064 202950 213184 202978
rect 213064 196026 213092 202950
rect 213052 196020 213104 196026
rect 213052 195962 213104 195968
rect 213432 195890 213460 203374
rect 213420 195884 213472 195890
rect 213420 195826 213472 195832
rect 212960 195816 213012 195822
rect 212960 195758 213012 195764
rect 191982 192792 192038 192801
rect 191982 192727 192038 192736
rect 183610 191976 183666 191985
rect 183610 191911 183666 191920
rect 209752 190846 209964 190874
rect 183518 189528 183574 189537
rect 183518 189463 183574 189472
rect 191982 188712 192038 188721
rect 191982 188647 192038 188656
rect 183334 188304 183390 188313
rect 191996 188274 192024 188647
rect 183334 188239 183390 188248
rect 187936 188268 187988 188274
rect 187936 188210 187988 188216
rect 191984 188268 192036 188274
rect 191984 188210 192036 188216
rect 183242 187080 183298 187089
rect 183242 187015 183298 187024
rect 183150 185856 183206 185865
rect 183150 185791 183206 185800
rect 183058 184632 183114 184641
rect 183058 184567 183114 184576
rect 187948 184058 187976 188210
rect 191154 186808 191210 186817
rect 191154 186743 191210 186752
rect 182876 184052 182928 184058
rect 182876 183994 182928 184000
rect 187936 184052 187988 184058
rect 187936 183994 187988 184000
rect 128502 183816 128558 183825
rect 128502 183751 128558 183760
rect 106988 183230 107200 183258
rect 104492 182760 104544 182766
rect 104492 182702 104544 182708
rect 104504 179910 104532 182702
rect 106988 182698 107016 183230
rect 107158 183136 107214 183145
rect 107158 183071 107214 183080
rect 107172 182766 107200 183071
rect 128516 182766 128544 183751
rect 182888 183417 182916 183994
rect 182874 183408 182930 183417
rect 182874 183343 182930 183352
rect 107160 182760 107212 182766
rect 107160 182702 107212 182708
rect 128504 182760 128556 182766
rect 128504 182702 128556 182708
rect 137520 182760 137572 182766
rect 137520 182702 137572 182708
rect 190602 182728 190658 182737
rect 106976 182692 107028 182698
rect 106976 182634 107028 182640
rect 106974 180824 107030 180833
rect 106974 180759 107030 180768
rect 106988 180386 107016 180759
rect 105136 180380 105188 180386
rect 105136 180322 105188 180328
rect 106976 180380 107028 180386
rect 106976 180322 107028 180328
rect 104492 179904 104544 179910
rect 104492 179846 104544 179852
rect 99524 179564 99576 179570
rect 99524 179506 99576 179512
rect 104400 179564 104452 179570
rect 104400 179506 104452 179512
rect 98418 179328 98474 179337
rect 98418 179263 98474 179272
rect 99522 177424 99578 177433
rect 105148 177394 105176 180322
rect 106790 178376 106846 178385
rect 106790 178311 106846 178320
rect 99522 177359 99524 177368
rect 99576 177359 99578 177368
rect 105136 177388 105188 177394
rect 99524 177330 99576 177336
rect 105136 177330 105188 177336
rect 106804 177190 106832 178311
rect 98604 177184 98656 177190
rect 98604 177126 98656 177132
rect 106792 177184 106844 177190
rect 106792 177126 106844 177132
rect 98616 176753 98644 177126
rect 98602 176744 98658 176753
rect 98602 176679 98658 176688
rect 106606 176064 106662 176073
rect 106606 175999 106662 176008
rect 106620 175830 106648 175999
rect 98236 175824 98288 175830
rect 98236 175766 98288 175772
rect 106608 175824 106660 175830
rect 106608 175766 106660 175772
rect 98248 175393 98276 175766
rect 98234 175384 98290 175393
rect 98234 175319 98290 175328
rect 137532 174441 137560 182702
rect 183152 182692 183204 182698
rect 191168 182698 191196 186743
rect 191982 184768 192038 184777
rect 191982 184703 192038 184712
rect 190602 182663 190658 182672
rect 191156 182692 191208 182698
rect 183152 182634 183204 182640
rect 183164 182193 183192 182634
rect 183150 182184 183206 182193
rect 183150 182119 183206 182128
rect 183704 181332 183756 181338
rect 183704 181274 183756 181280
rect 183716 181105 183744 181274
rect 183702 181096 183758 181105
rect 183702 181031 183758 181040
rect 182508 179904 182560 179910
rect 182508 179846 182560 179852
rect 183702 179872 183758 179881
rect 182520 178657 182548 179846
rect 190616 179842 190644 182663
rect 191156 182634 191208 182640
rect 191996 181338 192024 184703
rect 191984 181332 192036 181338
rect 191984 181274 192036 181280
rect 190694 180824 190750 180833
rect 190694 180759 190750 180768
rect 190708 179910 190736 180759
rect 190696 179904 190748 179910
rect 190696 179846 190748 179852
rect 183702 179807 183704 179816
rect 183756 179807 183758 179816
rect 190604 179836 190656 179842
rect 183704 179778 183756 179784
rect 190604 179778 190656 179784
rect 191982 178784 192038 178793
rect 191982 178719 192038 178728
rect 182506 178648 182562 178657
rect 182506 178583 182562 178592
rect 191996 178550 192024 178719
rect 182508 178544 182560 178550
rect 182508 178486 182560 178492
rect 191984 178544 192036 178550
rect 191984 178486 192036 178492
rect 182520 177433 182548 178486
rect 182506 177424 182562 177433
rect 182506 177359 182562 177368
rect 191982 176744 192038 176753
rect 191982 176679 192038 176688
rect 191996 176510 192024 176679
rect 183244 176504 183296 176510
rect 183244 176446 183296 176452
rect 191984 176504 192036 176510
rect 191984 176446 192036 176452
rect 183256 176209 183284 176446
rect 183242 176200 183298 176209
rect 183242 176135 183298 176144
rect 183704 175144 183756 175150
rect 183704 175086 183756 175092
rect 191524 175144 191576 175150
rect 191524 175086 191576 175092
rect 183716 174985 183744 175086
rect 183702 174976 183758 174985
rect 183702 174911 183758 174920
rect 191536 174849 191564 175086
rect 191522 174840 191578 174849
rect 191522 174775 191578 174784
rect 137518 174432 137574 174441
rect 137518 174367 137574 174376
rect 99522 173752 99578 173761
rect 99522 173687 99524 173696
rect 99576 173687 99578 173696
rect 106790 173752 106846 173761
rect 106790 173687 106792 173696
rect 99524 173658 99576 173664
rect 106844 173687 106846 173696
rect 183334 173752 183390 173761
rect 183334 173687 183390 173696
rect 106792 173658 106844 173664
rect 183348 173110 183376 173687
rect 183336 173104 183388 173110
rect 183336 173046 183388 173052
rect 191984 173104 192036 173110
rect 191984 173046 192036 173052
rect 191996 172809 192024 173046
rect 191982 172800 192038 172809
rect 191982 172735 192038 172744
rect 99522 172528 99578 172537
rect 99522 172463 99578 172472
rect 183518 172528 183574 172537
rect 183518 172463 183574 172472
rect 99536 171750 99564 172463
rect 183532 171750 183560 172463
rect 99524 171744 99576 171750
rect 99524 171686 99576 171692
rect 106792 171744 106844 171750
rect 106792 171686 106844 171692
rect 183520 171744 183572 171750
rect 183520 171686 183572 171692
rect 191156 171744 191208 171750
rect 191156 171686 191208 171692
rect 106804 171449 106832 171686
rect 106790 171440 106846 171449
rect 106790 171375 106846 171384
rect 99430 171304 99486 171313
rect 99430 171239 99486 171248
rect 182690 171304 182746 171313
rect 182690 171239 182692 171248
rect 99444 170322 99472 171239
rect 182744 171239 182746 171248
rect 185084 171268 185136 171274
rect 182692 171210 182744 171216
rect 185084 171210 185136 171216
rect 99432 170316 99484 170322
rect 99432 170258 99484 170264
rect 106792 170248 106844 170254
rect 106792 170190 106844 170196
rect 99522 170080 99578 170089
rect 99522 170015 99578 170024
rect 99536 168962 99564 170015
rect 106804 169001 106832 170190
rect 182506 170080 182562 170089
rect 182506 170015 182562 170024
rect 106790 168992 106846 169001
rect 99524 168956 99576 168962
rect 99524 168898 99576 168904
rect 106700 168956 106752 168962
rect 182520 168962 182548 170015
rect 106790 168927 106846 168936
rect 182508 168956 182560 168962
rect 106700 168898 106752 168904
rect 182508 168898 182560 168904
rect 99430 168856 99486 168865
rect 99430 168791 99486 168800
rect 99444 167602 99472 168791
rect 99522 167768 99578 167777
rect 99522 167703 99578 167712
rect 99536 167670 99564 167703
rect 99524 167664 99576 167670
rect 99524 167606 99576 167612
rect 99432 167596 99484 167602
rect 99432 167538 99484 167544
rect 106712 166689 106740 168898
rect 185096 168894 185124 171210
rect 191168 170769 191196 171686
rect 209752 171018 209780 190846
rect 209936 190761 209964 190846
rect 209922 190752 209978 190761
rect 209922 190687 209978 190696
rect 211948 190648 212000 190654
rect 211948 190590 212000 190596
rect 211960 190489 211988 190590
rect 211946 190480 212002 190489
rect 211946 190415 212002 190424
rect 212498 183816 212554 183825
rect 212498 183751 212554 183760
rect 212512 182766 212540 183751
rect 212500 182760 212552 182766
rect 212500 182702 212552 182708
rect 211762 177152 211818 177161
rect 211762 177087 211818 177096
rect 211776 176374 211804 177087
rect 211764 176368 211816 176374
rect 211764 176310 211816 176316
rect 209830 171032 209886 171041
rect 209752 170990 209830 171018
rect 209830 170967 209886 170976
rect 191154 170760 191210 170769
rect 191154 170695 191210 170704
rect 191892 168956 191944 168962
rect 191892 168898 191944 168904
rect 185084 168888 185136 168894
rect 183702 168856 183758 168865
rect 185084 168830 185136 168836
rect 183702 168791 183758 168800
rect 106884 167664 106936 167670
rect 106884 167606 106936 167612
rect 106792 167596 106844 167602
rect 106792 167538 106844 167544
rect 106698 166680 106754 166689
rect 106698 166615 106754 166624
rect 99522 166544 99578 166553
rect 99522 166479 99578 166488
rect 99536 166242 99564 166479
rect 99524 166236 99576 166242
rect 99524 166178 99576 166184
rect 99522 165320 99578 165329
rect 99522 165255 99578 165264
rect 99536 164814 99564 165255
rect 99524 164808 99576 164814
rect 99524 164750 99576 164756
rect 106804 164377 106832 167538
rect 106790 164368 106846 164377
rect 106790 164303 106846 164312
rect 99522 164096 99578 164105
rect 99522 164031 99578 164040
rect 99536 163454 99564 164031
rect 99524 163448 99576 163454
rect 99524 163390 99576 163396
rect 104400 163448 104452 163454
rect 104400 163390 104452 163396
rect 98970 162872 99026 162881
rect 98970 162807 99026 162816
rect 98786 154440 98842 154449
rect 98786 154375 98842 154384
rect 98236 151820 98288 151826
rect 98236 151762 98288 151768
rect 98248 151690 98276 151762
rect 98236 151684 98288 151690
rect 98236 151626 98288 151632
rect 98800 142986 98828 154375
rect 98880 151684 98932 151690
rect 98880 151626 98932 151632
rect 98788 142980 98840 142986
rect 98788 142922 98840 142928
rect 97868 137336 97920 137342
rect 97868 137278 97920 137284
rect 97880 137002 97908 137278
rect 97960 137268 98012 137274
rect 97960 137210 98012 137216
rect 97868 136996 97920 137002
rect 97868 136938 97920 136944
rect 97972 135710 98000 137210
rect 98052 135908 98104 135914
rect 98052 135850 98104 135856
rect 97960 135704 98012 135710
rect 97960 135646 98012 135652
rect 98064 134350 98092 135850
rect 98144 135840 98196 135846
rect 98144 135782 98196 135788
rect 98052 134344 98104 134350
rect 98052 134286 98104 134292
rect 98156 134282 98184 135782
rect 98144 134276 98196 134282
rect 98144 134218 98196 134224
rect 98052 126252 98104 126258
rect 98052 126194 98104 126200
rect 98064 124694 98092 126194
rect 98144 126184 98196 126190
rect 98144 126126 98196 126132
rect 98052 124688 98104 124694
rect 98052 124630 98104 124636
rect 98156 124626 98184 126126
rect 98144 124620 98196 124626
rect 98144 124562 98196 124568
rect 97868 120812 97920 120818
rect 97868 120754 97920 120760
rect 97684 119384 97736 119390
rect 97684 119326 97736 119332
rect 97696 117826 97724 119326
rect 97880 119118 97908 120754
rect 97960 120744 98012 120750
rect 97960 120686 98012 120692
rect 97972 119186 98000 120686
rect 98144 120676 98196 120682
rect 98144 120618 98196 120624
rect 98052 119316 98104 119322
rect 98052 119258 98104 119264
rect 97960 119180 98012 119186
rect 97960 119122 98012 119128
rect 97868 119112 97920 119118
rect 97868 119054 97920 119060
rect 97960 117956 98012 117962
rect 97960 117898 98012 117904
rect 97684 117820 97736 117826
rect 97684 117762 97736 117768
rect 97972 116398 98000 117898
rect 98064 117758 98092 119258
rect 98156 119254 98184 120618
rect 98144 119248 98196 119254
rect 98144 119190 98196 119196
rect 98144 117888 98196 117894
rect 98144 117830 98196 117836
rect 98052 117752 98104 117758
rect 98052 117694 98104 117700
rect 97960 116392 98012 116398
rect 97960 116334 98012 116340
rect 98156 116330 98184 117830
rect 98144 116324 98196 116330
rect 98144 116266 98196 116272
rect 98788 110272 98840 110278
rect 98788 110214 98840 110220
rect 98800 99777 98828 110214
rect 98786 99768 98842 99777
rect 98786 99703 98842 99712
rect 98788 97216 98840 97222
rect 98788 97158 98840 97164
rect 98696 93068 98748 93074
rect 98696 93010 98748 93016
rect 98708 87401 98736 93010
rect 98800 89985 98828 97158
rect 98786 89976 98842 89985
rect 98786 89911 98842 89920
rect 98694 87392 98750 87401
rect 98694 87327 98750 87336
rect 98234 75560 98290 75569
rect 98234 75495 98290 75504
rect 98248 75122 98276 75495
rect 98236 75116 98288 75122
rect 98236 75058 98288 75064
rect 98786 62776 98842 62785
rect 98786 62711 98842 62720
rect 98800 55062 98828 62711
rect 98892 58530 98920 151626
rect 98984 143394 99012 162807
rect 99062 161648 99118 161657
rect 99062 161583 99118 161592
rect 99076 143462 99104 161583
rect 99154 160424 99210 160433
rect 99154 160359 99210 160368
rect 99168 143530 99196 160359
rect 99246 159200 99302 159209
rect 99246 159135 99302 159144
rect 99260 143598 99288 159135
rect 99430 157976 99486 157985
rect 99430 157911 99486 157920
rect 99338 156752 99394 156761
rect 99338 156687 99394 156696
rect 99248 143592 99300 143598
rect 99248 143534 99300 143540
rect 99156 143524 99208 143530
rect 99156 143466 99208 143472
rect 99064 143456 99116 143462
rect 99064 143398 99116 143404
rect 98972 143388 99024 143394
rect 98972 143330 99024 143336
rect 99352 142850 99380 156687
rect 99444 142918 99472 157911
rect 99522 155528 99578 155537
rect 99522 155463 99578 155472
rect 99432 142912 99484 142918
rect 99432 142854 99484 142860
rect 99340 142844 99392 142850
rect 99340 142786 99392 142792
rect 99536 142782 99564 155463
rect 104412 155090 104440 163390
rect 106896 161929 106924 167606
rect 183716 167602 183744 168791
rect 183794 167768 183850 167777
rect 183794 167703 183850 167712
rect 183704 167596 183756 167602
rect 183704 167538 183756 167544
rect 182874 166544 182930 166553
rect 182874 166479 182876 166488
rect 182928 166479 182930 166488
rect 182876 166450 182928 166456
rect 107252 166236 107304 166242
rect 107252 166178 107304 166184
rect 107160 164808 107212 164814
rect 107160 164750 107212 164756
rect 106882 161920 106938 161929
rect 106882 161855 106938 161864
rect 107172 157305 107200 164750
rect 107264 159617 107292 166178
rect 183702 165320 183758 165329
rect 183702 165255 183758 165264
rect 183716 165018 183744 165255
rect 183704 165012 183756 165018
rect 183704 164954 183756 164960
rect 138162 164776 138218 164785
rect 138162 164711 138218 164720
rect 128502 163824 128558 163833
rect 128502 163759 128558 163768
rect 128516 163454 128544 163759
rect 138176 163454 138204 164711
rect 183058 164096 183114 164105
rect 183058 164031 183114 164040
rect 183072 163454 183100 164031
rect 128504 163448 128556 163454
rect 128504 163390 128556 163396
rect 138164 163448 138216 163454
rect 138164 163390 138216 163396
rect 183060 163448 183112 163454
rect 183060 163390 183112 163396
rect 138176 160569 138204 163390
rect 183808 163046 183836 167703
rect 191340 167596 191392 167602
rect 191340 167538 191392 167544
rect 187936 166508 187988 166514
rect 187936 166450 187988 166456
rect 183796 163040 183848 163046
rect 183796 162982 183848 162988
rect 183058 162872 183114 162881
rect 183058 162807 183114 162816
rect 138162 160560 138218 160569
rect 138162 160495 138218 160504
rect 107250 159608 107306 159617
rect 107250 159543 107306 159552
rect 107158 157296 107214 157305
rect 107158 157231 107214 157240
rect 182690 155528 182746 155537
rect 182690 155463 182692 155472
rect 182744 155463 182746 155472
rect 182692 155434 182744 155440
rect 104400 155084 104452 155090
rect 104400 155026 104452 155032
rect 106516 155084 106568 155090
rect 106516 155026 106568 155032
rect 106528 154993 106556 155026
rect 106514 154984 106570 154993
rect 106514 154919 106570 154928
rect 110116 152370 110144 153868
rect 109184 152364 109236 152370
rect 109184 152306 109236 152312
rect 110104 152364 110156 152370
rect 110104 152306 110156 152312
rect 106608 143592 106660 143598
rect 106608 143534 106660 143540
rect 103940 142980 103992 142986
rect 103940 142922 103992 142928
rect 99524 142776 99576 142782
rect 99524 142718 99576 142724
rect 103952 140826 103980 142922
rect 105596 142912 105648 142918
rect 105596 142854 105648 142860
rect 105136 142844 105188 142850
rect 105136 142786 105188 142792
rect 104584 142776 104636 142782
rect 104584 142718 104636 142724
rect 104596 140826 104624 142718
rect 105148 140826 105176 142786
rect 105608 140826 105636 142854
rect 103952 140798 104242 140826
rect 104596 140798 104794 140826
rect 105148 140798 105346 140826
rect 105608 140798 105990 140826
rect 106620 140690 106648 143534
rect 106792 143524 106844 143530
rect 106792 143466 106844 143472
rect 106804 140826 106832 143466
rect 107436 143456 107488 143462
rect 107436 143398 107488 143404
rect 107448 140826 107476 143398
rect 107988 143388 108040 143394
rect 107988 143330 108040 143336
rect 108000 140826 108028 143330
rect 106804 140798 107094 140826
rect 107448 140798 107738 140826
rect 108000 140798 108290 140826
rect 109196 140690 109224 152306
rect 110484 151010 110512 153868
rect 110668 153854 110866 153882
rect 110668 151026 110696 153854
rect 111312 151078 111340 153868
rect 109552 151004 109604 151010
rect 109552 150946 109604 150952
rect 110472 151004 110524 151010
rect 110472 150946 110524 150952
rect 110576 150998 110696 151026
rect 111300 151072 111352 151078
rect 111300 151014 111352 151020
rect 111680 151010 111708 153868
rect 112048 151026 112076 153868
rect 112508 151078 112536 153868
rect 111668 151004 111720 151010
rect 109564 140690 109592 150946
rect 110472 150868 110524 150874
rect 110472 150810 110524 150816
rect 110288 143252 110340 143258
rect 110288 143194 110340 143200
rect 110300 140690 110328 143194
rect 110484 140826 110512 150810
rect 110576 143258 110604 150998
rect 111668 150946 111720 150952
rect 111956 150998 112076 151026
rect 112496 151072 112548 151078
rect 112496 151014 112548 151020
rect 112876 151010 112904 153868
rect 112128 151004 112180 151010
rect 110656 150936 110708 150942
rect 110656 150878 110708 150884
rect 110564 143252 110616 143258
rect 110564 143194 110616 143200
rect 110484 140798 110590 140826
rect 106542 140662 106648 140690
rect 108842 140662 109224 140690
rect 109486 140662 109592 140690
rect 110038 140662 110328 140690
rect 110668 140690 110696 150878
rect 111956 140690 111984 150998
rect 112128 150946 112180 150952
rect 112864 151004 112916 151010
rect 112864 150946 112916 150952
rect 112036 150936 112088 150942
rect 112036 150878 112088 150884
rect 112048 140826 112076 150878
rect 112140 140962 112168 150946
rect 113244 142594 113272 153868
rect 113612 153854 113718 153882
rect 113244 142566 113456 142594
rect 112140 140934 112444 140962
rect 112048 140798 112338 140826
rect 110668 140662 111234 140690
rect 111786 140662 111984 140690
rect 112416 140690 112444 140934
rect 113428 140826 113456 142566
rect 113612 140826 113640 153854
rect 114072 141098 114100 153868
rect 114440 143666 114468 153868
rect 114428 143660 114480 143666
rect 114428 143602 114480 143608
rect 114900 143598 114928 153868
rect 115282 153854 115572 153882
rect 115544 150346 115572 153854
rect 115636 151010 115664 153868
rect 115912 153854 116110 153882
rect 115624 151004 115676 151010
rect 115624 150946 115676 150952
rect 115544 150318 115848 150346
rect 114980 143660 115032 143666
rect 114980 143602 115032 143608
rect 114888 143592 114940 143598
rect 114888 143534 114940 143540
rect 114072 141070 114192 141098
rect 114164 140826 114192 141070
rect 114992 140826 115020 143602
rect 115532 143592 115584 143598
rect 115532 143534 115584 143540
rect 115544 140826 115572 143534
rect 115820 142866 115848 150318
rect 115912 143598 115940 153854
rect 116464 151010 116492 153868
rect 115992 151004 116044 151010
rect 115992 150946 116044 150952
rect 116452 151004 116504 151010
rect 116452 150946 116504 150952
rect 116004 143666 116032 150946
rect 115992 143660 116044 143666
rect 115992 143602 116044 143608
rect 116636 143660 116688 143666
rect 116636 143602 116688 143608
rect 115900 143592 115952 143598
rect 115900 143534 115952 143540
rect 115820 142838 116216 142866
rect 116188 140826 116216 142838
rect 116648 140826 116676 143602
rect 116832 143122 116860 153868
rect 117292 143938 117320 153868
rect 117660 151010 117688 153868
rect 118120 151282 118148 153868
rect 118488 152302 118516 153868
rect 118476 152296 118528 152302
rect 118476 152238 118528 152244
rect 118856 152098 118884 153868
rect 118844 152092 118896 152098
rect 118844 152034 118896 152040
rect 119316 152030 119344 153868
rect 119684 152370 119712 153868
rect 119672 152364 119724 152370
rect 119672 152306 119724 152312
rect 120052 152166 120080 153868
rect 120512 152234 120540 153868
rect 120592 152296 120644 152302
rect 120592 152238 120644 152244
rect 120500 152228 120552 152234
rect 120500 152170 120552 152176
rect 120040 152160 120092 152166
rect 120040 152102 120092 152108
rect 119304 152024 119356 152030
rect 119304 151966 119356 151972
rect 118108 151276 118160 151282
rect 118108 151218 118160 151224
rect 120316 151276 120368 151282
rect 120316 151218 120368 151224
rect 117464 151004 117516 151010
rect 117464 150946 117516 150952
rect 117648 151004 117700 151010
rect 117648 150946 117700 150952
rect 118844 151004 118896 151010
rect 118844 150946 118896 150952
rect 117280 143932 117332 143938
rect 117280 143874 117332 143880
rect 117476 143666 117504 150946
rect 118856 144074 118884 150946
rect 118844 144068 118896 144074
rect 118844 144010 118896 144016
rect 119580 144068 119632 144074
rect 119580 144010 119632 144016
rect 119028 143932 119080 143938
rect 119028 143874 119080 143880
rect 117464 143660 117516 143666
rect 117464 143602 117516 143608
rect 117924 143660 117976 143666
rect 117924 143602 117976 143608
rect 117648 143592 117700 143598
rect 117648 143534 117700 143540
rect 116820 143116 116872 143122
rect 116820 143058 116872 143064
rect 113428 140798 113534 140826
rect 113612 140798 114086 140826
rect 114164 140798 114730 140826
rect 114992 140798 115282 140826
rect 115544 140798 115834 140826
rect 116188 140798 116478 140826
rect 116648 140798 117030 140826
rect 117660 140690 117688 143534
rect 117936 140826 117964 143602
rect 118476 143116 118528 143122
rect 118476 143058 118528 143064
rect 118488 140826 118516 143058
rect 119040 140826 119068 143874
rect 119592 140826 119620 144010
rect 120328 140826 120356 151218
rect 120604 140826 120632 152238
rect 120880 151078 120908 153868
rect 120960 152092 121012 152098
rect 120960 152034 121012 152040
rect 120868 151072 120920 151078
rect 120868 151014 120920 151020
rect 120972 144074 121000 152034
rect 121248 151282 121276 153868
rect 121708 151350 121736 153868
rect 121972 152364 122024 152370
rect 121972 152306 122024 152312
rect 121788 152024 121840 152030
rect 121788 151966 121840 151972
rect 121696 151344 121748 151350
rect 121696 151286 121748 151292
rect 121236 151276 121288 151282
rect 121236 151218 121288 151224
rect 120960 144068 121012 144074
rect 120960 144010 121012 144016
rect 121696 144068 121748 144074
rect 121696 144010 121748 144016
rect 121708 140962 121736 144010
rect 121800 141098 121828 151966
rect 121984 150890 122012 152306
rect 122076 151010 122104 153868
rect 122444 151486 122472 153868
rect 122904 151894 122932 153868
rect 123168 152228 123220 152234
rect 123168 152170 123220 152176
rect 123076 152160 123128 152166
rect 123076 152102 123128 152108
rect 122892 151888 122944 151894
rect 122892 151830 122944 151836
rect 122432 151480 122484 151486
rect 122432 151422 122484 151428
rect 122064 151004 122116 151010
rect 122064 150946 122116 150952
rect 121984 150862 122104 150890
rect 122076 150074 122104 150862
rect 122076 150046 122472 150074
rect 121800 141070 122012 141098
rect 121708 140934 121828 140962
rect 117936 140798 118226 140826
rect 118488 140798 118778 140826
rect 119040 140798 119330 140826
rect 119592 140798 119974 140826
rect 120328 140798 120526 140826
rect 120604 140798 121078 140826
rect 121800 140690 121828 140934
rect 121984 140826 122012 141070
rect 122444 140826 122472 150046
rect 123088 140826 123116 152102
rect 123180 140962 123208 152170
rect 123272 151894 123300 153868
rect 123640 152234 123668 153868
rect 123628 152228 123680 152234
rect 123628 152170 123680 152176
rect 123260 151888 123312 151894
rect 123260 151830 123312 151836
rect 124100 151554 124128 153868
rect 124468 152302 124496 153868
rect 124836 152370 124864 153868
rect 124824 152364 124876 152370
rect 124824 152306 124876 152312
rect 124456 152296 124508 152302
rect 124456 152238 124508 152244
rect 124088 151548 124140 151554
rect 124088 151490 124140 151496
rect 125100 151480 125152 151486
rect 125100 151422 125152 151428
rect 124640 151344 124692 151350
rect 124640 151286 124692 151292
rect 123720 151276 123772 151282
rect 123720 151218 123772 151224
rect 123732 144006 123760 151218
rect 123812 151072 123864 151078
rect 123812 151014 123864 151020
rect 123824 144074 123852 151014
rect 123812 144068 123864 144074
rect 123812 144010 123864 144016
rect 124456 144068 124508 144074
rect 124456 144010 124508 144016
rect 123720 144000 123772 144006
rect 123720 143942 123772 143948
rect 123180 140934 123760 140962
rect 123732 140826 123760 140934
rect 124468 140826 124496 144010
rect 124548 144000 124600 144006
rect 124548 143942 124600 143948
rect 124560 141098 124588 143942
rect 124652 143682 124680 151286
rect 125112 144006 125140 151422
rect 125296 151078 125324 153868
rect 125664 151350 125692 153868
rect 143250 153854 143724 153882
rect 129240 152364 129292 152370
rect 129240 152306 129292 152312
rect 128780 152296 128832 152302
rect 128780 152238 128832 152244
rect 127952 152228 128004 152234
rect 127952 152170 128004 152176
rect 127308 151956 127360 151962
rect 127308 151898 127360 151904
rect 127216 151888 127268 151894
rect 127216 151830 127268 151836
rect 125652 151344 125704 151350
rect 125652 151286 125704 151292
rect 125284 151072 125336 151078
rect 125284 151014 125336 151020
rect 125192 151004 125244 151010
rect 125192 150946 125244 150952
rect 125204 144074 125232 150946
rect 127228 146182 127256 151830
rect 127216 146176 127268 146182
rect 127216 146118 127268 146124
rect 125192 144068 125244 144074
rect 125192 144010 125244 144016
rect 126020 144068 126072 144074
rect 126020 144010 126072 144016
rect 125100 144000 125152 144006
rect 125100 143942 125152 143948
rect 124652 143654 125416 143682
rect 124560 141070 124772 141098
rect 121984 140798 122274 140826
rect 122444 140798 122826 140826
rect 123088 140798 123470 140826
rect 123732 140798 124022 140826
rect 124468 140798 124574 140826
rect 112416 140662 112982 140690
rect 117582 140662 117688 140690
rect 121722 140662 121828 140690
rect 124744 140690 124772 141070
rect 125388 140826 125416 143654
rect 126032 140826 126060 144010
rect 126572 144000 126624 144006
rect 126572 143942 126624 143948
rect 126584 140826 126612 143942
rect 127320 140826 127348 151898
rect 127860 151548 127912 151554
rect 127860 151490 127912 151496
rect 127676 146176 127728 146182
rect 127676 146118 127728 146124
rect 127688 140826 127716 146118
rect 127872 144006 127900 151490
rect 127964 144074 127992 152170
rect 127952 144068 128004 144074
rect 127952 144010 128004 144016
rect 128596 144068 128648 144074
rect 128596 144010 128648 144016
rect 127860 144000 127912 144006
rect 127860 143942 127912 143948
rect 128608 140826 128636 144010
rect 128688 144000 128740 144006
rect 128688 143942 128740 143948
rect 128700 141098 128728 143942
rect 128792 143682 128820 152238
rect 129252 144074 129280 152306
rect 131356 151344 131408 151350
rect 131356 151286 131408 151292
rect 129332 151072 129384 151078
rect 129332 151014 129384 151020
rect 129240 144068 129292 144074
rect 129240 144010 129292 144016
rect 129344 144006 129372 151014
rect 130068 144068 130120 144074
rect 130068 144010 130120 144016
rect 129332 144000 129384 144006
rect 129332 143942 129384 143948
rect 128792 143654 129464 143682
rect 128700 141070 128820 141098
rect 125388 140798 125770 140826
rect 126032 140798 126322 140826
rect 126584 140798 126966 140826
rect 127320 140798 127518 140826
rect 127688 140798 128070 140826
rect 128608 140798 128714 140826
rect 128792 140690 128820 141070
rect 129436 140826 129464 143654
rect 130080 140826 130108 144010
rect 130620 144000 130672 144006
rect 130620 143942 130672 143948
rect 130632 140826 130660 143942
rect 131368 140826 131396 151286
rect 129436 140798 129818 140826
rect 130080 140798 130462 140826
rect 130632 140798 131014 140826
rect 131368 140798 131566 140826
rect 124744 140662 125218 140690
rect 128792 140662 129266 140690
rect 134850 140568 134906 140577
rect 134850 140503 134906 140512
rect 100810 140160 100866 140169
rect 100810 140095 100866 140104
rect 100824 138566 100852 140095
rect 134864 140062 134892 140503
rect 134852 140056 134904 140062
rect 100902 140024 100958 140033
rect 143592 140056 143644 140062
rect 134852 139998 134904 140004
rect 135402 140024 135458 140033
rect 100902 139959 100958 139968
rect 143592 139998 143644 140004
rect 135402 139959 135404 139968
rect 100812 138560 100864 138566
rect 100812 138502 100864 138508
rect 100916 138498 100944 139959
rect 135456 139959 135458 139968
rect 143316 139988 143368 139994
rect 135404 139930 135456 139936
rect 143316 139930 143368 139936
rect 134666 139480 134722 139489
rect 134666 139415 134722 139424
rect 101178 138936 101234 138945
rect 101178 138871 101234 138880
rect 101086 138664 101142 138673
rect 101086 138599 101142 138608
rect 100904 138492 100956 138498
rect 100904 138434 100956 138440
rect 100994 137848 101050 137857
rect 100994 137783 101050 137792
rect 101008 137342 101036 137783
rect 100996 137336 101048 137342
rect 100996 137278 101048 137284
rect 101100 137070 101128 138599
rect 101192 137138 101220 138871
rect 134680 138634 134708 139415
rect 135402 138800 135458 138809
rect 135402 138735 135404 138744
rect 135456 138735 135458 138744
rect 139820 138764 139872 138770
rect 135404 138706 135456 138712
rect 139820 138706 139872 138712
rect 134668 138628 134720 138634
rect 134668 138570 134720 138576
rect 139636 138628 139688 138634
rect 139636 138570 139688 138576
rect 134666 138256 134722 138265
rect 134666 138191 134722 138200
rect 134680 137410 134708 138191
rect 135402 137712 135458 137721
rect 135402 137647 135458 137656
rect 134668 137404 134720 137410
rect 134668 137346 134720 137352
rect 101270 137304 101326 137313
rect 101270 137239 101272 137248
rect 101324 137239 101326 137248
rect 101272 137210 101324 137216
rect 135416 137206 135444 137647
rect 135404 137200 135456 137206
rect 135404 137142 135456 137148
rect 101180 137132 101232 137138
rect 101180 137074 101232 137080
rect 139648 137070 139676 138570
rect 139728 137404 139780 137410
rect 139728 137346 139780 137352
rect 101088 137064 101140 137070
rect 139636 137064 139688 137070
rect 101088 137006 101140 137012
rect 135034 137032 135090 137041
rect 139636 137006 139688 137012
rect 135034 136967 135090 136976
rect 101822 136624 101878 136633
rect 101822 136559 101878 136568
rect 101454 136216 101510 136225
rect 101454 136151 101510 136160
rect 101468 135914 101496 136151
rect 101730 135944 101786 135953
rect 101456 135908 101508 135914
rect 101730 135879 101786 135888
rect 101456 135850 101508 135856
rect 101744 135846 101772 135879
rect 101732 135840 101784 135846
rect 101732 135782 101784 135788
rect 101836 135778 101864 136559
rect 135048 135982 135076 136967
rect 139740 136662 139768 137346
rect 139832 137002 139860 138706
rect 143328 138265 143356 139930
rect 143604 138537 143632 139998
rect 143590 138528 143646 138537
rect 143590 138463 143646 138472
rect 143314 138256 143370 138265
rect 143314 138191 143370 138200
rect 143408 137200 143460 137206
rect 143408 137142 143460 137148
rect 143590 137168 143646 137177
rect 139820 136996 139872 137002
rect 139820 136938 139872 136944
rect 143132 136996 143184 137002
rect 143132 136938 143184 136944
rect 143144 136905 143172 136938
rect 143130 136896 143186 136905
rect 143130 136831 143186 136840
rect 139728 136656 139780 136662
rect 139728 136598 139780 136604
rect 135310 136488 135366 136497
rect 135310 136423 135366 136432
rect 135036 135976 135088 135982
rect 135036 135918 135088 135924
rect 135324 135914 135352 136423
rect 143316 135976 143368 135982
rect 135402 135944 135458 135953
rect 135312 135908 135364 135914
rect 143316 135918 143368 135924
rect 135402 135879 135458 135888
rect 135312 135850 135364 135856
rect 135416 135846 135444 135879
rect 135404 135840 135456 135846
rect 135404 135782 135456 135788
rect 143224 135840 143276 135846
rect 143224 135782 143276 135788
rect 101824 135772 101876 135778
rect 101824 135714 101876 135720
rect 134850 135400 134906 135409
rect 134850 135335 134906 135344
rect 101454 134856 101510 134865
rect 101454 134791 101510 134800
rect 100902 134448 100958 134457
rect 101468 134418 101496 134791
rect 134666 134720 134722 134729
rect 134666 134655 134722 134664
rect 134680 134622 134708 134655
rect 134668 134616 134720 134622
rect 134668 134558 134720 134564
rect 134864 134554 134892 135335
rect 136876 134616 136928 134622
rect 136876 134558 136928 134564
rect 134852 134548 134904 134554
rect 134852 134490 134904 134496
rect 100902 134383 100958 134392
rect 101456 134412 101508 134418
rect 100916 132922 100944 134383
rect 101456 134354 101508 134360
rect 135402 134176 135458 134185
rect 135402 134111 135458 134120
rect 101822 133768 101878 133777
rect 101822 133703 101878 133712
rect 101730 133088 101786 133097
rect 101730 133023 101786 133032
rect 100904 132916 100956 132922
rect 100904 132858 100956 132864
rect 101178 132000 101234 132009
rect 101178 131935 101234 131944
rect 101192 130270 101220 131935
rect 101546 131864 101602 131873
rect 101546 131799 101602 131808
rect 101362 130368 101418 130377
rect 101362 130303 101418 130312
rect 101180 130264 101232 130270
rect 101180 130206 101232 130212
rect 101270 129008 101326 129017
rect 101270 128943 101326 128952
rect 100994 128464 101050 128473
rect 100994 128399 101050 128408
rect 101008 127482 101036 128399
rect 101178 127920 101234 127929
rect 101178 127855 101234 127864
rect 101086 127784 101142 127793
rect 101086 127719 101142 127728
rect 100996 127476 101048 127482
rect 100996 127418 101048 127424
rect 101100 126122 101128 127719
rect 101088 126116 101140 126122
rect 101088 126058 101140 126064
rect 101192 126054 101220 127855
rect 101284 127414 101312 128943
rect 101376 128842 101404 130303
rect 101560 130202 101588 131799
rect 101744 131630 101772 133023
rect 101836 132990 101864 133703
rect 134114 133632 134170 133641
rect 134114 133567 134170 133576
rect 134128 133126 134156 133567
rect 134116 133120 134168 133126
rect 134116 133062 134168 133068
rect 135416 133058 135444 134111
rect 135404 133052 135456 133058
rect 135404 132994 135456 133000
rect 101824 132984 101876 132990
rect 101824 132926 101876 132932
rect 135126 132952 135182 132961
rect 135126 132887 135182 132896
rect 101822 132544 101878 132553
rect 101822 132479 101878 132488
rect 101732 131624 101784 131630
rect 101732 131566 101784 131572
rect 101836 131562 101864 132479
rect 134482 132408 134538 132417
rect 134482 132343 134538 132352
rect 134496 131970 134524 132343
rect 134484 131964 134536 131970
rect 134484 131906 134536 131912
rect 135140 131698 135168 132887
rect 136888 132854 136916 134558
rect 139636 134548 139688 134554
rect 139636 134490 139688 134496
rect 139648 133806 139676 134490
rect 143236 134049 143264 135782
rect 143328 135273 143356 135918
rect 143420 135817 143448 137142
rect 143590 137103 143646 137112
rect 143604 137070 143632 137103
rect 143592 137064 143644 137070
rect 143592 137006 143644 137012
rect 143500 136656 143552 136662
rect 143500 136598 143552 136604
rect 143512 136361 143540 136598
rect 143498 136352 143554 136361
rect 143498 136287 143554 136296
rect 143592 135908 143644 135914
rect 143592 135850 143644 135856
rect 143406 135808 143462 135817
rect 143406 135743 143462 135752
rect 143314 135264 143370 135273
rect 143314 135199 143370 135208
rect 143604 134321 143632 135850
rect 143590 134312 143646 134321
rect 143590 134247 143646 134256
rect 143222 134040 143278 134049
rect 143222 133975 143278 133984
rect 139636 133800 139688 133806
rect 139636 133742 139688 133748
rect 142948 133800 143000 133806
rect 142948 133742 143000 133748
rect 142960 133369 142988 133742
rect 142946 133360 143002 133369
rect 142946 133295 143002 133304
rect 138164 133120 138216 133126
rect 138164 133062 138216 133068
rect 136876 132848 136928 132854
rect 136876 132790 136928 132796
rect 137152 131964 137204 131970
rect 137152 131906 137204 131912
rect 135310 131864 135366 131873
rect 135310 131799 135366 131808
rect 135324 131766 135352 131799
rect 135312 131760 135364 131766
rect 135312 131702 135364 131708
rect 135128 131692 135180 131698
rect 135128 131634 135180 131640
rect 101824 131556 101876 131562
rect 101824 131498 101876 131504
rect 134850 131320 134906 131329
rect 134850 131255 134906 131264
rect 101822 130776 101878 130785
rect 101822 130711 101878 130720
rect 101548 130196 101600 130202
rect 101548 130138 101600 130144
rect 101730 129688 101786 129697
rect 101730 129623 101786 129632
rect 101364 128836 101416 128842
rect 101364 128778 101416 128784
rect 101744 128774 101772 129623
rect 101836 128910 101864 130711
rect 134666 130640 134722 130649
rect 134666 130575 134668 130584
rect 134720 130575 134722 130584
rect 134668 130546 134720 130552
rect 134864 130338 134892 131255
rect 134852 130332 134904 130338
rect 134852 130274 134904 130280
rect 137164 130270 137192 131906
rect 137980 131760 138032 131766
rect 137980 131702 138032 131708
rect 137612 130604 137664 130610
rect 137612 130546 137664 130552
rect 137428 130332 137480 130338
rect 137428 130274 137480 130280
rect 137152 130264 137204 130270
rect 137152 130206 137204 130212
rect 135402 130096 135458 130105
rect 135402 130031 135458 130040
rect 134666 129552 134722 129561
rect 134666 129487 134722 129496
rect 134680 129386 134708 129487
rect 134668 129380 134720 129386
rect 134668 129322 134720 129328
rect 135416 128978 135444 130031
rect 135404 128972 135456 128978
rect 135404 128914 135456 128920
rect 101824 128904 101876 128910
rect 101824 128846 101876 128852
rect 135402 128872 135458 128881
rect 137440 128842 137468 130274
rect 137520 129380 137572 129386
rect 137520 129322 137572 129328
rect 135402 128807 135458 128816
rect 137428 128836 137480 128842
rect 101732 128768 101784 128774
rect 101732 128710 101784 128716
rect 134666 128328 134722 128337
rect 134666 128263 134722 128272
rect 134680 127890 134708 128263
rect 134668 127884 134720 127890
rect 134668 127826 134720 127832
rect 134666 127784 134722 127793
rect 134666 127719 134668 127728
rect 134720 127719 134722 127728
rect 134668 127690 134720 127696
rect 135416 127550 135444 128807
rect 137428 128778 137480 128784
rect 136876 127748 136928 127754
rect 136876 127690 136928 127696
rect 135404 127544 135456 127550
rect 135404 127486 135456 127492
rect 101272 127408 101324 127414
rect 101272 127350 101324 127356
rect 135402 127240 135458 127249
rect 135458 127198 135628 127226
rect 135402 127175 135458 127184
rect 101822 126696 101878 126705
rect 101822 126631 101878 126640
rect 101730 126288 101786 126297
rect 101836 126258 101864 126631
rect 135402 126560 135458 126569
rect 135458 126518 135536 126546
rect 135402 126495 135458 126504
rect 101730 126223 101786 126232
rect 101824 126252 101876 126258
rect 101744 126190 101772 126223
rect 101824 126194 101876 126200
rect 101732 126184 101784 126190
rect 101732 126126 101784 126132
rect 101180 126048 101232 126054
rect 101180 125990 101232 125996
rect 135218 126016 135274 126025
rect 135218 125951 135274 125960
rect 101454 125608 101510 125617
rect 101454 125543 101510 125552
rect 101468 124762 101496 125543
rect 135034 125472 135090 125481
rect 135034 125407 135090 125416
rect 135048 125306 135076 125407
rect 135036 125300 135088 125306
rect 135036 125242 135088 125248
rect 101638 124928 101694 124937
rect 101638 124863 101694 124872
rect 101456 124756 101508 124762
rect 101456 124698 101508 124704
rect 101652 123334 101680 124863
rect 135232 124830 135260 125951
rect 135404 124892 135456 124898
rect 135404 124834 135456 124840
rect 135220 124824 135272 124830
rect 101730 124792 101786 124801
rect 135416 124801 135444 124834
rect 135220 124766 135272 124772
rect 135402 124792 135458 124801
rect 101730 124727 101786 124736
rect 135402 124727 135458 124736
rect 101640 123328 101692 123334
rect 101640 123270 101692 123276
rect 101744 123266 101772 124727
rect 135508 124422 135536 126518
rect 135600 124762 135628 127198
rect 136888 126054 136916 127690
rect 137532 127414 137560 129322
rect 137624 128774 137652 130546
rect 137992 130202 138020 131702
rect 138176 131562 138204 133062
rect 143224 132984 143276 132990
rect 143224 132926 143276 132932
rect 143236 132281 143264 132926
rect 143592 132848 143644 132854
rect 143590 132816 143592 132825
rect 143644 132816 143646 132825
rect 143590 132751 143646 132760
rect 143222 132272 143278 132281
rect 143222 132207 143278 132216
rect 142488 131624 142540 131630
rect 142488 131566 142540 131572
rect 138164 131556 138216 131562
rect 138164 131498 138216 131504
rect 142500 131057 142528 131566
rect 143592 131556 143644 131562
rect 143592 131498 143644 131504
rect 143604 131465 143632 131498
rect 143590 131456 143646 131465
rect 143590 131391 143646 131400
rect 142486 131048 142542 131057
rect 142486 130983 142542 130992
rect 143592 130264 143644 130270
rect 143590 130232 143592 130241
rect 143644 130232 143646 130241
rect 137980 130196 138032 130202
rect 137980 130138 138032 130144
rect 143040 130196 143092 130202
rect 143590 130167 143646 130176
rect 143040 130138 143092 130144
rect 143052 129969 143080 130138
rect 143038 129960 143094 129969
rect 143038 129895 143094 129904
rect 143132 128904 143184 128910
rect 142762 128872 142818 128881
rect 143132 128846 143184 128852
rect 142762 128807 142764 128816
rect 142816 128807 142818 128816
rect 142764 128778 142816 128784
rect 137612 128768 137664 128774
rect 137612 128710 137664 128716
rect 143144 128065 143172 128846
rect 143592 128768 143644 128774
rect 143590 128736 143592 128745
rect 143644 128736 143646 128745
rect 143590 128671 143646 128680
rect 143130 128056 143186 128065
rect 143130 127991 143186 128000
rect 137612 127884 137664 127890
rect 137612 127826 137664 127832
rect 137520 127408 137572 127414
rect 137520 127350 137572 127356
rect 137624 126122 137652 127826
rect 143316 127476 143368 127482
rect 143316 127418 143368 127424
rect 142488 127408 142540 127414
rect 142486 127376 142488 127385
rect 142540 127376 142542 127385
rect 142486 127311 142542 127320
rect 143328 126977 143356 127418
rect 143314 126968 143370 126977
rect 143314 126903 143370 126912
rect 137612 126116 137664 126122
rect 137612 126058 137664 126064
rect 143592 126116 143644 126122
rect 143592 126058 143644 126064
rect 136876 126048 136928 126054
rect 136876 125990 136928 125996
rect 143040 126048 143092 126054
rect 143604 126025 143632 126058
rect 143040 125990 143092 125996
rect 143590 126016 143646 126025
rect 143052 125753 143080 125990
rect 143590 125951 143646 125960
rect 143038 125744 143094 125753
rect 143038 125679 143094 125688
rect 137612 125300 137664 125306
rect 137612 125242 137664 125248
rect 136876 124892 136928 124898
rect 136876 124834 136928 124840
rect 135588 124756 135640 124762
rect 135588 124698 135640 124704
rect 135496 124416 135548 124422
rect 135496 124358 135548 124364
rect 134114 124248 134170 124257
rect 134114 124183 134170 124192
rect 101914 123840 101970 123849
rect 101914 123775 101970 123784
rect 101822 123432 101878 123441
rect 101822 123367 101878 123376
rect 101732 123260 101784 123266
rect 101732 123202 101784 123208
rect 101638 122616 101694 122625
rect 101638 122551 101694 122560
rect 101454 122072 101510 122081
rect 101454 122007 101510 122016
rect 101086 121120 101142 121129
rect 101086 121055 101142 121064
rect 101100 120750 101128 121055
rect 101088 120744 101140 120750
rect 101088 120686 101140 120692
rect 101468 120546 101496 122007
rect 101546 120712 101602 120721
rect 101546 120647 101548 120656
rect 101600 120647 101602 120656
rect 101548 120618 101600 120624
rect 101652 120614 101680 122551
rect 101836 121974 101864 123367
rect 101824 121968 101876 121974
rect 101824 121910 101876 121916
rect 101928 121906 101956 123775
rect 134128 123402 134156 124183
rect 134482 123704 134538 123713
rect 134482 123639 134538 123648
rect 134496 123538 134524 123639
rect 134484 123532 134536 123538
rect 134484 123474 134536 123480
rect 134116 123396 134168 123402
rect 134116 123338 134168 123344
rect 134482 123024 134538 123033
rect 134482 122959 134538 122968
rect 134496 122450 134524 122959
rect 136888 122926 136916 124834
rect 137624 123334 137652 125242
rect 142764 124824 142816 124830
rect 142764 124766 142816 124772
rect 142488 124416 142540 124422
rect 142486 124384 142488 124393
rect 142540 124384 142542 124393
rect 142486 124319 142542 124328
rect 142776 123985 142804 124766
rect 143592 124756 143644 124762
rect 143592 124698 143644 124704
rect 143604 124665 143632 124698
rect 143590 124656 143646 124665
rect 143590 124591 143646 124600
rect 142762 123976 142818 123985
rect 142762 123911 142818 123920
rect 137704 123532 137756 123538
rect 137704 123474 137756 123480
rect 137612 123328 137664 123334
rect 137612 123270 137664 123276
rect 136876 122920 136928 122926
rect 136876 122862 136928 122868
rect 134942 122480 134998 122489
rect 134484 122444 134536 122450
rect 134942 122415 134998 122424
rect 134484 122386 134536 122392
rect 134956 122314 134984 122415
rect 134944 122308 134996 122314
rect 134944 122250 134996 122256
rect 137244 122308 137296 122314
rect 137244 122250 137296 122256
rect 134482 121936 134538 121945
rect 101916 121900 101968 121906
rect 134482 121871 134538 121880
rect 101916 121842 101968 121848
rect 101730 121528 101786 121537
rect 101730 121463 101786 121472
rect 101744 120818 101772 121463
rect 134496 120818 134524 121871
rect 134666 121392 134722 121401
rect 134666 121327 134722 121336
rect 101732 120812 101784 120818
rect 101732 120754 101784 120760
rect 134484 120812 134536 120818
rect 134484 120754 134536 120760
rect 134680 120750 134708 121327
rect 134668 120744 134720 120750
rect 134668 120686 134720 120692
rect 135402 120712 135458 120721
rect 135402 120647 135404 120656
rect 135456 120647 135458 120656
rect 136876 120676 136928 120682
rect 135404 120618 135456 120624
rect 136876 120618 136928 120624
rect 101640 120608 101692 120614
rect 101640 120550 101692 120556
rect 101456 120540 101508 120546
rect 101456 120482 101508 120488
rect 134482 120168 134538 120177
rect 134482 120103 134538 120112
rect 101270 119760 101326 119769
rect 101270 119695 101326 119704
rect 101284 119390 101312 119695
rect 101272 119384 101324 119390
rect 101272 119326 101324 119332
rect 101362 119352 101418 119361
rect 134496 119322 134524 120103
rect 135402 119624 135458 119633
rect 135402 119559 135404 119568
rect 135456 119559 135458 119568
rect 135404 119530 135456 119536
rect 101362 119287 101364 119296
rect 101416 119287 101418 119296
rect 134484 119316 134536 119322
rect 101364 119258 101416 119264
rect 134484 119258 134536 119264
rect 136888 119186 136916 120618
rect 137256 120546 137284 122250
rect 137716 121974 137744 123474
rect 138164 123396 138216 123402
rect 138164 123338 138216 123344
rect 138072 122444 138124 122450
rect 138072 122386 138124 122392
rect 137704 121968 137756 121974
rect 137704 121910 137756 121916
rect 137428 120812 137480 120818
rect 137428 120754 137480 120760
rect 137244 120540 137296 120546
rect 137244 120482 137296 120488
rect 136968 119316 137020 119322
rect 136968 119258 137020 119264
rect 136876 119180 136928 119186
rect 136876 119122 136928 119128
rect 134666 118944 134722 118953
rect 134666 118879 134722 118888
rect 101362 118536 101418 118545
rect 134680 118506 134708 118879
rect 101362 118471 101418 118480
rect 134668 118500 134720 118506
rect 101376 117962 101404 118471
rect 134668 118442 134720 118448
rect 136876 118500 136928 118506
rect 136876 118442 136928 118448
rect 134666 118400 134722 118409
rect 134666 118335 134722 118344
rect 134680 118234 134708 118335
rect 134668 118228 134720 118234
rect 134668 118170 134720 118176
rect 101730 118128 101786 118137
rect 101730 118063 101786 118072
rect 101364 117956 101416 117962
rect 101364 117898 101416 117904
rect 101744 117894 101772 118063
rect 101732 117888 101784 117894
rect 101732 117830 101784 117836
rect 134850 117856 134906 117865
rect 134850 117791 134906 117800
rect 101178 117448 101234 117457
rect 101178 117383 101234 117392
rect 101086 116768 101142 116777
rect 101086 116703 101142 116712
rect 100994 116632 101050 116641
rect 101100 116602 101128 116703
rect 100994 116567 101050 116576
rect 101088 116596 101140 116602
rect 101008 116534 101036 116567
rect 101088 116538 101140 116544
rect 100996 116528 101048 116534
rect 100996 116470 101048 116476
rect 101192 116466 101220 117383
rect 134758 116632 134814 116641
rect 134758 116567 134814 116576
rect 101180 116460 101232 116466
rect 101180 116402 101232 116408
rect 101086 115680 101142 115689
rect 101086 115615 101142 115624
rect 100994 115272 101050 115281
rect 101100 115242 101128 115615
rect 100994 115207 101050 115216
rect 101088 115236 101140 115242
rect 101008 115174 101036 115207
rect 101088 115178 101140 115184
rect 100996 115168 101048 115174
rect 100996 115110 101048 115116
rect 101822 114456 101878 114465
rect 101822 114391 101878 114400
rect 101638 113776 101694 113785
rect 101638 113711 101694 113720
rect 100994 112552 101050 112561
rect 100994 112487 101050 112496
rect 101008 112386 101036 112487
rect 100996 112380 101048 112386
rect 100996 112322 101048 112328
rect 99524 110476 99576 110482
rect 99524 110418 99576 110424
rect 99432 110340 99484 110346
rect 99432 110282 99484 110288
rect 99248 109864 99300 109870
rect 99248 109806 99300 109812
rect 99156 109796 99208 109802
rect 99156 109738 99208 109744
rect 99064 109728 99116 109734
rect 99064 109670 99116 109676
rect 98972 109660 99024 109666
rect 98972 109602 99024 109608
rect 98984 91209 99012 109602
rect 99076 92433 99104 109670
rect 99168 93657 99196 109738
rect 99260 95561 99288 109806
rect 99340 109592 99392 109598
rect 99340 109534 99392 109540
rect 99246 95552 99302 95561
rect 99246 95487 99302 95496
rect 99352 94337 99380 109534
rect 99444 97057 99472 110282
rect 99536 98553 99564 110418
rect 101652 101982 101680 113711
rect 101836 102118 101864 114391
rect 102006 113912 102062 113921
rect 102006 113847 102062 113856
rect 101824 102112 101876 102118
rect 101824 102054 101876 102060
rect 102020 102050 102048 113847
rect 104136 109666 104164 112932
rect 104596 109734 104624 112932
rect 105148 109802 105176 112932
rect 105136 109796 105188 109802
rect 105136 109738 105188 109744
rect 104584 109728 104636 109734
rect 104584 109670 104636 109676
rect 104124 109660 104176 109666
rect 104124 109602 104176 109608
rect 105700 109598 105728 112932
rect 106252 109870 106280 112932
rect 106804 110346 106832 112932
rect 107356 110482 107384 112932
rect 107344 110476 107396 110482
rect 107344 110418 107396 110424
rect 106792 110340 106844 110346
rect 106792 110282 106844 110288
rect 107908 110278 107936 112932
rect 108460 111201 108488 112932
rect 108446 111192 108502 111201
rect 108446 111127 108502 111136
rect 109012 110958 109040 112932
rect 109000 110952 109052 110958
rect 109000 110894 109052 110900
rect 109564 110890 109592 112932
rect 109552 110884 109604 110890
rect 109552 110826 109604 110832
rect 107896 110272 107948 110278
rect 107896 110214 107948 110220
rect 106240 109864 106292 109870
rect 106240 109806 106292 109812
rect 105688 109592 105740 109598
rect 105688 109534 105740 109540
rect 102008 102044 102060 102050
rect 102008 101986 102060 101992
rect 101640 101976 101692 101982
rect 101640 101918 101692 101924
rect 110116 99740 110144 112932
rect 110668 110634 110696 112932
rect 110576 110606 110696 110634
rect 110576 99754 110604 110606
rect 111220 99754 111248 112932
rect 111772 102662 111800 112932
rect 111300 102656 111352 102662
rect 111300 102598 111352 102604
rect 111760 102656 111812 102662
rect 111760 102598 111812 102604
rect 110498 99726 110604 99754
rect 110866 99726 111248 99754
rect 111312 99740 111340 102598
rect 112324 102594 112352 112932
rect 112496 102656 112548 102662
rect 112496 102598 112548 102604
rect 111668 102588 111720 102594
rect 111668 102530 111720 102536
rect 112312 102588 112364 102594
rect 112312 102530 112364 102536
rect 111680 99740 111708 102530
rect 112036 101976 112088 101982
rect 112036 101918 112088 101924
rect 112048 99740 112076 101918
rect 112508 99740 112536 102598
rect 112876 101982 112904 112932
rect 113428 110634 113456 112932
rect 113232 110612 113284 110618
rect 113232 110554 113284 110560
rect 113336 110606 113456 110634
rect 113140 110544 113192 110550
rect 113140 110486 113192 110492
rect 112864 101976 112916 101982
rect 112864 101918 112916 101924
rect 113152 99754 113180 110486
rect 112890 99726 113180 99754
rect 113244 99740 113272 110554
rect 113336 102662 113364 110606
rect 113980 110550 114008 112932
rect 114532 110618 114560 112932
rect 115084 110634 115112 112932
rect 114520 110612 114572 110618
rect 114520 110554 114572 110560
rect 114716 110606 115112 110634
rect 113968 110544 114020 110550
rect 113968 110486 114020 110492
rect 114612 110544 114664 110550
rect 114612 110486 114664 110492
rect 113324 102656 113376 102662
rect 113324 102598 113376 102604
rect 113692 102656 113744 102662
rect 113692 102598 113744 102604
rect 113704 99740 113732 102598
rect 114624 102526 114652 110486
rect 114716 102662 114744 110606
rect 115636 110550 115664 112932
rect 115808 110612 115860 110618
rect 115808 110554 115860 110560
rect 115624 110544 115676 110550
rect 115624 110486 115676 110492
rect 115716 109864 115768 109870
rect 115716 109806 115768 109812
rect 114704 102656 114756 102662
rect 114704 102598 114756 102604
rect 114060 102520 114112 102526
rect 114060 102462 114112 102468
rect 114612 102520 114664 102526
rect 114612 102462 114664 102468
rect 115256 102520 115308 102526
rect 115256 102462 115308 102468
rect 114072 99740 114100 102462
rect 114428 102384 114480 102390
rect 114428 102326 114480 102332
rect 114440 99740 114468 102326
rect 114888 102044 114940 102050
rect 114888 101986 114940 101992
rect 114900 99740 114928 101986
rect 115268 99740 115296 102462
rect 115728 99754 115756 109806
rect 115650 99726 115756 99754
rect 115820 99754 115848 110554
rect 115900 110544 115952 110550
rect 115900 110486 115952 110492
rect 115912 102050 115940 110486
rect 115992 110340 116044 110346
rect 115992 110282 116044 110288
rect 116004 102526 116032 110282
rect 115992 102520 116044 102526
rect 115992 102462 116044 102468
rect 116188 102390 116216 112932
rect 116740 110550 116768 112932
rect 116728 110544 116780 110550
rect 116728 110486 116780 110492
rect 117292 110346 117320 112932
rect 117464 110544 117516 110550
rect 117464 110486 117516 110492
rect 117280 110340 117332 110346
rect 117280 110282 117332 110288
rect 116176 102384 116228 102390
rect 116176 102326 116228 102332
rect 115900 102044 115952 102050
rect 115900 101986 115952 101992
rect 117476 101846 117504 110486
rect 117844 109870 117872 112932
rect 118304 110618 118332 112932
rect 118292 110612 118344 110618
rect 118292 110554 118344 110560
rect 118856 110550 118884 112932
rect 118844 110544 118896 110550
rect 118844 110486 118896 110492
rect 117832 109864 117884 109870
rect 117832 109806 117884 109812
rect 118936 109864 118988 109870
rect 118936 109806 118988 109812
rect 116452 101840 116504 101846
rect 116452 101782 116504 101788
rect 117464 101840 117516 101846
rect 117464 101782 117516 101788
rect 115820 99726 116110 99754
rect 116464 99740 116492 101782
rect 116820 101704 116872 101710
rect 116820 101646 116872 101652
rect 116832 99740 116860 101646
rect 117648 101636 117700 101642
rect 117648 101578 117700 101584
rect 117280 101432 117332 101438
rect 117280 101374 117332 101380
rect 117292 99740 117320 101374
rect 117660 99740 117688 101578
rect 118476 101568 118528 101574
rect 118476 101510 118528 101516
rect 118108 101364 118160 101370
rect 118108 101306 118160 101312
rect 118120 99740 118148 101306
rect 118488 99740 118516 101510
rect 118844 101500 118896 101506
rect 118844 101442 118896 101448
rect 118856 99740 118884 101442
rect 118948 101438 118976 109806
rect 119408 101710 119436 112932
rect 119960 109870 119988 112932
rect 119948 109864 120000 109870
rect 119948 109806 120000 109812
rect 119580 109796 119632 109802
rect 119580 109738 119632 109744
rect 119396 101704 119448 101710
rect 119396 101646 119448 101652
rect 118936 101432 118988 101438
rect 118936 101374 118988 101380
rect 119304 101432 119356 101438
rect 119304 101374 119356 101380
rect 119316 99740 119344 101374
rect 119592 101370 119620 109738
rect 119948 109728 120000 109734
rect 119948 109670 120000 109676
rect 119856 109660 119908 109666
rect 119856 109602 119908 109608
rect 119764 109592 119816 109598
rect 119764 109534 119816 109540
rect 119672 102588 119724 102594
rect 119672 102530 119724 102536
rect 119580 101364 119632 101370
rect 119580 101306 119632 101312
rect 119684 99740 119712 102530
rect 119776 101642 119804 109534
rect 119764 101636 119816 101642
rect 119764 101578 119816 101584
rect 119868 101574 119896 109602
rect 119856 101568 119908 101574
rect 119856 101510 119908 101516
rect 119960 101506 119988 109670
rect 120512 109598 120540 112932
rect 121064 109802 121092 112932
rect 121052 109796 121104 109802
rect 121052 109738 121104 109744
rect 121616 109666 121644 112932
rect 122168 109734 122196 112932
rect 122156 109728 122208 109734
rect 122156 109670 122208 109676
rect 121604 109660 121656 109666
rect 121604 109602 121656 109608
rect 122720 109598 122748 112932
rect 120500 109592 120552 109598
rect 120500 109534 120552 109540
rect 120960 109592 121012 109598
rect 120960 109534 121012 109540
rect 122708 109592 122760 109598
rect 122708 109534 122760 109540
rect 120868 102520 120920 102526
rect 120868 102462 120920 102468
rect 120040 102452 120092 102458
rect 120040 102394 120092 102400
rect 119948 101500 120000 101506
rect 119948 101442 120000 101448
rect 120052 99740 120080 102394
rect 120500 102180 120552 102186
rect 120500 102122 120552 102128
rect 120512 99740 120540 102122
rect 120880 99740 120908 102462
rect 120972 101438 121000 109534
rect 123272 102594 123300 112932
rect 123260 102588 123312 102594
rect 123260 102530 123312 102536
rect 123824 102458 123852 112932
rect 123812 102452 123864 102458
rect 123812 102394 123864 102400
rect 122432 102384 122484 102390
rect 122432 102326 122484 102332
rect 122064 102316 122116 102322
rect 122064 102258 122116 102264
rect 121696 102248 121748 102254
rect 121696 102190 121748 102196
rect 121236 101772 121288 101778
rect 121236 101714 121288 101720
rect 120960 101432 121012 101438
rect 120960 101374 121012 101380
rect 121248 99740 121276 101714
rect 121708 99740 121736 102190
rect 122076 99740 122104 102258
rect 122444 99740 122472 102326
rect 124376 102186 124404 112932
rect 124928 102526 124956 112932
rect 124916 102520 124968 102526
rect 124916 102462 124968 102468
rect 124364 102180 124416 102186
rect 124364 102122 124416 102128
rect 122892 102112 122944 102118
rect 122892 102054 122944 102060
rect 122904 99740 122932 102054
rect 124456 101840 124508 101846
rect 124456 101782 124508 101788
rect 123260 101704 123312 101710
rect 123260 101646 123312 101652
rect 123272 99740 123300 101646
rect 123628 101568 123680 101574
rect 123628 101510 123680 101516
rect 123640 99740 123668 101510
rect 124088 101500 124140 101506
rect 124088 101442 124140 101448
rect 124100 99740 124128 101442
rect 124468 99740 124496 101782
rect 125480 101778 125508 112932
rect 126032 102254 126060 112932
rect 126584 109818 126612 112932
rect 126124 109790 126612 109818
rect 126664 109796 126716 109802
rect 126124 102322 126152 109790
rect 126664 109738 126716 109744
rect 126480 109660 126532 109666
rect 126480 109602 126532 109608
rect 126112 102316 126164 102322
rect 126112 102258 126164 102264
rect 126020 102248 126072 102254
rect 126020 102190 126072 102196
rect 125468 101772 125520 101778
rect 125468 101714 125520 101720
rect 124824 101636 124876 101642
rect 124824 101578 124876 101584
rect 124836 99740 124864 101578
rect 126492 101574 126520 109602
rect 126572 109592 126624 109598
rect 126572 109534 126624 109540
rect 126584 101710 126612 109534
rect 126572 101704 126624 101710
rect 126572 101646 126624 101652
rect 126480 101568 126532 101574
rect 126480 101510 126532 101516
rect 126676 101506 126704 109738
rect 127136 102390 127164 112932
rect 127124 102384 127176 102390
rect 127124 102326 127176 102332
rect 127688 102118 127716 112932
rect 128240 109598 128268 112932
rect 128792 109666 128820 112932
rect 129344 109802 129372 112932
rect 129332 109796 129384 109802
rect 129332 109738 129384 109744
rect 128780 109660 128832 109666
rect 128780 109602 128832 109608
rect 129332 109660 129384 109666
rect 129332 109602 129384 109608
rect 128228 109592 128280 109598
rect 128228 109534 128280 109540
rect 129240 109592 129292 109598
rect 129240 109534 129292 109540
rect 127676 102112 127728 102118
rect 127676 102054 127728 102060
rect 129252 101642 129280 109534
rect 129240 101636 129292 101642
rect 129240 101578 129292 101584
rect 126664 101500 126716 101506
rect 126664 101442 126716 101448
rect 125652 101432 125704 101438
rect 125652 101374 125704 101380
rect 125284 101364 125336 101370
rect 125284 101306 125336 101312
rect 125296 99740 125324 101306
rect 125664 99740 125692 101374
rect 129344 101370 129372 109602
rect 129896 101846 129924 112932
rect 129976 111632 130028 111638
rect 129976 111574 130028 111580
rect 129988 110958 130016 111574
rect 129976 110952 130028 110958
rect 129976 110894 130028 110900
rect 130448 109598 130476 112932
rect 131000 109666 131028 112932
rect 130988 109660 131040 109666
rect 130988 109602 131040 109608
rect 130436 109592 130488 109598
rect 130436 109534 130488 109540
rect 129884 101840 129936 101846
rect 129884 101782 129936 101788
rect 131552 101438 131580 112932
rect 134024 111700 134076 111706
rect 134024 111642 134076 111648
rect 134036 111201 134064 111642
rect 134022 111192 134078 111201
rect 134022 111127 134078 111136
rect 131540 101432 131592 101438
rect 131540 101374 131592 101380
rect 129332 101364 129384 101370
rect 129332 101306 129384 101312
rect 99522 98544 99578 98553
rect 99522 98479 99578 98488
rect 106790 98544 106846 98553
rect 106790 98479 106846 98488
rect 106804 97222 106832 98479
rect 106792 97216 106844 97222
rect 106792 97158 106844 97164
rect 99430 97048 99486 97057
rect 99430 96983 99486 96992
rect 106790 96232 106846 96241
rect 106790 96167 106846 96176
rect 106804 95862 106832 96167
rect 99524 95856 99576 95862
rect 99524 95798 99576 95804
rect 106792 95856 106844 95862
rect 106792 95798 106844 95804
rect 99338 94328 99394 94337
rect 99338 94263 99394 94272
rect 99154 93648 99210 93657
rect 99154 93583 99210 93592
rect 99062 92424 99118 92433
rect 99062 92359 99118 92368
rect 98970 91200 99026 91209
rect 98970 91135 99026 91144
rect 99536 88761 99564 95798
rect 106514 93920 106570 93929
rect 106514 93855 106570 93864
rect 106528 93074 106556 93855
rect 106516 93068 106568 93074
rect 106516 93010 106568 93016
rect 106790 91472 106846 91481
rect 106790 91407 106846 91416
rect 106804 90286 106832 91407
rect 105044 90280 105096 90286
rect 105044 90222 105096 90228
rect 106792 90280 106844 90286
rect 106792 90222 106844 90228
rect 104952 88920 105004 88926
rect 104952 88862 105004 88868
rect 99522 88752 99578 88761
rect 99522 88687 99578 88696
rect 99522 85352 99578 85361
rect 99522 85287 99578 85296
rect 99536 85254 99564 85287
rect 99524 85248 99576 85254
rect 99524 85190 99576 85196
rect 99432 84704 99484 84710
rect 99432 84646 99484 84652
rect 99522 84672 99578 84681
rect 99444 84001 99472 84646
rect 99522 84607 99578 84616
rect 99536 84506 99564 84607
rect 104964 84506 104992 88862
rect 105056 85254 105084 90222
rect 128502 89840 128558 89849
rect 128502 89775 128558 89784
rect 106790 89160 106846 89169
rect 106790 89095 106846 89104
rect 106804 88926 106832 89095
rect 128516 88926 128544 89775
rect 106792 88920 106844 88926
rect 106792 88862 106844 88868
rect 128504 88920 128556 88926
rect 128504 88862 128556 88868
rect 132000 88920 132052 88926
rect 132000 88862 132052 88868
rect 106790 86848 106846 86857
rect 106790 86783 106846 86792
rect 105044 85248 105096 85254
rect 105044 85190 105096 85196
rect 106804 84710 106832 86783
rect 106792 84704 106844 84710
rect 106792 84646 106844 84652
rect 99524 84500 99576 84506
rect 99524 84442 99576 84448
rect 104952 84500 105004 84506
rect 104952 84442 105004 84448
rect 107802 84400 107858 84409
rect 107802 84335 107858 84344
rect 99430 83992 99486 84001
rect 99430 83927 99486 83936
rect 107816 83350 107844 84335
rect 99524 83344 99576 83350
rect 99524 83286 99576 83292
rect 107804 83344 107856 83350
rect 107804 83286 107856 83292
rect 99536 82777 99564 83286
rect 99522 82768 99578 82777
rect 99522 82703 99578 82712
rect 106792 82120 106844 82126
rect 106790 82088 106792 82097
rect 106844 82088 106846 82097
rect 106790 82023 106846 82032
rect 99524 81984 99576 81990
rect 99524 81926 99576 81932
rect 99536 81553 99564 81926
rect 99522 81544 99578 81553
rect 99522 81479 99578 81488
rect 132012 80562 132040 88862
rect 132000 80556 132052 80562
rect 132000 80498 132052 80504
rect 99524 79876 99576 79882
rect 99524 79818 99576 79824
rect 106792 79876 106844 79882
rect 106792 79818 106844 79824
rect 99536 79785 99564 79818
rect 106804 79785 106832 79818
rect 99522 79776 99578 79785
rect 99522 79711 99578 79720
rect 106790 79776 106846 79785
rect 106790 79711 106846 79720
rect 99522 78008 99578 78017
rect 99522 77943 99578 77952
rect 99536 77910 99564 77943
rect 99524 77904 99576 77910
rect 99524 77846 99576 77852
rect 106516 77904 106568 77910
rect 106516 77846 106568 77852
rect 106528 77473 106556 77846
rect 106514 77464 106570 77473
rect 106514 77399 106570 77408
rect 99522 76784 99578 76793
rect 99522 76719 99578 76728
rect 99536 76482 99564 76719
rect 99524 76476 99576 76482
rect 99524 76418 99576 76424
rect 100996 76476 101048 76482
rect 100996 76418 101048 76424
rect 101008 75054 101036 76418
rect 100996 75048 101048 75054
rect 106792 75048 106844 75054
rect 100996 74990 101048 74996
rect 106790 75016 106792 75025
rect 106844 75016 106846 75025
rect 106790 74951 106846 74960
rect 100996 74912 101048 74918
rect 100996 74854 101048 74860
rect 99430 74336 99486 74345
rect 99430 74271 99486 74280
rect 99444 73762 99472 74271
rect 99524 73824 99576 73830
rect 99522 73792 99524 73801
rect 99576 73792 99578 73801
rect 99432 73756 99484 73762
rect 99522 73727 99578 73736
rect 99432 73698 99484 73704
rect 101008 73694 101036 74854
rect 105136 73824 105188 73830
rect 105136 73766 105188 73772
rect 100996 73688 101048 73694
rect 100996 73630 101048 73636
rect 99522 72568 99578 72577
rect 99522 72503 99578 72512
rect 99536 72402 99564 72503
rect 99524 72396 99576 72402
rect 99524 72338 99576 72344
rect 99522 71072 99578 71081
rect 99522 71007 99524 71016
rect 99576 71007 99578 71016
rect 104492 71036 104544 71042
rect 99524 70978 99576 70984
rect 104492 70978 104544 70984
rect 99522 69848 99578 69857
rect 99522 69783 99578 69792
rect 99536 69614 99564 69783
rect 99524 69608 99576 69614
rect 99524 69550 99576 69556
rect 104400 69608 104452 69614
rect 104400 69550 104452 69556
rect 98970 68352 99026 68361
rect 98970 68287 99026 68296
rect 98880 58524 98932 58530
rect 98880 58466 98932 58472
rect 98788 55056 98840 55062
rect 98788 54998 98840 55004
rect 98984 49554 99012 68287
rect 99062 67128 99118 67137
rect 99062 67063 99118 67072
rect 99076 49622 99104 67063
rect 99154 65904 99210 65913
rect 99154 65839 99210 65848
rect 99168 49758 99196 65839
rect 99246 64680 99302 64689
rect 99246 64615 99302 64624
rect 99260 50030 99288 64615
rect 99338 63456 99394 63465
rect 99338 63391 99394 63400
rect 99248 50024 99300 50030
rect 99248 49966 99300 49972
rect 99352 49962 99380 63391
rect 99522 61552 99578 61561
rect 99522 61487 99578 61496
rect 99536 61318 99564 61487
rect 99524 61312 99576 61318
rect 99524 61254 99576 61260
rect 103020 61312 103072 61318
rect 103020 61254 103072 61260
rect 99522 60056 99578 60065
rect 99522 59991 99578 60000
rect 99536 59958 99564 59991
rect 99524 59952 99576 59958
rect 99524 59894 99576 59900
rect 100352 59952 100404 59958
rect 100352 59894 100404 59900
rect 99524 55056 99576 55062
rect 99524 54998 99576 55004
rect 99536 50098 99564 54998
rect 99524 50092 99576 50098
rect 99524 50034 99576 50040
rect 99340 49956 99392 49962
rect 99340 49898 99392 49904
rect 99156 49752 99208 49758
rect 99156 49694 99208 49700
rect 99064 49616 99116 49622
rect 99064 49558 99116 49564
rect 98972 49548 99024 49554
rect 98972 49490 99024 49496
rect 100260 49072 100312 49078
rect 100260 49014 100312 49020
rect 96120 48868 96172 48874
rect 96120 48810 96172 48816
rect 80754 46864 80810 46873
rect 80754 46799 80810 46808
rect 77810 46728 77866 46737
rect 77810 46663 77866 46672
rect 74866 46456 74922 46465
rect 74866 46391 74922 46400
rect 73394 46320 73450 46329
rect 73394 46255 73450 46264
rect 73408 44810 73436 46255
rect 74880 44810 74908 46391
rect 76338 46184 76394 46193
rect 76338 46119 76394 46128
rect 76352 44810 76380 46119
rect 77824 44810 77852 46663
rect 79282 46592 79338 46601
rect 79282 46527 79338 46536
rect 79296 44810 79324 46527
rect 80768 44810 80796 46799
rect 93360 46352 93412 46358
rect 85722 46320 85778 46329
rect 93360 46294 93412 46300
rect 85722 46255 85778 46264
rect 82964 46216 83016 46222
rect 82964 46158 83016 46164
rect 82976 44810 83004 46158
rect 84068 46148 84120 46154
rect 84068 46090 84120 46096
rect 59044 44788 59096 44794
rect 61356 44782 61692 44810
rect 62828 44782 63164 44810
rect 64300 44782 64636 44810
rect 65772 44782 66108 44810
rect 67336 44782 67672 44810
rect 68808 44782 69144 44810
rect 70556 44782 70616 44810
rect 73408 44782 73652 44810
rect 74880 44782 75124 44810
rect 76352 44782 76688 44810
rect 77824 44782 78160 44810
rect 79296 44782 79632 44810
rect 80768 44782 81104 44810
rect 82668 44782 83004 44810
rect 84080 44810 84108 46090
rect 85736 44810 85764 46255
rect 87102 46184 87158 46193
rect 87102 46119 87158 46128
rect 88944 46148 88996 46154
rect 84080 44782 84140 44810
rect 85612 44782 85764 44810
rect 59044 44730 59096 44736
rect 58950 44416 59006 44425
rect 58950 44351 59006 44360
rect 58214 43872 58270 43881
rect 58214 43807 58270 43816
rect 58216 43292 58268 43298
rect 58216 43234 58268 43240
rect 58228 42657 58256 43234
rect 58308 43224 58360 43230
rect 59056 43201 59084 44730
rect 87116 44674 87144 46119
rect 88944 46090 88996 46096
rect 88956 44810 88984 46090
rect 88648 44782 88984 44810
rect 92808 44720 92860 44726
rect 87116 44646 87176 44674
rect 92808 44662 92860 44668
rect 92716 44652 92768 44658
rect 92716 44594 92768 44600
rect 90120 44510 90456 44538
rect 58308 43166 58360 43172
rect 59042 43192 59098 43201
rect 58214 42648 58270 42657
rect 58214 42583 58270 42592
rect 56284 42476 56336 42482
rect 56284 42418 56336 42424
rect 56296 41666 56324 42418
rect 56652 42340 56704 42346
rect 56652 42282 56704 42288
rect 56664 41938 56692 42282
rect 58320 42113 58348 43166
rect 59042 43127 59098 43136
rect 58306 42104 58362 42113
rect 58306 42039 58362 42048
rect 58400 42000 58452 42006
rect 58400 41942 58452 41948
rect 56652 41932 56704 41938
rect 56652 41874 56704 41880
rect 58216 41932 58268 41938
rect 58216 41874 58268 41880
rect 56284 41660 56336 41666
rect 56284 41602 56336 41608
rect 58228 41433 58256 41874
rect 58308 41660 58360 41666
rect 58308 41602 58360 41608
rect 58214 41424 58270 41433
rect 58214 41359 58270 41368
rect 58320 40889 58348 41602
rect 58306 40880 58362 40889
rect 58306 40815 58362 40824
rect 56652 40708 56704 40714
rect 56652 40650 56704 40656
rect 56560 40640 56612 40646
rect 56560 40582 56612 40588
rect 56572 40170 56600 40582
rect 56560 40164 56612 40170
rect 56560 40106 56612 40112
rect 56664 39082 56692 40650
rect 58412 40209 58440 41942
rect 58398 40200 58454 40209
rect 58216 40164 58268 40170
rect 58398 40135 58454 40144
rect 58216 40106 58268 40112
rect 58228 39665 58256 40106
rect 58214 39656 58270 39665
rect 58214 39591 58270 39600
rect 56744 39280 56796 39286
rect 56744 39222 56796 39228
rect 56652 39076 56704 39082
rect 56652 39018 56704 39024
rect 56756 38674 56784 39222
rect 58306 39112 58362 39121
rect 58306 39047 58308 39056
rect 58360 39047 58362 39056
rect 58308 39018 58360 39024
rect 58216 39008 58268 39014
rect 58216 38950 58268 38956
rect 56744 38668 56796 38674
rect 56744 38610 56796 38616
rect 58228 38441 58256 38950
rect 58400 38668 58452 38674
rect 58400 38610 58452 38616
rect 58214 38432 58270 38441
rect 58214 38367 58270 38376
rect 58308 37920 58360 37926
rect 58412 37897 58440 38610
rect 58308 37862 58360 37868
rect 58398 37888 58454 37897
rect 58216 37852 58268 37858
rect 58216 37794 58268 37800
rect 58228 37217 58256 37794
rect 58214 37208 58270 37217
rect 58214 37143 58270 37152
rect 58320 36673 58348 37862
rect 58398 37823 58454 37832
rect 58306 36664 58362 36673
rect 55548 36628 55600 36634
rect 58306 36599 58362 36608
rect 55548 36570 55600 36576
rect 55456 35404 55508 35410
rect 55456 35346 55508 35352
rect 55468 34798 55496 35346
rect 55560 35002 55588 36570
rect 58308 36560 58360 36566
rect 58308 36502 58360 36508
rect 58216 36492 58268 36498
rect 58216 36434 58268 36440
rect 58228 36129 58256 36434
rect 58214 36120 58270 36129
rect 58214 36055 58270 36064
rect 58320 35449 58348 36502
rect 58306 35440 58362 35449
rect 58306 35375 58362 35384
rect 59228 35132 59280 35138
rect 59228 35074 59280 35080
rect 55548 34996 55600 35002
rect 55548 34938 55600 34944
rect 58308 34996 58360 35002
rect 58308 34938 58360 34944
rect 58320 34905 58348 34938
rect 58306 34896 58362 34905
rect 58306 34831 58362 34840
rect 55456 34792 55508 34798
rect 55456 34734 55508 34740
rect 58216 34792 58268 34798
rect 58216 34734 58268 34740
rect 58228 34225 58256 34734
rect 58214 34216 58270 34225
rect 58214 34151 58270 34160
rect 56468 33772 56520 33778
rect 56468 33714 56520 33720
rect 56480 33098 56508 33714
rect 56744 33704 56796 33710
rect 59240 33681 59268 35074
rect 56744 33646 56796 33652
rect 59226 33672 59282 33681
rect 56756 33438 56784 33646
rect 59226 33607 59282 33616
rect 56744 33432 56796 33438
rect 56744 33374 56796 33380
rect 58216 33432 58268 33438
rect 58216 33374 58268 33380
rect 58228 33137 58256 33374
rect 58214 33128 58270 33137
rect 56468 33092 56520 33098
rect 58214 33063 58270 33072
rect 58308 33092 58360 33098
rect 56468 33034 56520 33040
rect 58308 33034 58360 33040
rect 58320 32457 58348 33034
rect 58306 32448 58362 32457
rect 58306 32383 58362 32392
rect 58216 32276 58268 32282
rect 58216 32218 58268 32224
rect 58228 31913 58256 32218
rect 58308 32208 58360 32214
rect 58308 32150 58360 32156
rect 58214 31904 58270 31913
rect 58214 31839 58270 31848
rect 56744 31324 56796 31330
rect 56744 31266 56796 31272
rect 56652 31188 56704 31194
rect 56652 31130 56704 31136
rect 56664 30922 56692 31130
rect 56652 30916 56704 30922
rect 56652 30858 56704 30864
rect 56756 30854 56784 31266
rect 58320 31233 58348 32150
rect 58306 31224 58362 31233
rect 58306 31159 58362 31168
rect 58400 30984 58452 30990
rect 58400 30926 58452 30932
rect 58216 30916 58268 30922
rect 58216 30858 58268 30864
rect 56744 30848 56796 30854
rect 56744 30790 56796 30796
rect 58228 30145 58256 30858
rect 58308 30848 58360 30854
rect 58308 30790 58360 30796
rect 58320 30689 58348 30790
rect 58306 30680 58362 30689
rect 58306 30615 58362 30624
rect 58214 30136 58270 30145
rect 58214 30071 58270 30080
rect 56008 29692 56060 29698
rect 56008 29634 56060 29640
rect 56020 28950 56048 29634
rect 58412 29465 58440 30926
rect 58398 29456 58454 29465
rect 58216 29420 58268 29426
rect 58398 29391 58454 29400
rect 58216 29362 58268 29368
rect 56008 28944 56060 28950
rect 58228 28921 58256 29362
rect 58308 28944 58360 28950
rect 56008 28886 56060 28892
rect 58214 28912 58270 28921
rect 58308 28886 58360 28892
rect 58214 28847 58270 28856
rect 56376 28332 56428 28338
rect 56376 28274 56428 28280
rect 56388 28066 56416 28274
rect 58320 28241 58348 28886
rect 58306 28232 58362 28241
rect 58306 28167 58362 28176
rect 56376 28060 56428 28066
rect 56376 28002 56428 28008
rect 58308 28060 58360 28066
rect 58308 28002 58360 28008
rect 58216 27992 58268 27998
rect 58216 27934 58268 27940
rect 58228 27153 58256 27934
rect 58320 27697 58348 28002
rect 58306 27688 58362 27697
rect 58306 27623 58362 27632
rect 58214 27144 58270 27153
rect 58214 27079 58270 27088
rect 59044 26972 59096 26978
rect 59044 26914 59096 26920
rect 58308 26904 58360 26910
rect 58308 26846 58360 26852
rect 58216 26836 58268 26842
rect 58216 26778 58268 26784
rect 58228 26473 58256 26778
rect 58214 26464 58270 26473
rect 58214 26399 58270 26408
rect 58320 25929 58348 26846
rect 58306 25920 58362 25929
rect 58306 25855 58362 25864
rect 59056 25249 59084 26914
rect 59412 25544 59464 25550
rect 59412 25486 59464 25492
rect 59042 25240 59098 25249
rect 59042 25175 59098 25184
rect 59424 24161 59452 25486
rect 59504 25476 59556 25482
rect 59504 25418 59556 25424
rect 59516 24705 59544 25418
rect 59502 24696 59558 24705
rect 59502 24631 59558 24640
rect 59410 24152 59466 24161
rect 56100 24116 56152 24122
rect 59410 24087 59466 24096
rect 56100 24058 56152 24064
rect 56112 23510 56140 24058
rect 58216 23980 58268 23986
rect 58216 23922 58268 23928
rect 56100 23504 56152 23510
rect 58228 23481 58256 23922
rect 58308 23504 58360 23510
rect 56100 23446 56152 23452
rect 58214 23472 58270 23481
rect 58308 23446 58360 23452
rect 58214 23407 58270 23416
rect 58320 22937 58348 23446
rect 58306 22928 58362 22937
rect 58306 22863 58362 22872
rect 53982 22792 54038 22801
rect 51224 22756 51276 22762
rect 53982 22727 54038 22736
rect 55732 22756 55784 22762
rect 51224 22698 51276 22704
rect 51038 20480 51094 20489
rect 51038 20415 51094 20424
rect 50762 19256 50818 19265
rect 50762 19191 50818 19200
rect 18104 18472 18156 18478
rect 18104 18414 18156 18420
rect 53996 18410 54024 22727
rect 55732 22698 55784 22704
rect 55744 22218 55772 22698
rect 90428 22626 90456 44510
rect 92728 44425 92756 44594
rect 92714 44416 92770 44425
rect 92714 44351 92770 44360
rect 92820 44289 92848 44662
rect 92806 44280 92862 44289
rect 92806 44215 92862 44224
rect 92716 43292 92768 43298
rect 92716 43234 92768 43240
rect 92728 43201 92756 43234
rect 92900 43224 92952 43230
rect 92714 43192 92770 43201
rect 92900 43166 92952 43172
rect 92714 43127 92770 43136
rect 92808 43156 92860 43162
rect 92808 43098 92860 43104
rect 92820 42521 92848 43098
rect 92912 42929 92940 43166
rect 92898 42920 92954 42929
rect 92898 42855 92954 42864
rect 92806 42512 92862 42521
rect 92806 42447 92862 42456
rect 92808 41932 92860 41938
rect 92808 41874 92860 41880
rect 92716 41864 92768 41870
rect 92716 41806 92768 41812
rect 92728 41705 92756 41806
rect 92714 41696 92770 41705
rect 92714 41631 92770 41640
rect 92820 41161 92848 41874
rect 92806 41152 92862 41161
rect 92806 41087 92862 41096
rect 92808 40572 92860 40578
rect 92808 40514 92860 40520
rect 92716 40504 92768 40510
rect 92716 40446 92768 40452
rect 92728 40209 92756 40446
rect 92714 40200 92770 40209
rect 92714 40135 92770 40144
rect 92820 40073 92848 40514
rect 92806 40064 92862 40073
rect 92806 39999 92862 40008
rect 92900 39144 92952 39150
rect 92714 39112 92770 39121
rect 92900 39086 92952 39092
rect 92714 39047 92770 39056
rect 92808 39076 92860 39082
rect 92728 39014 92756 39047
rect 92808 39018 92860 39024
rect 92716 39008 92768 39014
rect 92716 38950 92768 38956
rect 92820 38713 92848 39018
rect 92806 38704 92862 38713
rect 92806 38639 92862 38648
rect 92912 38305 92940 39086
rect 92898 38296 92954 38305
rect 92898 38231 92954 38240
rect 92808 37784 92860 37790
rect 92808 37726 92860 37732
rect 92716 37716 92768 37722
rect 92716 37658 92768 37664
rect 92728 37489 92756 37658
rect 92714 37480 92770 37489
rect 92714 37415 92770 37424
rect 92820 37081 92848 37726
rect 92806 37072 92862 37081
rect 92806 37007 92862 37016
rect 92808 36424 92860 36430
rect 92808 36366 92860 36372
rect 92716 36356 92768 36362
rect 92716 36298 92768 36304
rect 92728 36129 92756 36298
rect 92714 36120 92770 36129
rect 92714 36055 92770 36064
rect 92820 35993 92848 36366
rect 92806 35984 92862 35993
rect 92806 35919 92862 35928
rect 92808 35064 92860 35070
rect 92808 35006 92860 35012
rect 92716 34996 92768 35002
rect 92716 34938 92768 34944
rect 92728 34905 92756 34938
rect 92714 34896 92770 34905
rect 92714 34831 92770 34840
rect 92820 34633 92848 35006
rect 92806 34624 92862 34633
rect 92806 34559 92862 34568
rect 92714 33672 92770 33681
rect 92714 33607 92770 33616
rect 92808 33636 92860 33642
rect 92728 33506 92756 33607
rect 92808 33578 92860 33584
rect 92716 33500 92768 33506
rect 92716 33442 92768 33448
rect 92820 33409 92848 33578
rect 92900 33568 92952 33574
rect 92900 33510 92952 33516
rect 92806 33400 92862 33409
rect 92806 33335 92862 33344
rect 92912 33001 92940 33510
rect 92898 32992 92954 33001
rect 92898 32927 92954 32936
rect 92808 32276 92860 32282
rect 92808 32218 92860 32224
rect 92716 32208 92768 32214
rect 92716 32150 92768 32156
rect 92728 31913 92756 32150
rect 92714 31904 92770 31913
rect 92714 31839 92770 31848
rect 92820 31777 92848 32218
rect 92806 31768 92862 31777
rect 92806 31703 92862 31712
rect 92808 30916 92860 30922
rect 92808 30858 92860 30864
rect 92716 30848 92768 30854
rect 92716 30790 92768 30796
rect 92728 30689 92756 30790
rect 92714 30680 92770 30689
rect 92714 30615 92770 30624
rect 92820 30553 92848 30858
rect 92806 30544 92862 30553
rect 92806 30479 92862 30488
rect 92900 29488 92952 29494
rect 92714 29456 92770 29465
rect 92900 29430 92952 29436
rect 92714 29391 92770 29400
rect 92808 29420 92860 29426
rect 92728 29358 92756 29391
rect 92808 29362 92860 29368
rect 92716 29352 92768 29358
rect 92716 29294 92768 29300
rect 92820 28785 92848 29362
rect 92912 29193 92940 29430
rect 92898 29184 92954 29193
rect 92898 29119 92954 29128
rect 92806 28776 92862 28785
rect 92806 28711 92862 28720
rect 92900 28196 92952 28202
rect 92900 28138 92952 28144
rect 92808 28128 92860 28134
rect 92808 28070 92860 28076
rect 92716 28060 92768 28066
rect 92716 28002 92768 28008
rect 92728 27697 92756 28002
rect 92714 27688 92770 27697
rect 92714 27623 92770 27632
rect 92820 27425 92848 28070
rect 92806 27416 92862 27425
rect 92806 27351 92862 27360
rect 92716 26768 92768 26774
rect 92912 26745 92940 28138
rect 92716 26710 92768 26716
rect 92898 26736 92954 26745
rect 92728 26337 92756 26710
rect 92898 26671 92954 26680
rect 92714 26328 92770 26337
rect 92714 26263 92770 26272
rect 92900 25408 92952 25414
rect 92900 25350 92952 25356
rect 92808 25340 92860 25346
rect 92808 25282 92860 25288
rect 92716 25272 92768 25278
rect 92716 25214 92768 25220
rect 92728 24569 92756 25214
rect 92820 24977 92848 25282
rect 92912 25249 92940 25350
rect 92898 25240 92954 25249
rect 92898 25175 92954 25184
rect 92806 24968 92862 24977
rect 92806 24903 92862 24912
rect 92714 24560 92770 24569
rect 92714 24495 92770 24504
rect 92808 23980 92860 23986
rect 92808 23922 92860 23928
rect 92716 23912 92768 23918
rect 92716 23854 92768 23860
rect 92728 23753 92756 23854
rect 92714 23744 92770 23753
rect 92714 23679 92770 23688
rect 92820 23345 92848 23922
rect 92806 23336 92862 23345
rect 92806 23271 92862 23280
rect 58216 22620 58268 22626
rect 58216 22562 58268 22568
rect 90416 22620 90468 22626
rect 90416 22562 90468 22568
rect 58228 22257 58256 22562
rect 92808 22484 92860 22490
rect 92808 22426 92860 22432
rect 92716 22416 92768 22422
rect 92716 22358 92768 22364
rect 92728 22257 92756 22358
rect 58214 22248 58270 22257
rect 55732 22212 55784 22218
rect 92714 22248 92770 22257
rect 58214 22183 58270 22192
rect 58308 22212 58360 22218
rect 55732 22154 55784 22160
rect 92714 22183 92770 22192
rect 58308 22154 58360 22160
rect 58320 21713 58348 22154
rect 92820 22121 92848 22426
rect 92806 22112 92862 22121
rect 92806 22047 92862 22056
rect 58306 21704 58362 21713
rect 58306 21639 58362 21648
rect 58216 21260 58268 21266
rect 58216 21202 58268 21208
rect 92716 21260 92768 21266
rect 92716 21202 92768 21208
rect 58228 21169 58256 21202
rect 92728 21169 92756 21202
rect 58214 21160 58270 21169
rect 58214 21095 58270 21104
rect 92714 21160 92770 21169
rect 92714 21095 92770 21104
rect 61710 21024 61766 21033
rect 61416 20982 61710 21010
rect 61710 20959 61766 20968
rect 63274 21024 63330 21033
rect 64746 21024 64802 21033
rect 63330 20982 63440 21010
rect 64452 20982 64746 21010
rect 63274 20959 63330 20968
rect 65758 21024 65814 21033
rect 65464 20982 65758 21010
rect 64746 20959 64802 20968
rect 65758 20959 65814 20968
rect 62722 20888 62778 20897
rect 62428 20846 62722 20874
rect 66862 20888 66918 20897
rect 66568 20846 66862 20874
rect 62722 20823 62778 20832
rect 67580 20846 67824 20874
rect 66862 20823 66918 20832
rect 53984 18404 54036 18410
rect 53984 18346 54036 18352
rect 60792 18336 60844 18342
rect 60792 18278 60844 18284
rect 54812 18268 54864 18274
rect 54812 18210 54864 18216
rect 42852 18200 42904 18206
rect 42852 18142 42904 18148
rect 30800 18064 30852 18070
rect 30800 18006 30852 18012
rect 24820 17928 24872 17934
rect 24820 17870 24872 17876
rect 18840 17860 18892 17866
rect 18840 17802 18892 17808
rect 12860 17792 12912 17798
rect 12860 17734 12912 17740
rect 12872 9304 12900 17734
rect 18852 9304 18880 17802
rect 24832 9304 24860 17870
rect 30812 9304 30840 18006
rect 36780 17996 36832 18002
rect 36780 17938 36832 17944
rect 36792 9304 36820 17938
rect 42864 9304 42892 18142
rect 48832 18132 48884 18138
rect 48832 18074 48884 18080
rect 48844 9304 48872 18074
rect 54824 9304 54852 18210
rect 60804 9304 60832 18278
rect 67796 17118 67824 20846
rect 68256 20846 68592 20874
rect 69604 20846 69848 20874
rect 71720 20846 71964 20874
rect 68256 18478 68284 20846
rect 69820 18478 69848 20846
rect 68244 18472 68296 18478
rect 68244 18414 68296 18420
rect 69808 18472 69860 18478
rect 69808 18414 69860 18420
rect 71936 18410 71964 20846
rect 72396 20846 72732 20874
rect 73408 20846 73744 20874
rect 74788 20846 74848 20874
rect 75524 20846 75860 20874
rect 76536 20846 76872 20874
rect 77548 20846 77884 20874
rect 78928 20846 78988 20874
rect 79112 20846 80000 20874
rect 80676 20846 81012 20874
rect 81688 20846 82024 20874
rect 83068 20846 83128 20874
rect 83804 20846 84140 20874
rect 84448 20846 85152 20874
rect 85828 20846 86164 20874
rect 71924 18404 71976 18410
rect 71924 18346 71976 18352
rect 72396 18206 72424 20846
rect 72384 18200 72436 18206
rect 72384 18142 72436 18148
rect 73408 18002 73436 20846
rect 74788 18070 74816 20846
rect 74776 18064 74828 18070
rect 74776 18006 74828 18012
rect 73396 17996 73448 18002
rect 73396 17938 73448 17944
rect 75524 17934 75552 20846
rect 76156 18336 76208 18342
rect 76156 18278 76208 18284
rect 75512 17928 75564 17934
rect 75512 17870 75564 17876
rect 67784 17112 67836 17118
rect 67784 17054 67836 17060
rect 72844 12352 72896 12358
rect 72844 12294 72896 12300
rect 66864 12284 66916 12290
rect 66864 12226 66916 12232
rect 66876 9304 66904 12226
rect 72856 9304 72884 12294
rect 76168 12290 76196 18278
rect 76536 17866 76564 20846
rect 76524 17860 76576 17866
rect 76524 17802 76576 17808
rect 77548 17798 77576 20846
rect 78928 18290 78956 20846
rect 78836 18262 78956 18290
rect 77536 17792 77588 17798
rect 77536 17734 77588 17740
rect 76156 12284 76208 12290
rect 76156 12226 76208 12232
rect 78836 9304 78864 18262
rect 79112 12358 79140 20846
rect 80676 18342 80704 20846
rect 80664 18336 80716 18342
rect 80664 18278 80716 18284
rect 81688 18274 81716 20846
rect 81676 18268 81728 18274
rect 81676 18210 81728 18216
rect 83068 18070 83096 20846
rect 83804 18138 83832 20846
rect 83792 18132 83844 18138
rect 83792 18074 83844 18080
rect 83056 18064 83108 18070
rect 83056 18006 83108 18012
rect 79100 12352 79152 12358
rect 79100 12294 79152 12300
rect 84448 12290 84476 20846
rect 85828 12358 85856 20846
rect 87254 20602 87282 20860
rect 88280 20846 88524 20874
rect 89292 20846 89628 20874
rect 87254 20574 87328 20602
rect 87300 12426 87328 20574
rect 88496 18342 88524 20846
rect 88484 18336 88536 18342
rect 88484 18278 88536 18284
rect 89600 17594 89628 20846
rect 89968 20846 90304 20874
rect 89968 18290 89996 20846
rect 93372 19838 93400 46294
rect 94740 46216 94792 46222
rect 94740 46158 94792 46164
rect 93360 19832 93412 19838
rect 93360 19774 93412 19780
rect 94752 19770 94780 46158
rect 96120 46148 96172 46154
rect 96120 46090 96172 46096
rect 96132 22558 96160 46090
rect 98144 43496 98196 43502
rect 98144 43438 98196 43444
rect 98156 43162 98184 43438
rect 98144 43156 98196 43162
rect 98144 43098 98196 43104
rect 98972 38396 99024 38402
rect 98972 38338 99024 38344
rect 98880 38260 98932 38266
rect 98880 38202 98932 38208
rect 98892 37790 98920 38202
rect 98880 37784 98932 37790
rect 98880 37726 98932 37732
rect 98984 37722 99012 38338
rect 98972 37716 99024 37722
rect 98972 37658 99024 37664
rect 97684 23164 97736 23170
rect 97684 23106 97736 23112
rect 96120 22552 96172 22558
rect 96120 22494 96172 22500
rect 97696 22422 97724 23106
rect 98144 22688 98196 22694
rect 98144 22630 98196 22636
rect 98156 22490 98184 22630
rect 98144 22484 98196 22490
rect 98144 22426 98196 22432
rect 97684 22416 97736 22422
rect 97684 22358 97736 22364
rect 94740 19764 94792 19770
rect 94740 19706 94792 19712
rect 100272 18410 100300 49014
rect 100364 49010 100392 59894
rect 100352 49004 100404 49010
rect 100352 48946 100404 48952
rect 103032 48942 103060 61254
rect 104412 61250 104440 69550
rect 104504 63698 104532 70978
rect 105148 68186 105176 73766
rect 106700 73756 106752 73762
rect 106700 73698 106752 73704
rect 106516 72396 106568 72402
rect 106516 72338 106568 72344
rect 105136 68180 105188 68186
rect 105136 68122 105188 68128
rect 106528 65641 106556 72338
rect 106712 70401 106740 73698
rect 106792 73688 106844 73694
rect 106792 73630 106844 73636
rect 106804 72713 106832 73630
rect 106790 72704 106846 72713
rect 106790 72639 106846 72648
rect 106698 70392 106754 70401
rect 106698 70327 106754 70336
rect 134036 70226 134064 111127
rect 134772 102118 134800 116567
rect 134864 116534 134892 117791
rect 134942 117312 134998 117321
rect 134942 117247 134998 117256
rect 134852 116528 134904 116534
rect 134852 116470 134904 116476
rect 134850 115544 134906 115553
rect 134850 115479 134906 115488
rect 134864 102254 134892 115479
rect 134852 102248 134904 102254
rect 134852 102190 134904 102196
rect 134760 102112 134812 102118
rect 134760 102054 134812 102060
rect 134956 102050 134984 117247
rect 136888 116398 136916 118442
rect 136980 117826 137008 119258
rect 137440 119254 137468 120754
rect 137520 120744 137572 120750
rect 137520 120686 137572 120692
rect 137428 119248 137480 119254
rect 137428 119190 137480 119196
rect 137532 119118 137560 120686
rect 138084 120614 138112 122386
rect 138176 121906 138204 123338
rect 143592 123328 143644 123334
rect 143590 123296 143592 123305
rect 143644 123296 143646 123305
rect 143590 123231 143646 123240
rect 142856 122920 142908 122926
rect 142856 122862 142908 122868
rect 142868 122761 142896 122862
rect 142854 122752 142910 122761
rect 142854 122687 142910 122696
rect 142764 121968 142816 121974
rect 142764 121910 142816 121916
rect 138164 121900 138216 121906
rect 138164 121842 138216 121848
rect 142776 121537 142804 121910
rect 143040 121900 143092 121906
rect 143040 121842 143092 121848
rect 143052 121809 143080 121842
rect 143038 121800 143094 121809
rect 143038 121735 143094 121744
rect 142762 121528 142818 121537
rect 142762 121463 142818 121472
rect 138072 120608 138124 120614
rect 142948 120608 143000 120614
rect 138072 120550 138124 120556
rect 142946 120576 142948 120585
rect 143000 120576 143002 120585
rect 142946 120511 143002 120520
rect 143592 120540 143644 120546
rect 143592 120482 143644 120488
rect 143604 120313 143632 120482
rect 143590 120304 143646 120313
rect 143590 120239 143646 120248
rect 137612 119588 137664 119594
rect 137612 119530 137664 119536
rect 137520 119112 137572 119118
rect 137520 119054 137572 119060
rect 137520 118228 137572 118234
rect 137520 118170 137572 118176
rect 136968 117820 137020 117826
rect 136968 117762 137020 117768
rect 136876 116392 136928 116398
rect 136876 116334 136928 116340
rect 137532 116330 137560 118170
rect 137624 117758 137652 119530
rect 143592 119248 143644 119254
rect 143590 119216 143592 119225
rect 143644 119216 143646 119225
rect 142580 119180 142632 119186
rect 143590 119151 143646 119160
rect 142580 119122 142632 119128
rect 142592 118545 142620 119122
rect 143592 119112 143644 119118
rect 143590 119080 143592 119089
rect 143644 119080 143646 119089
rect 143590 119015 143646 119024
rect 142578 118536 142634 118545
rect 142578 118471 142634 118480
rect 142580 117820 142632 117826
rect 142580 117762 142632 117768
rect 137612 117752 137664 117758
rect 142592 117729 142620 117762
rect 143224 117752 143276 117758
rect 137612 117694 137664 117700
rect 142578 117720 142634 117729
rect 143224 117694 143276 117700
rect 142578 117655 142634 117664
rect 143236 117321 143264 117694
rect 143222 117312 143278 117321
rect 143222 117247 143278 117256
rect 142764 116460 142816 116466
rect 142764 116402 142816 116408
rect 137520 116324 137572 116330
rect 137520 116266 137572 116272
rect 135034 116088 135090 116097
rect 135034 116023 135090 116032
rect 135048 102186 135076 116023
rect 142776 115553 142804 116402
rect 142948 116392 143000 116398
rect 142946 116360 142948 116369
rect 143000 116360 143002 116369
rect 142946 116295 143002 116304
rect 143592 116324 143644 116330
rect 143592 116266 143644 116272
rect 143604 116097 143632 116266
rect 143590 116088 143646 116097
rect 143590 116023 143646 116032
rect 142762 115544 142818 115553
rect 142762 115479 142818 115488
rect 135126 114864 135182 114873
rect 135126 114799 135182 114808
rect 135140 102390 135168 114799
rect 135310 114320 135366 114329
rect 135310 114255 135366 114264
rect 135218 113232 135274 113241
rect 135218 113167 135274 113176
rect 135128 102384 135180 102390
rect 135128 102326 135180 102332
rect 135036 102180 135088 102186
rect 135036 102122 135088 102128
rect 134944 102044 134996 102050
rect 134944 101986 134996 101992
rect 135232 101370 135260 113167
rect 135324 101982 135352 114255
rect 135402 113776 135458 113785
rect 135402 113711 135404 113720
rect 135456 113711 135458 113720
rect 141568 113740 141620 113746
rect 135404 113682 135456 113688
rect 141568 113682 141620 113688
rect 135312 101976 135364 101982
rect 135312 101918 135364 101924
rect 135220 101364 135272 101370
rect 135220 101306 135272 101312
rect 140464 101364 140516 101370
rect 140464 101306 140516 101312
rect 140476 99740 140504 101306
rect 141580 99740 141608 113682
rect 143696 101982 143724 153854
rect 156576 151758 156604 153868
rect 156564 151752 156616 151758
rect 156564 151694 156616 151700
rect 163200 151690 163228 153868
rect 163188 151684 163240 151690
rect 163188 151626 163240 151632
rect 169916 142510 169944 153868
rect 183072 143462 183100 162807
rect 187948 162026 187976 166450
rect 190052 165012 190104 165018
rect 190052 164954 190104 164960
rect 189960 163448 190012 163454
rect 189960 163390 190012 163396
rect 187936 162020 187988 162026
rect 187936 161962 187988 161968
rect 183150 161648 183206 161657
rect 183150 161583 183206 161592
rect 183060 143456 183112 143462
rect 183060 143398 183112 143404
rect 183164 143394 183192 161583
rect 183242 160424 183298 160433
rect 183242 160359 183298 160368
rect 183256 143530 183284 160359
rect 183334 159200 183390 159209
rect 183334 159135 183390 159144
rect 183348 143870 183376 159135
rect 183518 157976 183574 157985
rect 183518 157911 183574 157920
rect 183426 156752 183482 156761
rect 183426 156687 183482 156696
rect 183440 144006 183468 156687
rect 183428 144000 183480 144006
rect 183428 143942 183480 143948
rect 183532 143938 183560 157911
rect 189972 156761 190000 163390
rect 190064 158801 190092 164954
rect 191352 164785 191380 167538
rect 191904 166825 191932 168898
rect 191984 168888 192036 168894
rect 191984 168830 192036 168836
rect 191996 168729 192024 168830
rect 191982 168720 192038 168729
rect 191982 168655 192038 168664
rect 191890 166816 191946 166825
rect 191890 166751 191946 166760
rect 212684 165284 212736 165290
rect 212684 165226 212736 165232
rect 212696 164921 212724 165226
rect 212682 164912 212738 164921
rect 212682 164847 212738 164856
rect 191338 164776 191394 164785
rect 191338 164711 191394 164720
rect 211762 163824 211818 163833
rect 211762 163759 211818 163768
rect 211776 163658 211804 163759
rect 211764 163652 211816 163658
rect 211764 163594 211816 163600
rect 191984 163040 192036 163046
rect 191984 162982 192036 162988
rect 191996 162745 192024 162982
rect 191982 162736 192038 162745
rect 191982 162671 192038 162680
rect 191340 162020 191392 162026
rect 191340 161962 191392 161968
rect 191352 160841 191380 161962
rect 191338 160832 191394 160841
rect 191338 160767 191394 160776
rect 190050 158792 190106 158801
rect 190050 158727 190106 158736
rect 211946 157160 212002 157169
rect 211946 157095 212002 157104
rect 189958 156752 190014 156761
rect 189958 156687 190014 156696
rect 211960 156518 211988 157095
rect 212696 156518 212724 164847
rect 211948 156512 212000 156518
rect 211948 156454 212000 156460
rect 212684 156512 212736 156518
rect 212684 156454 212736 156460
rect 188028 155492 188080 155498
rect 188028 155434 188080 155440
rect 183610 154440 183666 154449
rect 183610 154375 183666 154384
rect 183624 144074 183652 154375
rect 183612 144068 183664 144074
rect 183612 144010 183664 144016
rect 187936 144068 187988 144074
rect 187936 144010 187988 144016
rect 183520 143932 183572 143938
rect 183520 143874 183572 143880
rect 183336 143864 183388 143870
rect 183336 143806 183388 143812
rect 183244 143524 183296 143530
rect 183244 143466 183296 143472
rect 183152 143388 183204 143394
rect 183152 143330 183204 143336
rect 167696 142504 167748 142510
rect 167696 142446 167748 142452
rect 169904 142504 169956 142510
rect 169904 142446 169956 142452
rect 167708 138786 167736 142446
rect 187948 140826 187976 144010
rect 188040 140962 188068 155434
rect 191982 154848 192038 154857
rect 191982 154783 192038 154792
rect 189408 144000 189460 144006
rect 189408 143942 189460 143948
rect 188040 140934 188528 140962
rect 188500 140826 188528 140934
rect 187948 140798 188238 140826
rect 188500 140798 188790 140826
rect 189420 140690 189448 143942
rect 189500 143932 189552 143938
rect 189500 143874 189552 143880
rect 189512 140826 189540 143874
rect 190052 143864 190104 143870
rect 190052 143806 190104 143812
rect 190064 140826 190092 143806
rect 190788 143524 190840 143530
rect 190788 143466 190840 143472
rect 190800 140826 190828 143466
rect 191996 143394 192024 154783
rect 193272 152364 193324 152370
rect 193272 152306 193324 152312
rect 193088 144068 193140 144074
rect 193088 144010 193140 144016
rect 192076 143456 192128 143462
rect 192076 143398 192128 143404
rect 191340 143388 191392 143394
rect 191340 143330 191392 143336
rect 191984 143388 192036 143394
rect 191984 143330 192036 143336
rect 191352 140826 191380 143330
rect 192088 140826 192116 143398
rect 189512 140798 189894 140826
rect 190064 140798 190446 140826
rect 190800 140798 191090 140826
rect 191352 140798 191642 140826
rect 192088 140798 192194 140826
rect 193100 140690 193128 144010
rect 193284 140962 193312 152306
rect 194112 152302 194140 153868
rect 194480 152370 194508 153868
rect 194862 153854 195060 153882
rect 194468 152364 194520 152370
rect 194468 152306 194520 152312
rect 194928 152364 194980 152370
rect 194928 152306 194980 152312
rect 193364 152296 193416 152302
rect 193364 152238 193416 152244
rect 194100 152296 194152 152302
rect 194100 152238 194152 152244
rect 193376 144074 193404 152238
rect 194652 151276 194704 151282
rect 194652 151218 194704 151224
rect 193364 144068 193416 144074
rect 193364 144010 193416 144016
rect 194192 143456 194244 143462
rect 194192 143398 194244 143404
rect 193192 140934 193312 140962
rect 193192 140826 193220 140934
rect 193192 140798 193298 140826
rect 194204 140690 194232 143398
rect 194664 140690 194692 151218
rect 194744 151004 194796 151010
rect 194744 150946 194796 150952
rect 194756 143462 194784 150946
rect 194744 143456 194796 143462
rect 194744 143398 194796 143404
rect 194940 140826 194968 152306
rect 195032 151010 195060 153854
rect 195112 151548 195164 151554
rect 195112 151490 195164 151496
rect 195020 151004 195072 151010
rect 195020 150946 195072 150952
rect 195124 140826 195152 151490
rect 195308 151282 195336 153868
rect 195676 152370 195704 153868
rect 195664 152364 195716 152370
rect 195664 152306 195716 152312
rect 196044 151554 196072 153868
rect 196228 153854 196518 153882
rect 196228 152250 196256 153854
rect 196584 152364 196636 152370
rect 196584 152306 196636 152312
rect 196136 152222 196256 152250
rect 196032 151548 196084 151554
rect 196032 151490 196084 151496
rect 195296 151276 195348 151282
rect 195296 151218 195348 151224
rect 196136 140962 196164 152222
rect 196216 150936 196268 150942
rect 196216 150878 196268 150884
rect 196044 140934 196164 140962
rect 196044 140826 196072 140934
rect 196228 140826 196256 150878
rect 196596 146130 196624 152306
rect 196872 151078 196900 153868
rect 197240 152370 197268 153868
rect 197228 152364 197280 152370
rect 197228 152306 197280 152312
rect 197596 152364 197648 152370
rect 197596 152306 197648 152312
rect 196860 151072 196912 151078
rect 196860 151014 196912 151020
rect 197608 146182 197636 152306
rect 197596 146176 197648 146182
rect 196596 146102 196992 146130
rect 197596 146118 197648 146124
rect 196964 140826 196992 146102
rect 197700 140826 197728 153868
rect 198068 152370 198096 153868
rect 198056 152364 198108 152370
rect 198056 152306 198108 152312
rect 198148 146176 198200 146182
rect 198148 146118 198200 146124
rect 198160 140826 198188 146118
rect 198436 144074 198464 153868
rect 198424 144068 198476 144074
rect 198424 144010 198476 144016
rect 198896 144006 198924 153868
rect 199264 150890 199292 153868
rect 199632 151146 199660 153868
rect 200106 153854 200304 153882
rect 199620 151140 199672 151146
rect 199620 151082 199672 151088
rect 200172 151140 200224 151146
rect 200172 151082 200224 151088
rect 199264 150862 199752 150890
rect 199068 144068 199120 144074
rect 199068 144010 199120 144016
rect 198884 144000 198936 144006
rect 198884 143942 198936 143948
rect 194940 140798 195046 140826
rect 195124 140798 195598 140826
rect 196044 140798 196150 140826
rect 196228 140798 196794 140826
rect 196964 140798 197346 140826
rect 197700 140798 197898 140826
rect 198160 140798 198450 140826
rect 199080 140690 199108 144010
rect 199252 144000 199304 144006
rect 199252 143942 199304 143948
rect 199264 140826 199292 143942
rect 199724 140826 199752 150862
rect 200184 142764 200212 151082
rect 200276 142918 200304 153854
rect 200460 151690 200488 153868
rect 200448 151684 200500 151690
rect 200448 151626 200500 151632
rect 200828 143938 200856 153868
rect 201184 151684 201236 151690
rect 201184 151626 201236 151632
rect 201196 144074 201224 151626
rect 201184 144068 201236 144074
rect 201184 144010 201236 144016
rect 201288 144006 201316 153868
rect 201276 144000 201328 144006
rect 201276 143942 201328 143948
rect 200816 143932 200868 143938
rect 200816 143874 200868 143880
rect 201656 143870 201684 153868
rect 202116 152370 202144 153868
rect 202104 152364 202156 152370
rect 202104 152306 202156 152312
rect 201736 144068 201788 144074
rect 201736 144010 201788 144016
rect 201644 143864 201696 143870
rect 201644 143806 201696 143812
rect 200264 142912 200316 142918
rect 200264 142854 200316 142860
rect 200908 142912 200960 142918
rect 200908 142854 200960 142860
rect 200184 142736 200396 142764
rect 200368 140826 200396 142736
rect 200920 140826 200948 142854
rect 201748 140826 201776 144010
rect 202484 143938 202512 153868
rect 202866 153854 203064 153882
rect 202932 152364 202984 152370
rect 202932 152306 202984 152312
rect 202944 144074 202972 152306
rect 202932 144068 202984 144074
rect 202932 144010 202984 144016
rect 203036 144006 203064 153854
rect 203312 152302 203340 153868
rect 203680 152370 203708 153868
rect 203668 152364 203720 152370
rect 203668 152306 203720 152312
rect 203300 152296 203352 152302
rect 203300 152238 203352 152244
rect 204048 151010 204076 153868
rect 204508 152166 204536 153868
rect 204876 152234 204904 153868
rect 204864 152228 204916 152234
rect 204864 152170 204916 152176
rect 204496 152160 204548 152166
rect 204496 152102 204548 152108
rect 205244 152098 205272 153868
rect 205232 152092 205284 152098
rect 205232 152034 205284 152040
rect 205704 151690 205732 153868
rect 206086 153854 206376 153882
rect 205968 152364 206020 152370
rect 205968 152306 206020 152312
rect 205692 151684 205744 151690
rect 205692 151626 205744 151632
rect 204036 151004 204088 151010
rect 204036 150946 204088 150952
rect 203852 144068 203904 144074
rect 203852 144010 203904 144016
rect 202748 144000 202800 144006
rect 202748 143942 202800 143948
rect 203024 144000 203076 144006
rect 203024 143942 203076 143948
rect 202288 143932 202340 143938
rect 202288 143874 202340 143880
rect 202472 143932 202524 143938
rect 202472 143874 202524 143880
rect 202300 140826 202328 143874
rect 202760 140826 202788 143942
rect 203300 143864 203352 143870
rect 203300 143806 203352 143812
rect 203312 140826 203340 143806
rect 203864 140826 203892 144010
rect 204956 144000 205008 144006
rect 204956 143942 205008 143948
rect 204496 143932 204548 143938
rect 204496 143874 204548 143880
rect 204508 140826 204536 143874
rect 204968 140826 204996 143942
rect 205980 143666 206008 152306
rect 206060 152296 206112 152302
rect 206060 152238 206112 152244
rect 205968 143660 206020 143666
rect 205968 143602 206020 143608
rect 206072 140962 206100 152238
rect 206348 151894 206376 153854
rect 206440 151962 206468 153868
rect 206428 151956 206480 151962
rect 206428 151898 206480 151904
rect 206336 151888 206388 151894
rect 206336 151830 206388 151836
rect 206900 151214 206928 153868
rect 207282 153854 207572 153882
rect 207348 152228 207400 152234
rect 207348 152170 207400 152176
rect 207256 152160 207308 152166
rect 207256 152102 207308 152108
rect 206888 151208 206940 151214
rect 206888 151150 206940 151156
rect 206244 151004 206296 151010
rect 206244 150946 206296 150952
rect 206152 143660 206204 143666
rect 206152 143602 206204 143608
rect 205980 140934 206100 140962
rect 199264 140798 199646 140826
rect 199724 140798 200198 140826
rect 200368 140798 200750 140826
rect 200920 140798 201302 140826
rect 201748 140798 201854 140826
rect 202300 140798 202498 140826
rect 202760 140798 203050 140826
rect 203312 140798 203602 140826
rect 203864 140798 204154 140826
rect 204508 140798 204706 140826
rect 204968 140798 205350 140826
rect 205980 140690 206008 140934
rect 206164 140826 206192 143602
rect 206256 141098 206284 150946
rect 206256 141070 206560 141098
rect 206532 140826 206560 141070
rect 207268 140826 207296 152102
rect 207360 142186 207388 152170
rect 207544 151010 207572 153854
rect 207636 151826 207664 153868
rect 207992 152092 208044 152098
rect 207992 152034 208044 152040
rect 207624 151820 207676 151826
rect 207624 151762 207676 151768
rect 207900 151684 207952 151690
rect 207900 151626 207952 151632
rect 207532 151004 207584 151010
rect 207532 150946 207584 150952
rect 207912 143598 207940 151626
rect 208004 143666 208032 152034
rect 208096 151350 208124 153868
rect 208084 151344 208136 151350
rect 208084 151286 208136 151292
rect 208464 151078 208492 153868
rect 208832 152098 208860 153868
rect 208820 152092 208872 152098
rect 208820 152034 208872 152040
rect 208820 151888 208872 151894
rect 208820 151830 208872 151836
rect 208452 151072 208504 151078
rect 208452 151014 208504 151020
rect 208832 143666 208860 151830
rect 209292 151690 209320 153868
rect 209660 151758 209688 153868
rect 212868 152092 212920 152098
rect 212868 152034 212920 152040
rect 210016 151956 210068 151962
rect 210016 151898 210068 151904
rect 209648 151752 209700 151758
rect 209648 151694 209700 151700
rect 209280 151684 209332 151690
rect 209280 151626 209332 151632
rect 207992 143660 208044 143666
rect 207992 143602 208044 143608
rect 208636 143660 208688 143666
rect 208636 143602 208688 143608
rect 208820 143660 208872 143666
rect 208820 143602 208872 143608
rect 209556 143660 209608 143666
rect 209556 143602 209608 143608
rect 207900 143592 207952 143598
rect 207900 143534 207952 143540
rect 207360 142158 207940 142186
rect 207912 140826 207940 142158
rect 208648 140826 208676 143602
rect 209004 143592 209056 143598
rect 209004 143534 209056 143540
rect 209016 140826 209044 143534
rect 209568 140826 209596 143602
rect 210028 140826 210056 151898
rect 210936 151820 210988 151826
rect 210936 151762 210988 151768
rect 210752 151344 210804 151350
rect 210752 151286 210804 151292
rect 210108 151208 210160 151214
rect 210108 151150 210160 151156
rect 210120 140962 210148 151150
rect 210660 151072 210712 151078
rect 210660 151014 210712 151020
rect 210672 142986 210700 151014
rect 210660 142980 210712 142986
rect 210660 142922 210712 142928
rect 210764 142850 210792 151286
rect 210844 151004 210896 151010
rect 210844 150946 210896 150952
rect 210856 143666 210884 150946
rect 210844 143660 210896 143666
rect 210844 143602 210896 143608
rect 210948 143122 210976 151762
rect 211396 143660 211448 143666
rect 211396 143602 211448 143608
rect 210936 143116 210988 143122
rect 210936 143058 210988 143064
rect 210752 142844 210804 142850
rect 210752 142786 210804 142792
rect 210120 140934 210700 140962
rect 210672 140826 210700 140934
rect 211408 140826 211436 143602
rect 212880 143274 212908 152034
rect 214248 151752 214300 151758
rect 214248 151694 214300 151700
rect 214156 151684 214208 151690
rect 214156 151626 214208 151632
rect 212880 143246 213368 143274
rect 211764 143116 211816 143122
rect 211764 143058 211816 143064
rect 211776 140826 211804 143058
rect 212868 142980 212920 142986
rect 212868 142922 212920 142928
rect 212316 142844 212368 142850
rect 212316 142786 212368 142792
rect 212328 140826 212356 142786
rect 212880 140826 212908 142922
rect 206164 140798 206454 140826
rect 206532 140798 207006 140826
rect 207268 140798 207558 140826
rect 207912 140798 208202 140826
rect 208648 140798 208754 140826
rect 209016 140798 209306 140826
rect 209568 140798 209858 140826
rect 210028 140798 210410 140826
rect 210672 140798 211054 140826
rect 211408 140798 211606 140826
rect 211776 140798 212158 140826
rect 212328 140798 212710 140826
rect 212880 140798 213262 140826
rect 189342 140662 189448 140690
rect 192746 140662 193128 140690
rect 193942 140662 194232 140690
rect 194494 140662 194692 140690
rect 199002 140662 199108 140690
rect 205902 140662 206008 140690
rect 213340 140690 213368 143246
rect 214168 140826 214196 151626
rect 214260 143666 214288 151694
rect 214248 143660 214300 143666
rect 214248 143602 214300 143608
rect 214708 143660 214760 143666
rect 214708 143602 214760 143608
rect 214720 140826 214748 143602
rect 215628 143388 215680 143394
rect 215628 143330 215680 143336
rect 214168 140798 214458 140826
rect 214720 140798 215010 140826
rect 215640 140690 215668 143330
rect 213340 140662 213906 140690
rect 215562 140662 215668 140690
rect 184990 140160 185046 140169
rect 184990 140095 185046 140104
rect 167400 138758 167736 138786
rect 177632 138560 177684 138566
rect 177632 138502 177684 138508
rect 177722 138528 177778 138537
rect 177644 138265 177672 138502
rect 185004 138498 185032 140095
rect 185082 140024 185138 140033
rect 185082 139959 185138 139968
rect 185096 138566 185124 139959
rect 185358 138936 185414 138945
rect 185358 138871 185414 138880
rect 185266 138664 185322 138673
rect 185266 138599 185322 138608
rect 185084 138560 185136 138566
rect 185084 138502 185136 138508
rect 177722 138463 177724 138472
rect 177776 138463 177778 138472
rect 184992 138492 185044 138498
rect 177724 138434 177776 138440
rect 184992 138434 185044 138440
rect 177630 138256 177686 138265
rect 177630 138191 177686 138200
rect 185174 137848 185230 137857
rect 185174 137783 185230 137792
rect 185188 137274 185216 137783
rect 181588 137268 181640 137274
rect 181588 137210 181640 137216
rect 185176 137268 185228 137274
rect 185176 137210 185228 137216
rect 177632 137132 177684 137138
rect 177632 137074 177684 137080
rect 177644 136905 177672 137074
rect 177724 137064 177776 137070
rect 177722 137032 177724 137041
rect 177776 137032 177778 137041
rect 177722 136967 177778 136976
rect 177630 136896 177686 136905
rect 177630 136831 177686 136840
rect 181600 136662 181628 137210
rect 182232 137200 182284 137206
rect 182232 137142 182284 137148
rect 177724 136656 177776 136662
rect 177724 136598 177776 136604
rect 181588 136656 181640 136662
rect 181588 136598 181640 136604
rect 177736 136361 177764 136598
rect 177722 136352 177778 136361
rect 177722 136287 177778 136296
rect 181956 135840 182008 135846
rect 181956 135782 182008 135788
rect 177632 135772 177684 135778
rect 177632 135714 177684 135720
rect 177644 135273 177672 135714
rect 177724 135704 177776 135710
rect 177724 135646 177776 135652
rect 177736 135545 177764 135646
rect 177722 135536 177778 135545
rect 177722 135471 177778 135480
rect 177630 135264 177686 135273
rect 177630 135199 177686 135208
rect 177632 134412 177684 134418
rect 177632 134354 177684 134360
rect 177644 133505 177672 134354
rect 181968 134350 181996 135782
rect 182244 135710 182272 137142
rect 185280 137138 185308 138599
rect 185268 137132 185320 137138
rect 185268 137074 185320 137080
rect 185372 137070 185400 138871
rect 185450 137304 185506 137313
rect 185450 137239 185506 137248
rect 185464 137206 185492 137239
rect 185452 137200 185504 137206
rect 185452 137142 185504 137148
rect 185360 137064 185412 137070
rect 185360 137006 185412 137012
rect 185174 136624 185230 136633
rect 185174 136559 185230 136568
rect 182324 135908 182376 135914
rect 182324 135850 182376 135856
rect 182232 135704 182284 135710
rect 182232 135646 182284 135652
rect 177724 134344 177776 134350
rect 177722 134312 177724 134321
rect 181956 134344 182008 134350
rect 177776 134312 177778 134321
rect 181956 134286 182008 134292
rect 177722 134247 177778 134256
rect 182336 134078 182364 135850
rect 185188 135778 185216 136559
rect 185266 136080 185322 136089
rect 185266 136015 185322 136024
rect 185280 135846 185308 136015
rect 185358 135944 185414 135953
rect 185358 135879 185360 135888
rect 185412 135879 185414 135888
rect 185360 135850 185412 135856
rect 185268 135840 185320 135846
rect 185268 135782 185320 135788
rect 185176 135772 185228 135778
rect 185176 135714 185228 135720
rect 185174 134856 185230 134865
rect 185174 134791 185230 134800
rect 185082 134448 185138 134457
rect 185188 134418 185216 134791
rect 185082 134383 185138 134392
rect 185176 134412 185228 134418
rect 177724 134072 177776 134078
rect 177724 134014 177776 134020
rect 182324 134072 182376 134078
rect 182324 134014 182376 134020
rect 177736 133913 177764 134014
rect 177722 133904 177778 133913
rect 177722 133839 177778 133848
rect 177630 133496 177686 133505
rect 177630 133431 177686 133440
rect 177632 132984 177684 132990
rect 177632 132926 177684 132932
rect 177644 132281 177672 132926
rect 185096 132922 185124 134383
rect 185176 134354 185228 134360
rect 185174 133768 185230 133777
rect 185174 133703 185230 133712
rect 185188 132990 185216 133703
rect 185818 133088 185874 133097
rect 185818 133023 185874 133032
rect 185176 132984 185228 132990
rect 185176 132926 185228 132932
rect 177724 132916 177776 132922
rect 177724 132858 177776 132864
rect 185084 132916 185136 132922
rect 185084 132858 185136 132864
rect 177736 132689 177764 132858
rect 177722 132680 177778 132689
rect 177722 132615 177778 132624
rect 177630 132272 177686 132281
rect 177630 132207 177686 132216
rect 185726 132000 185782 132009
rect 185726 131935 185782 131944
rect 185542 131728 185598 131737
rect 185542 131663 185598 131672
rect 177632 131624 177684 131630
rect 177632 131566 177684 131572
rect 177644 131057 177672 131566
rect 177724 131556 177776 131562
rect 177724 131498 177776 131504
rect 177736 131329 177764 131498
rect 177722 131320 177778 131329
rect 177722 131255 177778 131264
rect 177630 131048 177686 131057
rect 177630 130983 177686 130992
rect 185358 130776 185414 130785
rect 185358 130711 185414 130720
rect 185266 130368 185322 130377
rect 185266 130303 185322 130312
rect 177632 130264 177684 130270
rect 177632 130206 177684 130212
rect 177722 130232 177778 130241
rect 177644 129833 177672 130206
rect 177722 130167 177724 130176
rect 177776 130167 177778 130176
rect 177724 130138 177776 130144
rect 177630 129824 177686 129833
rect 177630 129759 177686 129768
rect 185174 129688 185230 129697
rect 185174 129623 185230 129632
rect 185188 128910 185216 129623
rect 177356 128904 177408 128910
rect 177356 128846 177408 128852
rect 185176 128904 185228 128910
rect 185176 128846 185228 128852
rect 177368 128065 177396 128846
rect 185280 128842 185308 130303
rect 177632 128836 177684 128842
rect 177632 128778 177684 128784
rect 185268 128836 185320 128842
rect 185268 128778 185320 128784
rect 177644 128473 177672 128778
rect 185372 128774 185400 130711
rect 185556 130270 185584 131663
rect 185544 130264 185596 130270
rect 185544 130206 185596 130212
rect 185740 130202 185768 131935
rect 185832 131562 185860 133023
rect 185910 132544 185966 132553
rect 185910 132479 185966 132488
rect 185924 131630 185952 132479
rect 185912 131624 185964 131630
rect 185912 131566 185964 131572
rect 185820 131556 185872 131562
rect 185820 131498 185872 131504
rect 185728 130196 185780 130202
rect 185728 130138 185780 130144
rect 185450 129008 185506 129017
rect 185450 128943 185506 128952
rect 177724 128768 177776 128774
rect 177722 128736 177724 128745
rect 185360 128768 185412 128774
rect 177776 128736 177778 128745
rect 185360 128710 185412 128716
rect 177722 128671 177778 128680
rect 177630 128464 177686 128473
rect 177630 128399 177686 128408
rect 185174 128464 185230 128473
rect 185174 128399 185230 128408
rect 177354 128056 177410 128065
rect 177354 127991 177410 128000
rect 185188 127482 185216 128399
rect 185358 127920 185414 127929
rect 185358 127855 185414 127864
rect 185266 127648 185322 127657
rect 185266 127583 185322 127592
rect 177724 127476 177776 127482
rect 177724 127418 177776 127424
rect 185176 127476 185228 127482
rect 185176 127418 185228 127424
rect 177172 127408 177224 127414
rect 177172 127350 177224 127356
rect 177184 127249 177212 127350
rect 177170 127240 177226 127249
rect 177170 127175 177226 127184
rect 177736 126977 177764 127418
rect 177722 126968 177778 126977
rect 177722 126903 177778 126912
rect 185174 126288 185230 126297
rect 182232 126252 182284 126258
rect 185174 126223 185230 126232
rect 182232 126194 182284 126200
rect 177632 126116 177684 126122
rect 177632 126058 177684 126064
rect 177644 125617 177672 126058
rect 177724 126048 177776 126054
rect 177722 126016 177724 126025
rect 177776 126016 177778 126025
rect 177722 125951 177778 125960
rect 177630 125608 177686 125617
rect 177630 125543 177686 125552
rect 177632 124756 177684 124762
rect 177632 124698 177684 124704
rect 177172 124416 177224 124422
rect 177172 124358 177224 124364
rect 177184 124257 177212 124358
rect 177170 124248 177226 124257
rect 177170 124183 177226 124192
rect 177644 123985 177672 124698
rect 182244 124694 182272 126194
rect 185188 126190 185216 126223
rect 182324 126184 182376 126190
rect 182324 126126 182376 126132
rect 185176 126184 185228 126190
rect 185176 126126 185228 126132
rect 177724 124688 177776 124694
rect 177724 124630 177776 124636
rect 182232 124688 182284 124694
rect 182232 124630 182284 124636
rect 177736 124529 177764 124630
rect 177722 124520 177778 124529
rect 177722 124455 177778 124464
rect 182336 124422 182364 126126
rect 185280 126122 185308 127583
rect 185268 126116 185320 126122
rect 185268 126058 185320 126064
rect 185372 126054 185400 127855
rect 185464 127414 185492 128943
rect 185452 127408 185504 127414
rect 185452 127350 185504 127356
rect 185450 126696 185506 126705
rect 185450 126631 185506 126640
rect 185464 126258 185492 126631
rect 185452 126252 185504 126258
rect 185452 126194 185504 126200
rect 185360 126048 185412 126054
rect 185360 125990 185412 125996
rect 185174 125608 185230 125617
rect 185174 125543 185230 125552
rect 185188 124762 185216 125543
rect 185358 124928 185414 124937
rect 185358 124863 185414 124872
rect 185266 124792 185322 124801
rect 185176 124756 185228 124762
rect 185266 124727 185322 124736
rect 185176 124698 185228 124704
rect 182324 124416 182376 124422
rect 182324 124358 182376 124364
rect 177630 123976 177686 123985
rect 177630 123911 177686 123920
rect 185280 123334 185308 124727
rect 177632 123328 177684 123334
rect 177632 123270 177684 123276
rect 185268 123328 185320 123334
rect 185268 123270 185320 123276
rect 177644 122761 177672 123270
rect 185372 123266 185400 124863
rect 185910 123840 185966 123849
rect 185910 123775 185966 123784
rect 185726 123432 185782 123441
rect 185726 123367 185782 123376
rect 177724 123260 177776 123266
rect 177724 123202 177776 123208
rect 185360 123260 185412 123266
rect 185360 123202 185412 123208
rect 177736 123033 177764 123202
rect 177722 123024 177778 123033
rect 177722 122959 177778 122968
rect 177630 122752 177686 122761
rect 177630 122687 177686 122696
rect 185542 122208 185598 122217
rect 185542 122143 185598 122152
rect 177632 121968 177684 121974
rect 177632 121910 177684 121916
rect 177644 121537 177672 121910
rect 177724 121900 177776 121906
rect 177724 121842 177776 121848
rect 177736 121809 177764 121842
rect 177722 121800 177778 121809
rect 177722 121735 177778 121744
rect 177630 121528 177686 121537
rect 177630 121463 177686 121472
rect 185358 121528 185414 121537
rect 185358 121463 185414 121472
rect 185174 120848 185230 120857
rect 182048 120812 182100 120818
rect 185372 120818 185400 121463
rect 185174 120783 185230 120792
rect 185360 120812 185412 120818
rect 182048 120754 182100 120760
rect 181772 120676 181824 120682
rect 181772 120618 181824 120624
rect 177724 120608 177776 120614
rect 177722 120576 177724 120585
rect 177776 120576 177778 120585
rect 177632 120540 177684 120546
rect 177722 120511 177778 120520
rect 177632 120482 177684 120488
rect 177644 120177 177672 120482
rect 177630 120168 177686 120177
rect 177630 120103 177686 120112
rect 177724 119180 177776 119186
rect 177724 119122 177776 119128
rect 177736 119089 177764 119122
rect 177722 119080 177778 119089
rect 177722 119015 177778 119024
rect 181784 118982 181812 120618
rect 182060 119186 182088 120754
rect 182324 120744 182376 120750
rect 182324 120686 182376 120692
rect 182140 119384 182192 119390
rect 182140 119326 182192 119332
rect 182048 119180 182100 119186
rect 182048 119122 182100 119128
rect 177724 118976 177776 118982
rect 177724 118918 177776 118924
rect 181772 118976 181824 118982
rect 181772 118918 181824 118924
rect 177632 118840 177684 118846
rect 177736 118817 177764 118918
rect 177632 118782 177684 118788
rect 177722 118808 177778 118817
rect 177644 118545 177672 118782
rect 177722 118743 177778 118752
rect 177630 118536 177686 118545
rect 177630 118471 177686 118480
rect 181404 117956 181456 117962
rect 181404 117898 181456 117904
rect 177724 117752 177776 117758
rect 177724 117694 177776 117700
rect 177632 117616 177684 117622
rect 177736 117593 177764 117694
rect 177632 117558 177684 117564
rect 177722 117584 177778 117593
rect 177644 117321 177672 117558
rect 177722 117519 177778 117528
rect 177630 117312 177686 117321
rect 177630 117247 177686 117256
rect 178184 116596 178236 116602
rect 178184 116538 178236 116544
rect 176804 116528 176856 116534
rect 176804 116470 176856 116476
rect 175424 115236 175476 115242
rect 175424 115178 175476 115184
rect 174780 115168 174832 115174
rect 174780 115110 174832 115116
rect 145352 114822 145596 114850
rect 146976 114822 147312 114850
rect 145352 111706 145380 114822
rect 147284 113338 147312 114822
rect 148112 114822 148448 114850
rect 149308 114822 149828 114850
rect 150688 114822 151300 114850
rect 152068 114822 152680 114850
rect 153448 114822 154152 114850
rect 154828 114822 155532 114850
rect 156208 114822 157004 114850
rect 158048 114822 158384 114850
rect 159520 114822 159856 114850
rect 160900 114822 161236 114850
rect 161728 114822 162708 114850
rect 163752 114822 164088 114850
rect 164488 114822 165560 114850
rect 166604 114822 166940 114850
rect 168076 114822 168412 114850
rect 169456 114822 169792 114850
rect 170928 114822 171264 114850
rect 172644 114822 172704 114850
rect 147272 113332 147324 113338
rect 147272 113274 147324 113280
rect 145340 111700 145392 111706
rect 145340 111642 145392 111648
rect 148112 111638 148140 114822
rect 148100 111632 148152 111638
rect 148100 111574 148152 111580
rect 143776 102384 143828 102390
rect 143776 102326 143828 102332
rect 142672 101976 142724 101982
rect 142672 101918 142724 101924
rect 143684 101976 143736 101982
rect 143684 101918 143736 101924
rect 142684 99740 142712 101918
rect 143788 99740 143816 102326
rect 144880 102248 144932 102254
rect 144880 102190 144932 102196
rect 144892 99740 144920 102190
rect 145984 102180 146036 102186
rect 145984 102122 146036 102128
rect 145996 99740 146024 102122
rect 147088 102112 147140 102118
rect 147088 102054 147140 102060
rect 147100 99740 147128 102054
rect 148192 102044 148244 102050
rect 148192 101986 148244 101992
rect 148204 99740 148232 101986
rect 149308 99740 149336 114822
rect 150688 101386 150716 114822
rect 152068 101386 152096 114822
rect 150504 101358 150716 101386
rect 151976 101358 152096 101386
rect 153448 101370 153476 114822
rect 154828 101370 154856 114822
rect 156208 101438 156236 114822
rect 158048 111026 158076 114822
rect 158864 111088 158916 111094
rect 158864 111030 158916 111036
rect 156840 111020 156892 111026
rect 156840 110962 156892 110968
rect 158036 111020 158088 111026
rect 158036 110962 158088 110968
rect 158312 111020 158364 111026
rect 158312 110962 158364 110968
rect 154908 101432 154960 101438
rect 154908 101374 154960 101380
rect 156196 101432 156248 101438
rect 156196 101374 156248 101380
rect 152608 101364 152660 101370
rect 150504 99754 150532 101358
rect 151976 99754 152004 101358
rect 152608 101306 152660 101312
rect 153436 101364 153488 101370
rect 153436 101306 153488 101312
rect 153804 101364 153856 101370
rect 153804 101306 153856 101312
rect 154816 101364 154868 101370
rect 154816 101306 154868 101312
rect 150426 99726 150532 99754
rect 151530 99726 152004 99754
rect 152620 99740 152648 101306
rect 153816 99740 153844 101306
rect 154920 99740 154948 101374
rect 156852 101370 156880 110962
rect 158220 101432 158272 101438
rect 158220 101374 158272 101380
rect 156012 101364 156064 101370
rect 156012 101306 156064 101312
rect 156840 101364 156892 101370
rect 156840 101306 156892 101312
rect 157116 101364 157168 101370
rect 157116 101306 157168 101312
rect 156024 99740 156052 101306
rect 157128 99740 157156 101306
rect 158232 99740 158260 101374
rect 158324 101370 158352 110962
rect 158876 101438 158904 111030
rect 159520 111026 159548 114822
rect 160900 111094 160928 114822
rect 160888 111088 160940 111094
rect 160888 111030 160940 111036
rect 159508 111020 159560 111026
rect 159508 110962 159560 110968
rect 161624 111020 161676 111026
rect 161624 110962 161676 110968
rect 159324 102384 159376 102390
rect 159324 102326 159376 102332
rect 158864 101432 158916 101438
rect 158864 101374 158916 101380
rect 158312 101364 158364 101370
rect 158312 101306 158364 101312
rect 159336 99740 159364 102326
rect 161532 102044 161584 102050
rect 161532 101986 161584 101992
rect 160428 101364 160480 101370
rect 160428 101306 160480 101312
rect 160440 99740 160468 101306
rect 161544 99740 161572 101986
rect 161636 101370 161664 110962
rect 161728 102390 161756 114822
rect 163752 111026 163780 114822
rect 163832 111156 163884 111162
rect 163832 111098 163884 111104
rect 163740 111020 163792 111026
rect 163740 110962 163792 110968
rect 161716 102384 161768 102390
rect 161716 102326 161768 102332
rect 163740 101432 163792 101438
rect 163740 101374 163792 101380
rect 161624 101364 161676 101370
rect 161624 101306 161676 101312
rect 162636 101364 162688 101370
rect 162636 101306 162688 101312
rect 162648 99740 162676 101306
rect 163752 99740 163780 101374
rect 163844 101370 163872 111098
rect 164488 102050 164516 114822
rect 166604 111162 166632 114822
rect 166592 111156 166644 111162
rect 166592 111098 166644 111104
rect 167880 111156 167932 111162
rect 167880 111098 167932 111104
rect 166500 111088 166552 111094
rect 166500 111030 166552 111036
rect 165120 111020 165172 111026
rect 165120 110962 165172 110968
rect 164476 102044 164528 102050
rect 164476 101986 164528 101992
rect 165132 101438 165160 110962
rect 165120 101432 165172 101438
rect 165120 101374 165172 101380
rect 165948 101432 166000 101438
rect 165948 101374 166000 101380
rect 163832 101364 163884 101370
rect 163832 101306 163884 101312
rect 164844 101364 164896 101370
rect 164844 101306 164896 101312
rect 164856 99740 164884 101306
rect 165960 99740 165988 101374
rect 166512 101370 166540 111030
rect 167144 101976 167196 101982
rect 167144 101918 167196 101924
rect 166500 101364 166552 101370
rect 166500 101306 166552 101312
rect 167156 99740 167184 101918
rect 167892 101438 167920 111098
rect 168076 111026 168104 114822
rect 169456 111094 169484 114822
rect 169904 112380 169956 112386
rect 169904 112322 169956 112328
rect 169444 111088 169496 111094
rect 169444 111030 169496 111036
rect 168064 111020 168116 111026
rect 168064 110962 168116 110968
rect 167880 101432 167932 101438
rect 167880 101374 167932 101380
rect 169916 99890 169944 112322
rect 170928 111162 170956 114822
rect 170916 111156 170968 111162
rect 170916 111098 170968 111104
rect 172676 111026 172704 114822
rect 172664 111020 172716 111026
rect 172664 110962 172716 110968
rect 172664 102112 172716 102118
rect 172664 102054 172716 102060
rect 171560 102044 171612 102050
rect 171560 101986 171612 101992
rect 170456 101976 170508 101982
rect 170456 101918 170508 101924
rect 169732 99862 169944 99890
rect 169732 99754 169760 99862
rect 169378 99726 169760 99754
rect 170468 99740 170496 101918
rect 171572 99740 171600 101986
rect 172676 99740 172704 102054
rect 174792 101370 174820 115110
rect 173768 101364 173820 101370
rect 173768 101306 173820 101312
rect 174780 101364 174832 101370
rect 174780 101306 174832 101312
rect 173780 99740 173808 101306
rect 175436 99618 175464 115178
rect 176160 111020 176212 111026
rect 176160 110962 176212 110968
rect 176172 101438 176200 110962
rect 176160 101432 176212 101438
rect 176160 101374 176212 101380
rect 176816 101370 176844 116470
rect 177080 116460 177132 116466
rect 177080 116402 177132 116408
rect 177092 115553 177120 116402
rect 177724 116392 177776 116398
rect 177722 116360 177724 116369
rect 177776 116360 177778 116369
rect 177722 116295 177778 116304
rect 177724 116120 177776 116126
rect 177724 116062 177776 116068
rect 177736 115961 177764 116062
rect 177722 115952 177778 115961
rect 177722 115887 177778 115896
rect 177078 115544 177134 115553
rect 177078 115479 177134 115488
rect 178196 101370 178224 116538
rect 181416 116398 181444 117898
rect 182152 117758 182180 119326
rect 182232 119316 182284 119322
rect 182232 119258 182284 119264
rect 182140 117752 182192 117758
rect 182140 117694 182192 117700
rect 182244 117622 182272 119258
rect 182336 118846 182364 120686
rect 185188 120682 185216 120783
rect 185360 120754 185412 120760
rect 185268 120744 185320 120750
rect 185266 120712 185268 120721
rect 185320 120712 185322 120721
rect 185176 120676 185228 120682
rect 185266 120647 185322 120656
rect 185176 120618 185228 120624
rect 185556 120546 185584 122143
rect 185740 121974 185768 123367
rect 185818 122616 185874 122625
rect 185818 122551 185874 122560
rect 185728 121968 185780 121974
rect 185728 121910 185780 121916
rect 185832 120614 185860 122551
rect 185924 121906 185952 123775
rect 185912 121900 185964 121906
rect 185912 121842 185964 121848
rect 185820 120608 185872 120614
rect 185820 120550 185872 120556
rect 185544 120540 185596 120546
rect 185544 120482 185596 120488
rect 185266 119760 185322 119769
rect 185266 119695 185322 119704
rect 185280 119390 185308 119695
rect 185268 119384 185320 119390
rect 185174 119352 185230 119361
rect 185268 119326 185320 119332
rect 185174 119287 185176 119296
rect 185228 119287 185230 119296
rect 185176 119258 185228 119264
rect 182324 118840 182376 118846
rect 182324 118782 182376 118788
rect 185266 118536 185322 118545
rect 185266 118471 185322 118480
rect 185174 117992 185230 118001
rect 185280 117962 185308 118471
rect 185174 117927 185230 117936
rect 185268 117956 185320 117962
rect 185188 117894 185216 117927
rect 185268 117898 185320 117904
rect 182324 117888 182376 117894
rect 182324 117830 182376 117836
rect 185176 117888 185228 117894
rect 185176 117830 185228 117836
rect 182232 117616 182284 117622
rect 182232 117558 182284 117564
rect 181404 116392 181456 116398
rect 181404 116334 181456 116340
rect 182336 116126 182364 117830
rect 185358 117448 185414 117457
rect 185358 117383 185414 117392
rect 185266 116768 185322 116777
rect 185266 116703 185322 116712
rect 185280 116602 185308 116703
rect 185268 116596 185320 116602
rect 185268 116538 185320 116544
rect 185176 116528 185228 116534
rect 185174 116496 185176 116505
rect 185228 116496 185230 116505
rect 185372 116466 185400 117383
rect 185174 116431 185230 116440
rect 185360 116460 185412 116466
rect 185360 116402 185412 116408
rect 182324 116120 182376 116126
rect 182324 116062 182376 116068
rect 185266 115680 185322 115689
rect 185266 115615 185322 115624
rect 185174 115272 185230 115281
rect 185280 115242 185308 115615
rect 185174 115207 185230 115216
rect 185268 115236 185320 115242
rect 185188 115174 185216 115207
rect 185268 115178 185320 115184
rect 185176 115168 185228 115174
rect 185176 115110 185228 115116
rect 185818 114456 185874 114465
rect 185818 114391 185874 114400
rect 185174 112688 185230 112697
rect 185174 112623 185230 112632
rect 185188 112386 185216 112623
rect 185176 112380 185228 112386
rect 185176 112322 185228 112328
rect 183612 110408 183664 110414
rect 183612 110350 183664 110356
rect 183520 110272 183572 110278
rect 183520 110214 183572 110220
rect 183336 109864 183388 109870
rect 183336 109806 183388 109812
rect 183244 109796 183296 109802
rect 183244 109738 183296 109744
rect 183152 109728 183204 109734
rect 183152 109670 183204 109676
rect 183060 109660 183112 109666
rect 183060 109602 183112 109608
rect 179288 101432 179340 101438
rect 179288 101374 179340 101380
rect 175976 101364 176028 101370
rect 175976 101306 176028 101312
rect 176804 101364 176856 101370
rect 176804 101306 176856 101312
rect 177080 101364 177132 101370
rect 177080 101306 177132 101312
rect 178184 101364 178236 101370
rect 178184 101306 178236 101312
rect 175988 99740 176016 101306
rect 177092 99740 177120 101306
rect 179300 99740 179328 101374
rect 174898 99590 175464 99618
rect 183072 90665 183100 109602
rect 183164 91889 183192 109670
rect 183256 93113 183284 109738
rect 183348 95561 183376 109806
rect 183428 109592 183480 109598
rect 183428 109534 183480 109540
rect 183334 95552 183390 95561
rect 183334 95487 183390 95496
rect 183440 94337 183468 109534
rect 183532 96785 183560 110214
rect 183624 98009 183652 110350
rect 183704 110340 183756 110346
rect 183704 110282 183756 110288
rect 183716 99233 183744 110282
rect 185832 102118 185860 114391
rect 186002 113912 186058 113921
rect 186002 113847 186058 113856
rect 185820 102112 185872 102118
rect 185820 102054 185872 102060
rect 186016 102050 186044 113847
rect 186186 113776 186242 113785
rect 186186 113711 186242 113720
rect 186004 102044 186056 102050
rect 186004 101986 186056 101992
rect 186200 101982 186228 113711
rect 198068 113054 198450 113082
rect 207636 113054 208202 113082
rect 209384 113054 209858 113082
rect 188224 109666 188252 112932
rect 188776 109734 188804 112932
rect 189328 109802 189356 112932
rect 189316 109796 189368 109802
rect 189316 109738 189368 109744
rect 188764 109728 188816 109734
rect 188764 109670 188816 109676
rect 188212 109660 188264 109666
rect 188212 109602 188264 109608
rect 189880 109598 189908 112932
rect 190432 109870 190460 112932
rect 191076 110278 191104 112932
rect 191628 110414 191656 112932
rect 191616 110408 191668 110414
rect 191616 110350 191668 110356
rect 192180 110346 192208 112932
rect 192746 112918 193036 112946
rect 193298 112918 193404 112946
rect 193008 112538 193036 112918
rect 193008 112510 193312 112538
rect 192168 110340 192220 110346
rect 192168 110282 192220 110288
rect 191064 110272 191116 110278
rect 191064 110214 191116 110220
rect 191984 110272 192036 110278
rect 191984 110214 192036 110220
rect 190420 109864 190472 109870
rect 190420 109806 190472 109812
rect 189868 109592 189920 109598
rect 189868 109534 189920 109540
rect 186188 101976 186240 101982
rect 186188 101918 186240 101924
rect 183702 99224 183758 99233
rect 183702 99159 183758 99168
rect 191996 98825 192024 110214
rect 193284 102662 193312 112510
rect 193272 102656 193324 102662
rect 193272 102598 193324 102604
rect 193376 101438 193404 112918
rect 193928 109598 193956 112932
rect 194494 112918 194692 112946
rect 193916 109592 193968 109598
rect 193916 109534 193968 109540
rect 194100 102656 194152 102662
rect 194100 102598 194152 102604
rect 193364 101432 193416 101438
rect 193364 101374 193416 101380
rect 194112 99740 194140 102598
rect 194664 101506 194692 112918
rect 194940 112918 195046 112946
rect 195124 112918 195598 112946
rect 194744 109592 194796 109598
rect 194744 109534 194796 109540
rect 194652 101500 194704 101506
rect 194652 101442 194704 101448
rect 194756 101438 194784 109534
rect 194468 101432 194520 101438
rect 194468 101374 194520 101380
rect 194744 101432 194796 101438
rect 194744 101374 194796 101380
rect 194480 99740 194508 101374
rect 194940 101370 194968 112918
rect 195124 101438 195152 112918
rect 195296 101500 195348 101506
rect 195296 101442 195348 101448
rect 195020 101432 195072 101438
rect 195020 101374 195072 101380
rect 195112 101432 195164 101438
rect 195112 101374 195164 101380
rect 194928 101364 194980 101370
rect 194928 101306 194980 101312
rect 195032 99618 195060 101374
rect 195308 99740 195336 101442
rect 196032 101432 196084 101438
rect 196032 101374 196084 101380
rect 195664 101364 195716 101370
rect 195664 101306 195716 101312
rect 195676 99740 195704 101306
rect 196044 99740 196072 101374
rect 196136 101352 196164 112932
rect 196320 112918 196794 112946
rect 197056 112918 197346 112946
rect 197608 112918 197898 112946
rect 196320 102662 196348 112918
rect 196308 102656 196360 102662
rect 196308 102598 196360 102604
rect 196860 102656 196912 102662
rect 196860 102598 196912 102604
rect 196136 101324 196256 101352
rect 196228 99754 196256 101324
rect 196228 99726 196518 99754
rect 196872 99740 196900 102598
rect 197056 99754 197084 112918
rect 197608 99754 197636 112918
rect 198068 112674 198096 113054
rect 199002 112918 199200 112946
rect 197976 112646 198096 112674
rect 197976 99754 198004 112646
rect 199172 102662 199200 112918
rect 199264 112918 199646 112946
rect 199724 112918 200198 112946
rect 200368 112918 200750 112946
rect 201012 112918 201302 112946
rect 201748 112918 201854 112946
rect 198424 102656 198476 102662
rect 198424 102598 198476 102604
rect 199160 102656 199212 102662
rect 199160 102598 199212 102604
rect 197056 99726 197254 99754
rect 197608 99726 197714 99754
rect 197976 99726 198082 99754
rect 198436 99740 198464 102598
rect 199264 102202 199292 112918
rect 199620 102656 199672 102662
rect 199620 102598 199672 102604
rect 198896 102174 199292 102202
rect 198896 99740 198924 102174
rect 199252 102112 199304 102118
rect 199252 102054 199304 102060
rect 199264 99740 199292 102054
rect 199632 99740 199660 102598
rect 199724 102118 199752 112918
rect 200368 102662 200396 112918
rect 201012 112674 201040 112918
rect 200644 112646 201040 112674
rect 200356 102656 200408 102662
rect 200356 102598 200408 102604
rect 200644 102594 200672 112646
rect 201748 109682 201776 112918
rect 201460 109660 201512 109666
rect 201460 109602 201512 109608
rect 201564 109654 201776 109682
rect 202484 109666 202512 112932
rect 202472 109660 202524 109666
rect 201472 102746 201500 109602
rect 201380 102718 201500 102746
rect 201380 102662 201408 102718
rect 200816 102656 200868 102662
rect 200816 102598 200868 102604
rect 201368 102656 201420 102662
rect 201368 102598 201420 102604
rect 201460 102656 201512 102662
rect 201460 102598 201512 102604
rect 200080 102588 200132 102594
rect 200080 102530 200132 102536
rect 200632 102588 200684 102594
rect 200632 102530 200684 102536
rect 199712 102112 199764 102118
rect 199712 102054 199764 102060
rect 200092 99740 200120 102530
rect 200448 102248 200500 102254
rect 200448 102190 200500 102196
rect 200460 99740 200488 102190
rect 200828 99740 200856 102598
rect 201276 102588 201328 102594
rect 201276 102530 201328 102536
rect 201288 99740 201316 102530
rect 194862 99590 195060 99618
rect 201472 99618 201500 102598
rect 201564 102254 201592 109654
rect 202472 109602 202524 109608
rect 203036 109598 203064 112932
rect 203128 112918 203602 112946
rect 203772 112918 204154 112946
rect 201644 109592 201696 109598
rect 201644 109534 201696 109540
rect 203024 109592 203076 109598
rect 203024 109534 203076 109540
rect 201656 102594 201684 109534
rect 203128 102662 203156 112918
rect 203772 112674 203800 112918
rect 203220 112646 203800 112674
rect 203116 102656 203168 102662
rect 203116 102598 203168 102604
rect 201644 102588 201696 102594
rect 201644 102530 201696 102536
rect 202472 102452 202524 102458
rect 202472 102394 202524 102400
rect 201552 102248 201604 102254
rect 201552 102190 201604 102196
rect 202104 102112 202156 102118
rect 202104 102054 202156 102060
rect 202116 99740 202144 102054
rect 202484 99740 202512 102394
rect 203220 102118 203248 112646
rect 203760 109728 203812 109734
rect 203760 109670 203812 109676
rect 203300 102588 203352 102594
rect 203300 102530 203352 102536
rect 203208 102112 203260 102118
rect 203208 102054 203260 102060
rect 202840 101704 202892 101710
rect 202840 101646 202892 101652
rect 202852 99740 202880 101646
rect 203312 99740 203340 102530
rect 203772 101710 203800 109670
rect 204692 109598 204720 112932
rect 205232 109796 205284 109802
rect 205232 109738 205284 109744
rect 205140 109660 205192 109666
rect 205140 109602 205192 109608
rect 203852 109592 203904 109598
rect 203852 109534 203904 109540
rect 204680 109592 204732 109598
rect 204680 109534 204732 109540
rect 203864 102458 203892 109534
rect 204864 102656 204916 102662
rect 204864 102598 204916 102604
rect 203852 102452 203904 102458
rect 203852 102394 203904 102400
rect 204036 102112 204088 102118
rect 204036 102054 204088 102060
rect 203760 101704 203812 101710
rect 203760 101646 203812 101652
rect 203668 101500 203720 101506
rect 203668 101442 203720 101448
rect 203680 99740 203708 101442
rect 204048 99740 204076 102054
rect 204496 101704 204548 101710
rect 204496 101646 204548 101652
rect 204508 99740 204536 101646
rect 204876 99740 204904 102598
rect 205152 101506 205180 109602
rect 205244 102118 205272 109738
rect 205336 109734 205364 112932
rect 205324 109728 205376 109734
rect 205324 109670 205376 109676
rect 205888 109598 205916 112932
rect 206440 109666 206468 112932
rect 206992 109802 207020 112932
rect 207268 112918 207558 112946
rect 206980 109796 207032 109802
rect 206980 109738 207032 109744
rect 206428 109660 206480 109666
rect 206428 109602 206480 109608
rect 205416 109592 205468 109598
rect 205416 109534 205468 109540
rect 205876 109592 205928 109598
rect 205876 109534 205928 109540
rect 205428 102594 205456 109534
rect 205416 102588 205468 102594
rect 205416 102530 205468 102536
rect 206428 102588 206480 102594
rect 206428 102530 206480 102536
rect 206060 102384 206112 102390
rect 206060 102326 206112 102332
rect 205232 102112 205284 102118
rect 205232 102054 205284 102060
rect 205232 101840 205284 101846
rect 205232 101782 205284 101788
rect 205140 101500 205192 101506
rect 205140 101442 205192 101448
rect 205244 99740 205272 101782
rect 205692 101500 205744 101506
rect 205692 101442 205744 101448
rect 205704 99740 205732 101442
rect 206072 99740 206100 102326
rect 206440 99740 206468 102530
rect 206888 101772 206940 101778
rect 206888 101714 206940 101720
rect 206900 99740 206928 101714
rect 207268 101710 207296 112918
rect 207636 112674 207664 113054
rect 207360 112646 207664 112674
rect 207360 102662 207388 112646
rect 208268 110340 208320 110346
rect 208268 110282 208320 110288
rect 208176 109728 208228 109734
rect 208176 109670 208228 109676
rect 207348 102656 207400 102662
rect 207348 102598 207400 102604
rect 207256 101704 207308 101710
rect 207256 101646 207308 101652
rect 208188 101574 208216 109670
rect 207624 101568 207676 101574
rect 207624 101510 207676 101516
rect 208176 101568 208228 101574
rect 208176 101510 208228 101516
rect 207256 101432 207308 101438
rect 207256 101374 207308 101380
rect 207268 99740 207296 101374
rect 207636 99740 207664 101510
rect 208084 101364 208136 101370
rect 208084 101306 208136 101312
rect 208096 99740 208124 101306
rect 208280 99754 208308 110282
rect 208360 109660 208412 109666
rect 208360 109602 208412 109608
rect 208372 101370 208400 109602
rect 208544 109592 208596 109598
rect 208544 109534 208596 109540
rect 208556 101438 208584 109534
rect 208636 107552 208688 107558
rect 208636 107494 208688 107500
rect 208648 101506 208676 107494
rect 208740 101846 208768 112932
rect 209016 112918 209306 112946
rect 209016 107558 209044 112918
rect 209384 112674 209412 113054
rect 209108 112646 209412 112674
rect 210120 112918 210410 112946
rect 210672 112918 211054 112946
rect 209004 107552 209056 107558
rect 209004 107494 209056 107500
rect 209108 107370 209136 112646
rect 210016 107552 210068 107558
rect 210016 107494 210068 107500
rect 208832 107342 209136 107370
rect 208832 102390 208860 107342
rect 208820 102384 208872 102390
rect 208820 102326 208872 102332
rect 208820 102248 208872 102254
rect 208820 102190 208872 102196
rect 208728 101840 208780 101846
rect 208728 101782 208780 101788
rect 208636 101500 208688 101506
rect 208636 101442 208688 101448
rect 208544 101432 208596 101438
rect 208544 101374 208596 101380
rect 208360 101364 208412 101370
rect 208360 101306 208412 101312
rect 208280 99726 208478 99754
rect 208832 99740 208860 102190
rect 209280 102112 209332 102118
rect 209280 102054 209332 102060
rect 209292 99740 209320 102054
rect 209648 102044 209700 102050
rect 209648 101986 209700 101992
rect 209660 99740 209688 101986
rect 210028 101778 210056 107494
rect 210120 102594 210148 112918
rect 210672 107558 210700 112918
rect 211592 109598 211620 112932
rect 212144 109734 212172 112932
rect 212132 109728 212184 109734
rect 212132 109670 212184 109676
rect 212696 109666 212724 112932
rect 213248 110346 213276 112932
rect 213340 112918 213906 112946
rect 213236 110340 213288 110346
rect 213236 110282 213288 110288
rect 212684 109660 212736 109666
rect 212684 109602 212736 109608
rect 211580 109592 211632 109598
rect 211580 109534 211632 109540
rect 210660 107552 210712 107558
rect 213340 107506 213368 112918
rect 213512 109660 213564 109666
rect 213512 109602 213564 109608
rect 213420 109592 213472 109598
rect 213420 109534 213472 109540
rect 210660 107494 210712 107500
rect 212880 107478 213368 107506
rect 210108 102588 210160 102594
rect 210108 102530 210160 102536
rect 212880 102254 212908 107478
rect 212868 102248 212920 102254
rect 212868 102190 212920 102196
rect 213432 102118 213460 109534
rect 213420 102112 213472 102118
rect 213420 102054 213472 102060
rect 213524 102050 213552 109602
rect 214444 109598 214472 112932
rect 214996 109666 215024 112932
rect 215548 110278 215576 112932
rect 215536 110272 215588 110278
rect 215536 110214 215588 110220
rect 214984 109660 215036 109666
rect 214984 109602 215036 109608
rect 214432 109592 214484 109598
rect 214432 109534 214484 109540
rect 213512 102044 213564 102050
rect 213512 101986 213564 101992
rect 210016 101772 210068 101778
rect 210016 101714 210068 101720
rect 212040 99936 212092 99942
rect 212040 99878 212092 99884
rect 201472 99590 201670 99618
rect 191982 98816 192038 98825
rect 191982 98751 192038 98760
rect 183610 98000 183666 98009
rect 183610 97935 183666 97944
rect 211764 97148 211816 97154
rect 211764 97090 211816 97096
rect 209830 96912 209886 96921
rect 209752 96870 209830 96898
rect 183518 96776 183574 96785
rect 183518 96711 183574 96720
rect 191982 94736 192038 94745
rect 191982 94671 192038 94680
rect 191996 94434 192024 94671
rect 188580 94428 188632 94434
rect 188580 94370 188632 94376
rect 191984 94428 192036 94434
rect 191984 94370 192036 94376
rect 183426 94328 183482 94337
rect 183426 94263 183482 94272
rect 183242 93104 183298 93113
rect 183242 93039 183298 93048
rect 183150 91880 183206 91889
rect 183150 91815 183206 91824
rect 183058 90656 183114 90665
rect 183058 90591 183114 90600
rect 188592 90218 188620 94370
rect 191154 92832 191210 92841
rect 191154 92767 191210 92776
rect 190786 90792 190842 90801
rect 190786 90727 190842 90736
rect 182876 90212 182928 90218
rect 182876 90154 182928 90160
rect 188580 90212 188632 90218
rect 188580 90154 188632 90160
rect 182888 89441 182916 90154
rect 182874 89432 182930 89441
rect 182874 89367 182930 89376
rect 183520 88852 183572 88858
rect 183520 88794 183572 88800
rect 183532 88217 183560 88794
rect 183518 88208 183574 88217
rect 183518 88143 183574 88152
rect 190800 87498 190828 90727
rect 191168 88858 191196 92767
rect 191156 88852 191208 88858
rect 191156 88794 191208 88800
rect 191706 88752 191762 88761
rect 191706 88687 191762 88696
rect 183704 87492 183756 87498
rect 183704 87434 183756 87440
rect 190788 87492 190840 87498
rect 190788 87434 190840 87440
rect 183716 87129 183744 87434
rect 183702 87120 183758 87129
rect 183702 87055 183758 87064
rect 191614 86848 191670 86857
rect 191614 86783 191670 86792
rect 183704 86064 183756 86070
rect 183704 86006 183756 86012
rect 183716 85905 183744 86006
rect 183702 85896 183758 85905
rect 183702 85831 183758 85840
rect 182508 84704 182560 84710
rect 182508 84646 182560 84652
rect 183702 84672 183758 84681
rect 182520 83457 182548 84646
rect 191628 84642 191656 86783
rect 191720 86070 191748 88687
rect 191708 86064 191760 86070
rect 191708 86006 191760 86012
rect 191982 84808 192038 84817
rect 191982 84743 192038 84752
rect 191996 84710 192024 84743
rect 191984 84704 192036 84710
rect 191984 84646 192036 84652
rect 183702 84607 183704 84616
rect 183756 84607 183758 84616
rect 191616 84636 191668 84642
rect 183704 84578 183756 84584
rect 191616 84578 191668 84584
rect 182506 83448 182562 83457
rect 182506 83383 182562 83392
rect 191982 82768 192038 82777
rect 191982 82703 192038 82712
rect 191996 82670 192024 82703
rect 183704 82664 183756 82670
rect 183704 82606 183756 82612
rect 191984 82664 192036 82670
rect 191984 82606 192036 82612
rect 183716 82233 183744 82606
rect 183702 82224 183758 82233
rect 183702 82159 183758 82168
rect 183244 81304 183296 81310
rect 183244 81246 183296 81252
rect 191892 81304 191944 81310
rect 191892 81246 191944 81252
rect 183256 81009 183284 81246
rect 183242 81000 183298 81009
rect 183242 80935 183298 80944
rect 191904 80873 191932 81246
rect 191890 80864 191946 80873
rect 191890 80799 191946 80808
rect 136876 80556 136928 80562
rect 136876 80498 136928 80504
rect 136888 80465 136916 80498
rect 136874 80456 136930 80465
rect 136874 80391 136930 80400
rect 183702 79776 183758 79785
rect 183702 79711 183758 79720
rect 183716 79270 183744 79711
rect 183704 79264 183756 79270
rect 183704 79206 183756 79212
rect 191984 79196 192036 79202
rect 191984 79138 192036 79144
rect 191996 78833 192024 79138
rect 191982 78824 192038 78833
rect 191982 78759 192038 78768
rect 183518 78552 183574 78561
rect 183518 78487 183574 78496
rect 183532 77910 183560 78487
rect 183520 77904 183572 77910
rect 183520 77846 183572 77852
rect 191984 77904 192036 77910
rect 191984 77846 192036 77852
rect 183058 77328 183114 77337
rect 183058 77263 183114 77272
rect 183072 76482 183100 77263
rect 191996 76793 192024 77846
rect 209752 76906 209780 96870
rect 209830 96847 209886 96856
rect 211776 96513 211804 97090
rect 211762 96504 211818 96513
rect 211762 96439 211818 96448
rect 211856 90212 211908 90218
rect 211856 90154 211908 90160
rect 211868 89849 211896 90154
rect 211854 89840 211910 89849
rect 211854 89775 211910 89784
rect 212052 83185 212080 99878
rect 216192 97154 216220 204802
rect 217572 190654 217600 231050
rect 220318 215232 220374 215241
rect 220318 215167 220374 215176
rect 218294 209656 218350 209665
rect 218294 209591 218350 209600
rect 217560 190648 217612 190654
rect 217560 190590 217612 190596
rect 216272 176368 216324 176374
rect 216272 176310 216324 176316
rect 216284 127482 216312 176310
rect 218308 165290 218336 209591
rect 218296 165284 218348 165290
rect 218296 165226 218348 165232
rect 218296 163652 218348 163658
rect 218296 163594 218348 163600
rect 216916 156512 216968 156518
rect 216916 156454 216968 156460
rect 216272 127476 216324 127482
rect 216272 127418 216324 127424
rect 216928 117321 216956 156454
rect 218308 127385 218336 163594
rect 218386 135944 218442 135953
rect 218386 135879 218442 135888
rect 218294 127376 218350 127385
rect 218294 127311 218350 127320
rect 216914 117312 216970 117321
rect 216914 117247 216970 117256
rect 217558 117312 217614 117321
rect 217558 117247 217614 117256
rect 216180 97148 216232 97154
rect 216180 97090 216232 97096
rect 212038 83176 212094 83185
rect 212038 83111 212094 83120
rect 209830 76920 209886 76929
rect 209752 76878 209830 76906
rect 209830 76855 209886 76864
rect 191982 76784 192038 76793
rect 191982 76719 192038 76728
rect 183060 76476 183112 76482
rect 183060 76418 183112 76424
rect 185176 76476 185228 76482
rect 185176 76418 185228 76424
rect 183242 76104 183298 76113
rect 183242 76039 183298 76048
rect 183256 75122 183284 76039
rect 183244 75116 183296 75122
rect 183244 75058 183296 75064
rect 185188 75054 185216 76418
rect 186004 75116 186056 75122
rect 186004 75058 186056 75064
rect 185176 75048 185228 75054
rect 185176 74990 185228 74996
rect 183702 74880 183758 74889
rect 183702 74815 183758 74824
rect 183716 73898 183744 74815
rect 183704 73892 183756 73898
rect 183704 73834 183756 73840
rect 183702 73792 183758 73801
rect 183702 73727 183704 73736
rect 183756 73727 183758 73736
rect 183704 73698 183756 73704
rect 186016 73694 186044 75058
rect 191524 75048 191576 75054
rect 191524 74990 191576 74996
rect 191536 74753 191564 74990
rect 191522 74744 191578 74753
rect 191522 74679 191578 74688
rect 217572 73830 217600 117247
rect 218400 113338 218428 135879
rect 218388 113332 218440 113338
rect 218388 113274 218440 113280
rect 217560 73824 217612 73830
rect 217560 73766 217612 73772
rect 188488 73756 188540 73762
rect 188488 73698 188540 73704
rect 190788 73756 190840 73762
rect 190788 73698 190840 73704
rect 186004 73688 186056 73694
rect 186004 73630 186056 73636
rect 183702 72568 183758 72577
rect 183758 72526 183836 72554
rect 183702 72503 183758 72512
rect 183702 71344 183758 71353
rect 183702 71279 183758 71288
rect 183716 70974 183744 71279
rect 183704 70968 183756 70974
rect 183704 70910 183756 70916
rect 128504 70220 128556 70226
rect 128504 70162 128556 70168
rect 134024 70220 134076 70226
rect 134024 70162 134076 70168
rect 136876 70220 136928 70226
rect 136876 70162 136928 70168
rect 128516 69857 128544 70162
rect 128502 69848 128558 69857
rect 128502 69783 128558 69792
rect 106608 68180 106660 68186
rect 106608 68122 106660 68128
rect 106620 67953 106648 68122
rect 106606 67944 106662 67953
rect 106606 67879 106662 67888
rect 136888 66593 136916 70162
rect 182874 70120 182930 70129
rect 182874 70055 182930 70064
rect 182888 69954 182916 70055
rect 182876 69948 182928 69954
rect 182876 69890 182928 69896
rect 183058 68896 183114 68905
rect 183058 68831 183114 68840
rect 136874 66584 136930 66593
rect 136874 66519 136930 66528
rect 106514 65632 106570 65641
rect 106514 65567 106570 65576
rect 104492 63692 104544 63698
rect 104492 63634 104544 63640
rect 106608 63692 106660 63698
rect 106608 63634 106660 63640
rect 106620 63329 106648 63634
rect 106606 63320 106662 63329
rect 106606 63255 106662 63264
rect 104400 61244 104452 61250
rect 104400 61186 104452 61192
rect 107160 61244 107212 61250
rect 107160 61186 107212 61192
rect 107172 61017 107200 61186
rect 107158 61008 107214 61017
rect 107158 60943 107214 60952
rect 182690 60464 182746 60473
rect 182690 60399 182692 60408
rect 182744 60399 182746 60408
rect 182692 60370 182744 60376
rect 109092 57436 109144 57442
rect 109092 57378 109144 57384
rect 105320 50092 105372 50098
rect 105320 50034 105372 50040
rect 104216 49004 104268 49010
rect 104216 48946 104268 48952
rect 103020 48936 103072 48942
rect 103020 48878 103072 48884
rect 104228 46700 104256 48946
rect 104768 48936 104820 48942
rect 104768 48878 104820 48884
rect 104780 46700 104808 48878
rect 105332 46700 105360 50034
rect 106424 50024 106476 50030
rect 106424 49966 106476 49972
rect 105872 49956 105924 49962
rect 105872 49898 105924 49904
rect 105884 46700 105912 49898
rect 106436 46700 106464 49966
rect 106976 49752 107028 49758
rect 106976 49694 107028 49700
rect 106988 46700 107016 49694
rect 107528 49616 107580 49622
rect 107528 49558 107580 49564
rect 107540 46700 107568 49558
rect 108080 49548 108132 49554
rect 108080 49490 108132 49496
rect 108092 46700 108120 49490
rect 108632 49004 108684 49010
rect 108632 48946 108684 48952
rect 108644 46700 108672 48946
rect 109104 48346 109132 57378
rect 110116 57170 110144 59892
rect 110484 57442 110512 59892
rect 110668 59878 110866 59906
rect 110944 59878 111326 59906
rect 110472 57436 110524 57442
rect 110472 57378 110524 57384
rect 110668 57322 110696 59878
rect 110484 57294 110696 57322
rect 109184 57164 109236 57170
rect 109184 57106 109236 57112
rect 110104 57164 110156 57170
rect 110104 57106 110156 57112
rect 109196 49010 109224 57106
rect 110484 49010 110512 57294
rect 110944 57186 110972 59878
rect 110576 57158 110972 57186
rect 111680 57170 111708 59892
rect 111668 57164 111720 57170
rect 109184 49004 109236 49010
rect 109184 48946 109236 48952
rect 109736 49004 109788 49010
rect 109736 48946 109788 48952
rect 110472 49004 110524 49010
rect 110472 48946 110524 48952
rect 109104 48318 109224 48346
rect 109196 46700 109224 48318
rect 109748 46700 109776 48946
rect 110576 46714 110604 57158
rect 112048 57152 112076 59892
rect 111668 57106 111720 57112
rect 111956 57124 112076 57152
rect 112232 59878 112522 59906
rect 110656 57096 110708 57102
rect 110656 57038 110708 57044
rect 110314 46686 110604 46714
rect 110668 46714 110696 57038
rect 111956 46986 111984 57124
rect 111864 46958 111984 46986
rect 111864 46714 111892 46958
rect 112232 46714 112260 59878
rect 112876 57238 112904 59892
rect 112864 57232 112916 57238
rect 112864 57174 112916 57180
rect 113244 57170 113272 59892
rect 113428 59878 113718 59906
rect 112588 57164 112640 57170
rect 112588 57106 112640 57112
rect 112772 57164 112824 57170
rect 112772 57106 112824 57112
rect 113232 57164 113284 57170
rect 113232 57106 113284 57112
rect 112600 57050 112628 57106
rect 112508 57022 112628 57050
rect 112508 47514 112536 57022
rect 112496 47508 112548 47514
rect 112496 47450 112548 47456
rect 112588 47508 112640 47514
rect 112588 47450 112640 47456
rect 110668 46686 110866 46714
rect 111510 46686 111892 46714
rect 112062 46686 112260 46714
rect 112600 46700 112628 47450
rect 112784 46714 112812 57106
rect 113428 46714 113456 59878
rect 114072 57170 114100 59892
rect 114440 57170 114468 59892
rect 113508 57164 113560 57170
rect 113508 57106 113560 57112
rect 114060 57164 114112 57170
rect 114060 57106 114112 57112
rect 114428 57164 114480 57170
rect 114428 57106 114480 57112
rect 113520 46986 113548 57106
rect 114900 50370 114928 59892
rect 115282 59878 115480 59906
rect 114980 57164 115032 57170
rect 114980 57106 115032 57112
rect 114888 50364 114940 50370
rect 114888 50306 114940 50312
rect 114992 50302 115020 57106
rect 114980 50296 115032 50302
rect 114980 50238 115032 50244
rect 114980 50160 115032 50166
rect 114980 50102 115032 50108
rect 115072 50160 115124 50166
rect 115072 50102 115124 50108
rect 113520 46958 113916 46986
rect 113888 46714 113916 46958
rect 114992 46714 115020 50102
rect 112784 46686 113166 46714
rect 113428 46686 113718 46714
rect 113888 46686 114270 46714
rect 114822 46686 115020 46714
rect 115084 46714 115112 50102
rect 115452 46714 115480 59878
rect 115636 57170 115664 59892
rect 116096 57238 116124 59892
rect 116464 58122 116492 59892
rect 116452 58116 116504 58122
rect 116452 58058 116504 58064
rect 116084 57232 116136 57238
rect 116084 57174 116136 57180
rect 116636 57232 116688 57238
rect 116636 57174 116688 57180
rect 115624 57164 115676 57170
rect 115624 57106 115676 57112
rect 116268 57164 116320 57170
rect 116268 57106 116320 57112
rect 116280 46714 116308 57106
rect 116648 46714 116676 57174
rect 116832 57170 116860 59892
rect 117292 57646 117320 59892
rect 117674 59878 118056 59906
rect 117648 58116 117700 58122
rect 117648 58058 117700 58064
rect 117280 57640 117332 57646
rect 117280 57582 117332 57588
rect 116820 57164 116872 57170
rect 116820 57106 116872 57112
rect 117660 46714 117688 58058
rect 118028 57238 118056 59878
rect 118016 57232 118068 57238
rect 118016 57174 118068 57180
rect 118120 57170 118148 59892
rect 118292 57640 118344 57646
rect 118292 57582 118344 57588
rect 117740 57164 117792 57170
rect 117740 57106 117792 57112
rect 118108 57164 118160 57170
rect 118108 57106 118160 57112
rect 115084 46686 115374 46714
rect 115452 46686 115926 46714
rect 116280 46686 116478 46714
rect 116648 46686 117030 46714
rect 117582 46686 117688 46714
rect 117752 46714 117780 57106
rect 118304 46850 118332 57582
rect 118488 57374 118516 59892
rect 118476 57368 118528 57374
rect 118476 57310 118528 57316
rect 118856 57306 118884 59892
rect 119316 58190 119344 59892
rect 119304 58184 119356 58190
rect 119304 58126 119356 58132
rect 118844 57300 118896 57306
rect 118844 57242 118896 57248
rect 119684 57238 119712 59892
rect 119672 57232 119724 57238
rect 119672 57174 119724 57180
rect 120052 57170 120080 59892
rect 120512 57714 120540 59892
rect 120500 57708 120552 57714
rect 120500 57650 120552 57656
rect 120880 57374 120908 59892
rect 121144 58184 121196 58190
rect 121144 58126 121196 58132
rect 120500 57368 120552 57374
rect 120500 57310 120552 57316
rect 120868 57368 120920 57374
rect 120868 57310 120920 57316
rect 118660 57164 118712 57170
rect 118660 57106 118712 57112
rect 118844 57164 118896 57170
rect 118844 57106 118896 57112
rect 120040 57164 120092 57170
rect 120040 57106 120092 57112
rect 118672 50234 118700 57106
rect 118660 50228 118712 50234
rect 118660 50170 118712 50176
rect 118856 48890 118884 57106
rect 119856 50228 119908 50234
rect 119856 50170 119908 50176
rect 118856 48862 118976 48890
rect 118304 46822 118516 46850
rect 118488 46714 118516 46822
rect 118948 46714 118976 48862
rect 117752 46686 118226 46714
rect 118488 46686 118778 46714
rect 118948 46686 119330 46714
rect 119868 46700 119896 50170
rect 120512 46714 120540 57310
rect 120776 57300 120828 57306
rect 120776 57242 120828 57248
rect 120434 46686 120540 46714
rect 120788 46714 120816 57242
rect 120960 57232 121012 57238
rect 120960 57174 121012 57180
rect 120972 50234 121000 57174
rect 121052 57164 121104 57170
rect 121052 57106 121104 57112
rect 120960 50228 121012 50234
rect 120960 50170 121012 50176
rect 121064 49962 121092 57106
rect 121052 49956 121104 49962
rect 121052 49898 121104 49904
rect 121156 46714 121184 58126
rect 121248 57170 121276 59892
rect 121708 57306 121736 59892
rect 122076 58326 122104 59892
rect 122064 58320 122116 58326
rect 122064 58262 122116 58268
rect 122444 58054 122472 59892
rect 122432 58048 122484 58054
rect 122432 57990 122484 57996
rect 121696 57300 121748 57306
rect 121696 57242 121748 57248
rect 122904 57238 122932 59892
rect 123168 57708 123220 57714
rect 123168 57650 123220 57656
rect 122892 57232 122944 57238
rect 122892 57174 122944 57180
rect 121236 57164 121288 57170
rect 121236 57106 121288 57112
rect 122064 50228 122116 50234
rect 122064 50170 122116 50176
rect 120788 46686 120986 46714
rect 121156 46686 121538 46714
rect 122076 46700 122104 50170
rect 122616 49956 122668 49962
rect 122616 49898 122668 49904
rect 122628 46700 122656 49898
rect 123180 46700 123208 57650
rect 123272 57510 123300 59892
rect 123640 57850 123668 59892
rect 123628 57844 123680 57850
rect 123628 57786 123680 57792
rect 123260 57504 123312 57510
rect 123260 57446 123312 57452
rect 124100 57374 124128 59892
rect 124468 57986 124496 59892
rect 124548 58320 124600 58326
rect 124548 58262 124600 58268
rect 124456 57980 124508 57986
rect 124456 57922 124508 57928
rect 123352 57368 123404 57374
rect 123352 57310 123404 57316
rect 124088 57368 124140 57374
rect 124088 57310 124140 57316
rect 123364 46714 123392 57310
rect 124456 57300 124508 57306
rect 124456 57242 124508 57248
rect 123996 57164 124048 57170
rect 123996 57106 124048 57112
rect 124008 46714 124036 57106
rect 124468 46714 124496 57242
rect 124560 46986 124588 58262
rect 124836 57306 124864 59892
rect 125192 58048 125244 58054
rect 125192 57990 125244 57996
rect 124824 57300 124876 57306
rect 124824 57242 124876 57248
rect 125100 57232 125152 57238
rect 125100 57174 125152 57180
rect 125112 49622 125140 57174
rect 125204 50234 125232 57990
rect 125296 57170 125324 59892
rect 125664 57238 125692 59892
rect 156576 58326 156604 59892
rect 163200 58530 163228 59892
rect 163188 58524 163240 58530
rect 163188 58466 163240 58472
rect 156564 58320 156616 58326
rect 156564 58262 156616 58268
rect 128596 57980 128648 57986
rect 128596 57922 128648 57928
rect 127216 57844 127268 57850
rect 127216 57786 127268 57792
rect 126112 57504 126164 57510
rect 126112 57446 126164 57452
rect 125652 57232 125704 57238
rect 125652 57174 125704 57180
rect 125284 57164 125336 57170
rect 125284 57106 125336 57112
rect 125192 50228 125244 50234
rect 125192 50170 125244 50176
rect 126020 50228 126072 50234
rect 126020 50170 126072 50176
rect 125100 49616 125152 49622
rect 125100 49558 125152 49564
rect 124560 46958 125232 46986
rect 125204 46714 125232 46958
rect 123364 46686 123746 46714
rect 124008 46686 124298 46714
rect 124468 46686 124850 46714
rect 125204 46686 125494 46714
rect 126032 46700 126060 50170
rect 126124 49706 126152 57446
rect 126124 49678 126796 49706
rect 126572 49616 126624 49622
rect 126572 49558 126624 49564
rect 126584 46700 126612 49558
rect 126768 46714 126796 49678
rect 127228 46714 127256 57786
rect 127308 57368 127360 57374
rect 127308 57310 127360 57316
rect 127320 46986 127348 57310
rect 127320 46958 127900 46986
rect 127872 46714 127900 46958
rect 128608 46714 128636 57922
rect 169916 57850 169944 59892
rect 156104 57844 156156 57850
rect 156104 57786 156156 57792
rect 169904 57844 169956 57850
rect 169904 57786 169956 57792
rect 128872 57300 128924 57306
rect 128872 57242 128924 57248
rect 128884 46714 128912 57242
rect 130068 57232 130120 57238
rect 130068 57174 130120 57180
rect 128964 57164 129016 57170
rect 128964 57106 129016 57112
rect 128976 46986 129004 57106
rect 128976 46958 129556 46986
rect 129528 46714 129556 46958
rect 130080 46714 130108 57174
rect 130988 48936 131040 48942
rect 130988 48878 131040 48884
rect 126768 46686 127150 46714
rect 127228 46686 127702 46714
rect 127872 46686 128254 46714
rect 128608 46686 128806 46714
rect 128884 46686 129358 46714
rect 129528 46686 129910 46714
rect 130080 46686 130462 46714
rect 131000 46700 131028 48878
rect 101362 46592 101418 46601
rect 101362 46527 101418 46536
rect 135128 46556 135180 46562
rect 101270 44824 101326 44833
rect 101270 44759 101326 44768
rect 100810 43464 100866 43473
rect 100810 43399 100866 43408
rect 100824 41870 100852 43399
rect 101284 43230 101312 44759
rect 101376 44658 101404 46527
rect 135128 46498 135180 46504
rect 151320 46556 151372 46562
rect 151320 46498 151372 46504
rect 134760 46488 134812 46494
rect 134760 46430 134812 46436
rect 101730 45912 101786 45921
rect 101730 45847 101786 45856
rect 101744 44726 101772 45847
rect 101822 45232 101878 45241
rect 101822 45167 101878 45176
rect 101732 44720 101784 44726
rect 101732 44662 101784 44668
rect 101364 44652 101416 44658
rect 101364 44594 101416 44600
rect 101638 44008 101694 44017
rect 101638 43943 101694 43952
rect 101652 43502 101680 43943
rect 101640 43496 101692 43502
rect 101640 43438 101692 43444
rect 101836 43298 101864 45167
rect 101824 43292 101876 43298
rect 101824 43234 101876 43240
rect 101272 43224 101324 43230
rect 101272 43166 101324 43172
rect 101730 42784 101786 42793
rect 101730 42719 101786 42728
rect 100902 42240 100958 42249
rect 100902 42175 100958 42184
rect 100812 41864 100864 41870
rect 100812 41806 100864 41812
rect 100810 41016 100866 41025
rect 100810 40951 100866 40960
rect 100824 39014 100852 40951
rect 100916 40510 100944 42175
rect 101744 41938 101772 42719
rect 101732 41932 101784 41938
rect 101732 41874 101784 41880
rect 100994 41560 101050 41569
rect 100994 41495 101050 41504
rect 101008 40578 101036 41495
rect 100996 40572 101048 40578
rect 100996 40514 101048 40520
rect 100904 40504 100956 40510
rect 100904 40446 100956 40452
rect 101086 40336 101142 40345
rect 101086 40271 101142 40280
rect 100994 39792 101050 39801
rect 100994 39727 101050 39736
rect 101008 39150 101036 39727
rect 100996 39144 101048 39150
rect 100996 39086 101048 39092
rect 101100 39082 101128 40271
rect 101178 39112 101234 39121
rect 101088 39076 101140 39082
rect 101178 39047 101234 39056
rect 101088 39018 101140 39024
rect 100812 39008 100864 39014
rect 100812 38950 100864 38956
rect 100994 38568 101050 38577
rect 100994 38503 101050 38512
rect 101008 38266 101036 38503
rect 101192 38402 101220 39047
rect 101180 38396 101232 38402
rect 101180 38338 101232 38344
rect 100996 38260 101048 38266
rect 100996 38202 101048 38208
rect 100534 37888 100590 37897
rect 100534 37823 100590 37832
rect 100548 36362 100576 37823
rect 100994 37344 101050 37353
rect 100994 37279 101050 37288
rect 100902 36664 100958 36673
rect 100902 36599 100958 36608
rect 100536 36356 100588 36362
rect 100536 36298 100588 36304
rect 100718 35440 100774 35449
rect 100718 35375 100774 35384
rect 100732 33506 100760 35375
rect 100916 35002 100944 36599
rect 101008 36430 101036 37279
rect 134666 36664 134722 36673
rect 134666 36599 134668 36608
rect 134720 36599 134722 36608
rect 134668 36570 134720 36576
rect 100996 36424 101048 36430
rect 100996 36366 101048 36372
rect 100994 36120 101050 36129
rect 100994 36055 101050 36064
rect 101008 35070 101036 36055
rect 100996 35064 101048 35070
rect 100996 35006 101048 35012
rect 100904 34996 100956 35002
rect 100904 34938 100956 34944
rect 101086 34896 101142 34905
rect 101086 34831 101142 34840
rect 100994 34216 101050 34225
rect 100994 34151 101050 34160
rect 100810 33808 100866 33817
rect 100810 33743 100866 33752
rect 100720 33500 100772 33506
rect 100720 33442 100772 33448
rect 100824 32214 100852 33743
rect 101008 33574 101036 34151
rect 101100 33642 101128 34831
rect 134668 33840 134720 33846
rect 134666 33808 134668 33817
rect 134720 33808 134722 33817
rect 134666 33743 134722 33752
rect 101088 33636 101140 33642
rect 101088 33578 101140 33584
rect 100996 33568 101048 33574
rect 100996 33510 101048 33516
rect 100994 33128 101050 33137
rect 100994 33063 101050 33072
rect 100902 32448 100958 32457
rect 100902 32383 100958 32392
rect 100812 32208 100864 32214
rect 100812 32150 100864 32156
rect 100810 31224 100866 31233
rect 100810 31159 100866 31168
rect 100824 29358 100852 31159
rect 100916 30854 100944 32383
rect 101008 32282 101036 33063
rect 100996 32276 101048 32282
rect 100996 32218 101048 32224
rect 100994 31904 101050 31913
rect 100994 31839 101050 31848
rect 101008 30922 101036 31839
rect 100996 30916 101048 30922
rect 100996 30858 101048 30864
rect 100904 30848 100956 30854
rect 100904 30790 100956 30796
rect 101086 30680 101142 30689
rect 101086 30615 101142 30624
rect 100994 30000 101050 30009
rect 100994 29935 101050 29944
rect 101008 29426 101036 29935
rect 101100 29494 101128 30615
rect 101088 29488 101140 29494
rect 101088 29430 101140 29436
rect 101730 29456 101786 29465
rect 100996 29420 101048 29426
rect 101730 29391 101786 29400
rect 100996 29362 101048 29368
rect 100812 29352 100864 29358
rect 100812 29294 100864 29300
rect 100994 28232 101050 28241
rect 100994 28167 100996 28176
rect 101048 28167 101050 28176
rect 100996 28138 101048 28144
rect 101744 28066 101772 29391
rect 101914 28776 101970 28785
rect 101914 28711 101970 28720
rect 101928 28134 101956 28711
rect 101916 28128 101968 28134
rect 101916 28070 101968 28076
rect 101732 28060 101784 28066
rect 101732 28002 101784 28008
rect 100994 27552 101050 27561
rect 100994 27487 101050 27496
rect 101008 26842 101036 27487
rect 101178 27008 101234 27017
rect 101178 26943 101234 26952
rect 100996 26836 101048 26842
rect 100996 26778 101048 26784
rect 101086 26328 101142 26337
rect 101086 26263 101142 26272
rect 100994 25784 101050 25793
rect 100994 25719 101050 25728
rect 101008 25278 101036 25719
rect 101100 25346 101128 26263
rect 101192 25414 101220 26943
rect 101180 25408 101232 25414
rect 101180 25350 101232 25356
rect 101088 25340 101140 25346
rect 101088 25282 101140 25288
rect 100996 25272 101048 25278
rect 100996 25214 101048 25220
rect 101086 25104 101142 25113
rect 101086 25039 101142 25048
rect 134668 25068 134720 25074
rect 100994 24560 101050 24569
rect 100994 24495 101050 24504
rect 101008 23986 101036 24495
rect 100996 23980 101048 23986
rect 100996 23922 101048 23928
rect 101100 23918 101128 25039
rect 134668 25010 134720 25016
rect 101088 23912 101140 23918
rect 100994 23880 101050 23889
rect 101088 23854 101140 23860
rect 100994 23815 101050 23824
rect 101008 23170 101036 23815
rect 134482 23744 134538 23753
rect 134482 23679 134538 23688
rect 101086 23336 101142 23345
rect 101086 23271 101142 23280
rect 100996 23164 101048 23170
rect 100996 23106 101048 23112
rect 101100 22694 101128 23271
rect 134496 22762 134524 23679
rect 134484 22756 134536 22762
rect 134484 22698 134536 22704
rect 101088 22688 101140 22694
rect 101088 22630 101140 22636
rect 101178 22656 101234 22665
rect 100996 22620 101048 22626
rect 101178 22591 101234 22600
rect 100996 22562 101048 22568
rect 101008 22257 101036 22562
rect 101088 22552 101140 22558
rect 101088 22494 101140 22500
rect 100994 22248 101050 22257
rect 100994 22183 101050 22192
rect 101100 21577 101128 22494
rect 101086 21568 101142 21577
rect 101086 21503 101142 21512
rect 101192 21266 101220 22591
rect 101180 21260 101232 21266
rect 101180 21202 101232 21208
rect 101088 19832 101140 19838
rect 100994 19800 101050 19809
rect 134680 19809 134708 25010
rect 101088 19774 101140 19780
rect 134666 19800 134722 19809
rect 100994 19735 100996 19744
rect 101048 19735 101050 19744
rect 100996 19706 101048 19712
rect 101100 19265 101128 19774
rect 134666 19735 134722 19744
rect 134772 19537 134800 46430
rect 134944 46420 134996 46426
rect 134944 46362 134996 46368
rect 134852 46352 134904 46358
rect 134852 46294 134904 46300
rect 134864 20761 134892 46294
rect 134956 25074 134984 46362
rect 135036 46284 135088 46290
rect 135036 46226 135088 46232
rect 134944 25068 134996 25074
rect 134944 25010 134996 25016
rect 135048 24954 135076 46226
rect 134956 24926 135076 24954
rect 134956 21169 134984 24926
rect 135034 24832 135090 24841
rect 135034 24767 135090 24776
rect 135048 24054 135076 24767
rect 135036 24048 135088 24054
rect 135036 23990 135088 23996
rect 135036 22960 135088 22966
rect 135036 22902 135088 22908
rect 135048 22529 135076 22902
rect 135034 22520 135090 22529
rect 135034 22455 135090 22464
rect 135140 21985 135168 46498
rect 145340 46488 145392 46494
rect 145340 46430 145392 46436
rect 135402 46320 135458 46329
rect 135402 46255 135458 46264
rect 135416 46222 135444 46255
rect 135404 46216 135456 46222
rect 135404 46158 135456 46164
rect 140188 46216 140240 46222
rect 140188 46158 140240 46164
rect 135312 46148 135364 46154
rect 135312 46090 135364 46096
rect 135218 43464 135274 43473
rect 135218 43399 135220 43408
rect 135272 43399 135274 43408
rect 135220 43370 135272 43376
rect 135218 42240 135274 42249
rect 135218 42175 135220 42184
rect 135272 42175 135274 42184
rect 135220 42146 135272 42152
rect 135218 40880 135274 40889
rect 135218 40815 135220 40824
rect 135272 40815 135274 40824
rect 135220 40786 135272 40792
rect 135218 40064 135274 40073
rect 135218 39999 135274 40008
rect 135232 39286 135260 39999
rect 135220 39280 135272 39286
rect 135220 39222 135272 39228
rect 135218 38840 135274 38849
rect 135218 38775 135274 38784
rect 135232 37858 135260 38775
rect 135220 37852 135272 37858
rect 135220 37794 135272 37800
rect 135218 35304 135274 35313
rect 135218 35239 135220 35248
rect 135272 35239 135274 35248
rect 135220 35210 135272 35216
rect 135218 34488 135274 34497
rect 135218 34423 135274 34432
rect 135232 33778 135260 34423
rect 135220 33772 135272 33778
rect 135220 33714 135272 33720
rect 135218 32448 135274 32457
rect 135218 32383 135220 32392
rect 135272 32383 135274 32392
rect 135220 32354 135272 32360
rect 135218 31224 135274 31233
rect 135218 31159 135220 31168
rect 135272 31159 135274 31168
rect 135220 31130 135272 31136
rect 135218 30680 135274 30689
rect 135218 30615 135274 30624
rect 135232 29630 135260 30615
rect 135220 29624 135272 29630
rect 135220 29566 135272 29572
rect 135218 29320 135274 29329
rect 135218 29255 135274 29264
rect 135232 28202 135260 29255
rect 135220 28196 135272 28202
rect 135220 28138 135272 28144
rect 135218 27008 135274 27017
rect 135218 26943 135220 26952
rect 135272 26943 135274 26952
rect 135220 26914 135272 26920
rect 135218 26056 135274 26065
rect 135218 25991 135274 26000
rect 135232 25550 135260 25991
rect 135220 25544 135272 25550
rect 135220 25486 135272 25492
rect 135324 22966 135352 46090
rect 135402 45504 135458 45513
rect 135402 45439 135458 45448
rect 135416 45338 135444 45439
rect 135404 45332 135456 45338
rect 135404 45274 135456 45280
rect 135402 45096 135458 45105
rect 135402 45031 135404 45040
rect 135456 45031 135458 45040
rect 135404 45002 135456 45008
rect 135402 44824 135458 44833
rect 135402 44759 135404 44768
rect 135456 44759 135458 44768
rect 135404 44730 135456 44736
rect 140200 44726 140228 46158
rect 140280 45332 140332 45338
rect 140280 45274 140332 45280
rect 140188 44720 140240 44726
rect 140188 44662 140240 44668
rect 140292 44454 140320 45274
rect 142304 45060 142356 45066
rect 142304 45002 142356 45008
rect 142212 44788 142264 44794
rect 142212 44730 142264 44736
rect 140280 44448 140332 44454
rect 140280 44390 140332 44396
rect 135402 43736 135458 43745
rect 135402 43671 135458 43680
rect 135416 43366 135444 43671
rect 136968 43428 137020 43434
rect 136968 43370 137020 43376
rect 135404 43360 135456 43366
rect 135404 43302 135456 43308
rect 135402 42512 135458 42521
rect 135402 42447 135458 42456
rect 135416 42006 135444 42447
rect 136876 42204 136928 42210
rect 136876 42146 136928 42152
rect 135404 42000 135456 42006
rect 135404 41942 135456 41948
rect 135402 41288 135458 41297
rect 135402 41223 135458 41232
rect 135416 40646 135444 41223
rect 135404 40640 135456 40646
rect 135404 40582 135456 40588
rect 136888 40510 136916 42146
rect 136980 41870 137008 43370
rect 142224 43065 142252 44730
rect 142316 43337 142344 45002
rect 145352 44810 145380 46430
rect 146812 46420 146864 46426
rect 146812 46362 146864 46368
rect 146824 44810 146852 46362
rect 148284 46352 148336 46358
rect 148284 46294 148336 46300
rect 148296 44810 148324 46294
rect 149756 46284 149808 46290
rect 149756 46226 149808 46232
rect 149768 44810 149796 46226
rect 151332 44810 151360 46498
rect 154262 46184 154318 46193
rect 152792 46148 152844 46154
rect 154262 46119 154318 46128
rect 152792 46090 152844 46096
rect 152804 44810 152832 46090
rect 154276 44810 154304 46119
rect 156116 44810 156144 57786
rect 183072 49622 183100 68831
rect 183808 68186 183836 72526
rect 188500 69546 188528 73698
rect 190800 70809 190828 73698
rect 191984 73688 192036 73694
rect 191984 73630 192036 73636
rect 191996 72849 192024 73630
rect 191982 72840 192038 72849
rect 191982 72775 192038 72784
rect 191524 70968 191576 70974
rect 191524 70910 191576 70916
rect 190786 70800 190842 70809
rect 190786 70735 190842 70744
rect 189960 69948 190012 69954
rect 189960 69890 190012 69896
rect 188488 69540 188540 69546
rect 188488 69482 188540 69488
rect 183796 68180 183848 68186
rect 183796 68122 183848 68128
rect 183150 67672 183206 67681
rect 183150 67607 183206 67616
rect 183060 49616 183112 49622
rect 183060 49558 183112 49564
rect 183164 49554 183192 67607
rect 183242 66448 183298 66457
rect 183242 66383 183298 66392
rect 183256 49690 183284 66383
rect 183334 65224 183390 65233
rect 183334 65159 183390 65168
rect 183244 49684 183296 49690
rect 183244 49626 183296 49632
rect 183152 49548 183204 49554
rect 183152 49490 183204 49496
rect 183348 49146 183376 65159
rect 183426 64000 183482 64009
rect 183426 63935 183482 63944
rect 183440 49282 183468 63935
rect 189972 62785 190000 69890
rect 190972 69540 191024 69546
rect 190972 69482 191024 69488
rect 190984 68769 191012 69482
rect 190970 68760 191026 68769
rect 190970 68695 191026 68704
rect 191340 68180 191392 68186
rect 191340 68122 191392 68128
rect 191352 66865 191380 68122
rect 191338 66856 191394 66865
rect 191338 66791 191394 66800
rect 191536 64825 191564 70910
rect 191522 64816 191578 64825
rect 191522 64751 191578 64760
rect 217572 63222 217600 73766
rect 212684 63216 212736 63222
rect 212682 63184 212684 63193
rect 217560 63216 217612 63222
rect 212736 63184 212738 63193
rect 217560 63158 217612 63164
rect 212682 63119 212738 63128
rect 183610 62776 183666 62785
rect 183610 62711 183666 62720
rect 189958 62776 190014 62785
rect 189958 62711 190014 62720
rect 183624 50030 183652 62711
rect 183702 61552 183758 61561
rect 183702 61487 183704 61496
rect 183756 61487 183758 61496
rect 188028 61516 188080 61522
rect 183704 61458 183756 61464
rect 188028 61458 188080 61464
rect 184440 60428 184492 60434
rect 184440 60370 184492 60376
rect 184452 50234 184480 60370
rect 188040 55010 188068 61458
rect 191982 60872 192038 60881
rect 191982 60807 192038 60816
rect 188040 54982 188344 55010
rect 184440 50228 184492 50234
rect 184440 50170 184492 50176
rect 188212 50228 188264 50234
rect 188212 50170 188264 50176
rect 183612 50024 183664 50030
rect 183612 49966 183664 49972
rect 183428 49276 183480 49282
rect 183428 49218 183480 49224
rect 183336 49140 183388 49146
rect 183336 49082 183388 49088
rect 164750 47000 164806 47009
rect 164750 46935 164806 46944
rect 161898 46864 161954 46873
rect 161898 46799 161954 46808
rect 158954 46728 159010 46737
rect 158954 46663 159010 46672
rect 157574 46320 157630 46329
rect 157574 46255 157630 46264
rect 157588 44810 157616 46255
rect 158968 44810 158996 46663
rect 160334 46456 160390 46465
rect 160334 46391 160390 46400
rect 160348 44810 160376 46391
rect 161912 44810 161940 46799
rect 163278 46592 163334 46601
rect 163278 46527 163334 46536
rect 163292 44810 163320 46527
rect 164764 44810 164792 46935
rect 188224 46700 188252 50170
rect 188316 46714 188344 54982
rect 189316 50024 189368 50030
rect 189316 49966 189368 49972
rect 188316 46686 188790 46714
rect 189328 46700 189356 49966
rect 191064 49684 191116 49690
rect 191064 49626 191116 49632
rect 189868 49276 189920 49282
rect 189868 49218 189920 49224
rect 189880 46700 189908 49218
rect 190420 49140 190472 49146
rect 190420 49082 190472 49088
rect 190432 46700 190460 49082
rect 191076 46700 191104 49626
rect 191996 49554 192024 60807
rect 193272 57232 193324 57238
rect 193272 57174 193324 57180
rect 192168 49616 192220 49622
rect 192168 49558 192220 49564
rect 191616 49548 191668 49554
rect 191616 49490 191668 49496
rect 191984 49548 192036 49554
rect 191984 49490 192036 49496
rect 191628 46700 191656 49490
rect 192180 46700 192208 49558
rect 192720 48936 192772 48942
rect 192720 48878 192772 48884
rect 192732 46700 192760 48878
rect 193284 46700 193312 57174
rect 194112 57170 194140 59892
rect 194480 57238 194508 59892
rect 194862 59878 194968 59906
rect 194940 57458 194968 59878
rect 194664 57430 194968 57458
rect 195032 59878 195322 59906
rect 194468 57232 194520 57238
rect 194468 57174 194520 57180
rect 193364 57164 193416 57170
rect 193364 57106 193416 57112
rect 194100 57164 194152 57170
rect 194100 57106 194152 57112
rect 193376 48942 193404 57106
rect 194664 50234 194692 57430
rect 194928 57300 194980 57306
rect 194928 57242 194980 57248
rect 194744 57164 194796 57170
rect 194744 57106 194796 57112
rect 193916 50228 193968 50234
rect 193916 50170 193968 50176
rect 194652 50228 194704 50234
rect 194652 50170 194704 50176
rect 193364 48936 193416 48942
rect 193364 48878 193416 48884
rect 193928 46700 193956 50170
rect 194756 46714 194784 57106
rect 194494 46686 194784 46714
rect 194940 46714 194968 57242
rect 195032 57170 195060 59878
rect 195676 57306 195704 59892
rect 195664 57300 195716 57306
rect 195664 57242 195716 57248
rect 196044 57170 196072 59892
rect 196228 59878 196518 59906
rect 196228 57186 196256 59878
rect 195020 57164 195072 57170
rect 195020 57106 195072 57112
rect 195112 57164 195164 57170
rect 195112 57106 195164 57112
rect 196032 57164 196084 57170
rect 196032 57106 196084 57112
rect 196136 57158 196256 57186
rect 196872 57170 196900 59892
rect 196308 57164 196360 57170
rect 195124 46714 195152 57106
rect 194940 46686 195046 46714
rect 195124 46686 195598 46714
rect 196136 46700 196164 57158
rect 196308 57106 196360 57112
rect 196860 57164 196912 57170
rect 196860 57106 196912 57112
rect 196320 46850 196348 57106
rect 197240 47514 197268 59892
rect 197044 47508 197096 47514
rect 197044 47450 197096 47456
rect 197228 47508 197280 47514
rect 197228 47450 197280 47456
rect 196320 46822 196624 46850
rect 196596 46714 196624 46822
rect 197056 46714 197084 47450
rect 197700 46714 197728 59892
rect 198068 57102 198096 59892
rect 198450 59878 198832 59906
rect 198804 57170 198832 59878
rect 198792 57164 198844 57170
rect 198896 57152 198924 59892
rect 199080 59878 199278 59906
rect 199080 57306 199108 59878
rect 199632 57578 199660 59892
rect 200106 59878 200212 59906
rect 200474 59878 200764 59906
rect 199620 57572 199672 57578
rect 199620 57514 199672 57520
rect 199068 57300 199120 57306
rect 199068 57242 199120 57248
rect 199804 57300 199856 57306
rect 199804 57242 199856 57248
rect 198896 57124 199200 57152
rect 198792 57106 198844 57112
rect 198056 57096 198108 57102
rect 198056 57038 198108 57044
rect 199068 57028 199120 57034
rect 199068 56970 199120 56976
rect 198148 47508 198200 47514
rect 198148 47450 198200 47456
rect 198160 46714 198188 47450
rect 199080 46714 199108 56970
rect 196596 46686 196794 46714
rect 197056 46686 197346 46714
rect 197700 46686 197898 46714
rect 198160 46686 198450 46714
rect 199002 46686 199108 46714
rect 199172 46714 199200 57124
rect 199816 46714 199844 57242
rect 200184 57170 200212 59878
rect 200448 57572 200500 57578
rect 200448 57514 200500 57520
rect 200172 57164 200224 57170
rect 200172 57106 200224 57112
rect 200460 46714 200488 57514
rect 200736 57238 200764 59878
rect 200828 57646 200856 59892
rect 201302 59878 201592 59906
rect 201564 57918 201592 59878
rect 201552 57912 201604 57918
rect 201552 57854 201604 57860
rect 200816 57640 200868 57646
rect 200816 57582 200868 57588
rect 200724 57232 200776 57238
rect 200724 57174 200776 57180
rect 201656 57170 201684 59892
rect 202116 57238 202144 59892
rect 202196 57640 202248 57646
rect 202196 57582 202248 57588
rect 201828 57232 201880 57238
rect 201828 57174 201880 57180
rect 202104 57232 202156 57238
rect 202104 57174 202156 57180
rect 200908 57164 200960 57170
rect 200908 57106 200960 57112
rect 201644 57164 201696 57170
rect 201644 57106 201696 57112
rect 200920 46714 200948 57106
rect 199172 46686 199646 46714
rect 199816 46686 200198 46714
rect 200460 46686 200750 46714
rect 200920 46686 201302 46714
rect 201840 46700 201868 57174
rect 202208 46714 202236 57582
rect 202484 57306 202512 59892
rect 202748 57912 202800 57918
rect 202748 57854 202800 57860
rect 202472 57300 202524 57306
rect 202472 57242 202524 57248
rect 202380 57164 202432 57170
rect 202380 57106 202432 57112
rect 202392 50234 202420 57106
rect 202380 50228 202432 50234
rect 202380 50170 202432 50176
rect 202760 46714 202788 57854
rect 202852 57170 202880 59892
rect 203312 57238 203340 59892
rect 203680 57442 203708 59892
rect 203668 57436 203720 57442
rect 203668 57378 203720 57384
rect 204048 57374 204076 59892
rect 204508 57510 204536 59892
rect 204496 57504 204548 57510
rect 204496 57446 204548 57452
rect 204036 57368 204088 57374
rect 204036 57310 204088 57316
rect 204876 57306 204904 59892
rect 205244 57578 205272 59892
rect 205232 57572 205284 57578
rect 205232 57514 205284 57520
rect 205232 57436 205284 57442
rect 205232 57378 205284 57384
rect 204496 57300 204548 57306
rect 204496 57242 204548 57248
rect 204864 57300 204916 57306
rect 204864 57242 204916 57248
rect 203024 57232 203076 57238
rect 203024 57174 203076 57180
rect 203300 57232 203352 57238
rect 203300 57174 203352 57180
rect 202840 57164 202892 57170
rect 202840 57106 202892 57112
rect 203036 49146 203064 57174
rect 203576 50228 203628 50234
rect 203576 50170 203628 50176
rect 203024 49140 203076 49146
rect 203024 49082 203076 49088
rect 202208 46686 202498 46714
rect 202760 46686 203050 46714
rect 203588 46700 203616 50170
rect 204128 49140 204180 49146
rect 204128 49082 204180 49088
rect 204140 46700 204168 49082
rect 204508 46714 204536 57242
rect 205140 57232 205192 57238
rect 205140 57174 205192 57180
rect 204588 57164 204640 57170
rect 204588 57106 204640 57112
rect 204600 46986 204628 57106
rect 205152 50234 205180 57174
rect 205140 50228 205192 50234
rect 205140 50170 205192 50176
rect 205244 50166 205272 57378
rect 205324 57368 205376 57374
rect 205324 57310 205376 57316
rect 205232 50160 205284 50166
rect 205232 50102 205284 50108
rect 205336 50098 205364 57310
rect 205704 57238 205732 59892
rect 205692 57232 205744 57238
rect 205692 57174 205744 57180
rect 206072 57170 206100 59892
rect 206440 58054 206468 59892
rect 206900 58258 206928 59892
rect 206888 58252 206940 58258
rect 206888 58194 206940 58200
rect 207268 58190 207296 59892
rect 207636 58326 207664 59892
rect 208096 58530 208124 59892
rect 208084 58524 208136 58530
rect 208084 58466 208136 58472
rect 207624 58320 207676 58326
rect 207624 58262 207676 58268
rect 207256 58184 207308 58190
rect 207256 58126 207308 58132
rect 206428 58048 206480 58054
rect 206428 57990 206480 57996
rect 208464 57850 208492 59892
rect 208832 58122 208860 59892
rect 209292 58394 209320 59892
rect 209660 58462 209688 59892
rect 210660 58524 210712 58530
rect 210660 58466 210712 58472
rect 209648 58456 209700 58462
rect 209648 58398 209700 58404
rect 209280 58388 209332 58394
rect 209280 58330 209332 58336
rect 210016 58252 210068 58258
rect 210016 58194 210068 58200
rect 208820 58116 208872 58122
rect 208820 58058 208872 58064
rect 208452 57844 208504 57850
rect 208452 57786 208504 57792
rect 207992 57572 208044 57578
rect 207992 57514 208044 57520
rect 207348 57504 207400 57510
rect 207348 57446 207400 57452
rect 207256 57300 207308 57306
rect 207256 57242 207308 57248
rect 206060 57164 206112 57170
rect 206060 57106 206112 57112
rect 207164 57164 207216 57170
rect 207164 57106 207216 57112
rect 205876 50228 205928 50234
rect 205876 50170 205928 50176
rect 205324 50092 205376 50098
rect 205324 50034 205376 50040
rect 204600 46958 204996 46986
rect 204968 46714 204996 46958
rect 204508 46686 204706 46714
rect 204968 46686 205350 46714
rect 205888 46700 205916 50170
rect 206428 50160 206480 50166
rect 206428 50102 206480 50108
rect 206440 46700 206468 50102
rect 206980 50092 207032 50098
rect 206980 50034 207032 50040
rect 206992 46700 207020 50034
rect 207176 49214 207204 57106
rect 207268 50030 207296 57242
rect 207256 50024 207308 50030
rect 207256 49966 207308 49972
rect 207164 49208 207216 49214
rect 207164 49150 207216 49156
rect 207360 46714 207388 57446
rect 207900 57232 207952 57238
rect 207900 57174 207952 57180
rect 207912 50166 207940 57174
rect 208004 50234 208032 57514
rect 210028 50438 210056 58194
rect 210108 58048 210160 58054
rect 210108 57990 210160 57996
rect 210016 50432 210068 50438
rect 210016 50374 210068 50380
rect 207992 50228 208044 50234
rect 207992 50170 208044 50176
rect 208728 50228 208780 50234
rect 208728 50170 208780 50176
rect 207900 50160 207952 50166
rect 207900 50102 207952 50108
rect 207900 50024 207952 50030
rect 207900 49966 207952 49972
rect 207912 46714 207940 49966
rect 207360 46686 207558 46714
rect 207912 46686 208202 46714
rect 208740 46700 208768 50170
rect 209280 50160 209332 50166
rect 209280 50102 209332 50108
rect 209292 46700 209320 50102
rect 209832 49208 209884 49214
rect 209832 49150 209884 49156
rect 209844 46700 209872 49150
rect 210120 46714 210148 57990
rect 210672 50574 210700 58466
rect 212040 58456 212092 58462
rect 212040 58398 212092 58404
rect 210752 58320 210804 58326
rect 210752 58262 210804 58268
rect 210660 50568 210712 50574
rect 210660 50510 210712 50516
rect 210660 50432 210712 50438
rect 210660 50374 210712 50380
rect 210672 46714 210700 50374
rect 210764 49146 210792 58262
rect 210844 58184 210896 58190
rect 210844 58126 210896 58132
rect 210856 49554 210884 58126
rect 210936 50568 210988 50574
rect 210936 50510 210988 50516
rect 210948 50166 210976 50510
rect 212052 50234 212080 58398
rect 212132 58388 212184 58394
rect 212132 58330 212184 58336
rect 212040 50228 212092 50234
rect 212040 50170 212092 50176
rect 210936 50160 210988 50166
rect 210936 50102 210988 50108
rect 210844 49548 210896 49554
rect 210844 49490 210896 49496
rect 211580 49548 211632 49554
rect 211580 49490 211632 49496
rect 210752 49140 210804 49146
rect 210752 49082 210804 49088
rect 210120 46686 210410 46714
rect 210672 46686 211054 46714
rect 211592 46700 211620 49490
rect 212144 49282 212172 58330
rect 212224 58116 212276 58122
rect 212224 58058 212276 58064
rect 212236 49554 212264 58058
rect 212868 57844 212920 57850
rect 212868 57786 212920 57792
rect 212684 50160 212736 50166
rect 212684 50102 212736 50108
rect 212224 49548 212276 49554
rect 212224 49490 212276 49496
rect 212132 49276 212184 49282
rect 212132 49218 212184 49224
rect 212132 49140 212184 49146
rect 212132 49082 212184 49088
rect 212144 46700 212172 49082
rect 212696 46700 212724 50102
rect 212880 46714 212908 57786
rect 214984 50228 215036 50234
rect 214984 50170 215036 50176
rect 213880 49548 213932 49554
rect 213880 49490 213932 49496
rect 212880 46686 213262 46714
rect 213892 46700 213920 49490
rect 214432 49276 214484 49282
rect 214432 49218 214484 49224
rect 214444 46700 214472 49218
rect 214996 46700 215024 50170
rect 215536 49616 215588 49622
rect 215536 49558 215588 49564
rect 215548 46700 215576 49558
rect 166960 46216 167012 46222
rect 176160 46216 176212 46222
rect 166960 46158 167012 46164
rect 169902 46184 169958 46193
rect 166972 44810 167000 46158
rect 168432 46148 168484 46154
rect 176160 46158 176212 46164
rect 185910 46184 185966 46193
rect 169902 46119 169958 46128
rect 168432 46090 168484 46096
rect 168444 44810 168472 46090
rect 169916 44810 169944 46119
rect 171374 44824 171430 44833
rect 145352 44782 145688 44810
rect 146824 44782 147160 44810
rect 148296 44782 148632 44810
rect 149768 44782 150104 44810
rect 151332 44782 151668 44810
rect 152804 44782 153140 44810
rect 154276 44782 154612 44810
rect 156116 44782 156176 44810
rect 157588 44782 157648 44810
rect 158968 44782 159120 44810
rect 160348 44782 160684 44810
rect 161912 44782 162156 44810
rect 163292 44782 163628 44810
rect 164764 44782 165100 44810
rect 166664 44782 167000 44810
rect 168136 44782 168472 44810
rect 169608 44782 169944 44810
rect 171172 44782 171374 44810
rect 171374 44759 171430 44768
rect 143684 44720 143736 44726
rect 143682 44688 143684 44697
rect 143736 44688 143738 44697
rect 172938 44688 172994 44697
rect 172644 44646 172938 44674
rect 143682 44623 143738 44632
rect 172938 44623 172994 44632
rect 174116 44510 174452 44538
rect 143500 44448 143552 44454
rect 143500 44390 143552 44396
rect 143512 44153 143540 44390
rect 143498 44144 143554 44153
rect 143498 44079 143554 44088
rect 142302 43328 142358 43337
rect 142302 43263 142358 43272
rect 142764 43292 142816 43298
rect 142764 43234 142816 43240
rect 142210 43056 142266 43065
rect 142210 42991 142266 43000
rect 142776 42521 142804 43234
rect 142762 42512 142818 42521
rect 142762 42447 142818 42456
rect 143316 41932 143368 41938
rect 143316 41874 143368 41880
rect 136968 41864 137020 41870
rect 136968 41806 137020 41812
rect 143328 41297 143356 41874
rect 143408 41864 143460 41870
rect 143406 41832 143408 41841
rect 143460 41832 143462 41841
rect 143406 41767 143462 41776
rect 143314 41288 143370 41297
rect 143314 41223 143370 41232
rect 136968 40844 137020 40850
rect 136968 40786 137020 40792
rect 136876 40504 136928 40510
rect 136876 40446 136928 40452
rect 135402 39520 135458 39529
rect 135402 39455 135458 39464
rect 135416 39218 135444 39455
rect 135404 39212 135456 39218
rect 135404 39154 135456 39160
rect 136980 39014 137008 40786
rect 142488 40572 142540 40578
rect 142488 40514 142540 40520
rect 142500 40073 142528 40514
rect 143684 40504 143736 40510
rect 143682 40472 143684 40481
rect 143736 40472 143738 40481
rect 143682 40407 143738 40416
rect 142486 40064 142542 40073
rect 142486 39999 142542 40008
rect 142856 39144 142908 39150
rect 142856 39086 142908 39092
rect 143682 39112 143738 39121
rect 136968 39008 137020 39014
rect 142868 38985 142896 39086
rect 143408 39076 143460 39082
rect 143682 39047 143738 39056
rect 143408 39018 143460 39024
rect 136968 38950 137020 38956
rect 142854 38976 142910 38985
rect 142854 38911 142910 38920
rect 143420 38305 143448 39018
rect 143696 39014 143724 39047
rect 143684 39008 143736 39014
rect 143684 38950 143736 38956
rect 135402 38296 135458 38305
rect 143406 38296 143462 38305
rect 135402 38231 135404 38240
rect 135456 38231 135458 38240
rect 139636 38260 139688 38266
rect 135404 38202 135456 38208
rect 143406 38231 143462 38240
rect 139636 38202 139688 38208
rect 135404 37920 135456 37926
rect 135402 37888 135404 37897
rect 136876 37920 136928 37926
rect 135456 37888 135458 37897
rect 136876 37862 136928 37868
rect 135402 37823 135458 37832
rect 135402 36936 135458 36945
rect 135402 36871 135458 36880
rect 135416 36498 135444 36871
rect 136784 36628 136836 36634
rect 136784 36570 136836 36576
rect 135404 36492 135456 36498
rect 135404 36434 135456 36440
rect 135402 35712 135458 35721
rect 135402 35647 135458 35656
rect 135416 35138 135444 35647
rect 135404 35132 135456 35138
rect 135404 35074 135456 35080
rect 136796 35070 136824 36570
rect 136888 36294 136916 37862
rect 139648 37246 139676 38202
rect 143684 37512 143736 37518
rect 143682 37480 143684 37489
rect 143736 37480 143738 37489
rect 143682 37415 143738 37424
rect 139636 37240 139688 37246
rect 139636 37182 139688 37188
rect 143500 37240 143552 37246
rect 143500 37182 143552 37188
rect 143512 36945 143540 37182
rect 143498 36936 143554 36945
rect 143498 36871 143554 36880
rect 143040 36424 143092 36430
rect 143040 36366 143092 36372
rect 136876 36288 136928 36294
rect 136876 36230 136928 36236
rect 143052 35993 143080 36366
rect 143684 36288 143736 36294
rect 143684 36230 143736 36236
rect 143696 36129 143724 36230
rect 143682 36120 143738 36129
rect 143682 36055 143738 36064
rect 143038 35984 143094 35993
rect 143038 35919 143094 35928
rect 138164 35268 138216 35274
rect 138164 35210 138216 35216
rect 136784 35064 136836 35070
rect 136784 35006 136836 35012
rect 135402 33944 135458 33953
rect 135402 33879 135458 33888
rect 135416 33710 135444 33879
rect 136968 33840 137020 33846
rect 136968 33782 137020 33788
rect 135404 33704 135456 33710
rect 135404 33646 135456 33652
rect 135402 32720 135458 32729
rect 135402 32655 135458 32664
rect 135416 32350 135444 32655
rect 136876 32412 136928 32418
rect 136876 32354 136928 32360
rect 135404 32344 135456 32350
rect 135404 32286 135456 32292
rect 135402 31496 135458 31505
rect 135402 31431 135458 31440
rect 135416 30990 135444 31431
rect 135404 30984 135456 30990
rect 135404 30926 135456 30932
rect 136888 30854 136916 32354
rect 136980 32214 137008 33782
rect 138176 33506 138204 35210
rect 142396 35132 142448 35138
rect 142396 35074 142448 35080
rect 142408 34633 142436 35074
rect 143684 35064 143736 35070
rect 143684 35006 143736 35012
rect 143696 34905 143724 35006
rect 143682 34896 143738 34905
rect 143682 34831 143738 34840
rect 142394 34624 142450 34633
rect 142394 34559 142450 34568
rect 143682 33672 143738 33681
rect 143316 33636 143368 33642
rect 143682 33607 143738 33616
rect 143316 33578 143368 33584
rect 142764 33568 142816 33574
rect 142764 33510 142816 33516
rect 138164 33500 138216 33506
rect 138164 33442 138216 33448
rect 142776 33001 142804 33510
rect 143328 33409 143356 33578
rect 143696 33506 143724 33607
rect 143684 33500 143736 33506
rect 143684 33442 143736 33448
rect 143314 33400 143370 33409
rect 143314 33335 143370 33344
rect 142762 32992 142818 33001
rect 142762 32927 142818 32936
rect 142580 32276 142632 32282
rect 142580 32218 142632 32224
rect 136968 32208 137020 32214
rect 136968 32150 137020 32156
rect 142592 31777 142620 32218
rect 143684 32208 143736 32214
rect 143682 32176 143684 32185
rect 143736 32176 143738 32185
rect 143682 32111 143738 32120
rect 142578 31768 142634 31777
rect 142578 31703 142634 31712
rect 136968 31188 137020 31194
rect 136968 31130 137020 31136
rect 136876 30848 136928 30854
rect 136876 30790 136928 30796
rect 135402 29864 135458 29873
rect 135402 29799 135458 29808
rect 135416 29562 135444 29799
rect 135404 29556 135456 29562
rect 135404 29498 135456 29504
rect 136980 29358 137008 31130
rect 142764 30916 142816 30922
rect 142764 30858 142816 30864
rect 142776 30553 142804 30858
rect 143684 30848 143736 30854
rect 143684 30790 143736 30796
rect 143696 30689 143724 30790
rect 143682 30680 143738 30689
rect 143682 30615 143738 30624
rect 142762 30544 142818 30553
rect 142762 30479 142818 30488
rect 143592 29488 143644 29494
rect 143592 29430 143644 29436
rect 143682 29456 143738 29465
rect 142764 29420 142816 29426
rect 142764 29362 142816 29368
rect 136968 29352 137020 29358
rect 136968 29294 137020 29300
rect 142776 28785 142804 29362
rect 143604 29193 143632 29430
rect 143682 29391 143738 29400
rect 143696 29358 143724 29391
rect 143684 29352 143736 29358
rect 143684 29294 143736 29300
rect 143590 29184 143646 29193
rect 143590 29119 143646 29128
rect 142762 28776 142818 28785
rect 142762 28711 142818 28720
rect 135402 28504 135458 28513
rect 135402 28439 135404 28448
rect 135456 28439 135458 28448
rect 139636 28468 139688 28474
rect 135404 28410 135456 28416
rect 139636 28410 139688 28416
rect 135402 28368 135458 28377
rect 135402 28303 135404 28312
rect 135456 28303 135458 28312
rect 137336 28332 137388 28338
rect 135404 28274 135456 28280
rect 137336 28274 137388 28280
rect 135402 27280 135458 27289
rect 135402 27215 135458 27224
rect 135416 26842 135444 27215
rect 135404 26836 135456 26842
rect 135404 26778 135456 26784
rect 137348 26638 137376 28274
rect 139648 27590 139676 28410
rect 143684 27992 143736 27998
rect 143682 27960 143684 27969
rect 143736 27960 143738 27969
rect 143682 27895 143738 27904
rect 139636 27584 139688 27590
rect 143408 27584 143460 27590
rect 139636 27526 139688 27532
rect 143406 27552 143408 27561
rect 143460 27552 143462 27561
rect 143406 27487 143462 27496
rect 138164 26972 138216 26978
rect 138164 26914 138216 26920
rect 137336 26632 137388 26638
rect 137336 26574 137388 26580
rect 135402 25648 135458 25657
rect 135402 25583 135458 25592
rect 135416 25482 135444 25583
rect 135404 25476 135456 25482
rect 135404 25418 135456 25424
rect 138176 25278 138204 26914
rect 143592 26768 143644 26774
rect 143592 26710 143644 26716
rect 143604 26337 143632 26710
rect 143684 26632 143736 26638
rect 143684 26574 143736 26580
rect 143696 26473 143724 26574
rect 143682 26464 143738 26473
rect 143682 26399 143738 26408
rect 143590 26328 143646 26337
rect 143590 26263 143646 26272
rect 143684 25408 143736 25414
rect 143684 25350 143736 25356
rect 143500 25340 143552 25346
rect 143500 25282 143552 25288
rect 138164 25272 138216 25278
rect 143132 25272 143184 25278
rect 138164 25214 138216 25220
rect 143130 25240 143132 25249
rect 143184 25240 143186 25249
rect 143130 25175 143186 25184
rect 143512 24569 143540 25282
rect 143696 25113 143724 25350
rect 143682 25104 143738 25113
rect 143682 25039 143738 25048
rect 143498 24560 143554 24569
rect 143498 24495 143554 24504
rect 135402 24424 135458 24433
rect 135402 24359 135458 24368
rect 135416 24122 135444 24359
rect 135404 24116 135456 24122
rect 135404 24058 135456 24064
rect 143592 24116 143644 24122
rect 143592 24058 143644 24064
rect 143604 23345 143632 24058
rect 143684 24048 143736 24054
rect 143682 24016 143684 24025
rect 143736 24016 143738 24025
rect 143682 23951 143738 23960
rect 143590 23336 143646 23345
rect 143590 23271 143646 23280
rect 135402 23064 135458 23073
rect 135402 22999 135458 23008
rect 135312 22960 135364 22966
rect 135312 22902 135364 22908
rect 135312 22824 135364 22830
rect 135312 22766 135364 22772
rect 135324 22665 135352 22766
rect 135416 22694 135444 22999
rect 136876 22824 136928 22830
rect 136876 22766 136928 22772
rect 135404 22688 135456 22694
rect 135310 22656 135366 22665
rect 135404 22630 135456 22636
rect 135310 22591 135366 22600
rect 135126 21976 135182 21985
rect 135126 21911 135182 21920
rect 136888 21266 136916 22766
rect 142764 22620 142816 22626
rect 142764 22562 142816 22568
rect 142776 22529 142804 22562
rect 143316 22552 143368 22558
rect 142762 22520 142818 22529
rect 143316 22494 143368 22500
rect 142762 22455 142818 22464
rect 143328 22121 143356 22494
rect 174424 22490 174452 44510
rect 174412 22484 174464 22490
rect 174412 22426 174464 22432
rect 143314 22112 143370 22121
rect 143314 22047 143370 22056
rect 136876 21260 136928 21266
rect 136876 21202 136928 21208
rect 143684 21260 143736 21266
rect 143684 21202 143736 21208
rect 143696 21169 143724 21202
rect 134942 21160 134998 21169
rect 134942 21095 134998 21104
rect 143682 21160 143738 21169
rect 143682 21095 143738 21104
rect 146258 21024 146314 21033
rect 147730 21024 147786 21033
rect 146314 20982 146424 21010
rect 147436 20982 147730 21010
rect 146258 20959 146314 20968
rect 148742 21024 148798 21033
rect 148448 20982 148742 21010
rect 147730 20959 147786 20968
rect 148742 20959 148798 20968
rect 153540 20982 153600 21010
rect 166420 20982 167124 21010
rect 145706 20888 145762 20897
rect 145412 20846 145706 20874
rect 149460 20846 149796 20874
rect 145706 20823 145762 20832
rect 134850 20752 134906 20761
rect 134850 20687 134906 20696
rect 134758 19528 134814 19537
rect 134758 19463 134814 19472
rect 101086 19256 101142 19265
rect 101086 19191 101142 19200
rect 106712 18478 106740 18956
rect 106700 18472 106752 18478
rect 106700 18414 106752 18420
rect 112232 18410 112260 18956
rect 100260 18404 100312 18410
rect 100260 18346 100312 18352
rect 112220 18404 112272 18410
rect 112220 18346 112272 18352
rect 89876 18262 89996 18290
rect 92716 18336 92768 18342
rect 92716 18278 92768 18284
rect 89588 17588 89640 17594
rect 89588 17530 89640 17536
rect 87288 12420 87340 12426
rect 87288 12362 87340 12368
rect 85816 12352 85868 12358
rect 85816 12294 85868 12300
rect 84436 12284 84488 12290
rect 84436 12226 84488 12232
rect 89876 11882 89904 18262
rect 90784 17588 90836 17594
rect 90784 17530 90836 17536
rect 84804 11876 84856 11882
rect 84804 11818 84856 11824
rect 89864 11876 89916 11882
rect 89864 11818 89916 11824
rect 84816 9304 84844 11818
rect 90796 9304 90824 17530
rect 92728 12494 92756 18278
rect 117844 17118 117872 18956
rect 126848 17860 126900 17866
rect 126848 17802 126900 17808
rect 120868 17792 120920 17798
rect 120868 17734 120920 17740
rect 117832 17112 117884 17118
rect 117832 17054 117884 17060
rect 92716 12488 92768 12494
rect 92716 12430 92768 12436
rect 96856 12488 96908 12494
rect 96856 12430 96908 12436
rect 96868 9304 96896 12430
rect 102836 12420 102888 12426
rect 102836 12362 102888 12368
rect 102848 9304 102876 12362
rect 108816 12352 108868 12358
rect 108816 12294 108868 12300
rect 108828 9304 108856 12294
rect 114796 12284 114848 12290
rect 114796 12226 114848 12232
rect 114808 9304 114836 12226
rect 120880 9304 120908 17734
rect 126860 9304 126888 17802
rect 129068 17089 129096 18956
rect 149768 18313 149796 20846
rect 150550 20761 150578 20860
rect 151576 20846 151912 20874
rect 150536 20752 150592 20761
rect 150536 20687 150592 20696
rect 149754 18304 149810 18313
rect 149754 18239 149810 18248
rect 138808 17996 138860 18002
rect 138808 17938 138860 17944
rect 132828 17928 132880 17934
rect 132828 17870 132880 17876
rect 129054 17080 129110 17089
rect 129054 17015 129110 17024
rect 132840 9304 132868 17870
rect 138820 9304 138848 17938
rect 151884 17118 151912 20846
rect 152252 20846 152588 20874
rect 152252 18410 152280 20846
rect 153540 18478 153568 20982
rect 156208 20846 156728 20874
rect 157588 20846 157740 20874
rect 158508 20846 158844 20874
rect 159520 20846 159856 20874
rect 160532 20846 160868 20874
rect 161728 20846 161880 20874
rect 162648 20846 162984 20874
rect 163660 20846 163996 20874
rect 165008 20846 165344 20874
rect 166020 20846 166356 20874
rect 153528 18472 153580 18478
rect 153528 18414 153580 18420
rect 152240 18404 152292 18410
rect 152240 18346 152292 18352
rect 156012 18336 156064 18342
rect 156208 18290 156236 20846
rect 157588 18342 157616 20846
rect 156012 18278 156064 18284
rect 151872 17112 151924 17118
rect 151872 17054 151924 17060
rect 150860 12352 150912 12358
rect 150860 12294 150912 12300
rect 144788 12284 144840 12290
rect 144788 12226 144840 12232
rect 144800 9304 144828 12226
rect 150872 9304 150900 12294
rect 156024 12290 156052 18278
rect 156116 18262 156236 18290
rect 157576 18336 157628 18342
rect 157576 18278 157628 18284
rect 156116 12358 156144 18262
rect 158508 18002 158536 20846
rect 158496 17996 158548 18002
rect 158496 17938 158548 17944
rect 159520 17934 159548 20846
rect 159508 17928 159560 17934
rect 159508 17870 159560 17876
rect 160532 17866 160560 20846
rect 160520 17860 160572 17866
rect 160520 17802 160572 17808
rect 161728 17798 161756 20846
rect 162648 18342 162676 20846
rect 163660 18342 163688 20846
rect 161900 18336 161952 18342
rect 161900 18278 161952 18284
rect 162636 18336 162688 18342
rect 162636 18278 162688 18284
rect 163096 18336 163148 18342
rect 163096 18278 163148 18284
rect 163648 18336 163700 18342
rect 163648 18278 163700 18284
rect 161716 17792 161768 17798
rect 161716 17734 161768 17740
rect 161912 12562 161940 18278
rect 163108 12766 163136 18278
rect 165316 18002 165344 20846
rect 166328 18274 166356 20846
rect 166316 18268 166368 18274
rect 166316 18210 166368 18216
rect 166420 18154 166448 20982
rect 167800 20846 168136 20874
rect 168628 20846 169148 20874
rect 170100 20846 170160 20874
rect 170928 20846 171264 20874
rect 171940 20846 172276 20874
rect 172768 20846 173288 20874
rect 174148 20846 174300 20874
rect 167800 18342 167828 20846
rect 167144 18336 167196 18342
rect 167144 18278 167196 18284
rect 167788 18336 167840 18342
rect 167788 18278 167840 18284
rect 165868 18126 166448 18154
rect 165304 17996 165356 18002
rect 165304 17938 165356 17944
rect 163096 12760 163148 12766
rect 163096 12702 163148 12708
rect 161900 12556 161952 12562
rect 161900 12498 161952 12504
rect 165868 12358 165896 18126
rect 156104 12352 156156 12358
rect 156104 12294 156156 12300
rect 162820 12352 162872 12358
rect 162820 12294 162872 12300
rect 165856 12352 165908 12358
rect 165856 12294 165908 12300
rect 156012 12284 156064 12290
rect 156012 12226 156064 12232
rect 156840 12284 156892 12290
rect 156840 12226 156892 12232
rect 156852 9304 156880 12226
rect 162832 9304 162860 12294
rect 167156 12290 167184 18278
rect 168524 18268 168576 18274
rect 168524 18210 168576 18216
rect 168536 12306 168564 18210
rect 168628 12426 168656 20846
rect 168984 17996 169036 18002
rect 168984 17938 169036 17944
rect 168996 12698 169024 17938
rect 169996 17588 170048 17594
rect 169996 17530 170048 17536
rect 168984 12692 169036 12698
rect 168984 12634 169036 12640
rect 170008 12426 170036 17530
rect 168616 12420 168668 12426
rect 168616 12362 168668 12368
rect 169996 12420 170048 12426
rect 169996 12362 170048 12368
rect 170100 12358 170128 20846
rect 170928 17594 170956 20846
rect 171940 18342 171968 20846
rect 171376 18336 171428 18342
rect 171376 18278 171428 18284
rect 171928 18336 171980 18342
rect 171928 18278 171980 18284
rect 170916 17588 170968 17594
rect 170916 17530 170968 17536
rect 171388 12494 171416 18278
rect 172768 12630 172796 20846
rect 174148 12698 174176 20846
rect 176172 19838 176200 46158
rect 177540 46148 177592 46154
rect 185910 46119 185966 46128
rect 177540 46090 177592 46096
rect 177264 40572 177316 40578
rect 177264 40514 177316 40520
rect 177276 39665 177304 40514
rect 177262 39656 177318 39665
rect 177262 39591 177318 39600
rect 177262 39112 177318 39121
rect 177262 39047 177318 39056
rect 177356 39076 177408 39082
rect 177276 39014 177304 39047
rect 177356 39018 177408 39024
rect 177264 39008 177316 39014
rect 177264 38950 177316 38956
rect 177368 38441 177396 39018
rect 177354 38432 177410 38441
rect 177354 38367 177410 38376
rect 177448 36900 177500 36906
rect 177448 36842 177500 36848
rect 177460 36673 177488 36842
rect 177446 36664 177502 36673
rect 177446 36599 177502 36608
rect 177356 36424 177408 36430
rect 177356 36366 177408 36372
rect 177368 35449 177396 36366
rect 177448 36356 177500 36362
rect 177448 36298 177500 36304
rect 177460 36129 177488 36298
rect 177446 36120 177502 36129
rect 177446 36055 177502 36064
rect 177354 35440 177410 35449
rect 177354 35375 177410 35384
rect 177264 34996 177316 35002
rect 177264 34938 177316 34944
rect 177276 34905 177304 34938
rect 177262 34896 177318 34905
rect 177262 34831 177318 34840
rect 177448 30848 177500 30854
rect 177448 30790 177500 30796
rect 177460 30689 177488 30790
rect 177446 30680 177502 30689
rect 177446 30615 177502 30624
rect 177262 29456 177318 29465
rect 177262 29391 177318 29400
rect 177448 29420 177500 29426
rect 177276 29358 177304 29391
rect 177448 29362 177500 29368
rect 177264 29352 177316 29358
rect 177264 29294 177316 29300
rect 177460 28241 177488 29362
rect 177446 28232 177502 28241
rect 177446 28167 177502 28176
rect 177356 28128 177408 28134
rect 177356 28070 177408 28076
rect 177368 27153 177396 28070
rect 177354 27144 177410 27153
rect 177354 27079 177410 27088
rect 177356 25408 177408 25414
rect 177356 25350 177408 25356
rect 177368 24161 177396 25350
rect 177354 24152 177410 24161
rect 177354 24087 177410 24096
rect 177356 23912 177408 23918
rect 177356 23854 177408 23860
rect 177368 22937 177396 23854
rect 177354 22928 177410 22937
rect 177354 22863 177410 22872
rect 176160 19832 176212 19838
rect 176160 19774 176212 19780
rect 177552 19770 177580 46090
rect 185174 45504 185230 45513
rect 185174 45439 185230 45448
rect 185188 45338 185216 45439
rect 181036 45332 181088 45338
rect 181036 45274 181088 45280
rect 185176 45332 185228 45338
rect 185176 45274 185228 45280
rect 177724 44720 177776 44726
rect 177724 44662 177776 44668
rect 177736 44425 177764 44662
rect 177722 44416 177778 44425
rect 177722 44351 177778 44360
rect 181048 43910 181076 45274
rect 185818 44960 185874 44969
rect 185818 44895 185874 44904
rect 185450 44824 185506 44833
rect 185450 44759 185506 44768
rect 177724 43904 177776 43910
rect 177722 43872 177724 43881
rect 181036 43904 181088 43910
rect 177776 43872 177778 43881
rect 181036 43846 181088 43852
rect 177722 43807 177778 43816
rect 185174 43736 185230 43745
rect 185174 43671 185230 43680
rect 184990 43464 185046 43473
rect 184990 43399 185046 43408
rect 181864 43360 181916 43366
rect 181864 43302 181916 43308
rect 177816 43292 177868 43298
rect 177816 43234 177868 43240
rect 177724 43224 177776 43230
rect 177722 43192 177724 43201
rect 177776 43192 177778 43201
rect 177722 43127 177778 43136
rect 177828 42657 177856 43234
rect 177814 42648 177870 42657
rect 177814 42583 177870 42592
rect 181876 42414 181904 43302
rect 177724 42408 177776 42414
rect 177724 42350 177776 42356
rect 181864 42408 181916 42414
rect 181864 42350 181916 42356
rect 177736 42113 177764 42350
rect 177722 42104 177778 42113
rect 177722 42039 177778 42048
rect 177632 41932 177684 41938
rect 177632 41874 177684 41880
rect 177644 40889 177672 41874
rect 185004 41870 185032 43399
rect 185188 43366 185216 43671
rect 185176 43360 185228 43366
rect 185176 43302 185228 43308
rect 185464 43298 185492 44759
rect 185452 43292 185504 43298
rect 185452 43234 185504 43240
rect 185832 43230 185860 44895
rect 185924 44726 185952 46119
rect 185912 44720 185964 44726
rect 185912 44662 185964 44668
rect 185820 43224 185872 43230
rect 185820 43166 185872 43172
rect 185174 42512 185230 42521
rect 185174 42447 185230 42456
rect 185082 42104 185138 42113
rect 185082 42039 185138 42048
rect 177724 41864 177776 41870
rect 177724 41806 177776 41812
rect 184992 41864 185044 41870
rect 184992 41806 185044 41812
rect 177736 41433 177764 41806
rect 177722 41424 177778 41433
rect 177722 41359 177778 41368
rect 177630 40880 177686 40889
rect 177630 40815 177686 40824
rect 184990 40608 185046 40617
rect 184990 40543 185046 40552
rect 177724 40504 177776 40510
rect 177724 40446 177776 40452
rect 177736 40209 177764 40446
rect 177722 40200 177778 40209
rect 177722 40135 177778 40144
rect 177724 39144 177776 39150
rect 177724 39086 177776 39092
rect 177736 37897 177764 39086
rect 185004 39014 185032 40543
rect 185096 40510 185124 42039
rect 185188 41938 185216 42447
rect 185176 41932 185228 41938
rect 185176 41874 185228 41880
rect 185174 41288 185230 41297
rect 185174 41223 185230 41232
rect 185188 40578 185216 41223
rect 185176 40572 185228 40578
rect 185176 40514 185228 40520
rect 185084 40504 185136 40510
rect 185084 40446 185136 40452
rect 185266 40064 185322 40073
rect 185266 39999 185322 40008
rect 185174 39384 185230 39393
rect 185174 39319 185230 39328
rect 185188 39150 185216 39319
rect 185176 39144 185228 39150
rect 185176 39086 185228 39092
rect 185280 39082 185308 39999
rect 185268 39076 185320 39082
rect 185268 39018 185320 39024
rect 184992 39008 185044 39014
rect 184992 38950 185044 38956
rect 185266 38840 185322 38849
rect 185266 38775 185322 38784
rect 185174 38160 185230 38169
rect 183244 38124 183296 38130
rect 185280 38130 185308 38775
rect 185174 38095 185230 38104
rect 185268 38124 185320 38130
rect 183244 38066 183296 38072
rect 177722 37888 177778 37897
rect 177722 37823 177778 37832
rect 183256 37382 183284 38066
rect 184990 37888 185046 37897
rect 183704 37852 183756 37858
rect 185188 37858 185216 38095
rect 185268 38066 185320 38072
rect 184990 37823 185046 37832
rect 185176 37852 185228 37858
rect 183704 37794 183756 37800
rect 177724 37376 177776 37382
rect 177724 37318 177776 37324
rect 183244 37376 183296 37382
rect 183244 37318 183296 37324
rect 177736 37217 177764 37318
rect 177722 37208 177778 37217
rect 177722 37143 177778 37152
rect 183716 36906 183744 37794
rect 183704 36900 183756 36906
rect 183704 36842 183756 36848
rect 185004 36362 185032 37823
rect 185176 37794 185228 37800
rect 185174 36936 185230 36945
rect 185174 36871 185230 36880
rect 185082 36528 185138 36537
rect 185082 36463 185138 36472
rect 184992 36356 185044 36362
rect 184992 36298 185044 36304
rect 184898 35304 184954 35313
rect 184898 35239 184954 35248
rect 177724 35064 177776 35070
rect 177724 35006 177776 35012
rect 177736 34225 177764 35006
rect 177722 34216 177778 34225
rect 177722 34151 177778 34160
rect 177630 33672 177686 33681
rect 177630 33607 177686 33616
rect 177816 33636 177868 33642
rect 177644 33506 177672 33607
rect 177816 33578 177868 33584
rect 177724 33568 177776 33574
rect 177724 33510 177776 33516
rect 177632 33500 177684 33506
rect 177632 33442 177684 33448
rect 177736 33137 177764 33510
rect 177722 33128 177778 33137
rect 177722 33063 177778 33072
rect 177828 32457 177856 33578
rect 184912 33506 184940 35239
rect 185096 35002 185124 36463
rect 185188 36430 185216 36871
rect 185176 36424 185228 36430
rect 185176 36366 185228 36372
rect 185450 35712 185506 35721
rect 185450 35647 185506 35656
rect 185464 35070 185492 35647
rect 185452 35064 185504 35070
rect 185452 35006 185504 35012
rect 185084 34996 185136 35002
rect 185084 34938 185136 34944
rect 185266 34488 185322 34497
rect 185266 34423 185322 34432
rect 185174 33944 185230 33953
rect 185174 33879 185230 33888
rect 184990 33808 185046 33817
rect 184990 33743 185046 33752
rect 184900 33500 184952 33506
rect 184900 33442 184952 33448
rect 177814 32448 177870 32457
rect 177814 32383 177870 32392
rect 177632 32276 177684 32282
rect 177632 32218 177684 32224
rect 177644 31233 177672 32218
rect 185004 32214 185032 33743
rect 185188 33642 185216 33879
rect 185176 33636 185228 33642
rect 185176 33578 185228 33584
rect 185280 33574 185308 34423
rect 185268 33568 185320 33574
rect 185268 33510 185320 33516
rect 185174 32720 185230 32729
rect 185174 32655 185230 32664
rect 185082 32312 185138 32321
rect 185188 32282 185216 32655
rect 185082 32247 185138 32256
rect 185176 32276 185228 32282
rect 177724 32208 177776 32214
rect 177724 32150 177776 32156
rect 184992 32208 185044 32214
rect 184992 32150 185044 32156
rect 177736 31913 177764 32150
rect 177722 31904 177778 31913
rect 177722 31839 177778 31848
rect 177630 31224 177686 31233
rect 177630 31159 177686 31168
rect 184990 30952 185046 30961
rect 177724 30916 177776 30922
rect 184990 30887 185046 30896
rect 177724 30858 177776 30864
rect 177736 30145 177764 30858
rect 177722 30136 177778 30145
rect 177722 30071 177778 30080
rect 177724 29488 177776 29494
rect 177724 29430 177776 29436
rect 177736 28921 177764 29430
rect 185004 29358 185032 30887
rect 185096 30854 185124 32247
rect 185176 32218 185228 32224
rect 185174 31496 185230 31505
rect 185174 31431 185230 31440
rect 185188 30922 185216 31431
rect 185176 30916 185228 30922
rect 185176 30858 185228 30864
rect 185084 30848 185136 30854
rect 185084 30790 185136 30796
rect 185266 30272 185322 30281
rect 185266 30207 185322 30216
rect 185174 29728 185230 29737
rect 185174 29663 185230 29672
rect 185188 29426 185216 29663
rect 185280 29494 185308 30207
rect 185268 29488 185320 29494
rect 185268 29430 185320 29436
rect 185176 29420 185228 29426
rect 185176 29362 185228 29368
rect 184992 29352 185044 29358
rect 184992 29294 185044 29300
rect 185358 29048 185414 29057
rect 185358 28983 185414 28992
rect 177722 28912 177778 28921
rect 177722 28847 177778 28856
rect 185266 28504 185322 28513
rect 185266 28439 185322 28448
rect 185174 28232 185230 28241
rect 177632 28196 177684 28202
rect 185174 28167 185176 28176
rect 177632 28138 177684 28144
rect 185228 28167 185230 28176
rect 185176 28138 185228 28144
rect 177644 26473 177672 28138
rect 185280 28134 185308 28439
rect 185268 28128 185320 28134
rect 185268 28070 185320 28076
rect 185372 28066 185400 28983
rect 177724 28060 177776 28066
rect 177724 28002 177776 28008
rect 185360 28060 185412 28066
rect 185360 28002 185412 28008
rect 177736 27697 177764 28002
rect 177722 27688 177778 27697
rect 177722 27623 177778 27632
rect 185174 27280 185230 27289
rect 185174 27215 185230 27224
rect 185188 26842 185216 27215
rect 185818 26872 185874 26881
rect 185176 26836 185228 26842
rect 185818 26807 185874 26816
rect 185176 26778 185228 26784
rect 177724 26768 177776 26774
rect 177724 26710 177776 26716
rect 177630 26464 177686 26473
rect 177630 26399 177686 26408
rect 177736 25929 177764 26710
rect 185266 26056 185322 26065
rect 185266 25991 185322 26000
rect 177722 25920 177778 25929
rect 177722 25855 177778 25864
rect 185280 25346 185308 25991
rect 185726 25648 185782 25657
rect 185726 25583 185782 25592
rect 185740 25414 185768 25583
rect 185728 25408 185780 25414
rect 185728 25350 185780 25356
rect 177816 25340 177868 25346
rect 177816 25282 177868 25288
rect 185268 25340 185320 25346
rect 185268 25282 185320 25288
rect 177724 25272 177776 25278
rect 177722 25240 177724 25249
rect 177776 25240 177778 25249
rect 177722 25175 177778 25184
rect 177828 24705 177856 25282
rect 185832 25278 185860 26807
rect 185820 25272 185872 25278
rect 185820 25214 185872 25220
rect 185174 24832 185230 24841
rect 185174 24767 185230 24776
rect 177814 24696 177870 24705
rect 177814 24631 177870 24640
rect 185188 23986 185216 24767
rect 185266 24152 185322 24161
rect 185266 24087 185322 24096
rect 177632 23980 177684 23986
rect 177632 23922 177684 23928
rect 185176 23980 185228 23986
rect 185176 23922 185228 23928
rect 177644 23481 177672 23922
rect 185280 23918 185308 24087
rect 185268 23912 185320 23918
rect 185268 23854 185320 23860
rect 185266 23608 185322 23617
rect 185266 23543 185322 23552
rect 177630 23472 177686 23481
rect 177630 23407 177686 23416
rect 185174 22928 185230 22937
rect 185174 22863 185230 22872
rect 185188 22694 185216 22863
rect 185280 22830 185308 23543
rect 185268 22824 185320 22830
rect 185268 22766 185320 22772
rect 185176 22688 185228 22694
rect 185176 22630 185228 22636
rect 185266 22656 185322 22665
rect 177632 22620 177684 22626
rect 185266 22591 185322 22600
rect 177632 22562 177684 22568
rect 177644 22257 177672 22562
rect 177724 22552 177776 22558
rect 177724 22494 177776 22500
rect 177630 22248 177686 22257
rect 177630 22183 177686 22192
rect 177736 21713 177764 22494
rect 185176 22484 185228 22490
rect 185176 22426 185228 22432
rect 185188 22393 185216 22426
rect 185174 22384 185230 22393
rect 185174 22319 185230 22328
rect 177722 21704 177778 21713
rect 177722 21639 177778 21648
rect 185280 21266 185308 22591
rect 220332 21985 220360 215167
rect 222342 205440 222398 205449
rect 222342 205375 222398 205384
rect 222356 204866 222384 205375
rect 222344 204860 222396 204866
rect 222344 204802 222396 204808
rect 220412 182760 220464 182766
rect 220412 182702 220464 182708
rect 220424 179201 220452 182702
rect 220410 179192 220466 179201
rect 220410 179127 220466 179136
rect 221698 152944 221754 152953
rect 221698 152879 221754 152888
rect 221712 90218 221740 152879
rect 222344 127476 222396 127482
rect 222344 127418 222396 127424
rect 222356 126841 222384 127418
rect 222342 126832 222398 126841
rect 222342 126767 222398 126776
rect 222342 100584 222398 100593
rect 222342 100519 222398 100528
rect 222356 99942 222384 100519
rect 222344 99936 222396 99942
rect 222344 99878 222396 99884
rect 221700 90212 221752 90218
rect 221700 90154 221752 90160
rect 222342 74336 222398 74345
rect 222342 74271 222398 74280
rect 222356 73830 222384 74271
rect 222344 73824 222396 73830
rect 222344 73766 222396 73772
rect 222252 48868 222304 48874
rect 222252 48810 222304 48816
rect 222264 48097 222292 48810
rect 222250 48088 222306 48097
rect 222250 48023 222306 48032
rect 220318 21976 220374 21985
rect 220318 21911 220374 21920
rect 177724 21260 177776 21266
rect 177724 21202 177776 21208
rect 185268 21260 185320 21266
rect 185268 21202 185320 21208
rect 177736 21169 177764 21202
rect 177722 21160 177778 21169
rect 177722 21095 177778 21104
rect 185268 19832 185320 19838
rect 185174 19800 185230 19809
rect 177540 19764 177592 19770
rect 185268 19774 185320 19780
rect 185174 19735 185176 19744
rect 177540 19706 177592 19712
rect 185228 19735 185230 19744
rect 185176 19706 185228 19712
rect 185280 19537 185308 19774
rect 185266 19528 185322 19537
rect 185266 19463 185322 19472
rect 192548 18478 192576 18956
rect 192536 18472 192588 18478
rect 192536 18414 192588 18420
rect 201840 17089 201868 18956
rect 211132 17118 211160 18956
rect 211396 18472 211448 18478
rect 211394 18440 211396 18449
rect 211448 18440 211450 18449
rect 211394 18375 211450 18384
rect 211120 17112 211172 17118
rect 201826 17080 201882 17089
rect 211120 17054 211172 17060
rect 201826 17015 201882 17024
rect 180852 12896 180904 12902
rect 180852 12838 180904 12844
rect 174872 12760 174924 12766
rect 174872 12702 174924 12708
rect 174136 12692 174188 12698
rect 174136 12634 174188 12640
rect 172756 12624 172808 12630
rect 172756 12566 172808 12572
rect 171376 12488 171428 12494
rect 171376 12430 171428 12436
rect 170088 12352 170140 12358
rect 167144 12284 167196 12290
rect 168536 12278 168840 12306
rect 170088 12294 170140 12300
rect 167144 12226 167196 12232
rect 168812 9304 168840 12278
rect 174884 9304 174912 12702
rect 180864 9304 180892 12838
rect 192812 12692 192864 12698
rect 192812 12634 192864 12640
rect 186832 12556 186884 12562
rect 186832 12498 186884 12504
rect 186844 9304 186872 12498
rect 192824 9304 192852 12634
rect 198792 12624 198844 12630
rect 198792 12566 198844 12572
rect 198804 9304 198832 12566
rect 204864 12488 204916 12494
rect 204864 12430 204916 12436
rect 204876 9304 204904 12430
rect 210844 12420 210896 12426
rect 210844 12362 210896 12368
rect 210856 9304 210884 12362
rect 216824 12352 216876 12358
rect 216824 12294 216876 12300
rect 216836 9304 216864 12294
rect 222804 12284 222856 12290
rect 222804 12226 222856 12232
rect 222816 9304 222844 12226
rect 12858 8824 12914 9304
rect 18838 8824 18894 9304
rect 24818 8824 24874 9304
rect 30798 8824 30854 9304
rect 36778 8824 36834 9304
rect 42850 8824 42906 9304
rect 48830 8824 48886 9304
rect 54810 8824 54866 9304
rect 60790 8824 60846 9304
rect 66862 8824 66918 9304
rect 72842 8824 72898 9304
rect 78822 8824 78878 9304
rect 84802 8824 84858 9304
rect 90782 8824 90838 9304
rect 96854 8824 96910 9304
rect 102834 8824 102890 9304
rect 108814 8824 108870 9304
rect 114794 8824 114850 9304
rect 120866 8824 120922 9304
rect 126846 8824 126902 9304
rect 132826 8824 132882 9304
rect 138806 8824 138862 9304
rect 144786 8824 144842 9304
rect 150858 8824 150914 9304
rect 156838 8824 156894 9304
rect 162818 8824 162874 9304
rect 168798 8824 168854 9304
rect 174870 8824 174926 9304
rect 180850 8824 180906 9304
rect 186830 8824 186886 9304
rect 192810 8824 192866 9304
rect 198790 8824 198846 9304
rect 204862 8824 204918 9304
rect 210842 8824 210898 9304
rect 216822 8824 216878 9304
rect 222802 8824 222858 9304
<< via2 >>
rect 33374 236528 33430 236584
rect 13318 232856 13374 232912
rect 14698 209328 14754 209384
rect 13318 185664 13374 185720
rect 13410 162136 13466 162192
rect 13318 138472 13374 138528
rect 13318 114944 13374 115000
rect 13318 91280 13374 91336
rect 13318 67752 13374 67808
rect 13410 44088 13466 44144
rect 22794 190424 22850 190480
rect 41838 189200 41894 189256
rect 22334 183760 22390 183816
rect 23622 178728 23678 178784
rect 22334 177096 22390 177152
rect 23622 170432 23678 170488
rect 50578 234488 50634 234544
rect 50026 232856 50082 232912
rect 50118 231632 50174 231688
rect 50026 225920 50082 225976
rect 50394 215040 50450 215096
rect 50394 213952 50450 214008
rect 50486 207696 50542 207752
rect 51222 233964 51278 234000
rect 51222 233944 51224 233964
rect 51224 233944 51276 233964
rect 51276 233944 51278 233964
rect 51222 233400 51278 233456
rect 58122 232992 58178 233048
rect 79558 235168 79614 235224
rect 50762 232176 50818 232232
rect 58030 231904 58086 231960
rect 58122 231224 58178 231280
rect 51222 231088 51278 231144
rect 51130 230544 51186 230600
rect 51222 230000 51278 230056
rect 58214 230680 58270 230736
rect 58214 230136 58270 230192
rect 51130 229320 51186 229376
rect 58214 229456 58270 229512
rect 58214 228912 58270 228968
rect 51222 228776 51278 228832
rect 51038 228232 51094 228288
rect 50762 227688 50818 227744
rect 51222 227144 51278 227200
rect 51222 226464 51278 226520
rect 58306 228232 58362 228288
rect 58214 227688 58270 227744
rect 58306 227144 58362 227200
rect 58214 226464 58270 226520
rect 58214 225920 58270 225976
rect 51130 225376 51186 225432
rect 58214 225240 58270 225296
rect 51222 224832 51278 224888
rect 51130 224308 51186 224344
rect 51130 224288 51132 224308
rect 51132 224288 51184 224308
rect 51184 224288 51186 224308
rect 58306 224696 58362 224752
rect 51222 223608 51278 223664
rect 51130 223084 51186 223120
rect 51130 223064 51132 223084
rect 51132 223064 51184 223084
rect 51184 223064 51186 223084
rect 58398 224152 58454 224208
rect 51222 222520 51278 222576
rect 51130 221976 51186 222032
rect 51222 221432 51278 221488
rect 51222 220752 51278 220808
rect 51130 220208 51186 220264
rect 58306 223472 58362 223528
rect 58214 222928 58270 222984
rect 58214 222248 58270 222304
rect 58306 221704 58362 221760
rect 58214 221160 58270 221216
rect 58214 220480 58270 220536
rect 50854 219664 50910 219720
rect 51222 219120 51278 219176
rect 51222 218576 51278 218632
rect 58306 219936 58362 219992
rect 58214 219256 58270 219312
rect 50762 217896 50818 217952
rect 51222 217372 51278 217408
rect 51222 217352 51224 217372
rect 51224 217352 51276 217372
rect 51276 217352 51278 217372
rect 51130 216808 51186 216864
rect 51222 216264 51278 216320
rect 51222 215720 51278 215776
rect 51130 214532 51132 214552
rect 51132 214532 51184 214552
rect 51184 214532 51186 214552
rect 51130 214496 51186 214532
rect 58306 218712 58362 218768
rect 58214 218168 58270 218224
rect 58214 217488 58270 217544
rect 58214 216944 58270 217000
rect 58306 216264 58362 216320
rect 58214 215756 58216 215776
rect 58216 215756 58268 215776
rect 58268 215756 58270 215776
rect 58214 215720 58270 215756
rect 58306 215176 58362 215232
rect 51222 213428 51278 213464
rect 51222 213408 51224 213428
rect 51224 213408 51276 213428
rect 51276 213408 51278 213428
rect 58214 214496 58270 214552
rect 58214 213952 58270 214008
rect 51222 212864 51278 212920
rect 51130 212184 51186 212240
rect 51222 211640 51278 211696
rect 50854 211096 50910 211152
rect 50670 210552 50726 210608
rect 50762 210008 50818 210064
rect 58306 213272 58362 213328
rect 58214 212728 58270 212784
rect 58306 212184 58362 212240
rect 58214 211504 58270 211560
rect 58306 210960 58362 211016
rect 58398 210280 58454 210336
rect 58214 209736 58270 209792
rect 50946 209328 51002 209384
rect 58306 209192 58362 209248
rect 92714 232448 92770 232504
rect 94002 231904 94058 231960
rect 92714 231224 92770 231280
rect 93726 230680 93782 230736
rect 92714 230136 92770 230192
rect 92714 229456 92770 229512
rect 92806 228912 92862 228968
rect 92714 228232 92770 228288
rect 93174 227688 93230 227744
rect 92714 227144 92770 227200
rect 92714 226464 92770 226520
rect 92806 225920 92862 225976
rect 92714 225276 92716 225296
rect 92716 225276 92768 225296
rect 92768 225276 92770 225296
rect 92714 225240 92770 225276
rect 92806 224696 92862 224752
rect 93726 224152 93782 224208
rect 93726 223472 93782 223528
rect 93910 222928 93966 222984
rect 92714 222248 92770 222304
rect 92990 221704 93046 221760
rect 92714 221180 92770 221216
rect 92714 221160 92716 221180
rect 92716 221160 92768 221180
rect 92768 221160 92770 221180
rect 93726 220480 93782 220536
rect 92806 219936 92862 219992
rect 93726 219256 93782 219312
rect 93910 218712 93966 218768
rect 93174 218168 93230 218224
rect 93726 217488 93782 217544
rect 93542 216944 93598 217000
rect 92714 216264 92770 216320
rect 92714 215740 92770 215776
rect 92714 215720 92716 215740
rect 92716 215720 92768 215740
rect 92768 215720 92770 215740
rect 92806 215176 92862 215232
rect 93542 214496 93598 214552
rect 92714 213952 92770 214008
rect 93358 213272 93414 213328
rect 92714 212728 92770 212784
rect 93358 212184 93414 212240
rect 92714 211540 92716 211560
rect 92716 211540 92768 211560
rect 92768 211540 92770 211560
rect 92714 211504 92770 211540
rect 92806 210960 92862 211016
rect 51038 208784 51094 208840
rect 51222 208240 51278 208296
rect 51130 207152 51186 207208
rect 88758 208920 88814 208976
rect 92898 210280 92954 210336
rect 93174 209736 93230 209792
rect 92714 209192 92770 209248
rect 53338 173832 53394 173888
rect 44414 168664 44470 168720
rect 53338 163768 53394 163824
rect 53430 160504 53486 160560
rect 44506 158736 44562 158792
rect 51406 140376 51462 140432
rect 49934 140104 49990 140160
rect 50026 139016 50082 139072
rect 49934 138644 49936 138664
rect 49936 138644 49988 138664
rect 49988 138644 49990 138664
rect 49934 138608 49990 138644
rect 50026 137792 50082 137848
rect 49934 137384 49990 137440
rect 50394 136568 50450 136624
rect 18102 135888 18158 135944
rect 18010 126232 18066 126288
rect 18010 116984 18066 117040
rect 51222 136180 51278 136216
rect 51222 136160 51224 136180
rect 51224 136160 51276 136180
rect 51276 136160 51278 136180
rect 51222 136044 51278 136080
rect 51222 136024 51224 136044
rect 51224 136024 51276 136044
rect 51276 136024 51278 136044
rect 51222 134936 51278 134992
rect 51130 134548 51186 134584
rect 51130 134528 51132 134548
rect 51132 134528 51184 134548
rect 51184 134528 51186 134548
rect 58214 136024 58270 136080
rect 58398 137112 58454 137168
rect 59226 138508 59228 138528
rect 59228 138508 59280 138528
rect 59280 138508 59282 138528
rect 59226 138472 59282 138508
rect 92714 138508 92716 138528
rect 92716 138508 92768 138528
rect 92768 138508 92770 138528
rect 92714 138472 92770 138508
rect 58674 138200 58730 138256
rect 92806 138064 92862 138120
rect 92714 137132 92770 137168
rect 92714 137112 92716 137132
rect 92716 137112 92768 137132
rect 92768 137112 92770 137132
rect 58490 136568 58546 136624
rect 92806 136840 92862 136896
rect 92714 136432 92770 136488
rect 92714 135480 92770 135536
rect 58306 135344 58362 135400
rect 92806 135208 92862 135264
rect 58214 134800 58270 134856
rect 50210 133712 50266 133768
rect 50946 133168 51002 133224
rect 51222 132488 51278 132544
rect 50394 132080 50450 132136
rect 51222 131692 51278 131728
rect 51222 131672 51224 131692
rect 51224 131672 51276 131692
rect 51276 131672 51278 131692
rect 58214 134120 58270 134176
rect 58306 133576 58362 133632
rect 58214 133032 58270 133088
rect 92714 134292 92716 134312
rect 92716 134292 92768 134312
rect 92768 134292 92770 134312
rect 92714 134256 92770 134292
rect 92806 133848 92862 133904
rect 92898 133440 92954 133496
rect 92714 132624 92770 132680
rect 58214 132352 58270 132408
rect 51222 130740 51278 130776
rect 51222 130720 51224 130740
rect 51224 130720 51276 130740
rect 51276 130720 51278 130740
rect 51222 130332 51278 130368
rect 51222 130312 51224 130332
rect 51224 130312 51276 130332
rect 51276 130312 51278 130332
rect 50394 129632 50450 129688
rect 51222 128972 51278 129008
rect 51222 128952 51224 128972
rect 51224 128952 51276 128972
rect 51276 128952 51278 128972
rect 50946 128408 51002 128464
rect 51222 127864 51278 127920
rect 51222 127612 51278 127648
rect 51222 127592 51224 127612
rect 51224 127592 51276 127612
rect 51276 127592 51278 127612
rect 51222 126640 51278 126696
rect 51222 126096 51278 126152
rect 50210 125552 50266 125608
rect 51222 125028 51278 125064
rect 51222 125008 51224 125028
rect 51224 125008 51276 125028
rect 51276 125008 51278 125028
rect 51222 124892 51278 124928
rect 51222 124872 51224 124892
rect 51224 124872 51276 124892
rect 51276 124872 51278 124892
rect 92806 132216 92862 132272
rect 58306 131808 58362 131864
rect 92714 131400 92770 131456
rect 58214 131128 58270 131184
rect 92806 130992 92862 131048
rect 58306 130584 58362 130640
rect 92714 130212 92716 130232
rect 92716 130212 92768 130232
rect 92768 130212 92770 130232
rect 92714 130176 92770 130212
rect 58214 130040 58270 130096
rect 92806 129768 92862 129824
rect 58306 129360 58362 129416
rect 58214 128836 58270 128872
rect 92714 128852 92716 128872
rect 92716 128852 92768 128872
rect 92768 128852 92770 128872
rect 58214 128816 58216 128836
rect 58216 128816 58268 128836
rect 58268 128816 58270 128836
rect 92714 128816 92770 128852
rect 58306 128136 58362 128192
rect 92806 128408 92862 128464
rect 92714 128000 92770 128056
rect 58214 127592 58270 127648
rect 92714 127184 92770 127240
rect 58214 127048 58270 127104
rect 92806 126912 92862 126968
rect 58306 126368 58362 126424
rect 58214 125824 58270 125880
rect 92714 125996 92716 126016
rect 92716 125996 92768 126016
rect 92768 125996 92770 126016
rect 92714 125960 92770 125996
rect 92806 125552 92862 125608
rect 58306 125144 58362 125200
rect 50578 123784 50634 123840
rect 51130 123396 51186 123432
rect 51130 123376 51132 123396
rect 51132 123376 51184 123396
rect 51184 123376 51186 123396
rect 50854 122560 50910 122616
rect 50210 122288 50266 122344
rect 58214 124636 58216 124656
rect 58216 124636 58268 124656
rect 58268 124636 58270 124656
rect 58214 124600 58270 124636
rect 58306 124056 58362 124112
rect 92714 124636 92716 124656
rect 92716 124636 92768 124656
rect 92768 124636 92770 124656
rect 92714 124600 92770 124636
rect 92806 124328 92862 124384
rect 92898 123920 92954 123976
rect 58398 123376 58454 123432
rect 58214 122832 58270 122888
rect 50210 121472 50266 121528
rect 51222 120948 51278 120984
rect 51222 120928 51224 120948
rect 51224 120928 51276 120948
rect 51276 120928 51278 120948
rect 51222 120792 51278 120848
rect 51222 119704 51278 119760
rect 51222 119316 51278 119352
rect 51222 119296 51224 119316
rect 51224 119296 51276 119316
rect 51276 119296 51278 119316
rect 92714 123104 92770 123160
rect 92806 122696 92862 122752
rect 58306 122152 58362 122208
rect 58214 121608 58270 121664
rect 92714 121744 92770 121800
rect 92806 121472 92862 121528
rect 58306 121064 58362 121120
rect 51222 118480 51278 118536
rect 51222 117956 51278 117992
rect 51222 117936 51224 117956
rect 51224 117936 51276 117956
rect 51276 117936 51278 117956
rect 51222 117392 51278 117448
rect 50578 116712 50634 116768
rect 22334 96448 22390 96504
rect 50762 116440 50818 116496
rect 50670 115080 50726 115136
rect 92714 120556 92716 120576
rect 92716 120556 92768 120576
rect 92768 120556 92770 120576
rect 92714 120520 92770 120556
rect 58214 120384 58270 120440
rect 92806 120112 92862 120168
rect 58306 119840 58362 119896
rect 58214 119180 58270 119216
rect 58214 119160 58216 119180
rect 58216 119160 58268 119180
rect 58268 119160 58270 119180
rect 58306 118616 58362 118672
rect 92714 119160 92770 119216
rect 92806 118888 92862 118944
rect 92898 118480 92954 118536
rect 58398 118072 58454 118128
rect 58214 117392 58270 117448
rect 92714 117528 92770 117584
rect 92806 117256 92862 117312
rect 58306 116848 58362 116904
rect 58214 116168 58270 116224
rect 50854 115624 50910 115680
rect 58306 115624 58362 115680
rect 58398 115080 58454 115136
rect 50946 114400 51002 114456
rect 51130 113992 51186 114048
rect 51038 112768 51094 112824
rect 51222 113876 51278 113912
rect 51222 113856 51224 113876
rect 51224 113856 51276 113876
rect 51276 113856 51278 113876
rect 41838 95224 41894 95280
rect 22334 89784 22390 89840
rect 44414 84752 44470 84808
rect 22334 83120 22390 83176
rect 44414 76456 44470 76512
rect 61894 111136 61950 111192
rect 92714 116340 92716 116360
rect 92716 116340 92768 116360
rect 92768 116340 92770 116360
rect 92714 116304 92770 116340
rect 92806 115896 92862 115952
rect 92898 115488 92954 115544
rect 53338 79856 53394 79912
rect 44414 74688 44470 74744
rect 53338 69792 53394 69848
rect 53430 66528 53486 66584
rect 53982 66528 54038 66584
rect 44506 64760 44562 64816
rect 22334 63128 22390 63184
rect 49934 46264 49990 46320
rect 50026 43952 50082 44008
rect 49934 43544 49990 43600
rect 50026 42728 50082 42784
rect 49934 42476 49990 42512
rect 49934 42456 49936 42476
rect 49936 42456 49988 42476
rect 49988 42456 49990 42476
rect 49934 42048 49990 42104
rect 18102 41932 18158 41968
rect 18102 41912 18104 41932
rect 18104 41912 18156 41932
rect 18156 41912 18158 41932
rect 50026 40960 50082 41016
rect 49934 40708 49990 40744
rect 49934 40688 49936 40708
rect 49936 40688 49988 40708
rect 49988 40688 49990 40708
rect 50210 37288 50266 37344
rect 50026 33072 50082 33128
rect 18102 32392 18158 32448
rect 13318 20560 13374 20616
rect 50026 31848 50082 31904
rect 50026 27496 50082 27552
rect 50394 23280 50450 23336
rect 50302 21104 50358 21160
rect 50578 22056 50634 22112
rect 50486 19744 50542 19800
rect 50946 21920 51002 21976
rect 50854 20968 50910 21024
rect 53338 45176 53394 45232
rect 53246 44904 53302 44960
rect 51130 39736 51186 39792
rect 51222 39328 51278 39384
rect 51130 38512 51186 38568
rect 51222 38104 51278 38160
rect 51222 36744 51278 36800
rect 51130 36472 51186 36528
rect 51222 35656 51278 35712
rect 51222 35132 51278 35168
rect 51222 35112 51224 35132
rect 51224 35112 51276 35132
rect 51276 35112 51278 35132
rect 51130 34160 51186 34216
rect 51222 33888 51278 33944
rect 51222 32528 51278 32584
rect 51222 31440 51278 31496
rect 51222 30932 51224 30952
rect 51224 30932 51276 30952
rect 51276 30932 51278 30952
rect 51222 30896 51278 30932
rect 51130 29944 51186 30000
rect 51222 29692 51278 29728
rect 51222 29672 51224 29692
rect 51224 29672 51276 29692
rect 51276 29672 51278 29692
rect 51130 28720 51186 28776
rect 51222 28312 51278 28368
rect 51222 27088 51278 27144
rect 51130 26816 51186 26872
rect 51130 25728 51186 25784
rect 51222 25492 51224 25512
rect 51224 25492 51276 25512
rect 51276 25492 51278 25512
rect 51222 25456 51278 25492
rect 51130 24504 51186 24560
rect 51222 24232 51278 24288
rect 51222 22872 51278 22928
rect 59226 58368 59282 58424
rect 139450 235168 139506 235224
rect 134758 234508 134814 234544
rect 134758 234488 134760 234508
rect 134760 234488 134812 234508
rect 134812 234488 134814 234508
rect 101178 233944 101234 234000
rect 134758 233944 134814 234000
rect 134850 233400 134906 233456
rect 101362 233128 101418 233184
rect 101730 232856 101786 232912
rect 134758 232856 134814 232912
rect 142302 232992 142358 233048
rect 163554 235168 163610 235224
rect 185266 234488 185322 234544
rect 185174 233944 185230 234000
rect 177722 232720 177778 232776
rect 134850 232176 134906 232232
rect 101270 231904 101326 231960
rect 134758 231632 134814 231688
rect 101454 231496 101510 231552
rect 101730 231224 101786 231280
rect 134758 231108 134814 231144
rect 134758 231088 134760 231108
rect 134760 231088 134812 231108
rect 134812 231088 134814 231108
rect 134390 230544 134446 230600
rect 101730 230136 101786 230192
rect 101546 229728 101602 229784
rect 134298 230020 134354 230056
rect 134298 230000 134300 230020
rect 134300 230000 134352 230020
rect 134352 230000 134354 230020
rect 177722 232176 177778 232232
rect 142302 231904 142358 231960
rect 177722 231496 177778 231552
rect 142210 231224 142266 231280
rect 177722 230852 177724 230872
rect 177724 230852 177776 230872
rect 177776 230852 177778 230872
rect 177722 230816 177778 230852
rect 143682 230680 143738 230736
rect 177722 230408 177778 230464
rect 142946 230136 143002 230192
rect 177722 229592 177778 229648
rect 134390 229320 134446 229376
rect 101730 229184 101786 229240
rect 101454 228640 101510 228696
rect 134758 228776 134814 228832
rect 101730 228368 101786 228424
rect 134850 228268 134852 228288
rect 134852 228268 134904 228288
rect 134904 228268 134906 228288
rect 134850 228232 134906 228268
rect 143682 229492 143684 229512
rect 143684 229492 143736 229512
rect 143736 229492 143738 229512
rect 143682 229456 143738 229492
rect 177630 229184 177686 229240
rect 143590 228912 143646 228968
rect 176986 228504 177042 228560
rect 134758 227688 134814 227744
rect 101362 227416 101418 227472
rect 101454 227008 101510 227064
rect 135402 227144 135458 227200
rect 134390 226464 134446 226520
rect 101638 226328 101694 226384
rect 101546 225512 101602 225568
rect 101822 225648 101878 225704
rect 134758 225920 134814 225976
rect 143498 228232 143554 228288
rect 143682 227688 143738 227744
rect 177722 227960 177778 228016
rect 177630 227416 177686 227472
rect 143314 227144 143370 227200
rect 177170 226600 177226 226656
rect 143682 226464 143738 226520
rect 177722 226192 177778 226248
rect 143314 225920 143370 225976
rect 134666 225376 134722 225432
rect 134298 224832 134354 224888
rect 101086 224560 101142 224616
rect 100994 224424 101050 224480
rect 135402 224288 135458 224344
rect 177722 225412 177724 225432
rect 177724 225412 177776 225432
rect 177776 225412 177778 225432
rect 177722 225376 177778 225412
rect 143682 225240 143738 225296
rect 143314 224696 143370 224752
rect 177722 224968 177778 225024
rect 177170 224424 177226 224480
rect 101454 223472 101510 223528
rect 101362 222928 101418 222984
rect 100902 222792 100958 222848
rect 134482 223084 134538 223120
rect 134482 223064 134484 223084
rect 134484 223064 134536 223084
rect 134536 223064 134538 223084
rect 134666 221976 134722 222032
rect 101638 221840 101694 221896
rect 101546 221432 101602 221488
rect 101822 220616 101878 220672
rect 101270 220072 101326 220128
rect 100902 219936 100958 219992
rect 101362 218984 101418 219040
rect 101730 218848 101786 218904
rect 101178 217896 101234 217952
rect 100810 217352 100866 217408
rect 100718 215992 100774 216048
rect 100902 217216 100958 217272
rect 134482 217372 134538 217408
rect 134482 217352 134484 217372
rect 134484 217352 134536 217372
rect 134536 217352 134538 217372
rect 101362 216128 101418 216184
rect 100994 215040 101050 215096
rect 100810 214632 100866 214688
rect 100718 213408 100774 213464
rect 135402 223608 135458 223664
rect 142578 224152 142634 224208
rect 134850 222520 134906 222576
rect 135402 221432 135458 221488
rect 135402 220752 135458 220808
rect 135310 220208 135366 220264
rect 143682 223472 143738 223528
rect 177722 223744 177778 223800
rect 177630 223200 177686 223256
rect 143314 222928 143370 222984
rect 143682 222248 143738 222304
rect 177722 222384 177778 222440
rect 177630 221976 177686 222032
rect 143314 221704 143370 221760
rect 143682 221160 143738 221216
rect 143314 220480 143370 220536
rect 135402 219664 135458 219720
rect 135034 219120 135090 219176
rect 135310 218612 135312 218632
rect 135312 218612 135364 218632
rect 135364 218612 135366 218632
rect 135310 218576 135366 218612
rect 135402 217896 135458 217952
rect 135402 216808 135458 216864
rect 135494 216264 135550 216320
rect 135402 215720 135458 215776
rect 134850 215040 134906 215096
rect 135310 214532 135312 214552
rect 135312 214532 135364 214552
rect 135364 214532 135366 214552
rect 135310 214496 135366 214532
rect 177722 221024 177778 221080
rect 177630 220888 177686 220944
rect 177170 220208 177226 220264
rect 143682 219936 143738 219992
rect 143682 219256 143738 219312
rect 177722 219528 177778 219584
rect 177170 218984 177226 219040
rect 143130 218712 143186 218768
rect 143682 218168 143738 218224
rect 177722 218304 177778 218360
rect 177170 217896 177226 217952
rect 143498 217488 143554 217544
rect 143682 216944 143738 217000
rect 177998 217080 178054 217136
rect 177722 216672 177778 216728
rect 143130 216264 143186 216320
rect 143130 215740 143186 215776
rect 143130 215720 143132 215740
rect 143132 215720 143184 215740
rect 143184 215720 143186 215740
rect 142946 215176 143002 215232
rect 100994 213952 101050 214008
rect 134482 213952 134538 214008
rect 100902 213136 100958 213192
rect 134482 213408 134538 213464
rect 134482 212864 134538 212920
rect 100994 212320 101050 212376
rect 101270 211912 101326 211968
rect 134666 212184 134722 212240
rect 101178 211096 101234 211152
rect 101086 210688 101142 210744
rect 100994 210416 101050 210472
rect 134574 211640 134630 211696
rect 135034 211096 135090 211152
rect 134850 210552 134906 210608
rect 100994 209464 101050 209520
rect 101638 208920 101694 208976
rect 100994 206472 101050 206528
rect 99246 190696 99302 190752
rect 99154 189472 99210 189528
rect 101730 208376 101786 208432
rect 102098 207832 102154 207888
rect 101914 207560 101970 207616
rect 134206 207716 134262 207752
rect 134206 207696 134208 207716
rect 134208 207696 134260 207716
rect 134260 207696 134262 207716
rect 99522 193688 99578 193744
rect 134942 209328 134998 209384
rect 135126 210008 135182 210064
rect 135218 208240 135274 208296
rect 177722 215584 177778 215640
rect 177630 215448 177686 215504
rect 177170 214904 177226 214960
rect 143498 214496 143554 214552
rect 142946 213952 143002 214008
rect 177722 214088 177778 214144
rect 177630 213680 177686 213736
rect 143682 213272 143738 213328
rect 143682 212728 143738 212784
rect 177722 212864 177778 212920
rect 177170 212456 177226 212512
rect 143498 212184 143554 212240
rect 177722 211660 177778 211696
rect 177722 211640 177724 211660
rect 177724 211640 177776 211660
rect 177776 211640 177778 211660
rect 143682 211504 143738 211560
rect 177170 211232 177226 211288
rect 143682 210960 143738 211016
rect 177722 210552 177778 210608
rect 143590 210280 143646 210336
rect 142946 209736 143002 209792
rect 143682 209192 143738 209248
rect 135402 208784 135458 208840
rect 135310 207152 135366 207208
rect 167142 195184 167198 195240
rect 172294 208920 172350 208976
rect 177170 210008 177226 210064
rect 177722 209464 177778 209520
rect 185174 233400 185230 233456
rect 185174 232856 185230 232912
rect 185174 232312 185230 232368
rect 185266 231768 185322 231824
rect 185174 231224 185230 231280
rect 185266 230680 185322 230736
rect 185174 230000 185230 230056
rect 185174 229456 185230 229512
rect 185266 228912 185322 228968
rect 185174 228368 185230 228424
rect 185174 227824 185230 227880
rect 185266 227280 185322 227336
rect 185358 226736 185414 226792
rect 185266 226192 185322 226248
rect 185174 225512 185230 225568
rect 185266 224968 185322 225024
rect 185174 224424 185230 224480
rect 185266 223880 185322 223936
rect 185174 223336 185230 223392
rect 185082 222792 185138 222848
rect 185266 222248 185322 222304
rect 185174 221704 185230 221760
rect 185358 221160 185414 221216
rect 222342 231632 222398 231688
rect 215718 221160 215774 221216
rect 185174 220480 185230 220536
rect 185082 219936 185138 219992
rect 185818 219392 185874 219448
rect 185174 218848 185230 218904
rect 185174 218304 185230 218360
rect 184990 217760 185046 217816
rect 184806 215992 184862 216048
rect 185082 217216 185138 217272
rect 185174 216672 185230 216728
rect 185174 215448 185230 215504
rect 184898 214904 184954 214960
rect 185266 214360 185322 214416
rect 184990 213816 185046 213872
rect 185082 213272 185138 213328
rect 185174 212728 185230 212784
rect 185450 212184 185506 212240
rect 185358 211504 185414 211560
rect 185266 210960 185322 211016
rect 185174 210416 185230 210472
rect 185174 209872 185230 209928
rect 185726 209328 185782 209384
rect 185174 207152 185230 207208
rect 105778 192464 105834 192520
rect 99430 192328 99486 192384
rect 99338 188928 99394 188984
rect 99062 187704 99118 187760
rect 98970 186480 99026 186536
rect 98878 185256 98934 185312
rect 98602 182400 98658 182456
rect 99522 183624 99578 183680
rect 99430 181040 99486 181096
rect 99522 179816 99578 179872
rect 107158 190152 107214 190208
rect 106790 187840 106846 187896
rect 106790 185392 106846 185448
rect 183426 190696 183482 190752
rect 185910 208784 185966 208840
rect 186278 208240 186334 208296
rect 186094 207696 186150 207752
rect 183702 193144 183758 193200
rect 191982 192736 192038 192792
rect 183610 191920 183666 191976
rect 183518 189472 183574 189528
rect 191982 188656 192038 188712
rect 183334 188248 183390 188304
rect 183242 187024 183298 187080
rect 183150 185800 183206 185856
rect 183058 184576 183114 184632
rect 191154 186752 191210 186808
rect 128502 183760 128558 183816
rect 107158 183080 107214 183136
rect 182874 183352 182930 183408
rect 106974 180768 107030 180824
rect 98418 179272 98474 179328
rect 99522 177388 99578 177424
rect 106790 178320 106846 178376
rect 99522 177368 99524 177388
rect 99524 177368 99576 177388
rect 99576 177368 99578 177388
rect 98602 176688 98658 176744
rect 106606 176008 106662 176064
rect 98234 175328 98290 175384
rect 190602 182672 190658 182728
rect 191982 184712 192038 184768
rect 183150 182128 183206 182184
rect 183702 181040 183758 181096
rect 183702 179836 183758 179872
rect 190694 180768 190750 180824
rect 183702 179816 183704 179836
rect 183704 179816 183756 179836
rect 183756 179816 183758 179836
rect 191982 178728 192038 178784
rect 182506 178592 182562 178648
rect 182506 177368 182562 177424
rect 191982 176688 192038 176744
rect 183242 176144 183298 176200
rect 183702 174920 183758 174976
rect 191522 174784 191578 174840
rect 137518 174376 137574 174432
rect 99522 173716 99578 173752
rect 99522 173696 99524 173716
rect 99524 173696 99576 173716
rect 99576 173696 99578 173716
rect 106790 173716 106846 173752
rect 106790 173696 106792 173716
rect 106792 173696 106844 173716
rect 106844 173696 106846 173716
rect 183334 173696 183390 173752
rect 191982 172744 192038 172800
rect 99522 172472 99578 172528
rect 183518 172472 183574 172528
rect 106790 171384 106846 171440
rect 99430 171248 99486 171304
rect 182690 171268 182746 171304
rect 182690 171248 182692 171268
rect 182692 171248 182744 171268
rect 182744 171248 182746 171268
rect 99522 170024 99578 170080
rect 182506 170024 182562 170080
rect 106790 168936 106846 168992
rect 99430 168800 99486 168856
rect 99522 167712 99578 167768
rect 209922 190696 209978 190752
rect 211946 190424 212002 190480
rect 212498 183760 212554 183816
rect 211762 177096 211818 177152
rect 209830 170976 209886 171032
rect 191154 170704 191210 170760
rect 183702 168800 183758 168856
rect 106698 166624 106754 166680
rect 99522 166488 99578 166544
rect 99522 165264 99578 165320
rect 106790 164312 106846 164368
rect 99522 164040 99578 164096
rect 98970 162816 99026 162872
rect 98786 154384 98842 154440
rect 98786 99712 98842 99768
rect 98786 89920 98842 89976
rect 98694 87336 98750 87392
rect 98234 75504 98290 75560
rect 98786 62720 98842 62776
rect 99062 161592 99118 161648
rect 99154 160368 99210 160424
rect 99246 159144 99302 159200
rect 99430 157920 99486 157976
rect 99338 156696 99394 156752
rect 99522 155472 99578 155528
rect 183794 167712 183850 167768
rect 182874 166508 182930 166544
rect 182874 166488 182876 166508
rect 182876 166488 182928 166508
rect 182928 166488 182930 166508
rect 106882 161864 106938 161920
rect 183702 165264 183758 165320
rect 138162 164720 138218 164776
rect 128502 163768 128558 163824
rect 183058 164040 183114 164096
rect 183058 162816 183114 162872
rect 138162 160504 138218 160560
rect 107250 159552 107306 159608
rect 107158 157240 107214 157296
rect 182690 155492 182746 155528
rect 182690 155472 182692 155492
rect 182692 155472 182744 155492
rect 182744 155472 182746 155492
rect 106514 154928 106570 154984
rect 134850 140512 134906 140568
rect 100810 140104 100866 140160
rect 100902 139968 100958 140024
rect 135402 139988 135458 140024
rect 135402 139968 135404 139988
rect 135404 139968 135456 139988
rect 135456 139968 135458 139988
rect 134666 139424 134722 139480
rect 101178 138880 101234 138936
rect 101086 138608 101142 138664
rect 100994 137792 101050 137848
rect 135402 138764 135458 138800
rect 135402 138744 135404 138764
rect 135404 138744 135456 138764
rect 135456 138744 135458 138764
rect 134666 138200 134722 138256
rect 135402 137656 135458 137712
rect 101270 137268 101326 137304
rect 101270 137248 101272 137268
rect 101272 137248 101324 137268
rect 101324 137248 101326 137268
rect 135034 136976 135090 137032
rect 101822 136568 101878 136624
rect 101454 136160 101510 136216
rect 101730 135888 101786 135944
rect 143590 138472 143646 138528
rect 143314 138200 143370 138256
rect 143130 136840 143186 136896
rect 135310 136432 135366 136488
rect 135402 135888 135458 135944
rect 134850 135344 134906 135400
rect 101454 134800 101510 134856
rect 100902 134392 100958 134448
rect 134666 134664 134722 134720
rect 135402 134120 135458 134176
rect 101822 133712 101878 133768
rect 101730 133032 101786 133088
rect 101178 131944 101234 132000
rect 101546 131808 101602 131864
rect 101362 130312 101418 130368
rect 101270 128952 101326 129008
rect 100994 128408 101050 128464
rect 101178 127864 101234 127920
rect 101086 127728 101142 127784
rect 134114 133576 134170 133632
rect 135126 132896 135182 132952
rect 101822 132488 101878 132544
rect 134482 132352 134538 132408
rect 143590 137112 143646 137168
rect 143498 136296 143554 136352
rect 143406 135752 143462 135808
rect 143314 135208 143370 135264
rect 143590 134256 143646 134312
rect 143222 133984 143278 134040
rect 142946 133304 143002 133360
rect 135310 131808 135366 131864
rect 134850 131264 134906 131320
rect 101822 130720 101878 130776
rect 101730 129632 101786 129688
rect 134666 130604 134722 130640
rect 134666 130584 134668 130604
rect 134668 130584 134720 130604
rect 134720 130584 134722 130604
rect 135402 130040 135458 130096
rect 134666 129496 134722 129552
rect 135402 128816 135458 128872
rect 134666 128272 134722 128328
rect 134666 127748 134722 127784
rect 134666 127728 134668 127748
rect 134668 127728 134720 127748
rect 134720 127728 134722 127748
rect 135402 127184 135458 127240
rect 101822 126640 101878 126696
rect 101730 126232 101786 126288
rect 135402 126504 135458 126560
rect 135218 125960 135274 126016
rect 101454 125552 101510 125608
rect 135034 125416 135090 125472
rect 101638 124872 101694 124928
rect 101730 124736 101786 124792
rect 135402 124736 135458 124792
rect 143590 132796 143592 132816
rect 143592 132796 143644 132816
rect 143644 132796 143646 132816
rect 143590 132760 143646 132796
rect 143222 132216 143278 132272
rect 143590 131400 143646 131456
rect 142486 130992 142542 131048
rect 143590 130212 143592 130232
rect 143592 130212 143644 130232
rect 143644 130212 143646 130232
rect 143590 130176 143646 130212
rect 143038 129904 143094 129960
rect 142762 128836 142818 128872
rect 142762 128816 142764 128836
rect 142764 128816 142816 128836
rect 142816 128816 142818 128836
rect 143590 128716 143592 128736
rect 143592 128716 143644 128736
rect 143644 128716 143646 128736
rect 143590 128680 143646 128716
rect 143130 128000 143186 128056
rect 142486 127356 142488 127376
rect 142488 127356 142540 127376
rect 142540 127356 142542 127376
rect 142486 127320 142542 127356
rect 143314 126912 143370 126968
rect 143590 125960 143646 126016
rect 143038 125688 143094 125744
rect 134114 124192 134170 124248
rect 101914 123784 101970 123840
rect 101822 123376 101878 123432
rect 101638 122560 101694 122616
rect 101454 122016 101510 122072
rect 101086 121064 101142 121120
rect 101546 120676 101602 120712
rect 101546 120656 101548 120676
rect 101548 120656 101600 120676
rect 101600 120656 101602 120676
rect 134482 123648 134538 123704
rect 134482 122968 134538 123024
rect 142486 124364 142488 124384
rect 142488 124364 142540 124384
rect 142540 124364 142542 124384
rect 142486 124328 142542 124364
rect 143590 124600 143646 124656
rect 142762 123920 142818 123976
rect 134942 122424 134998 122480
rect 134482 121880 134538 121936
rect 101730 121472 101786 121528
rect 134666 121336 134722 121392
rect 135402 120676 135458 120712
rect 135402 120656 135404 120676
rect 135404 120656 135456 120676
rect 135456 120656 135458 120676
rect 134482 120112 134538 120168
rect 101270 119704 101326 119760
rect 101362 119316 101418 119352
rect 135402 119588 135458 119624
rect 135402 119568 135404 119588
rect 135404 119568 135456 119588
rect 135456 119568 135458 119588
rect 101362 119296 101364 119316
rect 101364 119296 101416 119316
rect 101416 119296 101418 119316
rect 134666 118888 134722 118944
rect 101362 118480 101418 118536
rect 134666 118344 134722 118400
rect 101730 118072 101786 118128
rect 134850 117800 134906 117856
rect 101178 117392 101234 117448
rect 101086 116712 101142 116768
rect 100994 116576 101050 116632
rect 134758 116576 134814 116632
rect 101086 115624 101142 115680
rect 100994 115216 101050 115272
rect 101822 114400 101878 114456
rect 101638 113720 101694 113776
rect 100994 112496 101050 112552
rect 99246 95496 99302 95552
rect 102006 113856 102062 113912
rect 108446 111136 108502 111192
rect 134022 111136 134078 111192
rect 99522 98488 99578 98544
rect 106790 98488 106846 98544
rect 99430 96992 99486 97048
rect 106790 96176 106846 96232
rect 99338 94272 99394 94328
rect 99154 93592 99210 93648
rect 99062 92368 99118 92424
rect 98970 91144 99026 91200
rect 106514 93864 106570 93920
rect 106790 91416 106846 91472
rect 99522 88696 99578 88752
rect 99522 85296 99578 85352
rect 99522 84616 99578 84672
rect 128502 89784 128558 89840
rect 106790 89104 106846 89160
rect 106790 86792 106846 86848
rect 107802 84344 107858 84400
rect 99430 83936 99486 83992
rect 99522 82712 99578 82768
rect 106790 82068 106792 82088
rect 106792 82068 106844 82088
rect 106844 82068 106846 82088
rect 106790 82032 106846 82068
rect 99522 81488 99578 81544
rect 99522 79720 99578 79776
rect 106790 79720 106846 79776
rect 99522 77952 99578 78008
rect 106514 77408 106570 77464
rect 99522 76728 99578 76784
rect 106790 74996 106792 75016
rect 106792 74996 106844 75016
rect 106844 74996 106846 75016
rect 106790 74960 106846 74996
rect 99430 74280 99486 74336
rect 99522 73772 99524 73792
rect 99524 73772 99576 73792
rect 99576 73772 99578 73792
rect 99522 73736 99578 73772
rect 99522 72512 99578 72568
rect 99522 71036 99578 71072
rect 99522 71016 99524 71036
rect 99524 71016 99576 71036
rect 99576 71016 99578 71036
rect 99522 69792 99578 69848
rect 98970 68296 99026 68352
rect 99062 67072 99118 67128
rect 99154 65848 99210 65904
rect 99246 64624 99302 64680
rect 99338 63400 99394 63456
rect 99522 61496 99578 61552
rect 99522 60000 99578 60056
rect 80754 46808 80810 46864
rect 77810 46672 77866 46728
rect 74866 46400 74922 46456
rect 73394 46264 73450 46320
rect 76338 46128 76394 46184
rect 79282 46536 79338 46592
rect 85722 46264 85778 46320
rect 87102 46128 87158 46184
rect 58950 44360 59006 44416
rect 58214 43816 58270 43872
rect 58214 42592 58270 42648
rect 59042 43136 59098 43192
rect 58306 42048 58362 42104
rect 58214 41368 58270 41424
rect 58306 40824 58362 40880
rect 58398 40144 58454 40200
rect 58214 39600 58270 39656
rect 58306 39076 58362 39112
rect 58306 39056 58308 39076
rect 58308 39056 58360 39076
rect 58360 39056 58362 39076
rect 58214 38376 58270 38432
rect 58214 37152 58270 37208
rect 58398 37832 58454 37888
rect 58306 36608 58362 36664
rect 58214 36064 58270 36120
rect 58306 35384 58362 35440
rect 58306 34840 58362 34896
rect 58214 34160 58270 34216
rect 59226 33616 59282 33672
rect 58214 33072 58270 33128
rect 58306 32392 58362 32448
rect 58214 31848 58270 31904
rect 58306 31168 58362 31224
rect 58306 30624 58362 30680
rect 58214 30080 58270 30136
rect 58398 29400 58454 29456
rect 58214 28856 58270 28912
rect 58306 28176 58362 28232
rect 58306 27632 58362 27688
rect 58214 27088 58270 27144
rect 58214 26408 58270 26464
rect 58306 25864 58362 25920
rect 59042 25184 59098 25240
rect 59502 24640 59558 24696
rect 59410 24096 59466 24152
rect 58214 23416 58270 23472
rect 58306 22872 58362 22928
rect 53982 22736 54038 22792
rect 51038 20424 51094 20480
rect 50762 19200 50818 19256
rect 92714 44360 92770 44416
rect 92806 44224 92862 44280
rect 92714 43136 92770 43192
rect 92898 42864 92954 42920
rect 92806 42456 92862 42512
rect 92714 41640 92770 41696
rect 92806 41096 92862 41152
rect 92714 40144 92770 40200
rect 92806 40008 92862 40064
rect 92714 39056 92770 39112
rect 92806 38648 92862 38704
rect 92898 38240 92954 38296
rect 92714 37424 92770 37480
rect 92806 37016 92862 37072
rect 92714 36064 92770 36120
rect 92806 35928 92862 35984
rect 92714 34840 92770 34896
rect 92806 34568 92862 34624
rect 92714 33616 92770 33672
rect 92806 33344 92862 33400
rect 92898 32936 92954 32992
rect 92714 31848 92770 31904
rect 92806 31712 92862 31768
rect 92714 30624 92770 30680
rect 92806 30488 92862 30544
rect 92714 29400 92770 29456
rect 92898 29128 92954 29184
rect 92806 28720 92862 28776
rect 92714 27632 92770 27688
rect 92806 27360 92862 27416
rect 92898 26680 92954 26736
rect 92714 26272 92770 26328
rect 92898 25184 92954 25240
rect 92806 24912 92862 24968
rect 92714 24504 92770 24560
rect 92714 23688 92770 23744
rect 92806 23280 92862 23336
rect 58214 22192 58270 22248
rect 92714 22192 92770 22248
rect 92806 22056 92862 22112
rect 58306 21648 58362 21704
rect 58214 21104 58270 21160
rect 92714 21104 92770 21160
rect 61710 20968 61766 21024
rect 63274 20968 63330 21024
rect 64746 20968 64802 21024
rect 65758 20968 65814 21024
rect 62722 20832 62778 20888
rect 66862 20832 66918 20888
rect 106790 72648 106846 72704
rect 106698 70336 106754 70392
rect 134942 117256 134998 117312
rect 134850 115488 134906 115544
rect 143590 123276 143592 123296
rect 143592 123276 143644 123296
rect 143644 123276 143646 123296
rect 143590 123240 143646 123276
rect 142854 122696 142910 122752
rect 143038 121744 143094 121800
rect 142762 121472 142818 121528
rect 142946 120556 142948 120576
rect 142948 120556 143000 120576
rect 143000 120556 143002 120576
rect 142946 120520 143002 120556
rect 143590 120248 143646 120304
rect 143590 119196 143592 119216
rect 143592 119196 143644 119216
rect 143644 119196 143646 119216
rect 143590 119160 143646 119196
rect 143590 119060 143592 119080
rect 143592 119060 143644 119080
rect 143644 119060 143646 119080
rect 143590 119024 143646 119060
rect 142578 118480 142634 118536
rect 142578 117664 142634 117720
rect 143222 117256 143278 117312
rect 135034 116032 135090 116088
rect 142946 116340 142948 116360
rect 142948 116340 143000 116360
rect 143000 116340 143002 116360
rect 142946 116304 143002 116340
rect 143590 116032 143646 116088
rect 142762 115488 142818 115544
rect 135126 114808 135182 114864
rect 135310 114264 135366 114320
rect 135218 113176 135274 113232
rect 135402 113740 135458 113776
rect 135402 113720 135404 113740
rect 135404 113720 135456 113740
rect 135456 113720 135458 113740
rect 183150 161592 183206 161648
rect 183242 160368 183298 160424
rect 183334 159144 183390 159200
rect 183518 157920 183574 157976
rect 183426 156696 183482 156752
rect 191982 168664 192038 168720
rect 191890 166760 191946 166816
rect 212682 164856 212738 164912
rect 191338 164720 191394 164776
rect 211762 163768 211818 163824
rect 191982 162680 192038 162736
rect 191338 160776 191394 160832
rect 190050 158736 190106 158792
rect 211946 157104 212002 157160
rect 189958 156696 190014 156752
rect 183610 154384 183666 154440
rect 191982 154792 192038 154848
rect 184990 140104 185046 140160
rect 177722 138492 177778 138528
rect 185082 139968 185138 140024
rect 185358 138880 185414 138936
rect 185266 138608 185322 138664
rect 177722 138472 177724 138492
rect 177724 138472 177776 138492
rect 177776 138472 177778 138492
rect 177630 138200 177686 138256
rect 185174 137792 185230 137848
rect 177722 137012 177724 137032
rect 177724 137012 177776 137032
rect 177776 137012 177778 137032
rect 177722 136976 177778 137012
rect 177630 136840 177686 136896
rect 177722 136296 177778 136352
rect 177722 135480 177778 135536
rect 177630 135208 177686 135264
rect 185450 137248 185506 137304
rect 185174 136568 185230 136624
rect 177722 134292 177724 134312
rect 177724 134292 177776 134312
rect 177776 134292 177778 134312
rect 177722 134256 177778 134292
rect 185266 136024 185322 136080
rect 185358 135908 185414 135944
rect 185358 135888 185360 135908
rect 185360 135888 185412 135908
rect 185412 135888 185414 135908
rect 185174 134800 185230 134856
rect 185082 134392 185138 134448
rect 177722 133848 177778 133904
rect 177630 133440 177686 133496
rect 185174 133712 185230 133768
rect 185818 133032 185874 133088
rect 177722 132624 177778 132680
rect 177630 132216 177686 132272
rect 185726 131944 185782 132000
rect 185542 131672 185598 131728
rect 177722 131264 177778 131320
rect 177630 130992 177686 131048
rect 185358 130720 185414 130776
rect 185266 130312 185322 130368
rect 177722 130196 177778 130232
rect 177722 130176 177724 130196
rect 177724 130176 177776 130196
rect 177776 130176 177778 130196
rect 177630 129768 177686 129824
rect 185174 129632 185230 129688
rect 185910 132488 185966 132544
rect 185450 128952 185506 129008
rect 177722 128716 177724 128736
rect 177724 128716 177776 128736
rect 177776 128716 177778 128736
rect 177722 128680 177778 128716
rect 177630 128408 177686 128464
rect 185174 128408 185230 128464
rect 177354 128000 177410 128056
rect 185358 127864 185414 127920
rect 185266 127592 185322 127648
rect 177170 127184 177226 127240
rect 177722 126912 177778 126968
rect 185174 126232 185230 126288
rect 177722 125996 177724 126016
rect 177724 125996 177776 126016
rect 177776 125996 177778 126016
rect 177722 125960 177778 125996
rect 177630 125552 177686 125608
rect 177170 124192 177226 124248
rect 177722 124464 177778 124520
rect 185450 126640 185506 126696
rect 185174 125552 185230 125608
rect 185358 124872 185414 124928
rect 185266 124736 185322 124792
rect 177630 123920 177686 123976
rect 185910 123784 185966 123840
rect 185726 123376 185782 123432
rect 177722 122968 177778 123024
rect 177630 122696 177686 122752
rect 185542 122152 185598 122208
rect 177722 121744 177778 121800
rect 177630 121472 177686 121528
rect 185358 121472 185414 121528
rect 185174 120792 185230 120848
rect 177722 120556 177724 120576
rect 177724 120556 177776 120576
rect 177776 120556 177778 120576
rect 177722 120520 177778 120556
rect 177630 120112 177686 120168
rect 177722 119024 177778 119080
rect 177722 118752 177778 118808
rect 177630 118480 177686 118536
rect 177722 117528 177778 117584
rect 177630 117256 177686 117312
rect 177722 116340 177724 116360
rect 177724 116340 177776 116360
rect 177776 116340 177778 116360
rect 177722 116304 177778 116340
rect 177722 115896 177778 115952
rect 177078 115488 177134 115544
rect 185266 120692 185268 120712
rect 185268 120692 185320 120712
rect 185320 120692 185322 120712
rect 185266 120656 185322 120692
rect 185818 122560 185874 122616
rect 185266 119704 185322 119760
rect 185174 119316 185230 119352
rect 185174 119296 185176 119316
rect 185176 119296 185228 119316
rect 185228 119296 185230 119316
rect 185266 118480 185322 118536
rect 185174 117936 185230 117992
rect 185358 117392 185414 117448
rect 185266 116712 185322 116768
rect 185174 116476 185176 116496
rect 185176 116476 185228 116496
rect 185228 116476 185230 116496
rect 185174 116440 185230 116476
rect 185266 115624 185322 115680
rect 185174 115216 185230 115272
rect 185818 114400 185874 114456
rect 185174 112632 185230 112688
rect 183334 95496 183390 95552
rect 186002 113856 186058 113912
rect 186186 113720 186242 113776
rect 183702 99168 183758 99224
rect 191982 98760 192038 98816
rect 183610 97944 183666 98000
rect 183518 96720 183574 96776
rect 191982 94680 192038 94736
rect 183426 94272 183482 94328
rect 183242 93048 183298 93104
rect 183150 91824 183206 91880
rect 183058 90600 183114 90656
rect 191154 92776 191210 92832
rect 190786 90736 190842 90792
rect 182874 89376 182930 89432
rect 183518 88152 183574 88208
rect 191706 88696 191762 88752
rect 183702 87064 183758 87120
rect 191614 86792 191670 86848
rect 183702 85840 183758 85896
rect 183702 84636 183758 84672
rect 191982 84752 192038 84808
rect 183702 84616 183704 84636
rect 183704 84616 183756 84636
rect 183756 84616 183758 84636
rect 182506 83392 182562 83448
rect 191982 82712 192038 82768
rect 183702 82168 183758 82224
rect 183242 80944 183298 81000
rect 191890 80808 191946 80864
rect 136874 80400 136930 80456
rect 183702 79720 183758 79776
rect 191982 78768 192038 78824
rect 183518 78496 183574 78552
rect 183058 77272 183114 77328
rect 209830 96856 209886 96912
rect 211762 96448 211818 96504
rect 211854 89784 211910 89840
rect 220318 215176 220374 215232
rect 218294 209600 218350 209656
rect 218386 135888 218442 135944
rect 218294 127320 218350 127376
rect 216914 117256 216970 117312
rect 217558 117256 217614 117312
rect 212038 83120 212094 83176
rect 209830 76864 209886 76920
rect 191982 76728 192038 76784
rect 183242 76048 183298 76104
rect 183702 74824 183758 74880
rect 183702 73756 183758 73792
rect 183702 73736 183704 73756
rect 183704 73736 183756 73756
rect 183756 73736 183758 73756
rect 191522 74688 191578 74744
rect 183702 72512 183758 72568
rect 183702 71288 183758 71344
rect 128502 69792 128558 69848
rect 106606 67888 106662 67944
rect 182874 70064 182930 70120
rect 183058 68840 183114 68896
rect 136874 66528 136930 66584
rect 106514 65576 106570 65632
rect 106606 63264 106662 63320
rect 107158 60952 107214 61008
rect 182690 60428 182746 60464
rect 182690 60408 182692 60428
rect 182692 60408 182744 60428
rect 182744 60408 182746 60428
rect 101362 46536 101418 46592
rect 101270 44768 101326 44824
rect 100810 43408 100866 43464
rect 101730 45856 101786 45912
rect 101822 45176 101878 45232
rect 101638 43952 101694 44008
rect 101730 42728 101786 42784
rect 100902 42184 100958 42240
rect 100810 40960 100866 41016
rect 100994 41504 101050 41560
rect 101086 40280 101142 40336
rect 100994 39736 101050 39792
rect 101178 39056 101234 39112
rect 100994 38512 101050 38568
rect 100534 37832 100590 37888
rect 100994 37288 101050 37344
rect 100902 36608 100958 36664
rect 100718 35384 100774 35440
rect 134666 36628 134722 36664
rect 134666 36608 134668 36628
rect 134668 36608 134720 36628
rect 134720 36608 134722 36628
rect 100994 36064 101050 36120
rect 101086 34840 101142 34896
rect 100994 34160 101050 34216
rect 100810 33752 100866 33808
rect 134666 33788 134668 33808
rect 134668 33788 134720 33808
rect 134720 33788 134722 33808
rect 134666 33752 134722 33788
rect 100994 33072 101050 33128
rect 100902 32392 100958 32448
rect 100810 31168 100866 31224
rect 100994 31848 101050 31904
rect 101086 30624 101142 30680
rect 100994 29944 101050 30000
rect 101730 29400 101786 29456
rect 100994 28196 101050 28232
rect 100994 28176 100996 28196
rect 100996 28176 101048 28196
rect 101048 28176 101050 28196
rect 101914 28720 101970 28776
rect 100994 27496 101050 27552
rect 101178 26952 101234 27008
rect 101086 26272 101142 26328
rect 100994 25728 101050 25784
rect 101086 25048 101142 25104
rect 100994 24504 101050 24560
rect 100994 23824 101050 23880
rect 134482 23688 134538 23744
rect 101086 23280 101142 23336
rect 101178 22600 101234 22656
rect 100994 22192 101050 22248
rect 101086 21512 101142 21568
rect 100994 19764 101050 19800
rect 100994 19744 100996 19764
rect 100996 19744 101048 19764
rect 101048 19744 101050 19764
rect 134666 19744 134722 19800
rect 135034 24776 135090 24832
rect 135034 22464 135090 22520
rect 135402 46264 135458 46320
rect 135218 43428 135274 43464
rect 135218 43408 135220 43428
rect 135220 43408 135272 43428
rect 135272 43408 135274 43428
rect 135218 42204 135274 42240
rect 135218 42184 135220 42204
rect 135220 42184 135272 42204
rect 135272 42184 135274 42204
rect 135218 40844 135274 40880
rect 135218 40824 135220 40844
rect 135220 40824 135272 40844
rect 135272 40824 135274 40844
rect 135218 40008 135274 40064
rect 135218 38784 135274 38840
rect 135218 35268 135274 35304
rect 135218 35248 135220 35268
rect 135220 35248 135272 35268
rect 135272 35248 135274 35268
rect 135218 34432 135274 34488
rect 135218 32412 135274 32448
rect 135218 32392 135220 32412
rect 135220 32392 135272 32412
rect 135272 32392 135274 32412
rect 135218 31188 135274 31224
rect 135218 31168 135220 31188
rect 135220 31168 135272 31188
rect 135272 31168 135274 31188
rect 135218 30624 135274 30680
rect 135218 29264 135274 29320
rect 135218 26972 135274 27008
rect 135218 26952 135220 26972
rect 135220 26952 135272 26972
rect 135272 26952 135274 26972
rect 135218 26000 135274 26056
rect 135402 45448 135458 45504
rect 135402 45060 135458 45096
rect 135402 45040 135404 45060
rect 135404 45040 135456 45060
rect 135456 45040 135458 45060
rect 135402 44788 135458 44824
rect 135402 44768 135404 44788
rect 135404 44768 135456 44788
rect 135456 44768 135458 44788
rect 135402 43680 135458 43736
rect 135402 42456 135458 42512
rect 135402 41232 135458 41288
rect 154262 46128 154318 46184
rect 191982 72784 192038 72840
rect 190786 70744 190842 70800
rect 183150 67616 183206 67672
rect 183242 66392 183298 66448
rect 183334 65168 183390 65224
rect 183426 63944 183482 64000
rect 190970 68704 191026 68760
rect 191338 66800 191394 66856
rect 191522 64760 191578 64816
rect 212682 63164 212684 63184
rect 212684 63164 212736 63184
rect 212736 63164 212738 63184
rect 212682 63128 212738 63164
rect 183610 62720 183666 62776
rect 189958 62720 190014 62776
rect 183702 61516 183758 61552
rect 183702 61496 183704 61516
rect 183704 61496 183756 61516
rect 183756 61496 183758 61516
rect 191982 60816 192038 60872
rect 164750 46944 164806 47000
rect 161898 46808 161954 46864
rect 158954 46672 159010 46728
rect 157574 46264 157630 46320
rect 160334 46400 160390 46456
rect 163278 46536 163334 46592
rect 169902 46128 169958 46184
rect 171374 44768 171430 44824
rect 143682 44668 143684 44688
rect 143684 44668 143736 44688
rect 143736 44668 143738 44688
rect 143682 44632 143738 44668
rect 172938 44632 172994 44688
rect 143498 44088 143554 44144
rect 142302 43272 142358 43328
rect 142210 43000 142266 43056
rect 142762 42456 142818 42512
rect 143406 41812 143408 41832
rect 143408 41812 143460 41832
rect 143460 41812 143462 41832
rect 143406 41776 143462 41812
rect 143314 41232 143370 41288
rect 135402 39464 135458 39520
rect 143682 40452 143684 40472
rect 143684 40452 143736 40472
rect 143736 40452 143738 40472
rect 143682 40416 143738 40452
rect 142486 40008 142542 40064
rect 143682 39056 143738 39112
rect 142854 38920 142910 38976
rect 135402 38260 135458 38296
rect 135402 38240 135404 38260
rect 135404 38240 135456 38260
rect 135456 38240 135458 38260
rect 143406 38240 143462 38296
rect 135402 37868 135404 37888
rect 135404 37868 135456 37888
rect 135456 37868 135458 37888
rect 135402 37832 135458 37868
rect 135402 36880 135458 36936
rect 135402 35656 135458 35712
rect 143682 37460 143684 37480
rect 143684 37460 143736 37480
rect 143736 37460 143738 37480
rect 143682 37424 143738 37460
rect 143498 36880 143554 36936
rect 143682 36064 143738 36120
rect 143038 35928 143094 35984
rect 135402 33888 135458 33944
rect 135402 32664 135458 32720
rect 135402 31440 135458 31496
rect 143682 34840 143738 34896
rect 142394 34568 142450 34624
rect 143682 33616 143738 33672
rect 143314 33344 143370 33400
rect 142762 32936 142818 32992
rect 143682 32156 143684 32176
rect 143684 32156 143736 32176
rect 143736 32156 143738 32176
rect 143682 32120 143738 32156
rect 142578 31712 142634 31768
rect 135402 29808 135458 29864
rect 143682 30624 143738 30680
rect 142762 30488 142818 30544
rect 143682 29400 143738 29456
rect 143590 29128 143646 29184
rect 142762 28720 142818 28776
rect 135402 28468 135458 28504
rect 135402 28448 135404 28468
rect 135404 28448 135456 28468
rect 135456 28448 135458 28468
rect 135402 28332 135458 28368
rect 135402 28312 135404 28332
rect 135404 28312 135456 28332
rect 135456 28312 135458 28332
rect 135402 27224 135458 27280
rect 143682 27940 143684 27960
rect 143684 27940 143736 27960
rect 143736 27940 143738 27960
rect 143682 27904 143738 27940
rect 143406 27532 143408 27552
rect 143408 27532 143460 27552
rect 143460 27532 143462 27552
rect 143406 27496 143462 27532
rect 135402 25592 135458 25648
rect 143682 26408 143738 26464
rect 143590 26272 143646 26328
rect 143130 25220 143132 25240
rect 143132 25220 143184 25240
rect 143184 25220 143186 25240
rect 143130 25184 143186 25220
rect 143682 25048 143738 25104
rect 143498 24504 143554 24560
rect 135402 24368 135458 24424
rect 143682 23996 143684 24016
rect 143684 23996 143736 24016
rect 143736 23996 143738 24016
rect 143682 23960 143738 23996
rect 143590 23280 143646 23336
rect 135402 23008 135458 23064
rect 135310 22600 135366 22656
rect 135126 21920 135182 21976
rect 142762 22464 142818 22520
rect 143314 22056 143370 22112
rect 134942 21104 134998 21160
rect 143682 21104 143738 21160
rect 146258 20968 146314 21024
rect 147730 20968 147786 21024
rect 148742 20968 148798 21024
rect 145706 20832 145762 20888
rect 134850 20696 134906 20752
rect 134758 19472 134814 19528
rect 101086 19200 101142 19256
rect 150536 20696 150592 20752
rect 149754 18248 149810 18304
rect 129054 17024 129110 17080
rect 185910 46128 185966 46184
rect 177262 39600 177318 39656
rect 177262 39056 177318 39112
rect 177354 38376 177410 38432
rect 177446 36608 177502 36664
rect 177446 36064 177502 36120
rect 177354 35384 177410 35440
rect 177262 34840 177318 34896
rect 177446 30624 177502 30680
rect 177262 29400 177318 29456
rect 177446 28176 177502 28232
rect 177354 27088 177410 27144
rect 177354 24096 177410 24152
rect 177354 22872 177410 22928
rect 185174 45448 185230 45504
rect 177722 44360 177778 44416
rect 185818 44904 185874 44960
rect 185450 44768 185506 44824
rect 177722 43852 177724 43872
rect 177724 43852 177776 43872
rect 177776 43852 177778 43872
rect 177722 43816 177778 43852
rect 185174 43680 185230 43736
rect 184990 43408 185046 43464
rect 177722 43172 177724 43192
rect 177724 43172 177776 43192
rect 177776 43172 177778 43192
rect 177722 43136 177778 43172
rect 177814 42592 177870 42648
rect 177722 42048 177778 42104
rect 185174 42456 185230 42512
rect 185082 42048 185138 42104
rect 177722 41368 177778 41424
rect 177630 40824 177686 40880
rect 184990 40552 185046 40608
rect 177722 40144 177778 40200
rect 185174 41232 185230 41288
rect 185266 40008 185322 40064
rect 185174 39328 185230 39384
rect 185266 38784 185322 38840
rect 185174 38104 185230 38160
rect 177722 37832 177778 37888
rect 184990 37832 185046 37888
rect 177722 37152 177778 37208
rect 185174 36880 185230 36936
rect 185082 36472 185138 36528
rect 184898 35248 184954 35304
rect 177722 34160 177778 34216
rect 177630 33616 177686 33672
rect 177722 33072 177778 33128
rect 185450 35656 185506 35712
rect 185266 34432 185322 34488
rect 185174 33888 185230 33944
rect 184990 33752 185046 33808
rect 177814 32392 177870 32448
rect 185174 32664 185230 32720
rect 185082 32256 185138 32312
rect 177722 31848 177778 31904
rect 177630 31168 177686 31224
rect 184990 30896 185046 30952
rect 177722 30080 177778 30136
rect 185174 31440 185230 31496
rect 185266 30216 185322 30272
rect 185174 29672 185230 29728
rect 185358 28992 185414 29048
rect 177722 28856 177778 28912
rect 185266 28448 185322 28504
rect 185174 28196 185230 28232
rect 185174 28176 185176 28196
rect 185176 28176 185228 28196
rect 185228 28176 185230 28196
rect 177722 27632 177778 27688
rect 185174 27224 185230 27280
rect 185818 26816 185874 26872
rect 177630 26408 177686 26464
rect 185266 26000 185322 26056
rect 177722 25864 177778 25920
rect 185726 25592 185782 25648
rect 177722 25220 177724 25240
rect 177724 25220 177776 25240
rect 177776 25220 177778 25240
rect 177722 25184 177778 25220
rect 185174 24776 185230 24832
rect 177814 24640 177870 24696
rect 185266 24096 185322 24152
rect 185266 23552 185322 23608
rect 177630 23416 177686 23472
rect 185174 22872 185230 22928
rect 185266 22600 185322 22656
rect 177630 22192 177686 22248
rect 185174 22328 185230 22384
rect 177722 21648 177778 21704
rect 222342 205384 222398 205440
rect 220410 179136 220466 179192
rect 221698 152888 221754 152944
rect 222342 126776 222398 126832
rect 222342 100528 222398 100584
rect 222342 74280 222398 74336
rect 222250 48032 222306 48088
rect 220318 21920 220374 21976
rect 177722 21104 177778 21160
rect 185174 19764 185230 19800
rect 185174 19744 185176 19764
rect 185176 19744 185228 19764
rect 185228 19744 185230 19764
rect 185266 19472 185322 19528
rect 211394 18420 211396 18440
rect 211396 18420 211448 18440
rect 211448 18420 211450 18440
rect 211394 18384 211450 18420
rect 201826 17024 201882 17080
<< metal3 >>
rect 23566 236524 23572 236588
rect 23636 236586 23642 236588
rect 33369 236586 33435 236589
rect 23636 236584 33435 236586
rect 23636 236528 33374 236584
rect 33430 236528 33435 236584
rect 23636 236526 33435 236528
rect 23636 236524 23642 236526
rect 33369 236523 33435 236526
rect 79553 235226 79619 235229
rect 139445 235228 139511 235229
rect 88518 235226 88524 235228
rect 79553 235224 88524 235226
rect 79553 235168 79558 235224
rect 79614 235168 88524 235224
rect 79553 235166 88524 235168
rect 79553 235163 79619 235166
rect 88518 235164 88524 235166
rect 88588 235164 88594 235228
rect 139445 235224 139492 235228
rect 139556 235226 139562 235228
rect 163549 235226 163615 235229
rect 171318 235226 171324 235228
rect 139445 235168 139450 235224
rect 139445 235164 139492 235168
rect 139556 235166 139602 235226
rect 163549 235224 171324 235226
rect 163549 235168 163554 235224
rect 163610 235168 171324 235224
rect 163549 235166 171324 235168
rect 139556 235164 139562 235166
rect 139445 235163 139511 235164
rect 163549 235163 163615 235166
rect 171318 235164 171324 235166
rect 171388 235164 171394 235228
rect 50573 234546 50639 234549
rect 134753 234546 134819 234549
rect 47524 234544 50639 234546
rect 47524 234488 50578 234544
rect 50634 234488 50639 234544
rect 47524 234486 50639 234488
rect 131796 234544 134819 234546
rect 131796 234488 134758 234544
rect 134814 234488 134819 234544
rect 131796 234486 134819 234488
rect 50573 234483 50639 234486
rect 134753 234483 134819 234486
rect 185261 234546 185327 234549
rect 185261 234544 187916 234546
rect 185261 234488 185266 234544
rect 185322 234488 187916 234544
rect 185261 234486 187916 234488
rect 185261 234483 185327 234486
rect 51217 234002 51283 234005
rect 47524 234000 51283 234002
rect 47524 233944 51222 234000
rect 51278 233944 51283 234000
rect 47524 233942 51283 233944
rect 51217 233939 51283 233942
rect 101173 234002 101239 234005
rect 134753 234002 134819 234005
rect 101173 234000 104012 234002
rect 101173 233944 101178 234000
rect 101234 233944 104012 234000
rect 101173 233942 104012 233944
rect 131796 234000 134819 234002
rect 131796 233944 134758 234000
rect 134814 233944 134819 234000
rect 131796 233942 134819 233944
rect 101173 233939 101239 233942
rect 134753 233939 134819 233942
rect 185169 234002 185235 234005
rect 185169 234000 187916 234002
rect 185169 233944 185174 234000
rect 185230 233944 187916 234000
rect 185169 233942 187916 233944
rect 185169 233939 185235 233942
rect 51217 233458 51283 233461
rect 134845 233458 134911 233461
rect 47524 233456 51283 233458
rect 47524 233400 51222 233456
rect 51278 233400 51283 233456
rect 47524 233398 51283 233400
rect 131796 233456 134911 233458
rect 131796 233400 134850 233456
rect 134906 233400 134911 233456
rect 131796 233398 134911 233400
rect 51217 233395 51283 233398
rect 134845 233395 134911 233398
rect 185169 233458 185235 233461
rect 185169 233456 187916 233458
rect 185169 233400 185174 233456
rect 185230 233400 187916 233456
rect 185169 233398 187916 233400
rect 185169 233395 185235 233398
rect 101357 233186 101423 233189
rect 103982 233186 104042 233360
rect 101357 233184 104042 233186
rect 101357 233128 101362 233184
rect 101418 233128 104042 233184
rect 101357 233126 104042 233128
rect 101357 233123 101423 233126
rect 58117 233050 58183 233053
rect 142297 233050 142363 233053
rect 58117 233048 60986 233050
rect 58117 232992 58122 233048
rect 58178 232992 60986 233048
rect 58117 232990 60986 232992
rect 58117 232987 58183 232990
rect 9896 232914 10376 232944
rect 13313 232914 13379 232917
rect 50021 232914 50087 232917
rect 9896 232912 13379 232914
rect 9896 232856 13318 232912
rect 13374 232856 13379 232912
rect 9896 232854 13379 232856
rect 47524 232912 50087 232914
rect 47524 232856 50026 232912
rect 50082 232856 50087 232912
rect 47524 232854 50087 232856
rect 9896 232824 10376 232854
rect 13313 232851 13379 232854
rect 50021 232851 50087 232854
rect 60926 232476 60986 232990
rect 142297 233048 145074 233050
rect 142297 232992 142302 233048
rect 142358 232992 145074 233048
rect 142297 232990 145074 232992
rect 142297 232987 142363 232990
rect 101725 232914 101791 232917
rect 134753 232914 134819 232917
rect 101725 232912 104012 232914
rect 101725 232856 101730 232912
rect 101786 232856 104012 232912
rect 101725 232854 104012 232856
rect 131796 232912 134819 232914
rect 131796 232856 134758 232912
rect 134814 232856 134819 232912
rect 131796 232854 134819 232856
rect 101725 232851 101791 232854
rect 134753 232851 134819 232854
rect 92709 232506 92775 232509
rect 90764 232504 92775 232506
rect 90764 232448 92714 232504
rect 92770 232448 92775 232504
rect 145014 232476 145074 232990
rect 185169 232914 185235 232917
rect 185169 232912 187916 232914
rect 185169 232856 185174 232912
rect 185230 232856 187916 232912
rect 185169 232854 187916 232856
rect 185169 232851 185235 232854
rect 177717 232778 177783 232781
rect 174822 232776 177783 232778
rect 174822 232720 177722 232776
rect 177778 232720 177783 232776
rect 174822 232718 177783 232720
rect 174822 232476 174882 232718
rect 177717 232715 177783 232718
rect 90764 232446 92775 232448
rect 92709 232443 92775 232446
rect 185169 232370 185235 232373
rect 185169 232368 187916 232370
rect 185169 232312 185174 232368
rect 185230 232312 187916 232368
rect 185169 232310 187916 232312
rect 185169 232307 185235 232310
rect 50757 232234 50823 232237
rect 47524 232232 50823 232234
rect 47524 232176 50762 232232
rect 50818 232176 50823 232232
rect 47524 232174 50823 232176
rect 50757 232171 50823 232174
rect 58025 231962 58091 231965
rect 93997 231962 94063 231965
rect 58025 231960 60956 231962
rect 58025 231904 58030 231960
rect 58086 231904 60956 231960
rect 58025 231902 60956 231904
rect 90764 231960 94063 231962
rect 90764 231904 94002 231960
rect 94058 231904 94063 231960
rect 90764 231902 94063 231904
rect 58025 231899 58091 231902
rect 93997 231899 94063 231902
rect 101265 231962 101331 231965
rect 103982 231962 104042 232272
rect 134845 232234 134911 232237
rect 177717 232234 177783 232237
rect 131796 232232 134911 232234
rect 131796 232176 134850 232232
rect 134906 232176 134911 232232
rect 131796 232174 134911 232176
rect 134845 232171 134911 232174
rect 174822 232232 177783 232234
rect 174822 232176 177722 232232
rect 177778 232176 177783 232232
rect 174822 232174 177783 232176
rect 101265 231960 104042 231962
rect 101265 231904 101270 231960
rect 101326 231904 104042 231960
rect 101265 231902 104042 231904
rect 142297 231962 142363 231965
rect 142297 231960 145044 231962
rect 142297 231904 142302 231960
rect 142358 231904 145044 231960
rect 174822 231932 174882 232174
rect 177717 232171 177783 232174
rect 142297 231902 145044 231904
rect 101265 231899 101331 231902
rect 142297 231899 142363 231902
rect 185261 231826 185327 231829
rect 185261 231824 187916 231826
rect 185261 231768 185266 231824
rect 185322 231768 187916 231824
rect 185261 231766 187916 231768
rect 185261 231763 185327 231766
rect 50113 231690 50179 231693
rect 47524 231688 50179 231690
rect 47524 231632 50118 231688
rect 50174 231632 50179 231688
rect 47524 231630 50179 231632
rect 50113 231627 50179 231630
rect 101449 231554 101515 231557
rect 103982 231554 104042 231728
rect 134753 231690 134819 231693
rect 131796 231688 134819 231690
rect 131796 231632 134758 231688
rect 134814 231632 134819 231688
rect 131796 231630 134819 231632
rect 134753 231627 134819 231630
rect 222337 231690 222403 231693
rect 225416 231690 225896 231720
rect 222337 231688 225896 231690
rect 222337 231632 222342 231688
rect 222398 231632 225896 231688
rect 222337 231630 225896 231632
rect 222337 231627 222403 231630
rect 225416 231600 225896 231630
rect 177717 231554 177783 231557
rect 101449 231552 104042 231554
rect 101449 231496 101454 231552
rect 101510 231496 104042 231552
rect 101449 231494 104042 231496
rect 174822 231552 177783 231554
rect 174822 231496 177722 231552
rect 177778 231496 177783 231552
rect 174822 231494 177783 231496
rect 101449 231491 101515 231494
rect 58117 231282 58183 231285
rect 92709 231282 92775 231285
rect 58117 231280 60956 231282
rect 58117 231224 58122 231280
rect 58178 231224 60956 231280
rect 58117 231222 60956 231224
rect 90764 231280 92775 231282
rect 90764 231224 92714 231280
rect 92770 231224 92775 231280
rect 90764 231222 92775 231224
rect 58117 231219 58183 231222
rect 92709 231219 92775 231222
rect 101725 231282 101791 231285
rect 142205 231282 142271 231285
rect 101725 231280 104012 231282
rect 101725 231224 101730 231280
rect 101786 231224 104012 231280
rect 101725 231222 104012 231224
rect 142205 231280 145044 231282
rect 142205 231224 142210 231280
rect 142266 231224 145044 231280
rect 174822 231252 174882 231494
rect 177717 231491 177783 231494
rect 185169 231282 185235 231285
rect 185169 231280 187916 231282
rect 142205 231222 145044 231224
rect 185169 231224 185174 231280
rect 185230 231224 187916 231280
rect 185169 231222 187916 231224
rect 101725 231219 101791 231222
rect 142205 231219 142271 231222
rect 185169 231219 185235 231222
rect 51217 231146 51283 231149
rect 134753 231146 134819 231149
rect 47524 231144 51283 231146
rect 47524 231088 51222 231144
rect 51278 231088 51283 231144
rect 47524 231086 51283 231088
rect 131796 231144 134819 231146
rect 131796 231088 134758 231144
rect 134814 231088 134819 231144
rect 131796 231086 134819 231088
rect 51217 231083 51283 231086
rect 134753 231083 134819 231086
rect 177717 230874 177783 230877
rect 174822 230872 177783 230874
rect 174822 230816 177722 230872
rect 177778 230816 177783 230872
rect 174822 230814 177783 230816
rect 58209 230738 58275 230741
rect 93721 230738 93787 230741
rect 58209 230736 60956 230738
rect 58209 230680 58214 230736
rect 58270 230680 60956 230736
rect 58209 230678 60956 230680
rect 90764 230736 93787 230738
rect 90764 230680 93726 230736
rect 93782 230680 93787 230736
rect 90764 230678 93787 230680
rect 58209 230675 58275 230678
rect 93721 230675 93787 230678
rect 143677 230738 143743 230741
rect 143677 230736 145044 230738
rect 143677 230680 143682 230736
rect 143738 230680 145044 230736
rect 174822 230708 174882 230814
rect 177717 230811 177783 230814
rect 185261 230738 185327 230741
rect 185261 230736 187916 230738
rect 143677 230678 145044 230680
rect 185261 230680 185266 230736
rect 185322 230680 187916 230736
rect 185261 230678 187916 230680
rect 143677 230675 143743 230678
rect 185261 230675 185327 230678
rect 51125 230602 51191 230605
rect 47524 230600 51191 230602
rect 47524 230544 51130 230600
rect 51186 230544 51191 230600
rect 47524 230542 51191 230544
rect 51125 230539 51191 230542
rect 58209 230194 58275 230197
rect 92709 230194 92775 230197
rect 58209 230192 60956 230194
rect 58209 230136 58214 230192
rect 58270 230136 60956 230192
rect 58209 230134 60956 230136
rect 90764 230192 92775 230194
rect 90764 230136 92714 230192
rect 92770 230136 92775 230192
rect 90764 230134 92775 230136
rect 58209 230131 58275 230134
rect 92709 230131 92775 230134
rect 101725 230194 101791 230197
rect 103982 230194 104042 230640
rect 134385 230602 134451 230605
rect 131796 230600 134451 230602
rect 131796 230544 134390 230600
rect 134446 230544 134451 230600
rect 131796 230542 134451 230544
rect 134385 230539 134451 230542
rect 177717 230466 177783 230469
rect 174822 230464 177783 230466
rect 174822 230408 177722 230464
rect 177778 230408 177783 230464
rect 174822 230406 177783 230408
rect 101725 230192 104042 230194
rect 101725 230136 101730 230192
rect 101786 230136 104042 230192
rect 101725 230134 104042 230136
rect 142941 230194 143007 230197
rect 142941 230192 145044 230194
rect 142941 230136 142946 230192
rect 143002 230136 145044 230192
rect 174822 230164 174882 230406
rect 177717 230403 177783 230406
rect 142941 230134 145044 230136
rect 101725 230131 101791 230134
rect 142941 230131 143007 230134
rect 51217 230058 51283 230061
rect 134293 230058 134359 230061
rect 47524 230056 51283 230058
rect 47524 230000 51222 230056
rect 51278 230000 51283 230056
rect 47524 229998 51283 230000
rect 131796 230056 134359 230058
rect 131796 230000 134298 230056
rect 134354 230000 134359 230056
rect 131796 229998 134359 230000
rect 51217 229995 51283 229998
rect 134293 229995 134359 229998
rect 185169 230058 185235 230061
rect 185169 230056 187916 230058
rect 185169 230000 185174 230056
rect 185230 230000 187916 230056
rect 185169 229998 187916 230000
rect 185169 229995 185235 229998
rect 101541 229786 101607 229789
rect 103982 229786 104042 229960
rect 101541 229784 104042 229786
rect 101541 229728 101546 229784
rect 101602 229728 104042 229784
rect 101541 229726 104042 229728
rect 101541 229723 101607 229726
rect 177717 229650 177783 229653
rect 174822 229648 177783 229650
rect 174822 229592 177722 229648
rect 177778 229592 177783 229648
rect 174822 229590 177783 229592
rect 58209 229514 58275 229517
rect 92709 229514 92775 229517
rect 58209 229512 60956 229514
rect 58209 229456 58214 229512
rect 58270 229456 60956 229512
rect 58209 229454 60956 229456
rect 90764 229512 92775 229514
rect 90764 229456 92714 229512
rect 92770 229456 92775 229512
rect 90764 229454 92775 229456
rect 58209 229451 58275 229454
rect 92709 229451 92775 229454
rect 143677 229514 143743 229517
rect 143677 229512 145044 229514
rect 143677 229456 143682 229512
rect 143738 229456 145044 229512
rect 174822 229484 174882 229590
rect 177717 229587 177783 229590
rect 185169 229514 185235 229517
rect 185169 229512 187916 229514
rect 143677 229454 145044 229456
rect 185169 229456 185174 229512
rect 185230 229456 187916 229512
rect 185169 229454 187916 229456
rect 143677 229451 143743 229454
rect 185169 229451 185235 229454
rect 51125 229378 51191 229381
rect 47524 229376 51191 229378
rect 47524 229320 51130 229376
rect 51186 229320 51191 229376
rect 47524 229318 51191 229320
rect 51125 229315 51191 229318
rect 101725 229242 101791 229245
rect 103982 229242 104042 229416
rect 134385 229378 134451 229381
rect 131796 229376 134451 229378
rect 131796 229320 134390 229376
rect 134446 229320 134451 229376
rect 131796 229318 134451 229320
rect 134385 229315 134451 229318
rect 177625 229242 177691 229245
rect 101725 229240 104042 229242
rect 101725 229184 101730 229240
rect 101786 229184 104042 229240
rect 101725 229182 104042 229184
rect 174822 229240 177691 229242
rect 174822 229184 177630 229240
rect 177686 229184 177691 229240
rect 174822 229182 177691 229184
rect 101725 229179 101791 229182
rect 58209 228970 58275 228973
rect 92801 228970 92867 228973
rect 58209 228968 60956 228970
rect 58209 228912 58214 228968
rect 58270 228912 60956 228968
rect 58209 228910 60956 228912
rect 90764 228968 92867 228970
rect 90764 228912 92806 228968
rect 92862 228912 92867 228968
rect 90764 228910 92867 228912
rect 58209 228907 58275 228910
rect 92801 228907 92867 228910
rect 143585 228970 143651 228973
rect 143585 228968 145044 228970
rect 143585 228912 143590 228968
rect 143646 228912 145044 228968
rect 174822 228940 174882 229182
rect 177625 229179 177691 229182
rect 185261 228970 185327 228973
rect 185261 228968 187916 228970
rect 143585 228910 145044 228912
rect 185261 228912 185266 228968
rect 185322 228912 187916 228968
rect 185261 228910 187916 228912
rect 143585 228907 143651 228910
rect 185261 228907 185327 228910
rect 51217 228834 51283 228837
rect 47524 228832 51283 228834
rect 47524 228776 51222 228832
rect 51278 228776 51283 228832
rect 47524 228774 51283 228776
rect 51217 228771 51283 228774
rect 101449 228698 101515 228701
rect 103982 228698 104042 228872
rect 134753 228834 134819 228837
rect 131796 228832 134819 228834
rect 131796 228776 134758 228832
rect 134814 228776 134819 228832
rect 131796 228774 134819 228776
rect 134753 228771 134819 228774
rect 101449 228696 104042 228698
rect 101449 228640 101454 228696
rect 101510 228640 104042 228696
rect 101449 228638 104042 228640
rect 101449 228635 101515 228638
rect 176981 228562 177047 228565
rect 174822 228560 177047 228562
rect 174822 228504 176986 228560
rect 177042 228504 177047 228560
rect 174822 228502 177047 228504
rect 101725 228426 101791 228429
rect 101725 228424 104012 228426
rect 101725 228368 101730 228424
rect 101786 228368 104012 228424
rect 101725 228366 104012 228368
rect 101725 228363 101791 228366
rect 51033 228290 51099 228293
rect 47524 228288 51099 228290
rect 47524 228232 51038 228288
rect 51094 228232 51099 228288
rect 47524 228230 51099 228232
rect 51033 228227 51099 228230
rect 58301 228290 58367 228293
rect 92709 228290 92775 228293
rect 134845 228290 134911 228293
rect 58301 228288 60956 228290
rect 58301 228232 58306 228288
rect 58362 228232 60956 228288
rect 58301 228230 60956 228232
rect 90764 228288 92775 228290
rect 90764 228232 92714 228288
rect 92770 228232 92775 228288
rect 90764 228230 92775 228232
rect 131796 228288 134911 228290
rect 131796 228232 134850 228288
rect 134906 228232 134911 228288
rect 131796 228230 134911 228232
rect 58301 228227 58367 228230
rect 92709 228227 92775 228230
rect 134845 228227 134911 228230
rect 143493 228290 143559 228293
rect 143493 228288 145044 228290
rect 143493 228232 143498 228288
rect 143554 228232 145044 228288
rect 174822 228260 174882 228502
rect 176981 228499 177047 228502
rect 185169 228426 185235 228429
rect 185169 228424 187916 228426
rect 185169 228368 185174 228424
rect 185230 228368 187916 228424
rect 185169 228366 187916 228368
rect 185169 228363 185235 228366
rect 143493 228230 145044 228232
rect 143493 228227 143559 228230
rect 177717 228018 177783 228021
rect 174822 228016 177783 228018
rect 174822 227960 177722 228016
rect 177778 227960 177783 228016
rect 174822 227958 177783 227960
rect 50757 227746 50823 227749
rect 47524 227744 50823 227746
rect 47524 227688 50762 227744
rect 50818 227688 50823 227744
rect 47524 227686 50823 227688
rect 50757 227683 50823 227686
rect 58209 227746 58275 227749
rect 93169 227746 93235 227749
rect 58209 227744 60956 227746
rect 58209 227688 58214 227744
rect 58270 227688 60956 227744
rect 58209 227686 60956 227688
rect 90764 227744 93235 227746
rect 90764 227688 93174 227744
rect 93230 227688 93235 227744
rect 90764 227686 93235 227688
rect 58209 227683 58275 227686
rect 93169 227683 93235 227686
rect 101357 227474 101423 227477
rect 103982 227474 104042 227784
rect 134753 227746 134819 227749
rect 131796 227744 134819 227746
rect 131796 227688 134758 227744
rect 134814 227688 134819 227744
rect 131796 227686 134819 227688
rect 134753 227683 134819 227686
rect 143677 227746 143743 227749
rect 143677 227744 145044 227746
rect 143677 227688 143682 227744
rect 143738 227688 145044 227744
rect 174822 227716 174882 227958
rect 177717 227955 177783 227958
rect 185169 227882 185235 227885
rect 185169 227880 187916 227882
rect 185169 227824 185174 227880
rect 185230 227824 187916 227880
rect 185169 227822 187916 227824
rect 185169 227819 185235 227822
rect 143677 227686 145044 227688
rect 143677 227683 143743 227686
rect 177625 227474 177691 227477
rect 101357 227472 104042 227474
rect 101357 227416 101362 227472
rect 101418 227416 104042 227472
rect 101357 227414 104042 227416
rect 174822 227472 177691 227474
rect 174822 227416 177630 227472
rect 177686 227416 177691 227472
rect 174822 227414 177691 227416
rect 101357 227411 101423 227414
rect 51217 227202 51283 227205
rect 47524 227200 51283 227202
rect 47524 227144 51222 227200
rect 51278 227144 51283 227200
rect 47524 227142 51283 227144
rect 51217 227139 51283 227142
rect 58301 227202 58367 227205
rect 92709 227202 92775 227205
rect 58301 227200 60956 227202
rect 58301 227144 58306 227200
rect 58362 227144 60956 227200
rect 58301 227142 60956 227144
rect 90764 227200 92775 227202
rect 90764 227144 92714 227200
rect 92770 227144 92775 227200
rect 90764 227142 92775 227144
rect 58301 227139 58367 227142
rect 92709 227139 92775 227142
rect 101449 227066 101515 227069
rect 103982 227066 104042 227240
rect 135397 227202 135463 227205
rect 131796 227200 135463 227202
rect 131796 227144 135402 227200
rect 135458 227144 135463 227200
rect 131796 227142 135463 227144
rect 135397 227139 135463 227142
rect 143309 227202 143375 227205
rect 143309 227200 145044 227202
rect 143309 227144 143314 227200
rect 143370 227144 145044 227200
rect 174822 227172 174882 227414
rect 177625 227411 177691 227414
rect 185261 227338 185327 227341
rect 185261 227336 187916 227338
rect 185261 227280 185266 227336
rect 185322 227280 187916 227336
rect 185261 227278 187916 227280
rect 185261 227275 185327 227278
rect 143309 227142 145044 227144
rect 143309 227139 143375 227142
rect 101449 227064 104042 227066
rect 101449 227008 101454 227064
rect 101510 227008 104042 227064
rect 101449 227006 104042 227008
rect 101449 227003 101515 227006
rect 185353 226794 185419 226797
rect 185353 226792 187916 226794
rect 185353 226736 185358 226792
rect 185414 226736 187916 226792
rect 185353 226734 187916 226736
rect 185353 226731 185419 226734
rect 51217 226522 51283 226525
rect 47524 226520 51283 226522
rect 47524 226464 51222 226520
rect 51278 226464 51283 226520
rect 47524 226462 51283 226464
rect 51217 226459 51283 226462
rect 58209 226522 58275 226525
rect 92709 226522 92775 226525
rect 58209 226520 60956 226522
rect 58209 226464 58214 226520
rect 58270 226464 60956 226520
rect 58209 226462 60956 226464
rect 90764 226520 92775 226522
rect 90764 226464 92714 226520
rect 92770 226464 92775 226520
rect 90764 226462 92775 226464
rect 58209 226459 58275 226462
rect 92709 226459 92775 226462
rect 101633 226386 101699 226389
rect 103982 226386 104042 226696
rect 177165 226658 177231 226661
rect 174822 226656 177231 226658
rect 174822 226600 177170 226656
rect 177226 226600 177231 226656
rect 174822 226598 177231 226600
rect 134385 226522 134451 226525
rect 131796 226520 134451 226522
rect 131796 226464 134390 226520
rect 134446 226464 134451 226520
rect 131796 226462 134451 226464
rect 134385 226459 134451 226462
rect 143677 226522 143743 226525
rect 143677 226520 145044 226522
rect 143677 226464 143682 226520
rect 143738 226464 145044 226520
rect 174822 226492 174882 226598
rect 177165 226595 177231 226598
rect 143677 226462 145044 226464
rect 143677 226459 143743 226462
rect 101633 226384 104042 226386
rect 101633 226328 101638 226384
rect 101694 226328 104042 226384
rect 101633 226326 104042 226328
rect 101633 226323 101699 226326
rect 177717 226250 177783 226253
rect 174822 226248 177783 226250
rect 174822 226192 177722 226248
rect 177778 226192 177783 226248
rect 174822 226190 177783 226192
rect 50021 225978 50087 225981
rect 47524 225976 50087 225978
rect 47524 225920 50026 225976
rect 50082 225920 50087 225976
rect 47524 225918 50087 225920
rect 50021 225915 50087 225918
rect 58209 225978 58275 225981
rect 92801 225978 92867 225981
rect 58209 225976 60956 225978
rect 58209 225920 58214 225976
rect 58270 225920 60956 225976
rect 58209 225918 60956 225920
rect 90764 225976 92867 225978
rect 90764 225920 92806 225976
rect 92862 225920 92867 225976
rect 90764 225918 92867 225920
rect 58209 225915 58275 225918
rect 92801 225915 92867 225918
rect 101817 225706 101883 225709
rect 103982 225706 104042 226152
rect 134753 225978 134819 225981
rect 131796 225976 134819 225978
rect 131796 225920 134758 225976
rect 134814 225920 134819 225976
rect 131796 225918 134819 225920
rect 134753 225915 134819 225918
rect 143309 225978 143375 225981
rect 143309 225976 145044 225978
rect 143309 225920 143314 225976
rect 143370 225920 145044 225976
rect 174822 225948 174882 226190
rect 177717 226187 177783 226190
rect 185261 226250 185327 226253
rect 185261 226248 187916 226250
rect 185261 226192 185266 226248
rect 185322 226192 187916 226248
rect 185261 226190 187916 226192
rect 185261 226187 185327 226190
rect 143309 225918 145044 225920
rect 143309 225915 143375 225918
rect 101817 225704 104042 225706
rect 101817 225648 101822 225704
rect 101878 225648 104042 225704
rect 101817 225646 104042 225648
rect 101817 225643 101883 225646
rect 101541 225570 101607 225573
rect 185169 225570 185235 225573
rect 101541 225568 104012 225570
rect 101541 225512 101546 225568
rect 101602 225512 104012 225568
rect 101541 225510 104012 225512
rect 185169 225568 187916 225570
rect 185169 225512 185174 225568
rect 185230 225512 187916 225568
rect 185169 225510 187916 225512
rect 101541 225507 101607 225510
rect 185169 225507 185235 225510
rect 51125 225434 51191 225437
rect 134661 225434 134727 225437
rect 177717 225434 177783 225437
rect 47524 225432 51191 225434
rect 47524 225376 51130 225432
rect 51186 225376 51191 225432
rect 47524 225374 51191 225376
rect 131796 225432 134727 225434
rect 131796 225376 134666 225432
rect 134722 225376 134727 225432
rect 131796 225374 134727 225376
rect 51125 225371 51191 225374
rect 134661 225371 134727 225374
rect 174822 225432 177783 225434
rect 174822 225376 177722 225432
rect 177778 225376 177783 225432
rect 174822 225374 177783 225376
rect 58209 225298 58275 225301
rect 92709 225298 92775 225301
rect 58209 225296 60956 225298
rect 58209 225240 58214 225296
rect 58270 225240 60956 225296
rect 58209 225238 60956 225240
rect 90764 225296 92775 225298
rect 90764 225240 92714 225296
rect 92770 225240 92775 225296
rect 90764 225238 92775 225240
rect 58209 225235 58275 225238
rect 92709 225235 92775 225238
rect 143677 225298 143743 225301
rect 143677 225296 145044 225298
rect 143677 225240 143682 225296
rect 143738 225240 145044 225296
rect 174822 225268 174882 225374
rect 177717 225371 177783 225374
rect 143677 225238 145044 225240
rect 143677 225235 143743 225238
rect 177717 225026 177783 225029
rect 174822 225024 177783 225026
rect 174822 224968 177722 225024
rect 177778 224968 177783 225024
rect 174822 224966 177783 224968
rect 51217 224890 51283 224893
rect 47524 224888 51283 224890
rect 47524 224832 51222 224888
rect 51278 224832 51283 224888
rect 47524 224830 51283 224832
rect 51217 224827 51283 224830
rect 58301 224754 58367 224757
rect 92801 224754 92867 224757
rect 58301 224752 60956 224754
rect 58301 224696 58306 224752
rect 58362 224696 60956 224752
rect 58301 224694 60956 224696
rect 90764 224752 92867 224754
rect 90764 224696 92806 224752
rect 92862 224696 92867 224752
rect 90764 224694 92867 224696
rect 58301 224691 58367 224694
rect 92801 224691 92867 224694
rect 101081 224618 101147 224621
rect 103982 224618 104042 224928
rect 134293 224890 134359 224893
rect 131796 224888 134359 224890
rect 131796 224832 134298 224888
rect 134354 224832 134359 224888
rect 131796 224830 134359 224832
rect 134293 224827 134359 224830
rect 143309 224754 143375 224757
rect 143309 224752 145044 224754
rect 143309 224696 143314 224752
rect 143370 224696 145044 224752
rect 174822 224724 174882 224966
rect 177717 224963 177783 224966
rect 185261 225026 185327 225029
rect 185261 225024 187916 225026
rect 185261 224968 185266 225024
rect 185322 224968 187916 225024
rect 185261 224966 187916 224968
rect 185261 224963 185327 224966
rect 143309 224694 145044 224696
rect 143309 224691 143375 224694
rect 101081 224616 104042 224618
rect 101081 224560 101086 224616
rect 101142 224560 104042 224616
rect 101081 224558 104042 224560
rect 101081 224555 101147 224558
rect 100989 224482 101055 224485
rect 177165 224482 177231 224485
rect 100989 224480 104012 224482
rect 100989 224424 100994 224480
rect 101050 224424 104012 224480
rect 100989 224422 104012 224424
rect 174822 224480 177231 224482
rect 174822 224424 177170 224480
rect 177226 224424 177231 224480
rect 174822 224422 177231 224424
rect 100989 224419 101055 224422
rect 51125 224346 51191 224349
rect 135397 224346 135463 224349
rect 47524 224344 51191 224346
rect 47524 224288 51130 224344
rect 51186 224288 51191 224344
rect 47524 224286 51191 224288
rect 131796 224344 135463 224346
rect 131796 224288 135402 224344
rect 135458 224288 135463 224344
rect 131796 224286 135463 224288
rect 51125 224283 51191 224286
rect 135397 224283 135463 224286
rect 58393 224210 58459 224213
rect 93721 224210 93787 224213
rect 58393 224208 60956 224210
rect 58393 224152 58398 224208
rect 58454 224152 60956 224208
rect 58393 224150 60956 224152
rect 90764 224208 93787 224210
rect 90764 224152 93726 224208
rect 93782 224152 93787 224208
rect 90764 224150 93787 224152
rect 58393 224147 58459 224150
rect 93721 224147 93787 224150
rect 142573 224210 142639 224213
rect 142573 224208 145044 224210
rect 142573 224152 142578 224208
rect 142634 224152 145044 224208
rect 174822 224180 174882 224422
rect 177165 224419 177231 224422
rect 185169 224482 185235 224485
rect 185169 224480 187916 224482
rect 185169 224424 185174 224480
rect 185230 224424 187916 224480
rect 185169 224422 187916 224424
rect 185169 224419 185235 224422
rect 142573 224150 145044 224152
rect 142573 224147 142639 224150
rect 185261 223938 185327 223941
rect 185261 223936 187916 223938
rect 185261 223880 185266 223936
rect 185322 223880 187916 223936
rect 185261 223878 187916 223880
rect 185261 223875 185327 223878
rect 51217 223666 51283 223669
rect 47524 223664 51283 223666
rect 47524 223608 51222 223664
rect 51278 223608 51283 223664
rect 47524 223606 51283 223608
rect 51217 223603 51283 223606
rect 58301 223530 58367 223533
rect 93721 223530 93787 223533
rect 58301 223528 60956 223530
rect 58301 223472 58306 223528
rect 58362 223472 60956 223528
rect 58301 223470 60956 223472
rect 90764 223528 93787 223530
rect 90764 223472 93726 223528
rect 93782 223472 93787 223528
rect 90764 223470 93787 223472
rect 58301 223467 58367 223470
rect 93721 223467 93787 223470
rect 101449 223530 101515 223533
rect 103982 223530 104042 223840
rect 177717 223802 177783 223805
rect 174822 223800 177783 223802
rect 174822 223744 177722 223800
rect 177778 223744 177783 223800
rect 174822 223742 177783 223744
rect 135397 223666 135463 223669
rect 131796 223664 135463 223666
rect 131796 223608 135402 223664
rect 135458 223608 135463 223664
rect 131796 223606 135463 223608
rect 135397 223603 135463 223606
rect 101449 223528 104042 223530
rect 101449 223472 101454 223528
rect 101510 223472 104042 223528
rect 101449 223470 104042 223472
rect 143677 223530 143743 223533
rect 143677 223528 145044 223530
rect 143677 223472 143682 223528
rect 143738 223472 145044 223528
rect 174822 223500 174882 223742
rect 177717 223739 177783 223742
rect 143677 223470 145044 223472
rect 101449 223467 101515 223470
rect 143677 223467 143743 223470
rect 185169 223394 185235 223397
rect 185169 223392 187916 223394
rect 185169 223336 185174 223392
rect 185230 223336 187916 223392
rect 185169 223334 187916 223336
rect 185169 223331 185235 223334
rect 51125 223122 51191 223125
rect 47524 223120 51191 223122
rect 47524 223064 51130 223120
rect 51186 223064 51191 223120
rect 47524 223062 51191 223064
rect 51125 223059 51191 223062
rect 58209 222986 58275 222989
rect 93905 222986 93971 222989
rect 58209 222984 60956 222986
rect 58209 222928 58214 222984
rect 58270 222928 60956 222984
rect 58209 222926 60956 222928
rect 90764 222984 93971 222986
rect 90764 222928 93910 222984
rect 93966 222928 93971 222984
rect 90764 222926 93971 222928
rect 58209 222923 58275 222926
rect 93905 222923 93971 222926
rect 101357 222986 101423 222989
rect 103982 222986 104042 223296
rect 177625 223258 177691 223261
rect 174822 223256 177691 223258
rect 174822 223200 177630 223256
rect 177686 223200 177691 223256
rect 174822 223198 177691 223200
rect 134477 223122 134543 223125
rect 131796 223120 134543 223122
rect 131796 223064 134482 223120
rect 134538 223064 134543 223120
rect 131796 223062 134543 223064
rect 134477 223059 134543 223062
rect 101357 222984 104042 222986
rect 101357 222928 101362 222984
rect 101418 222928 104042 222984
rect 101357 222926 104042 222928
rect 143309 222986 143375 222989
rect 143309 222984 145044 222986
rect 143309 222928 143314 222984
rect 143370 222928 145044 222984
rect 174822 222956 174882 223198
rect 177625 223195 177691 223198
rect 143309 222926 145044 222928
rect 101357 222923 101423 222926
rect 143309 222923 143375 222926
rect 100897 222850 100963 222853
rect 185077 222850 185143 222853
rect 100897 222848 104012 222850
rect 100897 222792 100902 222848
rect 100958 222792 104012 222848
rect 100897 222790 104012 222792
rect 185077 222848 187916 222850
rect 185077 222792 185082 222848
rect 185138 222792 187916 222848
rect 185077 222790 187916 222792
rect 100897 222787 100963 222790
rect 185077 222787 185143 222790
rect 51217 222578 51283 222581
rect 134845 222578 134911 222581
rect 47524 222576 51283 222578
rect 47524 222520 51222 222576
rect 51278 222520 51283 222576
rect 47524 222518 51283 222520
rect 131796 222576 134911 222578
rect 131796 222520 134850 222576
rect 134906 222520 134911 222576
rect 131796 222518 134911 222520
rect 51217 222515 51283 222518
rect 134845 222515 134911 222518
rect 177717 222442 177783 222445
rect 174822 222440 177783 222442
rect 174822 222384 177722 222440
rect 177778 222384 177783 222440
rect 174822 222382 177783 222384
rect 58209 222306 58275 222309
rect 92709 222306 92775 222309
rect 58209 222304 60956 222306
rect 58209 222248 58214 222304
rect 58270 222248 60956 222304
rect 58209 222246 60956 222248
rect 90764 222304 92775 222306
rect 90764 222248 92714 222304
rect 92770 222248 92775 222304
rect 90764 222246 92775 222248
rect 58209 222243 58275 222246
rect 92709 222243 92775 222246
rect 143677 222306 143743 222309
rect 143677 222304 145044 222306
rect 143677 222248 143682 222304
rect 143738 222248 145044 222304
rect 174822 222276 174882 222382
rect 177717 222379 177783 222382
rect 185261 222306 185327 222309
rect 185261 222304 187916 222306
rect 143677 222246 145044 222248
rect 185261 222248 185266 222304
rect 185322 222248 187916 222304
rect 185261 222246 187916 222248
rect 143677 222243 143743 222246
rect 185261 222243 185327 222246
rect 51125 222034 51191 222037
rect 47524 222032 51191 222034
rect 47524 221976 51130 222032
rect 51186 221976 51191 222032
rect 47524 221974 51191 221976
rect 51125 221971 51191 221974
rect 101633 221898 101699 221901
rect 103982 221898 104042 222208
rect 134661 222034 134727 222037
rect 177625 222034 177691 222037
rect 131796 222032 134727 222034
rect 131796 221976 134666 222032
rect 134722 221976 134727 222032
rect 131796 221974 134727 221976
rect 134661 221971 134727 221974
rect 174822 222032 177691 222034
rect 174822 221976 177630 222032
rect 177686 221976 177691 222032
rect 174822 221974 177691 221976
rect 101633 221896 104042 221898
rect 101633 221840 101638 221896
rect 101694 221840 104042 221896
rect 101633 221838 104042 221840
rect 101633 221835 101699 221838
rect 58301 221762 58367 221765
rect 92985 221762 93051 221765
rect 58301 221760 60956 221762
rect 58301 221704 58306 221760
rect 58362 221704 60956 221760
rect 58301 221702 60956 221704
rect 90764 221760 93051 221762
rect 90764 221704 92990 221760
rect 93046 221704 93051 221760
rect 90764 221702 93051 221704
rect 58301 221699 58367 221702
rect 92985 221699 93051 221702
rect 143309 221762 143375 221765
rect 143309 221760 145044 221762
rect 143309 221704 143314 221760
rect 143370 221704 145044 221760
rect 174822 221732 174882 221974
rect 177625 221971 177691 221974
rect 185169 221762 185235 221765
rect 185169 221760 187916 221762
rect 143309 221702 145044 221704
rect 185169 221704 185174 221760
rect 185230 221704 187916 221760
rect 185169 221702 187916 221704
rect 143309 221699 143375 221702
rect 185169 221699 185235 221702
rect 51217 221490 51283 221493
rect 47524 221488 51283 221490
rect 47524 221432 51222 221488
rect 51278 221432 51283 221488
rect 47524 221430 51283 221432
rect 51217 221427 51283 221430
rect 101541 221490 101607 221493
rect 103982 221490 104042 221664
rect 135397 221490 135463 221493
rect 101541 221488 104042 221490
rect 101541 221432 101546 221488
rect 101602 221432 104042 221488
rect 101541 221430 104042 221432
rect 131796 221488 135463 221490
rect 131796 221432 135402 221488
rect 135458 221432 135463 221488
rect 131796 221430 135463 221432
rect 101541 221427 101607 221430
rect 135397 221427 135463 221430
rect 58209 221218 58275 221221
rect 92709 221218 92775 221221
rect 58209 221216 60956 221218
rect 58209 221160 58214 221216
rect 58270 221160 60956 221216
rect 58209 221158 60956 221160
rect 90764 221216 92775 221218
rect 90764 221160 92714 221216
rect 92770 221160 92775 221216
rect 90764 221158 92775 221160
rect 58209 221155 58275 221158
rect 92709 221155 92775 221158
rect 143677 221218 143743 221221
rect 185353 221218 185419 221221
rect 215713 221218 215779 221221
rect 143677 221216 145044 221218
rect 143677 221160 143682 221216
rect 143738 221160 145044 221216
rect 185353 221216 187916 221218
rect 143677 221158 145044 221160
rect 143677 221155 143743 221158
rect 51217 220810 51283 220813
rect 47524 220808 51283 220810
rect 47524 220752 51222 220808
rect 51278 220752 51283 220808
rect 47524 220750 51283 220752
rect 51217 220747 51283 220750
rect 101817 220674 101883 220677
rect 103982 220674 104042 221120
rect 174822 221082 174882 221188
rect 185353 221160 185358 221216
rect 185414 221160 187916 221216
rect 185353 221158 187916 221160
rect 215670 221216 215779 221218
rect 215670 221160 215718 221216
rect 215774 221160 215779 221216
rect 185353 221155 185419 221158
rect 215670 221155 215779 221160
rect 177717 221082 177783 221085
rect 174822 221080 177783 221082
rect 174822 221024 177722 221080
rect 177778 221024 177783 221080
rect 174822 221022 177783 221024
rect 177717 221019 177783 221022
rect 177625 220946 177691 220949
rect 174822 220944 177691 220946
rect 174822 220888 177630 220944
rect 177686 220888 177691 220944
rect 174822 220886 177691 220888
rect 135397 220810 135463 220813
rect 131796 220808 135463 220810
rect 131796 220752 135402 220808
rect 135458 220752 135463 220808
rect 131796 220750 135463 220752
rect 135397 220747 135463 220750
rect 101817 220672 104042 220674
rect 101817 220616 101822 220672
rect 101878 220616 104042 220672
rect 101817 220614 104042 220616
rect 101817 220611 101883 220614
rect 58209 220538 58275 220541
rect 93721 220538 93787 220541
rect 58209 220536 60956 220538
rect 58209 220480 58214 220536
rect 58270 220480 60956 220536
rect 58209 220478 60956 220480
rect 90764 220536 93787 220538
rect 90764 220480 93726 220536
rect 93782 220480 93787 220536
rect 90764 220478 93787 220480
rect 58209 220475 58275 220478
rect 93721 220475 93787 220478
rect 143309 220538 143375 220541
rect 143309 220536 145044 220538
rect 143309 220480 143314 220536
rect 143370 220480 145044 220536
rect 174822 220508 174882 220886
rect 177625 220883 177691 220886
rect 215670 220780 215730 221155
rect 185169 220538 185235 220541
rect 185169 220536 187916 220538
rect 143309 220478 145044 220480
rect 185169 220480 185174 220536
rect 185230 220480 187916 220536
rect 185169 220478 187916 220480
rect 143309 220475 143375 220478
rect 185169 220475 185235 220478
rect 51125 220266 51191 220269
rect 47524 220264 51191 220266
rect 47524 220208 51130 220264
rect 51186 220208 51191 220264
rect 47524 220206 51191 220208
rect 51125 220203 51191 220206
rect 101265 220130 101331 220133
rect 103982 220130 104042 220440
rect 135305 220266 135371 220269
rect 177165 220266 177231 220269
rect 131796 220264 135371 220266
rect 131796 220208 135310 220264
rect 135366 220208 135371 220264
rect 131796 220206 135371 220208
rect 135305 220203 135371 220206
rect 174822 220264 177231 220266
rect 174822 220208 177170 220264
rect 177226 220208 177231 220264
rect 174822 220206 177231 220208
rect 101265 220128 104042 220130
rect 101265 220072 101270 220128
rect 101326 220072 104042 220128
rect 101265 220070 104042 220072
rect 101265 220067 101331 220070
rect 58301 219994 58367 219997
rect 92801 219994 92867 219997
rect 58301 219992 60956 219994
rect 58301 219936 58306 219992
rect 58362 219936 60956 219992
rect 58301 219934 60956 219936
rect 90764 219992 92867 219994
rect 90764 219936 92806 219992
rect 92862 219936 92867 219992
rect 90764 219934 92867 219936
rect 58301 219931 58367 219934
rect 92801 219931 92867 219934
rect 100897 219994 100963 219997
rect 143677 219994 143743 219997
rect 100897 219992 104012 219994
rect 100897 219936 100902 219992
rect 100958 219936 104012 219992
rect 100897 219934 104012 219936
rect 143677 219992 145044 219994
rect 143677 219936 143682 219992
rect 143738 219936 145044 219992
rect 174822 219964 174882 220206
rect 177165 220203 177231 220206
rect 185077 219994 185143 219997
rect 185077 219992 187916 219994
rect 143677 219934 145044 219936
rect 185077 219936 185082 219992
rect 185138 219936 187916 219992
rect 185077 219934 187916 219936
rect 100897 219931 100963 219934
rect 143677 219931 143743 219934
rect 185077 219931 185143 219934
rect 50849 219722 50915 219725
rect 135397 219722 135463 219725
rect 47524 219720 50915 219722
rect 47524 219664 50854 219720
rect 50910 219664 50915 219720
rect 47524 219662 50915 219664
rect 131796 219720 135463 219722
rect 131796 219664 135402 219720
rect 135458 219664 135463 219720
rect 131796 219662 135463 219664
rect 50849 219659 50915 219662
rect 135397 219659 135463 219662
rect 177717 219586 177783 219589
rect 174822 219584 177783 219586
rect 174822 219528 177722 219584
rect 177778 219528 177783 219584
rect 174822 219526 177783 219528
rect 58209 219314 58275 219317
rect 93721 219314 93787 219317
rect 58209 219312 60956 219314
rect 58209 219256 58214 219312
rect 58270 219256 60956 219312
rect 58209 219254 60956 219256
rect 90764 219312 93787 219314
rect 90764 219256 93726 219312
rect 93782 219256 93787 219312
rect 90764 219254 93787 219256
rect 58209 219251 58275 219254
rect 93721 219251 93787 219254
rect 51217 219178 51283 219181
rect 47524 219176 51283 219178
rect 47524 219120 51222 219176
rect 51278 219120 51283 219176
rect 47524 219118 51283 219120
rect 51217 219115 51283 219118
rect 101357 219042 101423 219045
rect 103982 219042 104042 219352
rect 143677 219314 143743 219317
rect 143677 219312 145044 219314
rect 143677 219256 143682 219312
rect 143738 219256 145044 219312
rect 174822 219284 174882 219526
rect 177717 219523 177783 219526
rect 185813 219450 185879 219453
rect 185813 219448 187916 219450
rect 185813 219392 185818 219448
rect 185874 219392 187916 219448
rect 185813 219390 187916 219392
rect 185813 219387 185879 219390
rect 143677 219254 145044 219256
rect 143677 219251 143743 219254
rect 135029 219178 135095 219181
rect 131796 219176 135095 219178
rect 131796 219120 135034 219176
rect 135090 219120 135095 219176
rect 131796 219118 135095 219120
rect 135029 219115 135095 219118
rect 177165 219042 177231 219045
rect 101357 219040 104042 219042
rect 101357 218984 101362 219040
rect 101418 218984 104042 219040
rect 101357 218982 104042 218984
rect 174822 219040 177231 219042
rect 174822 218984 177170 219040
rect 177226 218984 177231 219040
rect 174822 218982 177231 218984
rect 101357 218979 101423 218982
rect 101725 218906 101791 218909
rect 101725 218904 104012 218906
rect 101725 218848 101730 218904
rect 101786 218848 104012 218904
rect 101725 218846 104012 218848
rect 101725 218843 101791 218846
rect 58301 218770 58367 218773
rect 93905 218770 93971 218773
rect 58301 218768 60956 218770
rect 58301 218712 58306 218768
rect 58362 218712 60956 218768
rect 58301 218710 60956 218712
rect 90764 218768 93971 218770
rect 90764 218712 93910 218768
rect 93966 218712 93971 218768
rect 90764 218710 93971 218712
rect 58301 218707 58367 218710
rect 93905 218707 93971 218710
rect 143125 218770 143191 218773
rect 143125 218768 145044 218770
rect 143125 218712 143130 218768
rect 143186 218712 145044 218768
rect 174822 218740 174882 218982
rect 177165 218979 177231 218982
rect 185169 218906 185235 218909
rect 185169 218904 187916 218906
rect 185169 218848 185174 218904
rect 185230 218848 187916 218904
rect 185169 218846 187916 218848
rect 185169 218843 185235 218846
rect 143125 218710 145044 218712
rect 143125 218707 143191 218710
rect 51217 218634 51283 218637
rect 135305 218634 135371 218637
rect 47524 218632 51283 218634
rect 47524 218576 51222 218632
rect 51278 218576 51283 218632
rect 47524 218574 51283 218576
rect 131796 218632 135371 218634
rect 131796 218576 135310 218632
rect 135366 218576 135371 218632
rect 131796 218574 135371 218576
rect 51217 218571 51283 218574
rect 135305 218571 135371 218574
rect 177717 218362 177783 218365
rect 174822 218360 177783 218362
rect 174822 218304 177722 218360
rect 177778 218304 177783 218360
rect 174822 218302 177783 218304
rect 58209 218226 58275 218229
rect 93169 218226 93235 218229
rect 58209 218224 60956 218226
rect 58209 218168 58214 218224
rect 58270 218168 60956 218224
rect 58209 218166 60956 218168
rect 90764 218224 93235 218226
rect 90764 218168 93174 218224
rect 93230 218168 93235 218224
rect 90764 218166 93235 218168
rect 58209 218163 58275 218166
rect 93169 218163 93235 218166
rect 50757 217954 50823 217957
rect 47524 217952 50823 217954
rect 47524 217896 50762 217952
rect 50818 217896 50823 217952
rect 47524 217894 50823 217896
rect 50757 217891 50823 217894
rect 101173 217954 101239 217957
rect 103982 217954 104042 218264
rect 143677 218226 143743 218229
rect 143677 218224 145044 218226
rect 143677 218168 143682 218224
rect 143738 218168 145044 218224
rect 174822 218196 174882 218302
rect 177717 218299 177783 218302
rect 185169 218362 185235 218365
rect 185169 218360 187916 218362
rect 185169 218304 185174 218360
rect 185230 218304 187916 218360
rect 185169 218302 187916 218304
rect 185169 218299 185235 218302
rect 143677 218166 145044 218168
rect 143677 218163 143743 218166
rect 135397 217954 135463 217957
rect 177165 217954 177231 217957
rect 101173 217952 104042 217954
rect 101173 217896 101178 217952
rect 101234 217896 104042 217952
rect 101173 217894 104042 217896
rect 131796 217952 135463 217954
rect 131796 217896 135402 217952
rect 135458 217896 135463 217952
rect 131796 217894 135463 217896
rect 101173 217891 101239 217894
rect 135397 217891 135463 217894
rect 174822 217952 177231 217954
rect 174822 217896 177170 217952
rect 177226 217896 177231 217952
rect 174822 217894 177231 217896
rect 58209 217546 58275 217549
rect 93721 217546 93787 217549
rect 58209 217544 60956 217546
rect 58209 217488 58214 217544
rect 58270 217488 60956 217544
rect 58209 217486 60956 217488
rect 90764 217544 93787 217546
rect 90764 217488 93726 217544
rect 93782 217488 93787 217544
rect 90764 217486 93787 217488
rect 58209 217483 58275 217486
rect 93721 217483 93787 217486
rect 51217 217410 51283 217413
rect 47524 217408 51283 217410
rect 47524 217352 51222 217408
rect 51278 217352 51283 217408
rect 47524 217350 51283 217352
rect 51217 217347 51283 217350
rect 100805 217410 100871 217413
rect 103982 217410 104042 217720
rect 143493 217546 143559 217549
rect 143493 217544 145044 217546
rect 143493 217488 143498 217544
rect 143554 217488 145044 217544
rect 174822 217516 174882 217894
rect 177165 217891 177231 217894
rect 184985 217818 185051 217821
rect 184985 217816 187916 217818
rect 184985 217760 184990 217816
rect 185046 217760 187916 217816
rect 184985 217758 187916 217760
rect 184985 217755 185051 217758
rect 143493 217486 145044 217488
rect 143493 217483 143559 217486
rect 134477 217410 134543 217413
rect 100805 217408 104042 217410
rect 100805 217352 100810 217408
rect 100866 217352 104042 217408
rect 100805 217350 104042 217352
rect 131796 217408 134543 217410
rect 131796 217352 134482 217408
rect 134538 217352 134543 217408
rect 131796 217350 134543 217352
rect 100805 217347 100871 217350
rect 134477 217347 134543 217350
rect 100897 217274 100963 217277
rect 185077 217274 185143 217277
rect 100897 217272 104012 217274
rect 100897 217216 100902 217272
rect 100958 217216 104012 217272
rect 100897 217214 104012 217216
rect 185077 217272 187916 217274
rect 185077 217216 185082 217272
rect 185138 217216 187916 217272
rect 185077 217214 187916 217216
rect 100897 217211 100963 217214
rect 185077 217211 185143 217214
rect 177993 217138 178059 217141
rect 174822 217136 178059 217138
rect 174822 217080 177998 217136
rect 178054 217080 178059 217136
rect 174822 217078 178059 217080
rect 58209 217002 58275 217005
rect 93537 217002 93603 217005
rect 58209 217000 60956 217002
rect 58209 216944 58214 217000
rect 58270 216944 60956 217000
rect 58209 216942 60956 216944
rect 90764 217000 93603 217002
rect 90764 216944 93542 217000
rect 93598 216944 93603 217000
rect 90764 216942 93603 216944
rect 58209 216939 58275 216942
rect 93537 216939 93603 216942
rect 143677 217002 143743 217005
rect 143677 217000 145044 217002
rect 143677 216944 143682 217000
rect 143738 216944 145044 217000
rect 174822 216972 174882 217078
rect 177993 217075 178059 217078
rect 143677 216942 145044 216944
rect 143677 216939 143743 216942
rect 51125 216866 51191 216869
rect 135397 216866 135463 216869
rect 47524 216864 51191 216866
rect 47524 216808 51130 216864
rect 51186 216808 51191 216864
rect 47524 216806 51191 216808
rect 131796 216864 135463 216866
rect 131796 216808 135402 216864
rect 135458 216808 135463 216864
rect 131796 216806 135463 216808
rect 51125 216803 51191 216806
rect 135397 216803 135463 216806
rect 177717 216730 177783 216733
rect 174822 216728 177783 216730
rect 174822 216672 177722 216728
rect 177778 216672 177783 216728
rect 174822 216670 177783 216672
rect 51217 216322 51283 216325
rect 47524 216320 51283 216322
rect 47524 216264 51222 216320
rect 51278 216264 51283 216320
rect 47524 216262 51283 216264
rect 51217 216259 51283 216262
rect 58301 216322 58367 216325
rect 92709 216322 92775 216325
rect 58301 216320 60956 216322
rect 58301 216264 58306 216320
rect 58362 216264 60956 216320
rect 58301 216262 60956 216264
rect 90764 216320 92775 216322
rect 90764 216264 92714 216320
rect 92770 216264 92775 216320
rect 90764 216262 92775 216264
rect 58301 216259 58367 216262
rect 92709 216259 92775 216262
rect 101357 216186 101423 216189
rect 103982 216186 104042 216632
rect 135489 216322 135555 216325
rect 131796 216320 135555 216322
rect 131796 216264 135494 216320
rect 135550 216264 135555 216320
rect 131796 216262 135555 216264
rect 135489 216259 135555 216262
rect 143125 216322 143191 216325
rect 143125 216320 145044 216322
rect 143125 216264 143130 216320
rect 143186 216264 145044 216320
rect 174822 216292 174882 216670
rect 177717 216667 177783 216670
rect 185169 216730 185235 216733
rect 185169 216728 187916 216730
rect 185169 216672 185174 216728
rect 185230 216672 187916 216728
rect 185169 216670 187916 216672
rect 185169 216667 185235 216670
rect 143125 216262 145044 216264
rect 143125 216259 143191 216262
rect 101357 216184 104042 216186
rect 101357 216128 101362 216184
rect 101418 216128 104042 216184
rect 101357 216126 104042 216128
rect 101357 216123 101423 216126
rect 100713 216050 100779 216053
rect 184801 216050 184867 216053
rect 100713 216048 104012 216050
rect 100713 215992 100718 216048
rect 100774 215992 104012 216048
rect 100713 215990 104012 215992
rect 184801 216048 187916 216050
rect 184801 215992 184806 216048
rect 184862 215992 187916 216048
rect 184801 215990 187916 215992
rect 100713 215987 100779 215990
rect 184801 215987 184867 215990
rect 51217 215778 51283 215781
rect 47524 215776 51283 215778
rect 47524 215720 51222 215776
rect 51278 215720 51283 215776
rect 47524 215718 51283 215720
rect 51217 215715 51283 215718
rect 58209 215778 58275 215781
rect 92709 215778 92775 215781
rect 135397 215778 135463 215781
rect 58209 215776 60956 215778
rect 58209 215720 58214 215776
rect 58270 215720 60956 215776
rect 58209 215718 60956 215720
rect 90764 215776 92775 215778
rect 90764 215720 92714 215776
rect 92770 215720 92775 215776
rect 90764 215718 92775 215720
rect 131796 215776 135463 215778
rect 131796 215720 135402 215776
rect 135458 215720 135463 215776
rect 131796 215718 135463 215720
rect 58209 215715 58275 215718
rect 92709 215715 92775 215718
rect 135397 215715 135463 215718
rect 143125 215778 143191 215781
rect 143125 215776 145044 215778
rect 143125 215720 143130 215776
rect 143186 215720 145044 215776
rect 143125 215718 145044 215720
rect 143125 215715 143191 215718
rect 174822 215642 174882 215748
rect 177717 215642 177783 215645
rect 174822 215640 177783 215642
rect 174822 215584 177722 215640
rect 177778 215584 177783 215640
rect 174822 215582 177783 215584
rect 177717 215579 177783 215582
rect 177625 215506 177691 215509
rect 174822 215504 177691 215506
rect 174822 215448 177630 215504
rect 177686 215448 177691 215504
rect 174822 215446 177691 215448
rect 58301 215234 58367 215237
rect 92801 215234 92867 215237
rect 58301 215232 60956 215234
rect 58301 215176 58306 215232
rect 58362 215176 60956 215232
rect 58301 215174 60956 215176
rect 90764 215232 92867 215234
rect 90764 215176 92806 215232
rect 92862 215176 92867 215232
rect 90764 215174 92867 215176
rect 58301 215171 58367 215174
rect 92801 215171 92867 215174
rect 50389 215098 50455 215101
rect 47524 215096 50455 215098
rect 47524 215040 50394 215096
rect 50450 215040 50455 215096
rect 47524 215038 50455 215040
rect 50389 215035 50455 215038
rect 100989 215098 101055 215101
rect 103982 215098 104042 215408
rect 142941 215234 143007 215237
rect 142941 215232 145044 215234
rect 142941 215176 142946 215232
rect 143002 215176 145044 215232
rect 174822 215204 174882 215446
rect 177625 215443 177691 215446
rect 185169 215506 185235 215509
rect 185169 215504 187916 215506
rect 185169 215448 185174 215504
rect 185230 215448 187916 215504
rect 185169 215446 187916 215448
rect 185169 215443 185235 215446
rect 220313 215234 220379 215237
rect 215884 215232 220379 215234
rect 142941 215174 145044 215176
rect 215884 215176 220318 215232
rect 220374 215176 220379 215232
rect 215884 215174 220379 215176
rect 142941 215171 143007 215174
rect 220313 215171 220379 215174
rect 134845 215098 134911 215101
rect 100989 215096 104042 215098
rect 100989 215040 100994 215096
rect 101050 215040 104042 215096
rect 100989 215038 104042 215040
rect 131796 215096 134911 215098
rect 131796 215040 134850 215096
rect 134906 215040 134911 215096
rect 131796 215038 134911 215040
rect 100989 215035 101055 215038
rect 134845 215035 134911 215038
rect 177165 214962 177231 214965
rect 174822 214960 177231 214962
rect 174822 214904 177170 214960
rect 177226 214904 177231 214960
rect 174822 214902 177231 214904
rect 100805 214690 100871 214693
rect 103982 214690 104042 214864
rect 100805 214688 104042 214690
rect 100805 214632 100810 214688
rect 100866 214632 104042 214688
rect 100805 214630 104042 214632
rect 100805 214627 100871 214630
rect 51125 214554 51191 214557
rect 47524 214552 51191 214554
rect 47524 214496 51130 214552
rect 51186 214496 51191 214552
rect 47524 214494 51191 214496
rect 51125 214491 51191 214494
rect 58209 214554 58275 214557
rect 93537 214554 93603 214557
rect 135305 214554 135371 214557
rect 58209 214552 60956 214554
rect 58209 214496 58214 214552
rect 58270 214496 60956 214552
rect 58209 214494 60956 214496
rect 90764 214552 93603 214554
rect 90764 214496 93542 214552
rect 93598 214496 93603 214552
rect 90764 214494 93603 214496
rect 131796 214552 135371 214554
rect 131796 214496 135310 214552
rect 135366 214496 135371 214552
rect 131796 214494 135371 214496
rect 58209 214491 58275 214494
rect 93537 214491 93603 214494
rect 135305 214491 135371 214494
rect 143493 214554 143559 214557
rect 143493 214552 145044 214554
rect 143493 214496 143498 214552
rect 143554 214496 145044 214552
rect 174822 214524 174882 214902
rect 177165 214899 177231 214902
rect 184893 214962 184959 214965
rect 184893 214960 187916 214962
rect 184893 214904 184898 214960
rect 184954 214904 187916 214960
rect 184893 214902 187916 214904
rect 184893 214899 184959 214902
rect 143493 214494 145044 214496
rect 143493 214491 143559 214494
rect 185261 214418 185327 214421
rect 185261 214416 187916 214418
rect 185261 214360 185266 214416
rect 185322 214360 187916 214416
rect 185261 214358 187916 214360
rect 185261 214355 185327 214358
rect 50389 214010 50455 214013
rect 47524 214008 50455 214010
rect 47524 213952 50394 214008
rect 50450 213952 50455 214008
rect 47524 213950 50455 213952
rect 50389 213947 50455 213950
rect 58209 214010 58275 214013
rect 92709 214010 92775 214013
rect 58209 214008 60956 214010
rect 58209 213952 58214 214008
rect 58270 213952 60956 214008
rect 58209 213950 60956 213952
rect 90764 214008 92775 214010
rect 90764 213952 92714 214008
rect 92770 213952 92775 214008
rect 90764 213950 92775 213952
rect 58209 213947 58275 213950
rect 92709 213947 92775 213950
rect 100989 214010 101055 214013
rect 103982 214010 104042 214320
rect 177717 214146 177783 214149
rect 174822 214144 177783 214146
rect 174822 214088 177722 214144
rect 177778 214088 177783 214144
rect 174822 214086 177783 214088
rect 134477 214010 134543 214013
rect 100989 214008 104042 214010
rect 100989 213952 100994 214008
rect 101050 213952 104042 214008
rect 100989 213950 104042 213952
rect 131796 214008 134543 214010
rect 131796 213952 134482 214008
rect 134538 213952 134543 214008
rect 131796 213950 134543 213952
rect 100989 213947 101055 213950
rect 134477 213947 134543 213950
rect 142941 214010 143007 214013
rect 142941 214008 145044 214010
rect 142941 213952 142946 214008
rect 143002 213952 145044 214008
rect 174822 213980 174882 214086
rect 177717 214083 177783 214086
rect 142941 213950 145044 213952
rect 142941 213947 143007 213950
rect 184985 213874 185051 213877
rect 184985 213872 187916 213874
rect 184985 213816 184990 213872
rect 185046 213816 187916 213872
rect 184985 213814 187916 213816
rect 184985 213811 185051 213814
rect 51217 213466 51283 213469
rect 47524 213464 51283 213466
rect 47524 213408 51222 213464
rect 51278 213408 51283 213464
rect 47524 213406 51283 213408
rect 51217 213403 51283 213406
rect 100713 213466 100779 213469
rect 103982 213466 104042 213776
rect 177625 213738 177691 213741
rect 174822 213736 177691 213738
rect 174822 213680 177630 213736
rect 177686 213680 177691 213736
rect 174822 213678 177691 213680
rect 134477 213466 134543 213469
rect 100713 213464 104042 213466
rect 100713 213408 100718 213464
rect 100774 213408 104042 213464
rect 100713 213406 104042 213408
rect 131796 213464 134543 213466
rect 131796 213408 134482 213464
rect 134538 213408 134543 213464
rect 131796 213406 134543 213408
rect 100713 213403 100779 213406
rect 134477 213403 134543 213406
rect 58301 213330 58367 213333
rect 93353 213330 93419 213333
rect 58301 213328 60956 213330
rect 58301 213272 58306 213328
rect 58362 213272 60956 213328
rect 58301 213270 60956 213272
rect 90764 213328 93419 213330
rect 90764 213272 93358 213328
rect 93414 213272 93419 213328
rect 90764 213270 93419 213272
rect 58301 213267 58367 213270
rect 93353 213267 93419 213270
rect 143677 213330 143743 213333
rect 143677 213328 145044 213330
rect 143677 213272 143682 213328
rect 143738 213272 145044 213328
rect 174822 213300 174882 213678
rect 177625 213675 177691 213678
rect 185077 213330 185143 213333
rect 185077 213328 187916 213330
rect 143677 213270 145044 213272
rect 185077 213272 185082 213328
rect 185138 213272 187916 213328
rect 185077 213270 187916 213272
rect 143677 213267 143743 213270
rect 185077 213267 185143 213270
rect 103614 213202 104012 213262
rect 100897 213194 100963 213197
rect 103614 213194 103674 213202
rect 100897 213192 103674 213194
rect 100897 213136 100902 213192
rect 100958 213136 103674 213192
rect 100897 213134 103674 213136
rect 100897 213131 100963 213134
rect 51217 212922 51283 212925
rect 134477 212922 134543 212925
rect 177717 212922 177783 212925
rect 47524 212920 51283 212922
rect 47524 212864 51222 212920
rect 51278 212864 51283 212920
rect 47524 212862 51283 212864
rect 131796 212920 134543 212922
rect 131796 212864 134482 212920
rect 134538 212864 134543 212920
rect 131796 212862 134543 212864
rect 51217 212859 51283 212862
rect 134477 212859 134543 212862
rect 174822 212920 177783 212922
rect 174822 212864 177722 212920
rect 177778 212864 177783 212920
rect 174822 212862 177783 212864
rect 58209 212786 58275 212789
rect 92709 212786 92775 212789
rect 58209 212784 60956 212786
rect 58209 212728 58214 212784
rect 58270 212728 60956 212784
rect 58209 212726 60956 212728
rect 90764 212784 92775 212786
rect 90764 212728 92714 212784
rect 92770 212728 92775 212784
rect 90764 212726 92775 212728
rect 58209 212723 58275 212726
rect 92709 212723 92775 212726
rect 143677 212786 143743 212789
rect 143677 212784 145044 212786
rect 143677 212728 143682 212784
rect 143738 212728 145044 212784
rect 174822 212756 174882 212862
rect 177717 212859 177783 212862
rect 185169 212786 185235 212789
rect 185169 212784 187916 212786
rect 143677 212726 145044 212728
rect 185169 212728 185174 212784
rect 185230 212728 187916 212784
rect 185169 212726 187916 212728
rect 143677 212723 143743 212726
rect 185169 212723 185235 212726
rect 100989 212378 101055 212381
rect 103982 212378 104042 212688
rect 177165 212514 177231 212517
rect 100989 212376 104042 212378
rect 100989 212320 100994 212376
rect 101050 212320 104042 212376
rect 100989 212318 104042 212320
rect 174822 212512 177231 212514
rect 174822 212456 177170 212512
rect 177226 212456 177231 212512
rect 174822 212454 177231 212456
rect 100989 212315 101055 212318
rect 51125 212242 51191 212245
rect 47524 212240 51191 212242
rect 47524 212184 51130 212240
rect 51186 212184 51191 212240
rect 47524 212182 51191 212184
rect 51125 212179 51191 212182
rect 58301 212242 58367 212245
rect 93353 212242 93419 212245
rect 134661 212242 134727 212245
rect 58301 212240 60956 212242
rect 58301 212184 58306 212240
rect 58362 212184 60956 212240
rect 58301 212182 60956 212184
rect 90764 212240 93419 212242
rect 90764 212184 93358 212240
rect 93414 212184 93419 212240
rect 90764 212182 93419 212184
rect 131796 212240 134727 212242
rect 131796 212184 134666 212240
rect 134722 212184 134727 212240
rect 131796 212182 134727 212184
rect 58301 212179 58367 212182
rect 93353 212179 93419 212182
rect 134661 212179 134727 212182
rect 143493 212242 143559 212245
rect 143493 212240 145044 212242
rect 143493 212184 143498 212240
rect 143554 212184 145044 212240
rect 174822 212212 174882 212454
rect 177165 212451 177231 212454
rect 185445 212242 185511 212245
rect 185445 212240 187916 212242
rect 143493 212182 145044 212184
rect 185445 212184 185450 212240
rect 185506 212184 187916 212240
rect 185445 212182 187916 212184
rect 143493 212179 143559 212182
rect 185445 212179 185511 212182
rect 101265 211970 101331 211973
rect 103982 211970 104042 212144
rect 101265 211968 104042 211970
rect 101265 211912 101270 211968
rect 101326 211912 104042 211968
rect 101265 211910 104042 211912
rect 101265 211907 101331 211910
rect 51217 211698 51283 211701
rect 134569 211698 134635 211701
rect 177717 211698 177783 211701
rect 47524 211696 51283 211698
rect 47524 211640 51222 211696
rect 51278 211640 51283 211696
rect 47524 211638 51283 211640
rect 131796 211696 134635 211698
rect 131796 211640 134574 211696
rect 134630 211640 134635 211696
rect 131796 211638 134635 211640
rect 51217 211635 51283 211638
rect 134569 211635 134635 211638
rect 174822 211696 177783 211698
rect 174822 211640 177722 211696
rect 177778 211640 177783 211696
rect 174822 211638 177783 211640
rect 58209 211562 58275 211565
rect 92709 211562 92775 211565
rect 58209 211560 60956 211562
rect 58209 211504 58214 211560
rect 58270 211504 60956 211560
rect 58209 211502 60956 211504
rect 90764 211560 92775 211562
rect 90764 211504 92714 211560
rect 92770 211504 92775 211560
rect 90764 211502 92775 211504
rect 58209 211499 58275 211502
rect 92709 211499 92775 211502
rect 143677 211562 143743 211565
rect 143677 211560 145044 211562
rect 143677 211504 143682 211560
rect 143738 211504 145044 211560
rect 174822 211532 174882 211638
rect 177717 211635 177783 211638
rect 185353 211562 185419 211565
rect 185353 211560 187916 211562
rect 143677 211502 145044 211504
rect 185353 211504 185358 211560
rect 185414 211504 187916 211560
rect 185353 211502 187916 211504
rect 143677 211499 143743 211502
rect 185353 211499 185419 211502
rect 50849 211154 50915 211157
rect 47524 211152 50915 211154
rect 47524 211096 50854 211152
rect 50910 211096 50915 211152
rect 47524 211094 50915 211096
rect 50849 211091 50915 211094
rect 101173 211154 101239 211157
rect 103982 211154 104042 211464
rect 177165 211290 177231 211293
rect 174822 211288 177231 211290
rect 174822 211232 177170 211288
rect 177226 211232 177231 211288
rect 174822 211230 177231 211232
rect 135029 211154 135095 211157
rect 101173 211152 104042 211154
rect 101173 211096 101178 211152
rect 101234 211096 104042 211152
rect 101173 211094 104042 211096
rect 131796 211152 135095 211154
rect 131796 211096 135034 211152
rect 135090 211096 135095 211152
rect 131796 211094 135095 211096
rect 101173 211091 101239 211094
rect 135029 211091 135095 211094
rect 58301 211018 58367 211021
rect 92801 211018 92867 211021
rect 58301 211016 60956 211018
rect 58301 210960 58306 211016
rect 58362 210960 60956 211016
rect 58301 210958 60956 210960
rect 90764 211016 92867 211018
rect 90764 210960 92806 211016
rect 92862 210960 92867 211016
rect 90764 210958 92867 210960
rect 58301 210955 58367 210958
rect 92801 210955 92867 210958
rect 143677 211018 143743 211021
rect 143677 211016 145044 211018
rect 143677 210960 143682 211016
rect 143738 210960 145044 211016
rect 174822 210988 174882 211230
rect 177165 211227 177231 211230
rect 185261 211018 185327 211021
rect 185261 211016 187916 211018
rect 143677 210958 145044 210960
rect 185261 210960 185266 211016
rect 185322 210960 187916 211016
rect 185261 210958 187916 210960
rect 143677 210955 143743 210958
rect 185261 210955 185327 210958
rect 101081 210746 101147 210749
rect 103982 210746 104042 210920
rect 101081 210744 104042 210746
rect 101081 210688 101086 210744
rect 101142 210688 104042 210744
rect 101081 210686 104042 210688
rect 101081 210683 101147 210686
rect 50665 210610 50731 210613
rect 134845 210610 134911 210613
rect 177717 210610 177783 210613
rect 47524 210608 50731 210610
rect 47524 210552 50670 210608
rect 50726 210552 50731 210608
rect 47524 210550 50731 210552
rect 131796 210608 134911 210610
rect 131796 210552 134850 210608
rect 134906 210552 134911 210608
rect 131796 210550 134911 210552
rect 50665 210547 50731 210550
rect 134845 210547 134911 210550
rect 174822 210608 177783 210610
rect 174822 210552 177722 210608
rect 177778 210552 177783 210608
rect 174822 210550 177783 210552
rect 100989 210474 101055 210477
rect 100989 210472 104012 210474
rect 100989 210416 100994 210472
rect 101050 210416 104012 210472
rect 100989 210414 104012 210416
rect 100989 210411 101055 210414
rect 58393 210338 58459 210341
rect 92893 210338 92959 210341
rect 58393 210336 60956 210338
rect 58393 210280 58398 210336
rect 58454 210280 60956 210336
rect 58393 210278 60956 210280
rect 90764 210336 92959 210338
rect 90764 210280 92898 210336
rect 92954 210280 92959 210336
rect 90764 210278 92959 210280
rect 58393 210275 58459 210278
rect 92893 210275 92959 210278
rect 143585 210338 143651 210341
rect 143585 210336 145044 210338
rect 143585 210280 143590 210336
rect 143646 210280 145044 210336
rect 174822 210308 174882 210550
rect 177717 210547 177783 210550
rect 185169 210474 185235 210477
rect 185169 210472 187916 210474
rect 185169 210416 185174 210472
rect 185230 210416 187916 210472
rect 185169 210414 187916 210416
rect 185169 210411 185235 210414
rect 143585 210278 145044 210280
rect 143585 210275 143651 210278
rect 50757 210066 50823 210069
rect 135121 210066 135187 210069
rect 177165 210066 177231 210069
rect 47524 210064 50823 210066
rect 47524 210008 50762 210064
rect 50818 210008 50823 210064
rect 47524 210006 50823 210008
rect 131796 210064 135187 210066
rect 131796 210008 135126 210064
rect 135182 210008 135187 210064
rect 131796 210006 135187 210008
rect 50757 210003 50823 210006
rect 135121 210003 135187 210006
rect 174822 210064 177231 210066
rect 174822 210008 177170 210064
rect 177226 210008 177231 210064
rect 174822 210006 177231 210008
rect 58209 209794 58275 209797
rect 93169 209794 93235 209797
rect 58209 209792 60956 209794
rect 58209 209736 58214 209792
rect 58270 209736 60956 209792
rect 58209 209734 60956 209736
rect 90764 209792 93235 209794
rect 90764 209736 93174 209792
rect 93230 209736 93235 209792
rect 90764 209734 93235 209736
rect 58209 209731 58275 209734
rect 93169 209731 93235 209734
rect 100989 209522 101055 209525
rect 103982 209522 104042 209832
rect 142941 209794 143007 209797
rect 142941 209792 145044 209794
rect 142941 209736 142946 209792
rect 143002 209736 145044 209792
rect 174822 209764 174882 210006
rect 177165 210003 177231 210006
rect 185169 209930 185235 209933
rect 185169 209928 187916 209930
rect 185169 209872 185174 209928
rect 185230 209872 187916 209928
rect 185169 209870 187916 209872
rect 185169 209867 185235 209870
rect 142941 209734 145044 209736
rect 142941 209731 143007 209734
rect 218289 209658 218355 209661
rect 215884 209656 218355 209658
rect 215884 209600 218294 209656
rect 218350 209600 218355 209656
rect 215884 209598 218355 209600
rect 218289 209595 218355 209598
rect 177717 209522 177783 209525
rect 100989 209520 104042 209522
rect 100989 209464 100994 209520
rect 101050 209464 104042 209520
rect 100989 209462 104042 209464
rect 174822 209520 177783 209522
rect 174822 209464 177722 209520
rect 177778 209464 177783 209520
rect 174822 209462 177783 209464
rect 100989 209459 101055 209462
rect 9896 209386 10376 209416
rect 14693 209386 14759 209389
rect 50941 209386 51007 209389
rect 134937 209386 135003 209389
rect 9896 209384 14759 209386
rect 9896 209328 14698 209384
rect 14754 209328 14759 209384
rect 9896 209326 14759 209328
rect 47524 209384 51007 209386
rect 47524 209328 50946 209384
rect 51002 209328 51007 209384
rect 47524 209326 51007 209328
rect 131796 209384 135003 209386
rect 131796 209328 134942 209384
rect 134998 209328 135003 209384
rect 131796 209326 135003 209328
rect 9896 209296 10376 209326
rect 14693 209323 14759 209326
rect 50941 209323 51007 209326
rect 134937 209323 135003 209326
rect 58301 209250 58367 209253
rect 92709 209250 92775 209253
rect 58301 209248 60956 209250
rect 58301 209192 58306 209248
rect 58362 209192 60956 209248
rect 58301 209190 60956 209192
rect 90764 209248 92775 209250
rect 90764 209192 92714 209248
rect 92770 209192 92775 209248
rect 90764 209190 92775 209192
rect 58301 209187 58367 209190
rect 92709 209187 92775 209190
rect 88518 208916 88524 208980
rect 88588 208978 88594 208980
rect 88753 208978 88819 208981
rect 88588 208976 88819 208978
rect 88588 208920 88758 208976
rect 88814 208920 88819 208976
rect 88588 208918 88819 208920
rect 88588 208916 88594 208918
rect 88753 208915 88819 208918
rect 101633 208978 101699 208981
rect 103982 208978 104042 209288
rect 143677 209250 143743 209253
rect 143677 209248 145044 209250
rect 143677 209192 143682 209248
rect 143738 209192 145044 209248
rect 174822 209220 174882 209462
rect 177717 209459 177783 209462
rect 185721 209386 185787 209389
rect 185721 209384 187916 209386
rect 185721 209328 185726 209384
rect 185782 209328 187916 209384
rect 185721 209326 187916 209328
rect 185721 209323 185787 209326
rect 143677 209190 145044 209192
rect 143677 209187 143743 209190
rect 101633 208976 104042 208978
rect 101633 208920 101638 208976
rect 101694 208920 104042 208976
rect 101633 208918 104042 208920
rect 101633 208915 101699 208918
rect 171318 208916 171324 208980
rect 171388 208978 171394 208980
rect 172289 208978 172355 208981
rect 171388 208976 172355 208978
rect 171388 208920 172294 208976
rect 172350 208920 172355 208976
rect 171388 208918 172355 208920
rect 171388 208916 171394 208918
rect 172289 208915 172355 208918
rect 51033 208842 51099 208845
rect 135397 208842 135463 208845
rect 47524 208840 51099 208842
rect 47524 208784 51038 208840
rect 51094 208784 51099 208840
rect 47524 208782 51099 208784
rect 131796 208840 135463 208842
rect 131796 208784 135402 208840
rect 135458 208784 135463 208840
rect 131796 208782 135463 208784
rect 51033 208779 51099 208782
rect 135397 208779 135463 208782
rect 185905 208842 185971 208845
rect 185905 208840 187916 208842
rect 185905 208784 185910 208840
rect 185966 208784 187916 208840
rect 185905 208782 187916 208784
rect 185905 208779 185971 208782
rect 101725 208434 101791 208437
rect 103982 208434 104042 208744
rect 101725 208432 104042 208434
rect 101725 208376 101730 208432
rect 101786 208376 104042 208432
rect 101725 208374 104042 208376
rect 101725 208371 101791 208374
rect 51217 208298 51283 208301
rect 135213 208298 135279 208301
rect 47524 208296 51283 208298
rect 47524 208240 51222 208296
rect 51278 208240 51283 208296
rect 47524 208238 51283 208240
rect 131796 208296 135279 208298
rect 131796 208240 135218 208296
rect 135274 208240 135279 208296
rect 131796 208238 135279 208240
rect 51217 208235 51283 208238
rect 135213 208235 135279 208238
rect 186273 208298 186339 208301
rect 186273 208296 187916 208298
rect 186273 208240 186278 208296
rect 186334 208240 187916 208296
rect 186273 208238 187916 208240
rect 186273 208235 186339 208238
rect 102093 207890 102159 207893
rect 103982 207890 104042 208200
rect 102093 207888 104042 207890
rect 102093 207832 102098 207888
rect 102154 207832 104042 207888
rect 102093 207830 104042 207832
rect 102093 207827 102159 207830
rect 50481 207754 50547 207757
rect 134201 207754 134267 207757
rect 47524 207752 50547 207754
rect 47524 207696 50486 207752
rect 50542 207696 50547 207752
rect 47524 207694 50547 207696
rect 131796 207752 134267 207754
rect 131796 207696 134206 207752
rect 134262 207696 134267 207752
rect 131796 207694 134267 207696
rect 50481 207691 50547 207694
rect 134201 207691 134267 207694
rect 186089 207754 186155 207757
rect 186089 207752 187916 207754
rect 186089 207696 186094 207752
rect 186150 207696 187916 207752
rect 186089 207694 187916 207696
rect 186089 207691 186155 207694
rect 103614 207626 104012 207686
rect 101909 207618 101975 207621
rect 103614 207618 103674 207626
rect 101909 207616 103674 207618
rect 101909 207560 101914 207616
rect 101970 207560 103674 207616
rect 101909 207558 103674 207560
rect 101909 207555 101975 207558
rect 51125 207210 51191 207213
rect 135305 207210 135371 207213
rect 47524 207208 51191 207210
rect 47524 207152 51130 207208
rect 51186 207152 51191 207208
rect 47524 207150 51191 207152
rect 131796 207208 135371 207210
rect 131796 207152 135310 207208
rect 135366 207152 135371 207208
rect 131796 207150 135371 207152
rect 51125 207147 51191 207150
rect 135305 207147 135371 207150
rect 185169 207210 185235 207213
rect 185169 207208 187916 207210
rect 185169 207152 185174 207208
rect 185230 207152 187916 207208
rect 185169 207150 187916 207152
rect 185169 207147 185235 207150
rect 100989 206530 101055 206533
rect 103982 206530 104042 207112
rect 100989 206528 104042 206530
rect 100989 206472 100994 206528
rect 101050 206472 104042 206528
rect 100989 206470 104042 206472
rect 100989 206467 101055 206470
rect 222337 205442 222403 205445
rect 225416 205442 225896 205472
rect 222337 205440 225896 205442
rect 222337 205384 222342 205440
rect 222398 205384 225896 205440
rect 222337 205382 225896 205384
rect 222337 205379 222403 205382
rect 225416 205352 225896 205382
rect 140222 195180 140228 195244
rect 140292 195242 140298 195244
rect 167137 195242 167203 195245
rect 140292 195240 167203 195242
rect 140292 195184 167142 195240
rect 167198 195184 167203 195240
rect 140292 195182 167203 195184
rect 140292 195180 140298 195182
rect 167137 195179 167203 195182
rect 99517 193746 99583 193749
rect 95702 193744 99583 193746
rect 95702 193688 99522 193744
rect 99578 193688 99583 193744
rect 95702 193686 99583 193688
rect 95702 193240 95762 193686
rect 99517 193683 99583 193686
rect 183697 193202 183763 193205
rect 179820 193200 183763 193202
rect 179820 193144 183702 193200
rect 183758 193144 183763 193200
rect 179820 193142 183763 193144
rect 183697 193139 183763 193142
rect 191977 192794 192043 192797
rect 191977 192792 193988 192794
rect 191977 192736 191982 192792
rect 192038 192736 193988 192792
rect 191977 192734 193988 192736
rect 191977 192731 192043 192734
rect 105773 192522 105839 192525
rect 105773 192520 109900 192522
rect 105773 192464 105778 192520
rect 105834 192464 109900 192520
rect 105773 192462 109900 192464
rect 105773 192459 105839 192462
rect 99425 192386 99491 192389
rect 95702 192384 99491 192386
rect 95702 192328 99430 192384
rect 99486 192328 99491 192384
rect 95702 192326 99491 192328
rect 95702 192016 95762 192326
rect 99425 192323 99491 192326
rect 183605 191978 183671 191981
rect 179820 191976 183671 191978
rect 179820 191920 183610 191976
rect 183666 191920 183671 191976
rect 179820 191918 183671 191920
rect 183605 191915 183671 191918
rect 99241 190754 99307 190757
rect 183421 190754 183487 190757
rect 209917 190756 209983 190757
rect 209917 190754 209964 190756
rect 95732 190752 99307 190754
rect 95732 190696 99246 190752
rect 99302 190696 99307 190752
rect 95732 190694 99307 190696
rect 179820 190752 183487 190754
rect 179820 190696 183426 190752
rect 183482 190696 183487 190752
rect 209876 190752 209964 190754
rect 210028 190754 210034 190756
rect 179820 190694 183487 190696
rect 99241 190691 99307 190694
rect 183421 190691 183487 190694
rect 193958 190620 194018 190724
rect 209876 190696 209922 190752
rect 209876 190694 209964 190696
rect 209917 190692 209964 190694
rect 210028 190694 210110 190754
rect 210028 190692 210034 190694
rect 209917 190691 209983 190692
rect 193950 190556 193956 190620
rect 194020 190556 194026 190620
rect 22789 190482 22855 190485
rect 211941 190482 212007 190485
rect 22789 190480 25996 190482
rect 22789 190424 22794 190480
rect 22850 190424 25996 190480
rect 22789 190422 25996 190424
rect 209812 190480 212007 190482
rect 209812 190424 211946 190480
rect 212002 190424 212007 190480
rect 209812 190422 212007 190424
rect 22789 190419 22855 190422
rect 211941 190419 212007 190422
rect 107153 190210 107219 190213
rect 107153 190208 109900 190210
rect 107153 190152 107158 190208
rect 107214 190152 109900 190208
rect 107153 190150 109900 190152
rect 107153 190147 107219 190150
rect 99149 189530 99215 189533
rect 183513 189530 183579 189533
rect 95732 189528 99215 189530
rect 95732 189472 99154 189528
rect 99210 189472 99215 189528
rect 95732 189470 99215 189472
rect 179820 189528 183579 189530
rect 179820 189472 183518 189528
rect 183574 189472 183579 189528
rect 179820 189470 183579 189472
rect 99149 189467 99215 189470
rect 183513 189467 183579 189470
rect 41833 189258 41899 189261
rect 41790 189256 41899 189258
rect 41790 189200 41838 189256
rect 41894 189200 41899 189256
rect 41790 189195 41899 189200
rect 41790 188684 41850 189195
rect 99333 188986 99399 188989
rect 95702 188984 99399 188986
rect 95702 188928 99338 188984
rect 99394 188928 99399 188984
rect 95702 188926 99399 188928
rect 95702 188344 95762 188926
rect 99333 188923 99399 188926
rect 191977 188714 192043 188717
rect 191977 188712 193988 188714
rect 191977 188656 191982 188712
rect 192038 188656 193988 188712
rect 191977 188654 193988 188656
rect 191977 188651 192043 188654
rect 183329 188306 183395 188309
rect 179820 188304 183395 188306
rect 179820 188248 183334 188304
rect 183390 188248 183395 188304
rect 179820 188246 183395 188248
rect 183329 188243 183395 188246
rect 106785 187898 106851 187901
rect 106785 187896 109900 187898
rect 106785 187840 106790 187896
rect 106846 187840 109900 187896
rect 106785 187838 109900 187840
rect 106785 187835 106851 187838
rect 99057 187762 99123 187765
rect 95702 187760 99123 187762
rect 95702 187704 99062 187760
rect 99118 187704 99123 187760
rect 95702 187702 99123 187704
rect 95702 187120 95762 187702
rect 99057 187699 99123 187702
rect 183237 187082 183303 187085
rect 179820 187080 183303 187082
rect 179820 187024 183242 187080
rect 183298 187024 183303 187080
rect 179820 187022 183303 187024
rect 183237 187019 183303 187022
rect 191149 186810 191215 186813
rect 191149 186808 193988 186810
rect 191149 186752 191154 186808
rect 191210 186752 193988 186808
rect 191149 186750 193988 186752
rect 191149 186747 191215 186750
rect 98965 186538 99031 186541
rect 95702 186536 99031 186538
rect 95702 186480 98970 186536
rect 99026 186480 99031 186536
rect 95702 186478 99031 186480
rect 95702 185896 95762 186478
rect 98965 186475 99031 186478
rect 183145 185858 183211 185861
rect 179820 185856 183211 185858
rect 179820 185800 183150 185856
rect 183206 185800 183211 185856
rect 179820 185798 183211 185800
rect 183145 185795 183211 185798
rect 9896 185722 10376 185752
rect 13313 185722 13379 185725
rect 9896 185720 13379 185722
rect 9896 185664 13318 185720
rect 13374 185664 13379 185720
rect 9896 185662 13379 185664
rect 9896 185632 10376 185662
rect 13313 185659 13379 185662
rect 106785 185450 106851 185453
rect 106785 185448 109900 185450
rect 106785 185392 106790 185448
rect 106846 185392 109900 185448
rect 106785 185390 109900 185392
rect 106785 185387 106851 185390
rect 98873 185314 98939 185317
rect 95702 185312 98939 185314
rect 95702 185256 98878 185312
rect 98934 185256 98939 185312
rect 95702 185254 98939 185256
rect 95702 184672 95762 185254
rect 98873 185251 98939 185254
rect 191977 184770 192043 184773
rect 191977 184768 193988 184770
rect 191977 184712 191982 184768
rect 192038 184712 193988 184768
rect 191977 184710 193988 184712
rect 191977 184707 192043 184710
rect 183053 184634 183119 184637
rect 179820 184632 183119 184634
rect 179820 184576 183058 184632
rect 183114 184576 183119 184632
rect 179820 184574 183119 184576
rect 183053 184571 183119 184574
rect 22329 183818 22395 183821
rect 128497 183818 128563 183821
rect 212493 183818 212559 183821
rect 22329 183816 25996 183818
rect 22329 183760 22334 183816
rect 22390 183760 25996 183816
rect 22329 183758 25996 183760
rect 125724 183816 128563 183818
rect 125724 183760 128502 183816
rect 128558 183760 128563 183816
rect 125724 183758 128563 183760
rect 209812 183816 212559 183818
rect 209812 183760 212498 183816
rect 212554 183760 212559 183816
rect 209812 183758 212559 183760
rect 22329 183755 22395 183758
rect 128497 183755 128563 183758
rect 212493 183755 212559 183758
rect 99517 183682 99583 183685
rect 95702 183680 99583 183682
rect 95702 183624 99522 183680
rect 99578 183624 99583 183680
rect 95702 183622 99583 183624
rect 95702 183448 95762 183622
rect 99517 183619 99583 183622
rect 182869 183410 182935 183413
rect 179820 183408 182935 183410
rect 179820 183352 182874 183408
rect 182930 183352 182935 183408
rect 179820 183350 182935 183352
rect 182869 183347 182935 183350
rect 107153 183138 107219 183141
rect 107153 183136 109900 183138
rect 107153 183080 107158 183136
rect 107214 183080 109900 183136
rect 107153 183078 109900 183080
rect 107153 183075 107219 183078
rect 190597 182730 190663 182733
rect 190597 182728 193988 182730
rect 190597 182672 190602 182728
rect 190658 182672 193988 182728
rect 190597 182670 193988 182672
rect 190597 182667 190663 182670
rect 98597 182458 98663 182461
rect 95702 182456 98663 182458
rect 95702 182400 98602 182456
rect 98658 182400 98663 182456
rect 95702 182398 98663 182400
rect 95702 182224 95762 182398
rect 98597 182395 98663 182398
rect 183145 182186 183211 182189
rect 179820 182184 183211 182186
rect 179820 182128 183150 182184
rect 183206 182128 183211 182184
rect 179820 182126 183211 182128
rect 183145 182123 183211 182126
rect 99425 181098 99491 181101
rect 183697 181098 183763 181101
rect 95732 181096 99491 181098
rect 95732 181040 99430 181096
rect 99486 181040 99491 181096
rect 95732 181038 99491 181040
rect 179820 181096 183763 181098
rect 179820 181040 183702 181096
rect 183758 181040 183763 181096
rect 179820 181038 183763 181040
rect 99425 181035 99491 181038
rect 183697 181035 183763 181038
rect 106969 180826 107035 180829
rect 190689 180826 190755 180829
rect 106969 180824 109900 180826
rect 106969 180768 106974 180824
rect 107030 180768 109900 180824
rect 106969 180766 109900 180768
rect 190689 180824 193988 180826
rect 190689 180768 190694 180824
rect 190750 180768 193988 180824
rect 190689 180766 193988 180768
rect 106969 180763 107035 180766
rect 190689 180763 190755 180766
rect 99517 179874 99583 179877
rect 183697 179874 183763 179877
rect 95732 179872 99583 179874
rect 95732 179816 99522 179872
rect 99578 179816 99583 179872
rect 95732 179814 99583 179816
rect 179820 179872 183763 179874
rect 179820 179816 183702 179872
rect 183758 179816 183763 179872
rect 179820 179814 183763 179816
rect 99517 179811 99583 179814
rect 183697 179811 183763 179814
rect 98413 179330 98479 179333
rect 95702 179328 98479 179330
rect 95702 179272 98418 179328
rect 98474 179272 98479 179328
rect 95702 179270 98479 179272
rect 23617 178786 23683 178789
rect 25774 178786 25780 178788
rect 23617 178784 25780 178786
rect 23617 178728 23622 178784
rect 23678 178728 25780 178784
rect 23617 178726 25780 178728
rect 23617 178723 23683 178726
rect 25774 178724 25780 178726
rect 25844 178724 25850 178788
rect 41790 178650 41850 178756
rect 95702 178688 95762 179270
rect 98413 179267 98479 179270
rect 220405 179194 220471 179197
rect 225416 179194 225896 179224
rect 220405 179192 225896 179194
rect 220405 179136 220410 179192
rect 220466 179136 225896 179192
rect 220405 179134 225896 179136
rect 220405 179131 220471 179134
rect 225416 179104 225896 179134
rect 191977 178786 192043 178789
rect 191977 178784 193988 178786
rect 191977 178728 191982 178784
rect 192038 178728 193988 178784
rect 191977 178726 193988 178728
rect 191977 178723 192043 178726
rect 41966 178650 41972 178652
rect 41790 178590 41972 178650
rect 41966 178588 41972 178590
rect 42036 178588 42042 178652
rect 182501 178650 182567 178653
rect 179820 178648 182567 178650
rect 179820 178592 182506 178648
rect 182562 178592 182567 178648
rect 179820 178590 182567 178592
rect 182501 178587 182567 178590
rect 106785 178378 106851 178381
rect 106785 178376 109900 178378
rect 106785 178320 106790 178376
rect 106846 178320 109900 178376
rect 106785 178318 109900 178320
rect 106785 178315 106851 178318
rect 99517 177426 99583 177429
rect 182501 177426 182567 177429
rect 95732 177424 99583 177426
rect 95732 177368 99522 177424
rect 99578 177368 99583 177424
rect 95732 177366 99583 177368
rect 179820 177424 182567 177426
rect 179820 177368 182506 177424
rect 182562 177368 182567 177424
rect 179820 177366 182567 177368
rect 99517 177363 99583 177366
rect 182501 177363 182567 177366
rect 22329 177154 22395 177157
rect 211757 177154 211823 177157
rect 22329 177152 25996 177154
rect 22329 177096 22334 177152
rect 22390 177096 25996 177152
rect 22329 177094 25996 177096
rect 209812 177152 211823 177154
rect 209812 177096 211762 177152
rect 211818 177096 211823 177152
rect 209812 177094 211823 177096
rect 22329 177091 22395 177094
rect 211757 177091 211823 177094
rect 98597 176746 98663 176749
rect 95702 176744 98663 176746
rect 95702 176688 98602 176744
rect 98658 176688 98663 176744
rect 95702 176686 98663 176688
rect 95702 176240 95762 176686
rect 98597 176683 98663 176686
rect 191977 176746 192043 176749
rect 191977 176744 193988 176746
rect 191977 176688 191982 176744
rect 192038 176688 193988 176744
rect 191977 176686 193988 176688
rect 191977 176683 192043 176686
rect 183237 176202 183303 176205
rect 179820 176200 183303 176202
rect 179820 176144 183242 176200
rect 183298 176144 183303 176200
rect 179820 176142 183303 176144
rect 183237 176139 183303 176142
rect 106601 176066 106667 176069
rect 106601 176064 109900 176066
rect 106601 176008 106606 176064
rect 106662 176008 109900 176064
rect 106601 176006 109900 176008
rect 106601 176003 106667 176006
rect 98229 175386 98295 175389
rect 95702 175384 98295 175386
rect 95702 175328 98234 175384
rect 98290 175328 98295 175384
rect 95702 175326 98295 175328
rect 95702 175016 95762 175326
rect 98229 175323 98295 175326
rect 183697 174978 183763 174981
rect 179820 174976 183763 174978
rect 179820 174920 183702 174976
rect 183758 174920 183763 174976
rect 179820 174918 183763 174920
rect 183697 174915 183763 174918
rect 191517 174842 191583 174845
rect 191517 174840 193988 174842
rect 191517 174784 191522 174840
rect 191578 174784 193988 174840
rect 191517 174782 193988 174784
rect 191517 174779 191583 174782
rect 137513 174434 137579 174437
rect 137513 174432 140106 174434
rect 137513 174376 137518 174432
rect 137574 174376 140106 174432
rect 137513 174374 140106 174376
rect 137513 174371 137579 174374
rect 140046 173928 140106 174374
rect 53333 173890 53399 173893
rect 53333 173888 55988 173890
rect 53333 173832 53338 173888
rect 53394 173832 55988 173888
rect 53333 173830 55988 173832
rect 53333 173827 53399 173830
rect 99517 173754 99583 173757
rect 95732 173752 99583 173754
rect 95732 173696 99522 173752
rect 99578 173696 99583 173752
rect 95732 173694 99583 173696
rect 99517 173691 99583 173694
rect 106785 173754 106851 173757
rect 183329 173754 183395 173757
rect 106785 173752 109900 173754
rect 106785 173696 106790 173752
rect 106846 173696 109900 173752
rect 106785 173694 109900 173696
rect 179820 173752 183395 173754
rect 179820 173696 183334 173752
rect 183390 173696 183395 173752
rect 179820 173694 183395 173696
rect 106785 173691 106851 173694
rect 183329 173691 183395 173694
rect 191977 172802 192043 172805
rect 191977 172800 193988 172802
rect 191977 172744 191982 172800
rect 192038 172744 193988 172800
rect 191977 172742 193988 172744
rect 191977 172739 192043 172742
rect 99517 172530 99583 172533
rect 183513 172530 183579 172533
rect 95732 172528 99583 172530
rect 95732 172472 99522 172528
rect 99578 172472 99583 172528
rect 95732 172470 99583 172472
rect 179820 172528 183579 172530
rect 179820 172472 183518 172528
rect 183574 172472 183579 172528
rect 179820 172470 183579 172472
rect 99517 172467 99583 172470
rect 183513 172467 183579 172470
rect 106785 171442 106851 171445
rect 106785 171440 109900 171442
rect 106785 171384 106790 171440
rect 106846 171384 109900 171440
rect 106785 171382 109900 171384
rect 106785 171379 106851 171382
rect 99425 171306 99491 171309
rect 182685 171306 182751 171309
rect 95732 171304 99491 171306
rect 95732 171248 99430 171304
rect 99486 171248 99491 171304
rect 95732 171246 99491 171248
rect 179820 171304 182751 171306
rect 179820 171248 182690 171304
rect 182746 171248 182751 171304
rect 179820 171246 182751 171248
rect 99425 171243 99491 171246
rect 182685 171243 182751 171246
rect 209825 171034 209891 171037
rect 209782 171032 209891 171034
rect 209782 170976 209830 171032
rect 209886 170976 209891 171032
rect 209782 170971 209891 170976
rect 191149 170762 191215 170765
rect 191149 170760 193988 170762
rect 191149 170704 191154 170760
rect 191210 170704 193988 170760
rect 191149 170702 193988 170704
rect 191149 170699 191215 170702
rect 23617 170490 23683 170493
rect 23617 170488 25996 170490
rect 23617 170432 23622 170488
rect 23678 170432 25996 170488
rect 209782 170460 209842 170971
rect 23617 170430 25996 170432
rect 23617 170427 23683 170430
rect 99517 170082 99583 170085
rect 182501 170082 182567 170085
rect 95732 170080 99583 170082
rect 95732 170024 99522 170080
rect 99578 170024 99583 170080
rect 95732 170022 99583 170024
rect 179820 170080 182567 170082
rect 179820 170024 182506 170080
rect 182562 170024 182567 170080
rect 179820 170022 182567 170024
rect 99517 170019 99583 170022
rect 182501 170019 182567 170022
rect 106785 168994 106851 168997
rect 106785 168992 109900 168994
rect 106785 168936 106790 168992
rect 106846 168936 109900 168992
rect 106785 168934 109900 168936
rect 106785 168931 106851 168934
rect 99425 168858 99491 168861
rect 183697 168858 183763 168861
rect 95732 168856 99491 168858
rect 95732 168800 99430 168856
rect 99486 168800 99491 168856
rect 95732 168798 99491 168800
rect 179820 168856 183763 168858
rect 179820 168800 183702 168856
rect 183758 168800 183763 168856
rect 179820 168798 183763 168800
rect 99425 168795 99491 168798
rect 183697 168795 183763 168798
rect 44409 168722 44475 168725
rect 41820 168720 44475 168722
rect 41820 168664 44414 168720
rect 44470 168664 44475 168720
rect 41820 168662 44475 168664
rect 44409 168659 44475 168662
rect 191977 168722 192043 168725
rect 191977 168720 193988 168722
rect 191977 168664 191982 168720
rect 192038 168664 193988 168720
rect 191977 168662 193988 168664
rect 191977 168659 192043 168662
rect 99517 167770 99583 167773
rect 183789 167770 183855 167773
rect 95732 167768 99583 167770
rect 95732 167712 99522 167768
rect 99578 167712 99583 167768
rect 95732 167710 99583 167712
rect 179820 167768 183855 167770
rect 179820 167712 183794 167768
rect 183850 167712 183855 167768
rect 179820 167710 183855 167712
rect 99517 167707 99583 167710
rect 183789 167707 183855 167710
rect 191885 166818 191951 166821
rect 191885 166816 193988 166818
rect 191885 166760 191890 166816
rect 191946 166760 193988 166816
rect 191885 166758 193988 166760
rect 191885 166755 191951 166758
rect 106693 166682 106759 166685
rect 106693 166680 109900 166682
rect 106693 166624 106698 166680
rect 106754 166624 109900 166680
rect 106693 166622 109900 166624
rect 106693 166619 106759 166622
rect 99517 166546 99583 166549
rect 182869 166546 182935 166549
rect 95732 166544 99583 166546
rect 95732 166488 99522 166544
rect 99578 166488 99583 166544
rect 95732 166486 99583 166488
rect 179820 166544 182935 166546
rect 179820 166488 182874 166544
rect 182930 166488 182935 166544
rect 179820 166486 182935 166488
rect 99517 166483 99583 166486
rect 182869 166483 182935 166486
rect 99517 165322 99583 165325
rect 183697 165322 183763 165325
rect 95732 165320 99583 165322
rect 95732 165264 99522 165320
rect 99578 165264 99583 165320
rect 95732 165262 99583 165264
rect 179820 165320 183763 165322
rect 179820 165264 183702 165320
rect 183758 165264 183763 165320
rect 179820 165262 183763 165264
rect 99517 165259 99583 165262
rect 183697 165259 183763 165262
rect 212534 164852 212540 164916
rect 212604 164914 212610 164916
rect 212677 164914 212743 164917
rect 212604 164912 212743 164914
rect 212604 164856 212682 164912
rect 212738 164856 212743 164912
rect 212604 164854 212743 164856
rect 212604 164852 212610 164854
rect 212677 164851 212743 164854
rect 138157 164778 138223 164781
rect 139486 164778 139492 164780
rect 138157 164776 139492 164778
rect 138157 164720 138162 164776
rect 138218 164720 139492 164776
rect 138157 164718 139492 164720
rect 138157 164715 138223 164718
rect 139486 164716 139492 164718
rect 139556 164716 139562 164780
rect 191333 164778 191399 164781
rect 191333 164776 193988 164778
rect 191333 164720 191338 164776
rect 191394 164720 193988 164776
rect 191333 164718 193988 164720
rect 191333 164715 191399 164718
rect 106785 164370 106851 164373
rect 106785 164368 109900 164370
rect 106785 164312 106790 164368
rect 106846 164312 109900 164368
rect 106785 164310 109900 164312
rect 106785 164307 106851 164310
rect 99517 164098 99583 164101
rect 183053 164098 183119 164101
rect 95732 164096 99583 164098
rect 95732 164040 99522 164096
rect 99578 164040 99583 164096
rect 95732 164038 99583 164040
rect 179820 164096 183119 164098
rect 179820 164040 183058 164096
rect 183114 164040 183119 164096
rect 179820 164038 183119 164040
rect 99517 164035 99583 164038
rect 183053 164035 183119 164038
rect 25774 163628 25780 163692
rect 25844 163690 25850 163692
rect 25966 163690 26026 163796
rect 41782 163764 41788 163828
rect 41852 163826 41858 163828
rect 53333 163826 53399 163829
rect 128497 163826 128563 163829
rect 211757 163826 211823 163829
rect 41852 163824 53399 163826
rect 41852 163768 53338 163824
rect 53394 163768 53399 163824
rect 41852 163766 53399 163768
rect 125724 163824 128563 163826
rect 125724 163768 128502 163824
rect 128558 163768 128563 163824
rect 125724 163766 128563 163768
rect 209812 163824 211823 163826
rect 209812 163768 211762 163824
rect 211818 163768 211823 163824
rect 209812 163766 211823 163768
rect 41852 163764 41858 163766
rect 53333 163763 53399 163766
rect 128497 163763 128563 163766
rect 211757 163763 211823 163766
rect 25844 163630 26026 163690
rect 25844 163628 25850 163630
rect 98965 162874 99031 162877
rect 183053 162874 183119 162877
rect 95732 162872 99031 162874
rect 95732 162816 98970 162872
rect 99026 162816 99031 162872
rect 95732 162814 99031 162816
rect 179820 162872 183119 162874
rect 179820 162816 183058 162872
rect 183114 162816 183119 162872
rect 179820 162814 183119 162816
rect 98965 162811 99031 162814
rect 183053 162811 183119 162814
rect 191977 162738 192043 162741
rect 191977 162736 193988 162738
rect 191977 162680 191982 162736
rect 192038 162680 193988 162736
rect 191977 162678 193988 162680
rect 191977 162675 192043 162678
rect 9896 162194 10376 162224
rect 13405 162194 13471 162197
rect 9896 162192 13471 162194
rect 9896 162136 13410 162192
rect 13466 162136 13471 162192
rect 9896 162134 13471 162136
rect 9896 162104 10376 162134
rect 13405 162131 13471 162134
rect 106877 161922 106943 161925
rect 106877 161920 109900 161922
rect 106877 161864 106882 161920
rect 106938 161864 109900 161920
rect 106877 161862 109900 161864
rect 106877 161859 106943 161862
rect 99057 161650 99123 161653
rect 183145 161650 183211 161653
rect 95732 161648 99123 161650
rect 95732 161592 99062 161648
rect 99118 161592 99123 161648
rect 95732 161590 99123 161592
rect 179820 161648 183211 161650
rect 179820 161592 183150 161648
rect 183206 161592 183211 161648
rect 179820 161590 183211 161592
rect 99057 161587 99123 161590
rect 183145 161587 183211 161590
rect 191333 160834 191399 160837
rect 191333 160832 193988 160834
rect 191333 160776 191338 160832
rect 191394 160776 193988 160832
rect 191333 160774 193988 160776
rect 191333 160771 191399 160774
rect 53425 160562 53491 160565
rect 138157 160562 138223 160565
rect 53425 160560 55988 160562
rect 53425 160504 53430 160560
rect 53486 160504 55988 160560
rect 53425 160502 55988 160504
rect 138157 160560 140076 160562
rect 138157 160504 138162 160560
rect 138218 160504 140076 160560
rect 138157 160502 140076 160504
rect 53425 160499 53491 160502
rect 138157 160499 138223 160502
rect 99149 160426 99215 160429
rect 183237 160426 183303 160429
rect 95732 160424 99215 160426
rect 95732 160368 99154 160424
rect 99210 160368 99215 160424
rect 95732 160366 99215 160368
rect 179820 160424 183303 160426
rect 179820 160368 183242 160424
rect 183298 160368 183303 160424
rect 179820 160366 183303 160368
rect 99149 160363 99215 160366
rect 183237 160363 183303 160366
rect 107245 159610 107311 159613
rect 107245 159608 109900 159610
rect 107245 159552 107250 159608
rect 107306 159552 109900 159608
rect 107245 159550 109900 159552
rect 107245 159547 107311 159550
rect 99241 159202 99307 159205
rect 183329 159202 183395 159205
rect 95732 159200 99307 159202
rect 95732 159144 99246 159200
rect 99302 159144 99307 159200
rect 95732 159142 99307 159144
rect 179820 159200 183395 159202
rect 179820 159144 183334 159200
rect 183390 159144 183395 159200
rect 179820 159142 183395 159144
rect 99241 159139 99307 159142
rect 183329 159139 183395 159142
rect 44501 158794 44567 158797
rect 41820 158792 44567 158794
rect 41820 158736 44506 158792
rect 44562 158736 44567 158792
rect 41820 158734 44567 158736
rect 44501 158731 44567 158734
rect 190045 158794 190111 158797
rect 190045 158792 193988 158794
rect 190045 158736 190050 158792
rect 190106 158736 193988 158792
rect 190045 158734 193988 158736
rect 190045 158731 190111 158734
rect 99425 157978 99491 157981
rect 183513 157978 183579 157981
rect 95732 157976 99491 157978
rect 95732 157920 99430 157976
rect 99486 157920 99491 157976
rect 95732 157918 99491 157920
rect 179820 157976 183579 157978
rect 179820 157920 183518 157976
rect 183574 157920 183579 157976
rect 179820 157918 183579 157920
rect 99425 157915 99491 157918
rect 183513 157915 183579 157918
rect 107153 157298 107219 157301
rect 107153 157296 109900 157298
rect 107153 157240 107158 157296
rect 107214 157240 109900 157296
rect 107153 157238 109900 157240
rect 107153 157235 107219 157238
rect 23566 157100 23572 157164
rect 23636 157162 23642 157164
rect 211941 157162 212007 157165
rect 23636 157102 25996 157162
rect 209812 157160 212007 157162
rect 209812 157104 211946 157160
rect 212002 157104 212007 157160
rect 209812 157102 212007 157104
rect 23636 157100 23642 157102
rect 211941 157099 212007 157102
rect 99333 156754 99399 156757
rect 183421 156754 183487 156757
rect 95732 156752 99399 156754
rect 95732 156696 99338 156752
rect 99394 156696 99399 156752
rect 95732 156694 99399 156696
rect 179820 156752 183487 156754
rect 179820 156696 183426 156752
rect 183482 156696 183487 156752
rect 179820 156694 183487 156696
rect 99333 156691 99399 156694
rect 183421 156691 183487 156694
rect 189953 156754 190019 156757
rect 189953 156752 193988 156754
rect 189953 156696 189958 156752
rect 190014 156696 193988 156752
rect 189953 156694 193988 156696
rect 189953 156691 190019 156694
rect 99517 155530 99583 155533
rect 182685 155530 182751 155533
rect 95732 155528 99583 155530
rect 95732 155472 99522 155528
rect 99578 155472 99583 155528
rect 95732 155470 99583 155472
rect 179820 155528 182751 155530
rect 179820 155472 182690 155528
rect 182746 155472 182751 155528
rect 179820 155470 182751 155472
rect 99517 155467 99583 155470
rect 182685 155467 182751 155470
rect 106509 154986 106575 154989
rect 106509 154984 109900 154986
rect 106509 154928 106514 154984
rect 106570 154928 109900 154984
rect 106509 154926 109900 154928
rect 106509 154923 106575 154926
rect 191977 154850 192043 154853
rect 191977 154848 193988 154850
rect 191977 154792 191982 154848
rect 192038 154792 193988 154848
rect 191977 154790 193988 154792
rect 191977 154787 192043 154790
rect 98781 154442 98847 154445
rect 183605 154442 183671 154445
rect 95732 154440 98847 154442
rect 95732 154384 98786 154440
rect 98842 154384 98847 154440
rect 95732 154382 98847 154384
rect 179820 154440 183671 154442
rect 179820 154384 183610 154440
rect 183666 154384 183671 154440
rect 179820 154382 183671 154384
rect 98781 154379 98847 154382
rect 183605 154379 183671 154382
rect 221693 152946 221759 152949
rect 225416 152946 225896 152976
rect 221693 152944 225896 152946
rect 221693 152888 221698 152944
rect 221754 152888 225896 152944
rect 221693 152886 225896 152888
rect 221693 152883 221759 152886
rect 225416 152856 225896 152886
rect 134845 140570 134911 140573
rect 131796 140568 134911 140570
rect 47862 140434 47922 140540
rect 131796 140512 134850 140568
rect 134906 140512 134911 140568
rect 131796 140510 134911 140512
rect 134845 140507 134911 140510
rect 51401 140434 51467 140437
rect 47862 140432 51467 140434
rect 47862 140376 51406 140432
rect 51462 140376 51467 140432
rect 47862 140374 51467 140376
rect 51401 140371 51467 140374
rect 49929 140162 49995 140165
rect 47678 140160 49995 140162
rect 47678 140104 49934 140160
rect 49990 140104 49995 140160
rect 47678 140102 49995 140104
rect 47678 139996 47738 140102
rect 49929 140099 49995 140102
rect 100805 140162 100871 140165
rect 103982 140162 104042 140472
rect 100805 140160 104042 140162
rect 100805 140104 100810 140160
rect 100866 140104 104042 140160
rect 100805 140102 104042 140104
rect 184985 140162 185051 140165
rect 187886 140162 187946 140540
rect 184985 140160 187946 140162
rect 184985 140104 184990 140160
rect 185046 140104 187946 140160
rect 184985 140102 187946 140104
rect 100805 140099 100871 140102
rect 184985 140099 185051 140102
rect 100897 140026 100963 140029
rect 135397 140026 135463 140029
rect 100897 140024 104012 140026
rect 100897 139968 100902 140024
rect 100958 139968 104012 140024
rect 100897 139966 104012 139968
rect 131796 140024 135463 140026
rect 131796 139968 135402 140024
rect 135458 139968 135463 140024
rect 131796 139966 135463 139968
rect 100897 139963 100963 139966
rect 135397 139963 135463 139966
rect 185077 140026 185143 140029
rect 185077 140024 187762 140026
rect 185077 139968 185082 140024
rect 185138 139968 187762 140024
rect 185077 139966 187762 139968
rect 185077 139963 185143 139966
rect 187702 139890 187762 139966
rect 187886 139890 187946 139996
rect 187702 139830 187946 139890
rect 134661 139482 134727 139485
rect 131796 139480 134727 139482
rect 47862 139074 47922 139452
rect 131796 139424 134666 139480
rect 134722 139424 134727 139480
rect 131796 139422 134727 139424
rect 134661 139419 134727 139422
rect 50021 139074 50087 139077
rect 47862 139072 50087 139074
rect 47862 139016 50026 139072
rect 50082 139016 50087 139072
rect 47862 139014 50087 139016
rect 50021 139011 50087 139014
rect 101173 138938 101239 138941
rect 103982 138938 104042 139384
rect 101173 138936 104042 138938
rect 101173 138880 101178 138936
rect 101234 138880 104042 138936
rect 101173 138878 104042 138880
rect 185353 138938 185419 138941
rect 187886 138938 187946 139452
rect 185353 138936 187946 138938
rect 185353 138880 185358 138936
rect 185414 138880 187946 138936
rect 185353 138878 187946 138880
rect 101173 138875 101239 138878
rect 185353 138875 185419 138878
rect 135397 138802 135463 138805
rect 131796 138800 135463 138802
rect 47862 138666 47922 138772
rect 131796 138744 135402 138800
rect 135458 138744 135463 138800
rect 131796 138742 135463 138744
rect 135397 138739 135463 138742
rect 103614 138674 104012 138734
rect 49929 138666 49995 138669
rect 47862 138664 49995 138666
rect 47862 138608 49934 138664
rect 49990 138608 49995 138664
rect 47862 138606 49995 138608
rect 49929 138603 49995 138606
rect 101081 138666 101147 138669
rect 103614 138666 103674 138674
rect 101081 138664 103674 138666
rect 101081 138608 101086 138664
rect 101142 138608 103674 138664
rect 101081 138606 103674 138608
rect 185261 138666 185327 138669
rect 187886 138666 187946 138772
rect 185261 138664 187946 138666
rect 185261 138608 185266 138664
rect 185322 138608 187946 138664
rect 185261 138606 187946 138608
rect 101081 138603 101147 138606
rect 185261 138603 185327 138606
rect 9896 138530 10376 138560
rect 13313 138530 13379 138533
rect 9896 138528 13379 138530
rect 9896 138472 13318 138528
rect 13374 138472 13379 138528
rect 9896 138470 13379 138472
rect 9896 138440 10376 138470
rect 13313 138467 13379 138470
rect 59221 138530 59287 138533
rect 92709 138530 92775 138533
rect 59221 138528 60986 138530
rect 59221 138472 59226 138528
rect 59282 138472 60986 138528
rect 59221 138470 60986 138472
rect 59221 138467 59287 138470
rect 60926 138364 60986 138470
rect 90734 138528 92775 138530
rect 90734 138472 92714 138528
rect 92770 138472 92775 138528
rect 90734 138470 92775 138472
rect 90734 138432 90794 138470
rect 92709 138467 92775 138470
rect 143585 138530 143651 138533
rect 177717 138530 177783 138533
rect 143585 138528 145074 138530
rect 143585 138472 143590 138528
rect 143646 138472 145074 138528
rect 143585 138470 145074 138472
rect 143585 138467 143651 138470
rect 145014 138432 145074 138470
rect 174822 138528 177783 138530
rect 174822 138472 177722 138528
rect 177778 138472 177783 138528
rect 174822 138470 177783 138472
rect 174822 138364 174882 138470
rect 177717 138467 177783 138470
rect 58669 138258 58735 138261
rect 134661 138258 134727 138261
rect 58669 138256 60986 138258
rect 47862 137850 47922 138228
rect 58669 138200 58674 138256
rect 58730 138200 60986 138256
rect 58669 138198 60986 138200
rect 131796 138256 134727 138258
rect 131796 138200 134666 138256
rect 134722 138200 134727 138256
rect 131796 138198 134727 138200
rect 58669 138195 58735 138198
rect 50021 137850 50087 137853
rect 47862 137848 50087 137850
rect 47862 137792 50026 137848
rect 50082 137792 50087 137848
rect 60926 137820 60986 138198
rect 134661 138195 134727 138198
rect 143309 138258 143375 138261
rect 177625 138258 177691 138261
rect 143309 138256 145074 138258
rect 143309 138200 143314 138256
rect 143370 138200 145074 138256
rect 143309 138198 145074 138200
rect 143309 138195 143375 138198
rect 92801 138122 92867 138125
rect 90734 138120 92867 138122
rect 90734 138064 92806 138120
rect 92862 138064 92867 138120
rect 90734 138062 92867 138064
rect 90734 137888 90794 138062
rect 92801 138059 92867 138062
rect 100989 137850 101055 137853
rect 103982 137850 104042 138160
rect 145014 137888 145074 138198
rect 174822 138256 177691 138258
rect 174822 138200 177630 138256
rect 177686 138200 177691 138256
rect 174822 138198 177691 138200
rect 100989 137848 104042 137850
rect 47862 137790 50087 137792
rect 50021 137787 50087 137790
rect 100989 137792 100994 137848
rect 101050 137792 104042 137848
rect 174822 137820 174882 138198
rect 177625 138195 177691 138198
rect 185169 137850 185235 137853
rect 187886 137850 187946 138228
rect 185169 137848 187946 137850
rect 100989 137790 104042 137792
rect 185169 137792 185174 137848
rect 185230 137792 187946 137848
rect 185169 137790 187946 137792
rect 100989 137787 101055 137790
rect 185169 137787 185235 137790
rect 135397 137714 135463 137717
rect 131796 137712 135463 137714
rect 47862 137442 47922 137684
rect 131796 137656 135402 137712
rect 135458 137656 135463 137712
rect 131796 137654 135463 137656
rect 135397 137651 135463 137654
rect 49929 137442 49995 137445
rect 47862 137440 49995 137442
rect 47862 137384 49934 137440
rect 49990 137384 49995 137440
rect 47862 137382 49995 137384
rect 49929 137379 49995 137382
rect 101265 137306 101331 137309
rect 103982 137306 104042 137616
rect 101265 137304 104042 137306
rect 101265 137248 101270 137304
rect 101326 137248 104042 137304
rect 101265 137246 104042 137248
rect 185445 137306 185511 137309
rect 187886 137306 187946 137684
rect 185445 137304 187946 137306
rect 185445 137248 185450 137304
rect 185506 137248 187946 137304
rect 185445 137246 187946 137248
rect 101265 137243 101331 137246
rect 185445 137243 185511 137246
rect 58393 137170 58459 137173
rect 92709 137170 92775 137173
rect 58393 137168 60956 137170
rect 58393 137112 58398 137168
rect 58454 137112 60956 137168
rect 58393 137110 60956 137112
rect 90764 137168 92775 137170
rect 90764 137112 92714 137168
rect 92770 137112 92775 137168
rect 90764 137110 92775 137112
rect 58393 137107 58459 137110
rect 92709 137107 92775 137110
rect 143585 137170 143651 137173
rect 143585 137168 145044 137170
rect 143585 137112 143590 137168
rect 143646 137112 145044 137168
rect 143585 137110 145044 137112
rect 143585 137107 143651 137110
rect 135029 137034 135095 137037
rect 131796 137032 135095 137034
rect 47862 136626 47922 137004
rect 131796 136976 135034 137032
rect 135090 136976 135095 137032
rect 131796 136974 135095 136976
rect 174822 137034 174882 137140
rect 177717 137034 177783 137037
rect 174822 137032 177783 137034
rect 174822 136976 177722 137032
rect 177778 136976 177783 137032
rect 174822 136974 177783 136976
rect 135029 136971 135095 136974
rect 177717 136971 177783 136974
rect 92801 136898 92867 136901
rect 90734 136896 92867 136898
rect 90734 136840 92806 136896
rect 92862 136840 92867 136896
rect 90734 136838 92867 136840
rect 90734 136664 90794 136838
rect 92801 136835 92867 136838
rect 50389 136626 50455 136629
rect 47862 136624 50455 136626
rect 47862 136568 50394 136624
rect 50450 136568 50455 136624
rect 47862 136566 50455 136568
rect 50389 136563 50455 136566
rect 58485 136626 58551 136629
rect 101817 136626 101883 136629
rect 103982 136626 104042 136936
rect 143125 136898 143191 136901
rect 177625 136898 177691 136901
rect 143125 136896 145074 136898
rect 143125 136840 143130 136896
rect 143186 136840 145074 136896
rect 143125 136838 145074 136840
rect 143125 136835 143191 136838
rect 145014 136664 145074 136838
rect 174822 136896 177691 136898
rect 174822 136840 177630 136896
rect 177686 136840 177691 136896
rect 174822 136838 177691 136840
rect 58485 136624 60956 136626
rect 58485 136568 58490 136624
rect 58546 136568 60956 136624
rect 58485 136566 60956 136568
rect 101817 136624 104042 136626
rect 101817 136568 101822 136624
rect 101878 136568 104042 136624
rect 174822 136596 174882 136838
rect 177625 136835 177691 136838
rect 185169 136626 185235 136629
rect 187886 136626 187946 137004
rect 185169 136624 187946 136626
rect 101817 136566 104042 136568
rect 185169 136568 185174 136624
rect 185230 136568 187946 136624
rect 185169 136566 187946 136568
rect 58485 136563 58551 136566
rect 101817 136563 101883 136566
rect 185169 136563 185235 136566
rect 92709 136490 92775 136493
rect 135305 136490 135371 136493
rect 90734 136488 92775 136490
rect 47862 136218 47922 136460
rect 90734 136432 92714 136488
rect 92770 136432 92775 136488
rect 90734 136430 92775 136432
rect 131796 136488 135371 136490
rect 131796 136432 135310 136488
rect 135366 136432 135371 136488
rect 131796 136430 135371 136432
rect 51217 136218 51283 136221
rect 47862 136216 51283 136218
rect 18097 135946 18163 135949
rect 19894 135946 19954 136188
rect 47862 136160 51222 136216
rect 51278 136160 51283 136216
rect 47862 136158 51283 136160
rect 51217 136155 51283 136158
rect 90734 136120 90794 136430
rect 92709 136427 92775 136430
rect 135305 136427 135371 136430
rect 101449 136218 101515 136221
rect 103982 136218 104042 136392
rect 143493 136354 143559 136357
rect 177717 136354 177783 136357
rect 143493 136352 145074 136354
rect 143493 136296 143498 136352
rect 143554 136296 145074 136352
rect 143493 136294 145074 136296
rect 143493 136291 143559 136294
rect 101449 136216 104042 136218
rect 101449 136160 101454 136216
rect 101510 136160 104042 136216
rect 101449 136158 104042 136160
rect 101449 136155 101515 136158
rect 145014 136120 145074 136294
rect 174822 136352 177783 136354
rect 174822 136296 177722 136352
rect 177778 136296 177783 136352
rect 174822 136294 177783 136296
rect 51217 136082 51283 136085
rect 18097 135944 19954 135946
rect 18097 135888 18102 135944
rect 18158 135888 19954 135944
rect 47678 136080 51283 136082
rect 47678 136024 51222 136080
rect 51278 136024 51283 136080
rect 47678 136022 51283 136024
rect 47678 135916 47738 136022
rect 51217 136019 51283 136022
rect 58209 136082 58275 136085
rect 58209 136080 60956 136082
rect 58209 136024 58214 136080
rect 58270 136024 60956 136080
rect 174822 136052 174882 136294
rect 177717 136291 177783 136294
rect 185261 136082 185327 136085
rect 187886 136082 187946 136460
rect 185261 136080 187946 136082
rect 58209 136022 60956 136024
rect 185261 136024 185266 136080
rect 185322 136024 187946 136080
rect 185261 136022 187946 136024
rect 58209 136019 58275 136022
rect 185261 136019 185327 136022
rect 101725 135946 101791 135949
rect 135397 135946 135463 135949
rect 101725 135944 104012 135946
rect 18097 135886 19954 135888
rect 101725 135888 101730 135944
rect 101786 135888 104012 135944
rect 101725 135886 104012 135888
rect 131796 135944 135463 135946
rect 131796 135888 135402 135944
rect 135458 135888 135463 135944
rect 131796 135886 135463 135888
rect 18097 135883 18163 135886
rect 101725 135883 101791 135886
rect 135397 135883 135463 135886
rect 185353 135946 185419 135949
rect 215854 135946 215914 136188
rect 218381 135946 218447 135949
rect 185353 135944 187762 135946
rect 185353 135888 185358 135944
rect 185414 135888 187762 135944
rect 215854 135944 218447 135946
rect 185353 135886 187762 135888
rect 185353 135883 185419 135886
rect 143401 135810 143467 135813
rect 187702 135810 187762 135886
rect 187886 135810 187946 135916
rect 215854 135888 218386 135944
rect 218442 135888 218447 135944
rect 215854 135886 218447 135888
rect 218381 135883 218447 135886
rect 143401 135808 145074 135810
rect 143401 135752 143406 135808
rect 143462 135752 145074 135808
rect 143401 135750 145074 135752
rect 187702 135750 187946 135810
rect 143401 135747 143467 135750
rect 92709 135538 92775 135541
rect 90734 135536 92775 135538
rect 90734 135480 92714 135536
rect 92770 135480 92775 135536
rect 90734 135478 92775 135480
rect 90734 135440 90794 135478
rect 92709 135475 92775 135478
rect 145014 135440 145074 135750
rect 177717 135538 177783 135541
rect 174822 135536 177783 135538
rect 174822 135480 177722 135536
rect 177778 135480 177783 135536
rect 174822 135478 177783 135480
rect 58301 135402 58367 135405
rect 134845 135402 134911 135405
rect 58301 135400 60956 135402
rect 47862 134994 47922 135372
rect 58301 135344 58306 135400
rect 58362 135344 60956 135400
rect 58301 135342 60956 135344
rect 131796 135400 134911 135402
rect 131796 135344 134850 135400
rect 134906 135344 134911 135400
rect 174822 135372 174882 135478
rect 177717 135475 177783 135478
rect 131796 135342 134911 135344
rect 58301 135339 58367 135342
rect 134845 135339 134911 135342
rect 92801 135266 92867 135269
rect 90734 135264 92867 135266
rect 90734 135208 92806 135264
rect 92862 135208 92867 135264
rect 90734 135206 92867 135208
rect 51217 134994 51283 134997
rect 47862 134992 51283 134994
rect 47862 134936 51222 134992
rect 51278 134936 51283 134992
rect 47862 134934 51283 134936
rect 51217 134931 51283 134934
rect 90734 134896 90794 135206
rect 92801 135203 92867 135206
rect 58209 134858 58275 134861
rect 101449 134858 101515 134861
rect 103982 134858 104042 135304
rect 143309 135266 143375 135269
rect 177625 135266 177691 135269
rect 143309 135264 145074 135266
rect 143309 135208 143314 135264
rect 143370 135208 145074 135264
rect 143309 135206 145074 135208
rect 143309 135203 143375 135206
rect 145014 134896 145074 135206
rect 174822 135264 177691 135266
rect 174822 135208 177630 135264
rect 177686 135208 177691 135264
rect 174822 135206 177691 135208
rect 58209 134856 60956 134858
rect 58209 134800 58214 134856
rect 58270 134800 60956 134856
rect 58209 134798 60956 134800
rect 101449 134856 104042 134858
rect 101449 134800 101454 134856
rect 101510 134800 104042 134856
rect 174822 134828 174882 135206
rect 177625 135203 177691 135206
rect 185169 134858 185235 134861
rect 187886 134858 187946 135372
rect 185169 134856 187946 134858
rect 101449 134798 104042 134800
rect 185169 134800 185174 134856
rect 185230 134800 187946 134856
rect 185169 134798 187946 134800
rect 58209 134795 58275 134798
rect 101449 134795 101515 134798
rect 185169 134795 185235 134798
rect 134661 134722 134727 134725
rect 131796 134720 134727 134722
rect 47862 134586 47922 134692
rect 131796 134664 134666 134720
rect 134722 134664 134727 134720
rect 131796 134662 134727 134664
rect 134661 134659 134727 134662
rect 51125 134586 51191 134589
rect 47862 134584 51191 134586
rect 47862 134528 51130 134584
rect 51186 134528 51191 134584
rect 47862 134526 51191 134528
rect 51125 134523 51191 134526
rect 100897 134450 100963 134453
rect 103982 134450 104042 134624
rect 100897 134448 104042 134450
rect 100897 134392 100902 134448
rect 100958 134392 104042 134448
rect 100897 134390 104042 134392
rect 185077 134450 185143 134453
rect 187886 134450 187946 134692
rect 185077 134448 187946 134450
rect 185077 134392 185082 134448
rect 185138 134392 187946 134448
rect 185077 134390 187946 134392
rect 100897 134387 100963 134390
rect 185077 134387 185143 134390
rect 92709 134314 92775 134317
rect 90734 134312 92775 134314
rect 90734 134256 92714 134312
rect 92770 134256 92775 134312
rect 90734 134254 92775 134256
rect 90734 134216 90794 134254
rect 92709 134251 92775 134254
rect 143585 134314 143651 134317
rect 177717 134314 177783 134317
rect 143585 134312 145074 134314
rect 143585 134256 143590 134312
rect 143646 134256 145074 134312
rect 143585 134254 145074 134256
rect 143585 134251 143651 134254
rect 145014 134216 145074 134254
rect 174822 134312 177783 134314
rect 174822 134256 177722 134312
rect 177778 134256 177783 134312
rect 174822 134254 177783 134256
rect 58209 134178 58275 134181
rect 135397 134178 135463 134181
rect 58209 134176 60956 134178
rect 47862 133770 47922 134148
rect 58209 134120 58214 134176
rect 58270 134120 60956 134176
rect 58209 134118 60956 134120
rect 131796 134176 135463 134178
rect 131796 134120 135402 134176
rect 135458 134120 135463 134176
rect 174822 134148 174882 134254
rect 177717 134251 177783 134254
rect 131796 134118 135463 134120
rect 58209 134115 58275 134118
rect 135397 134115 135463 134118
rect 92801 133906 92867 133909
rect 90734 133904 92867 133906
rect 90734 133848 92806 133904
rect 92862 133848 92867 133904
rect 90734 133846 92867 133848
rect 50205 133770 50271 133773
rect 47862 133768 50271 133770
rect 47862 133712 50210 133768
rect 50266 133712 50271 133768
rect 47862 133710 50271 133712
rect 50205 133707 50271 133710
rect 90734 133672 90794 133846
rect 92801 133843 92867 133846
rect 101817 133770 101883 133773
rect 103982 133770 104042 134080
rect 143217 134042 143283 134045
rect 143217 134040 145074 134042
rect 143217 133984 143222 134040
rect 143278 133984 145074 134040
rect 143217 133982 145074 133984
rect 143217 133979 143283 133982
rect 101817 133768 104042 133770
rect 101817 133712 101822 133768
rect 101878 133712 104042 133768
rect 101817 133710 104042 133712
rect 101817 133707 101883 133710
rect 145014 133672 145074 133982
rect 177717 133906 177783 133909
rect 174822 133904 177783 133906
rect 174822 133848 177722 133904
rect 177778 133848 177783 133904
rect 174822 133846 177783 133848
rect 58301 133634 58367 133637
rect 134109 133634 134175 133637
rect 58301 133632 60956 133634
rect 47862 133226 47922 133604
rect 58301 133576 58306 133632
rect 58362 133576 60956 133632
rect 58301 133574 60956 133576
rect 131796 133632 134175 133634
rect 131796 133576 134114 133632
rect 134170 133576 134175 133632
rect 174822 133604 174882 133846
rect 177717 133843 177783 133846
rect 185169 133770 185235 133773
rect 187886 133770 187946 134148
rect 185169 133768 187946 133770
rect 185169 133712 185174 133768
rect 185230 133712 187946 133768
rect 185169 133710 187946 133712
rect 185169 133707 185235 133710
rect 131796 133574 134175 133576
rect 58301 133571 58367 133574
rect 134109 133571 134175 133574
rect 92893 133498 92959 133501
rect 90734 133496 92959 133498
rect 90734 133440 92898 133496
rect 92954 133440 92959 133496
rect 90734 133438 92959 133440
rect 50941 133226 51007 133229
rect 47862 133224 51007 133226
rect 47862 133168 50946 133224
rect 51002 133168 51007 133224
rect 47862 133166 51007 133168
rect 50941 133163 51007 133166
rect 90734 133128 90794 133438
rect 92893 133435 92959 133438
rect 58209 133090 58275 133093
rect 101725 133090 101791 133093
rect 103982 133090 104042 133536
rect 177625 133498 177691 133501
rect 174822 133496 177691 133498
rect 174822 133440 177630 133496
rect 177686 133440 177691 133496
rect 174822 133438 177691 133440
rect 142941 133362 143007 133365
rect 142941 133360 145074 133362
rect 142941 133304 142946 133360
rect 143002 133304 145074 133360
rect 142941 133302 145074 133304
rect 142941 133299 143007 133302
rect 145014 133128 145074 133302
rect 58209 133088 60956 133090
rect 58209 133032 58214 133088
rect 58270 133032 60956 133088
rect 58209 133030 60956 133032
rect 101725 133088 104042 133090
rect 101725 133032 101730 133088
rect 101786 133032 104042 133088
rect 174822 133060 174882 133438
rect 177625 133435 177691 133438
rect 185813 133090 185879 133093
rect 187886 133090 187946 133604
rect 185813 133088 187946 133090
rect 101725 133030 104042 133032
rect 185813 133032 185818 133088
rect 185874 133032 187946 133088
rect 185813 133030 187946 133032
rect 58209 133027 58275 133030
rect 101725 133027 101791 133030
rect 185813 133027 185879 133030
rect 135121 132954 135187 132957
rect 131796 132952 135187 132954
rect 47862 132546 47922 132924
rect 131796 132896 135126 132952
rect 135182 132896 135187 132952
rect 131796 132894 135187 132896
rect 135121 132891 135187 132894
rect 92709 132682 92775 132685
rect 90734 132680 92775 132682
rect 90734 132624 92714 132680
rect 92770 132624 92775 132680
rect 90734 132622 92775 132624
rect 51217 132546 51283 132549
rect 47862 132544 51283 132546
rect 47862 132488 51222 132544
rect 51278 132488 51283 132544
rect 47862 132486 51283 132488
rect 51217 132483 51283 132486
rect 90734 132448 90794 132622
rect 92709 132619 92775 132622
rect 101817 132546 101883 132549
rect 103982 132546 104042 132856
rect 143585 132818 143651 132821
rect 143585 132816 145074 132818
rect 143585 132760 143590 132816
rect 143646 132760 145074 132816
rect 143585 132758 145074 132760
rect 143585 132755 143651 132758
rect 101817 132544 104042 132546
rect 101817 132488 101822 132544
rect 101878 132488 104042 132544
rect 101817 132486 104042 132488
rect 101817 132483 101883 132486
rect 145014 132448 145074 132758
rect 177717 132682 177783 132685
rect 174822 132680 177783 132682
rect 174822 132624 177722 132680
rect 177778 132624 177783 132680
rect 174822 132622 177783 132624
rect 58209 132410 58275 132413
rect 134477 132410 134543 132413
rect 58209 132408 60956 132410
rect 47862 132138 47922 132380
rect 58209 132352 58214 132408
rect 58270 132352 60956 132408
rect 58209 132350 60956 132352
rect 131796 132408 134543 132410
rect 131796 132352 134482 132408
rect 134538 132352 134543 132408
rect 174822 132380 174882 132622
rect 177717 132619 177783 132622
rect 185905 132546 185971 132549
rect 187886 132546 187946 132924
rect 185905 132544 187946 132546
rect 185905 132488 185910 132544
rect 185966 132488 187946 132544
rect 185905 132486 187946 132488
rect 185905 132483 185971 132486
rect 131796 132350 134543 132352
rect 58209 132347 58275 132350
rect 134477 132347 134543 132350
rect 92801 132274 92867 132277
rect 90734 132272 92867 132274
rect 90734 132216 92806 132272
rect 92862 132216 92867 132272
rect 90734 132214 92867 132216
rect 50389 132138 50455 132141
rect 47862 132136 50455 132138
rect 47862 132080 50394 132136
rect 50450 132080 50455 132136
rect 47862 132078 50455 132080
rect 50389 132075 50455 132078
rect 90734 131904 90794 132214
rect 92801 132211 92867 132214
rect 101173 132002 101239 132005
rect 103982 132002 104042 132312
rect 143217 132274 143283 132277
rect 177625 132274 177691 132277
rect 143217 132272 145074 132274
rect 143217 132216 143222 132272
rect 143278 132216 145074 132272
rect 143217 132214 145074 132216
rect 143217 132211 143283 132214
rect 101173 132000 104042 132002
rect 101173 131944 101178 132000
rect 101234 131944 104042 132000
rect 101173 131942 104042 131944
rect 101173 131939 101239 131942
rect 145014 131904 145074 132214
rect 174822 132272 177691 132274
rect 174822 132216 177630 132272
rect 177686 132216 177691 132272
rect 174822 132214 177691 132216
rect 58301 131866 58367 131869
rect 101541 131866 101607 131869
rect 135305 131866 135371 131869
rect 58301 131864 60956 131866
rect 47862 131730 47922 131836
rect 58301 131808 58306 131864
rect 58362 131808 60956 131864
rect 58301 131806 60956 131808
rect 101541 131864 104012 131866
rect 101541 131808 101546 131864
rect 101602 131808 104012 131864
rect 101541 131806 104012 131808
rect 131796 131864 135371 131866
rect 131796 131808 135310 131864
rect 135366 131808 135371 131864
rect 174822 131836 174882 132214
rect 177625 132211 177691 132214
rect 185721 132002 185787 132005
rect 187886 132002 187946 132380
rect 185721 132000 187946 132002
rect 185721 131944 185726 132000
rect 185782 131944 187946 132000
rect 185721 131942 187946 131944
rect 185721 131939 185787 131942
rect 131796 131806 135371 131808
rect 58301 131803 58367 131806
rect 101541 131803 101607 131806
rect 135305 131803 135371 131806
rect 51217 131730 51283 131733
rect 47862 131728 51283 131730
rect 47862 131672 51222 131728
rect 51278 131672 51283 131728
rect 47862 131670 51283 131672
rect 51217 131667 51283 131670
rect 185537 131730 185603 131733
rect 187886 131730 187946 131836
rect 185537 131728 187946 131730
rect 185537 131672 185542 131728
rect 185598 131672 187946 131728
rect 185537 131670 187946 131672
rect 185537 131667 185603 131670
rect 92709 131458 92775 131461
rect 90734 131456 92775 131458
rect 90734 131400 92714 131456
rect 92770 131400 92775 131456
rect 90734 131398 92775 131400
rect 47862 130778 47922 131292
rect 90734 131224 90794 131398
rect 92709 131395 92775 131398
rect 143585 131458 143651 131461
rect 143585 131456 145074 131458
rect 143585 131400 143590 131456
rect 143646 131400 145074 131456
rect 143585 131398 145074 131400
rect 143585 131395 143651 131398
rect 134845 131322 134911 131325
rect 131796 131320 134911 131322
rect 131796 131264 134850 131320
rect 134906 131264 134911 131320
rect 131796 131262 134911 131264
rect 134845 131259 134911 131262
rect 145014 131224 145074 131398
rect 177717 131322 177783 131325
rect 174822 131320 177783 131322
rect 174822 131264 177722 131320
rect 177778 131264 177783 131320
rect 174822 131262 177783 131264
rect 58209 131186 58275 131189
rect 58209 131184 60956 131186
rect 58209 131128 58214 131184
rect 58270 131128 60956 131184
rect 58209 131126 60956 131128
rect 58209 131123 58275 131126
rect 92801 131050 92867 131053
rect 90734 131048 92867 131050
rect 90734 130992 92806 131048
rect 92862 130992 92867 131048
rect 90734 130990 92867 130992
rect 51217 130778 51283 130781
rect 47862 130776 51283 130778
rect 47862 130720 51222 130776
rect 51278 130720 51283 130776
rect 47862 130718 51283 130720
rect 51217 130715 51283 130718
rect 90734 130680 90794 130990
rect 92801 130987 92867 130990
rect 101817 130778 101883 130781
rect 103982 130778 104042 131224
rect 174822 131156 174882 131262
rect 177717 131259 177783 131262
rect 142481 131050 142547 131053
rect 177625 131050 177691 131053
rect 142481 131048 145074 131050
rect 142481 130992 142486 131048
rect 142542 130992 145074 131048
rect 142481 130990 145074 130992
rect 142481 130987 142547 130990
rect 101817 130776 104042 130778
rect 101817 130720 101822 130776
rect 101878 130720 104042 130776
rect 101817 130718 104042 130720
rect 101817 130715 101883 130718
rect 145014 130680 145074 130990
rect 174822 131048 177691 131050
rect 174822 130992 177630 131048
rect 177686 130992 177691 131048
rect 174822 130990 177691 130992
rect 58301 130642 58367 130645
rect 134661 130642 134727 130645
rect 58301 130640 60956 130642
rect 47862 130370 47922 130612
rect 58301 130584 58306 130640
rect 58362 130584 60956 130640
rect 58301 130582 60956 130584
rect 131796 130640 134727 130642
rect 131796 130584 134666 130640
rect 134722 130584 134727 130640
rect 174822 130612 174882 130990
rect 177625 130987 177691 130990
rect 185353 130778 185419 130781
rect 187886 130778 187946 131292
rect 185353 130776 187946 130778
rect 185353 130720 185358 130776
rect 185414 130720 187946 130776
rect 185353 130718 187946 130720
rect 185353 130715 185419 130718
rect 131796 130582 134727 130584
rect 58301 130579 58367 130582
rect 134661 130579 134727 130582
rect 51217 130370 51283 130373
rect 47862 130368 51283 130370
rect 47862 130312 51222 130368
rect 51278 130312 51283 130368
rect 47862 130310 51283 130312
rect 51217 130307 51283 130310
rect 101357 130370 101423 130373
rect 103982 130370 104042 130544
rect 101357 130368 104042 130370
rect 101357 130312 101362 130368
rect 101418 130312 104042 130368
rect 101357 130310 104042 130312
rect 185261 130370 185327 130373
rect 187886 130370 187946 130612
rect 185261 130368 187946 130370
rect 185261 130312 185266 130368
rect 185322 130312 187946 130368
rect 185261 130310 187946 130312
rect 101357 130307 101423 130310
rect 185261 130307 185327 130310
rect 92709 130234 92775 130237
rect 90734 130232 92775 130234
rect 90734 130176 92714 130232
rect 92770 130176 92775 130232
rect 90734 130174 92775 130176
rect 90734 130136 90794 130174
rect 92709 130171 92775 130174
rect 143585 130234 143651 130237
rect 177717 130234 177783 130237
rect 143585 130232 145074 130234
rect 143585 130176 143590 130232
rect 143646 130176 145074 130232
rect 143585 130174 145074 130176
rect 143585 130171 143651 130174
rect 145014 130136 145074 130174
rect 174822 130232 177783 130234
rect 174822 130176 177722 130232
rect 177778 130176 177783 130232
rect 174822 130174 177783 130176
rect 58209 130098 58275 130101
rect 135397 130098 135463 130101
rect 58209 130096 60956 130098
rect 47862 129690 47922 130068
rect 58209 130040 58214 130096
rect 58270 130040 60956 130096
rect 58209 130038 60956 130040
rect 131796 130096 135463 130098
rect 131796 130040 135402 130096
rect 135458 130040 135463 130096
rect 174822 130068 174882 130174
rect 177717 130171 177783 130174
rect 131796 130038 135463 130040
rect 58209 130035 58275 130038
rect 135397 130035 135463 130038
rect 92801 129826 92867 129829
rect 90734 129824 92867 129826
rect 90734 129768 92806 129824
rect 92862 129768 92867 129824
rect 90734 129766 92867 129768
rect 50389 129690 50455 129693
rect 47862 129688 50455 129690
rect 47862 129632 50394 129688
rect 50450 129632 50455 129688
rect 47862 129630 50455 129632
rect 50389 129627 50455 129630
rect 47862 129010 47922 129524
rect 90734 129456 90794 129766
rect 92801 129763 92867 129766
rect 101725 129690 101791 129693
rect 103982 129690 104042 130000
rect 143033 129962 143099 129965
rect 143033 129960 145074 129962
rect 143033 129904 143038 129960
rect 143094 129904 145074 129960
rect 143033 129902 145074 129904
rect 143033 129899 143099 129902
rect 101725 129688 104042 129690
rect 101725 129632 101730 129688
rect 101786 129632 104042 129688
rect 101725 129630 104042 129632
rect 101725 129627 101791 129630
rect 134661 129554 134727 129557
rect 131796 129552 134727 129554
rect 131796 129496 134666 129552
rect 134722 129496 134727 129552
rect 131796 129494 134727 129496
rect 134661 129491 134727 129494
rect 145014 129456 145074 129902
rect 177625 129826 177691 129829
rect 174822 129824 177691 129826
rect 174822 129768 177630 129824
rect 177686 129768 177691 129824
rect 174822 129766 177691 129768
rect 58301 129418 58367 129421
rect 58301 129416 60956 129418
rect 58301 129360 58306 129416
rect 58362 129360 60956 129416
rect 58301 129358 60956 129360
rect 58301 129355 58367 129358
rect 51217 129010 51283 129013
rect 47862 129008 51283 129010
rect 47862 128952 51222 129008
rect 51278 128952 51283 129008
rect 47862 128950 51283 128952
rect 51217 128947 51283 128950
rect 101265 129010 101331 129013
rect 103982 129010 104042 129456
rect 174822 129388 174882 129766
rect 177625 129763 177691 129766
rect 185169 129690 185235 129693
rect 187886 129690 187946 130068
rect 185169 129688 187946 129690
rect 185169 129632 185174 129688
rect 185230 129632 187946 129688
rect 185169 129630 187946 129632
rect 185169 129627 185235 129630
rect 101265 129008 104042 129010
rect 101265 128952 101270 129008
rect 101326 128952 104042 129008
rect 101265 128950 104042 128952
rect 185445 129010 185511 129013
rect 187886 129010 187946 129524
rect 185445 129008 187946 129010
rect 185445 128952 185450 129008
rect 185506 128952 187946 129008
rect 185445 128950 187946 128952
rect 101265 128947 101331 128950
rect 185445 128947 185511 128950
rect 58209 128874 58275 128877
rect 92709 128874 92775 128877
rect 135397 128874 135463 128877
rect 58209 128872 60956 128874
rect 47862 128466 47922 128844
rect 58209 128816 58214 128872
rect 58270 128816 60956 128872
rect 58209 128814 60956 128816
rect 90764 128872 92775 128874
rect 90764 128816 92714 128872
rect 92770 128816 92775 128872
rect 90764 128814 92775 128816
rect 131796 128872 135463 128874
rect 131796 128816 135402 128872
rect 135458 128816 135463 128872
rect 131796 128814 135463 128816
rect 58209 128811 58275 128814
rect 92709 128811 92775 128814
rect 135397 128811 135463 128814
rect 142757 128874 142823 128877
rect 142757 128872 145044 128874
rect 142757 128816 142762 128872
rect 142818 128816 145044 128872
rect 142757 128814 145044 128816
rect 142757 128811 142823 128814
rect 50941 128466 51007 128469
rect 92801 128466 92867 128469
rect 47862 128464 51007 128466
rect 47862 128408 50946 128464
rect 51002 128408 51007 128464
rect 47862 128406 51007 128408
rect 50941 128403 51007 128406
rect 90734 128464 92867 128466
rect 90734 128408 92806 128464
rect 92862 128408 92867 128464
rect 90734 128406 92867 128408
rect 47862 127922 47922 128300
rect 90734 128232 90794 128406
rect 92801 128403 92867 128406
rect 100989 128466 101055 128469
rect 103982 128466 104042 128776
rect 143585 128738 143651 128741
rect 174822 128738 174882 128844
rect 177717 128738 177783 128741
rect 143585 128736 145074 128738
rect 143585 128680 143590 128736
rect 143646 128680 145074 128736
rect 143585 128678 145074 128680
rect 174822 128736 177783 128738
rect 174822 128680 177722 128736
rect 177778 128680 177783 128736
rect 174822 128678 177783 128680
rect 143585 128675 143651 128678
rect 100989 128464 104042 128466
rect 100989 128408 100994 128464
rect 101050 128408 104042 128464
rect 100989 128406 104042 128408
rect 100989 128403 101055 128406
rect 134661 128330 134727 128333
rect 131796 128328 134727 128330
rect 131796 128272 134666 128328
rect 134722 128272 134727 128328
rect 131796 128270 134727 128272
rect 134661 128267 134727 128270
rect 145014 128232 145074 128678
rect 177717 128675 177783 128678
rect 177625 128466 177691 128469
rect 174822 128464 177691 128466
rect 174822 128408 177630 128464
rect 177686 128408 177691 128464
rect 174822 128406 177691 128408
rect 58301 128194 58367 128197
rect 58301 128192 60956 128194
rect 58301 128136 58306 128192
rect 58362 128136 60956 128192
rect 58301 128134 60956 128136
rect 58301 128131 58367 128134
rect 92709 128058 92775 128061
rect 90734 128056 92775 128058
rect 90734 128000 92714 128056
rect 92770 128000 92775 128056
rect 90734 127998 92775 128000
rect 51217 127922 51283 127925
rect 47862 127920 51283 127922
rect 47862 127864 51222 127920
rect 51278 127864 51283 127920
rect 47862 127862 51283 127864
rect 51217 127859 51283 127862
rect 47862 127650 47922 127756
rect 90734 127688 90794 127998
rect 92709 127995 92775 127998
rect 101173 127922 101239 127925
rect 103982 127922 104042 128232
rect 174822 128164 174882 128406
rect 177625 128403 177691 128406
rect 185169 128466 185235 128469
rect 187886 128466 187946 128844
rect 185169 128464 187946 128466
rect 185169 128408 185174 128464
rect 185230 128408 187946 128464
rect 185169 128406 187946 128408
rect 185169 128403 185235 128406
rect 143125 128058 143191 128061
rect 177349 128058 177415 128061
rect 143125 128056 145074 128058
rect 143125 128000 143130 128056
rect 143186 128000 145074 128056
rect 143125 127998 145074 128000
rect 143125 127995 143191 127998
rect 101173 127920 104042 127922
rect 101173 127864 101178 127920
rect 101234 127864 104042 127920
rect 101173 127862 104042 127864
rect 101173 127859 101239 127862
rect 101081 127786 101147 127789
rect 134661 127786 134727 127789
rect 101081 127784 104012 127786
rect 101081 127728 101086 127784
rect 101142 127728 104012 127784
rect 101081 127726 104012 127728
rect 131796 127784 134727 127786
rect 131796 127728 134666 127784
rect 134722 127728 134727 127784
rect 131796 127726 134727 127728
rect 101081 127723 101147 127726
rect 134661 127723 134727 127726
rect 145014 127688 145074 127998
rect 174822 128056 177415 128058
rect 174822 128000 177354 128056
rect 177410 128000 177415 128056
rect 174822 127998 177415 128000
rect 51217 127650 51283 127653
rect 47862 127648 51283 127650
rect 47862 127592 51222 127648
rect 51278 127592 51283 127648
rect 47862 127590 51283 127592
rect 51217 127587 51283 127590
rect 58209 127650 58275 127653
rect 58209 127648 60956 127650
rect 58209 127592 58214 127648
rect 58270 127592 60956 127648
rect 174822 127620 174882 127998
rect 177349 127995 177415 127998
rect 185353 127922 185419 127925
rect 187886 127922 187946 128300
rect 185353 127920 187946 127922
rect 185353 127864 185358 127920
rect 185414 127864 187946 127920
rect 185353 127862 187946 127864
rect 185353 127859 185419 127862
rect 185261 127650 185327 127653
rect 187886 127650 187946 127756
rect 185261 127648 187946 127650
rect 58209 127590 60956 127592
rect 185261 127592 185266 127648
rect 185322 127592 187946 127648
rect 185261 127590 187946 127592
rect 58209 127587 58275 127590
rect 185261 127587 185327 127590
rect 142481 127378 142547 127381
rect 218289 127378 218355 127381
rect 142481 127376 145074 127378
rect 142481 127320 142486 127376
rect 142542 127320 145074 127376
rect 142481 127318 145074 127320
rect 142481 127315 142547 127318
rect 92709 127242 92775 127245
rect 135397 127242 135463 127245
rect 90734 127240 92775 127242
rect 18005 126290 18071 126293
rect 19894 126290 19954 126804
rect 47862 126698 47922 127212
rect 90734 127184 92714 127240
rect 92770 127184 92775 127240
rect 90734 127182 92775 127184
rect 131796 127240 135463 127242
rect 131796 127184 135402 127240
rect 135458 127184 135463 127240
rect 131796 127182 135463 127184
rect 90734 127144 90794 127182
rect 92709 127179 92775 127182
rect 135397 127179 135463 127182
rect 145014 127144 145074 127318
rect 215670 127376 218355 127378
rect 215670 127320 218294 127376
rect 218350 127320 218355 127376
rect 215670 127318 218355 127320
rect 177165 127242 177231 127245
rect 174822 127240 177231 127242
rect 174822 127184 177170 127240
rect 177226 127184 177231 127240
rect 174822 127182 177231 127184
rect 58209 127106 58275 127109
rect 58209 127104 60956 127106
rect 58209 127048 58214 127104
rect 58270 127048 60956 127104
rect 58209 127046 60956 127048
rect 58209 127043 58275 127046
rect 92801 126970 92867 126973
rect 90734 126968 92867 126970
rect 90734 126912 92806 126968
rect 92862 126912 92867 126968
rect 90734 126910 92867 126912
rect 51217 126698 51283 126701
rect 47862 126696 51283 126698
rect 47862 126640 51222 126696
rect 51278 126640 51283 126696
rect 47862 126638 51283 126640
rect 51217 126635 51283 126638
rect 18005 126288 19954 126290
rect 18005 126232 18010 126288
rect 18066 126232 19954 126288
rect 18005 126230 19954 126232
rect 18005 126227 18071 126230
rect 47862 126154 47922 126532
rect 90734 126464 90794 126910
rect 92801 126907 92867 126910
rect 101817 126698 101883 126701
rect 103982 126698 104042 127144
rect 174822 127076 174882 127182
rect 177165 127179 177231 127182
rect 143309 126970 143375 126973
rect 177717 126970 177783 126973
rect 143309 126968 145074 126970
rect 143309 126912 143314 126968
rect 143370 126912 145074 126968
rect 143309 126910 145074 126912
rect 143309 126907 143375 126910
rect 101817 126696 104042 126698
rect 101817 126640 101822 126696
rect 101878 126640 104042 126696
rect 101817 126638 104042 126640
rect 101817 126635 101883 126638
rect 135397 126562 135463 126565
rect 131796 126560 135463 126562
rect 131796 126504 135402 126560
rect 135458 126504 135463 126560
rect 131796 126502 135463 126504
rect 135397 126499 135463 126502
rect 145014 126464 145074 126910
rect 174822 126968 177783 126970
rect 174822 126912 177722 126968
rect 177778 126912 177783 126968
rect 174822 126910 177783 126912
rect 58301 126426 58367 126429
rect 58301 126424 60956 126426
rect 58301 126368 58306 126424
rect 58362 126368 60956 126424
rect 58301 126366 60956 126368
rect 58301 126363 58367 126366
rect 101725 126290 101791 126293
rect 103982 126290 104042 126464
rect 174822 126396 174882 126910
rect 177717 126907 177783 126910
rect 185445 126698 185511 126701
rect 187886 126698 187946 127212
rect 215670 126804 215730 127318
rect 218289 127315 218355 127318
rect 222337 126834 222403 126837
rect 225416 126834 225896 126864
rect 222337 126832 225896 126834
rect 222337 126776 222342 126832
rect 222398 126776 225896 126832
rect 222337 126774 225896 126776
rect 222337 126771 222403 126774
rect 225416 126744 225896 126774
rect 185445 126696 187946 126698
rect 185445 126640 185450 126696
rect 185506 126640 187946 126696
rect 185445 126638 187946 126640
rect 185445 126635 185511 126638
rect 101725 126288 104042 126290
rect 101725 126232 101730 126288
rect 101786 126232 104042 126288
rect 101725 126230 104042 126232
rect 185169 126290 185235 126293
rect 187886 126290 187946 126532
rect 185169 126288 187946 126290
rect 185169 126232 185174 126288
rect 185230 126232 187946 126288
rect 185169 126230 187946 126232
rect 101725 126227 101791 126230
rect 185169 126227 185235 126230
rect 51217 126154 51283 126157
rect 47862 126152 51283 126154
rect 47862 126096 51222 126152
rect 51278 126096 51283 126152
rect 47862 126094 51283 126096
rect 51217 126091 51283 126094
rect 92709 126018 92775 126021
rect 135213 126018 135279 126021
rect 90734 126016 92775 126018
rect 47862 125610 47922 125988
rect 90734 125960 92714 126016
rect 92770 125960 92775 126016
rect 90734 125958 92775 125960
rect 131796 126016 135279 126018
rect 131796 125960 135218 126016
rect 135274 125960 135279 126016
rect 131796 125958 135279 125960
rect 90734 125920 90794 125958
rect 92709 125955 92775 125958
rect 135213 125955 135279 125958
rect 143585 126018 143651 126021
rect 177717 126018 177783 126021
rect 143585 126016 145074 126018
rect 143585 125960 143590 126016
rect 143646 125960 145074 126016
rect 143585 125958 145074 125960
rect 143585 125955 143651 125958
rect 145014 125920 145074 125958
rect 174822 126016 177783 126018
rect 174822 125960 177722 126016
rect 177778 125960 177783 126016
rect 174822 125958 177783 125960
rect 58209 125882 58275 125885
rect 58209 125880 60956 125882
rect 58209 125824 58214 125880
rect 58270 125824 60956 125880
rect 58209 125822 60956 125824
rect 58209 125819 58275 125822
rect 50205 125610 50271 125613
rect 92801 125610 92867 125613
rect 47862 125608 50271 125610
rect 47862 125552 50210 125608
rect 50266 125552 50271 125608
rect 47862 125550 50271 125552
rect 50205 125547 50271 125550
rect 90734 125608 92867 125610
rect 90734 125552 92806 125608
rect 92862 125552 92867 125608
rect 90734 125550 92867 125552
rect 47862 125066 47922 125444
rect 90734 125240 90794 125550
rect 92801 125547 92867 125550
rect 101449 125610 101515 125613
rect 103982 125610 104042 125920
rect 174822 125852 174882 125958
rect 177717 125955 177783 125958
rect 143033 125746 143099 125749
rect 143033 125744 145074 125746
rect 143033 125688 143038 125744
rect 143094 125688 145074 125744
rect 143033 125686 145074 125688
rect 143033 125683 143099 125686
rect 101449 125608 104042 125610
rect 101449 125552 101454 125608
rect 101510 125552 104042 125608
rect 101449 125550 104042 125552
rect 101449 125547 101515 125550
rect 135029 125474 135095 125477
rect 131796 125472 135095 125474
rect 131796 125416 135034 125472
rect 135090 125416 135095 125472
rect 131796 125414 135095 125416
rect 135029 125411 135095 125414
rect 58301 125202 58367 125205
rect 58301 125200 60956 125202
rect 58301 125144 58306 125200
rect 58362 125144 60956 125200
rect 58301 125142 60956 125144
rect 58301 125139 58367 125142
rect 51217 125066 51283 125069
rect 47862 125064 51283 125066
rect 47862 125008 51222 125064
rect 51278 125008 51283 125064
rect 47862 125006 51283 125008
rect 51217 125003 51283 125006
rect 51217 124930 51283 124933
rect 47678 124928 51283 124930
rect 47678 124872 51222 124928
rect 51278 124872 51283 124928
rect 47678 124870 51283 124872
rect 47678 124764 47738 124870
rect 51217 124867 51283 124870
rect 101633 124930 101699 124933
rect 103982 124930 104042 125376
rect 145014 125240 145074 125686
rect 177625 125610 177691 125613
rect 174822 125608 177691 125610
rect 174822 125552 177630 125608
rect 177686 125552 177691 125608
rect 174822 125550 177691 125552
rect 174822 125172 174882 125550
rect 177625 125547 177691 125550
rect 185169 125610 185235 125613
rect 187886 125610 187946 125988
rect 185169 125608 187946 125610
rect 185169 125552 185174 125608
rect 185230 125552 187946 125608
rect 185169 125550 187946 125552
rect 185169 125547 185235 125550
rect 101633 124928 104042 124930
rect 101633 124872 101638 124928
rect 101694 124872 104042 124928
rect 101633 124870 104042 124872
rect 185353 124930 185419 124933
rect 187886 124930 187946 125444
rect 185353 124928 187946 124930
rect 185353 124872 185358 124928
rect 185414 124872 187946 124928
rect 185353 124870 187946 124872
rect 101633 124867 101699 124870
rect 185353 124867 185419 124870
rect 101725 124794 101791 124797
rect 135397 124794 135463 124797
rect 101725 124792 104012 124794
rect 101725 124736 101730 124792
rect 101786 124736 104012 124792
rect 101725 124734 104012 124736
rect 131796 124792 135463 124794
rect 131796 124736 135402 124792
rect 135458 124736 135463 124792
rect 131796 124734 135463 124736
rect 101725 124731 101791 124734
rect 135397 124731 135463 124734
rect 185261 124794 185327 124797
rect 185261 124792 187762 124794
rect 185261 124736 185266 124792
rect 185322 124736 187762 124792
rect 185261 124734 187762 124736
rect 185261 124731 185327 124734
rect 58209 124658 58275 124661
rect 92709 124658 92775 124661
rect 58209 124656 60956 124658
rect 58209 124600 58214 124656
rect 58270 124600 60956 124656
rect 58209 124598 60956 124600
rect 90764 124656 92775 124658
rect 90764 124600 92714 124656
rect 92770 124600 92775 124656
rect 90764 124598 92775 124600
rect 58209 124595 58275 124598
rect 92709 124595 92775 124598
rect 143585 124658 143651 124661
rect 187702 124658 187762 124734
rect 187886 124658 187946 124764
rect 143585 124656 145044 124658
rect 143585 124600 143590 124656
rect 143646 124600 145044 124656
rect 143585 124598 145044 124600
rect 143585 124595 143651 124598
rect 174822 124522 174882 124628
rect 187702 124598 187946 124658
rect 177717 124522 177783 124525
rect 174822 124520 177783 124522
rect 174822 124464 177722 124520
rect 177778 124464 177783 124520
rect 174822 124462 177783 124464
rect 177717 124459 177783 124462
rect 92801 124386 92867 124389
rect 90734 124384 92867 124386
rect 90734 124328 92806 124384
rect 92862 124328 92867 124384
rect 90734 124326 92867 124328
rect 47862 123842 47922 124220
rect 90734 124152 90794 124326
rect 92801 124323 92867 124326
rect 142481 124386 142547 124389
rect 142481 124384 145074 124386
rect 142481 124328 142486 124384
rect 142542 124328 145074 124384
rect 142481 124326 145074 124328
rect 142481 124323 142547 124326
rect 134109 124250 134175 124253
rect 131796 124248 134175 124250
rect 131796 124192 134114 124248
rect 134170 124192 134175 124248
rect 131796 124190 134175 124192
rect 134109 124187 134175 124190
rect 145014 124152 145074 124326
rect 177165 124250 177231 124253
rect 174822 124248 177231 124250
rect 174822 124192 177170 124248
rect 177226 124192 177231 124248
rect 174822 124190 177231 124192
rect 58301 124114 58367 124117
rect 58301 124112 60956 124114
rect 58301 124056 58306 124112
rect 58362 124056 60956 124112
rect 58301 124054 60956 124056
rect 58301 124051 58367 124054
rect 92893 123978 92959 123981
rect 90734 123976 92959 123978
rect 90734 123920 92898 123976
rect 92954 123920 92959 123976
rect 90734 123918 92959 123920
rect 50573 123842 50639 123845
rect 47862 123840 50639 123842
rect 47862 123784 50578 123840
rect 50634 123784 50639 123840
rect 47862 123782 50639 123784
rect 50573 123779 50639 123782
rect 47862 123434 47922 123676
rect 90734 123472 90794 123918
rect 92893 123915 92959 123918
rect 101909 123842 101975 123845
rect 103982 123842 104042 124152
rect 174822 124084 174882 124190
rect 177165 124187 177231 124190
rect 142757 123978 142823 123981
rect 177625 123978 177691 123981
rect 142757 123976 145074 123978
rect 142757 123920 142762 123976
rect 142818 123920 145074 123976
rect 142757 123918 145074 123920
rect 142757 123915 142823 123918
rect 101909 123840 104042 123842
rect 101909 123784 101914 123840
rect 101970 123784 104042 123840
rect 101909 123782 104042 123784
rect 101909 123779 101975 123782
rect 134477 123706 134543 123709
rect 131796 123704 134543 123706
rect 131796 123648 134482 123704
rect 134538 123648 134543 123704
rect 131796 123646 134543 123648
rect 134477 123643 134543 123646
rect 51125 123434 51191 123437
rect 47862 123432 51191 123434
rect 47862 123376 51130 123432
rect 51186 123376 51191 123432
rect 47862 123374 51191 123376
rect 51125 123371 51191 123374
rect 58393 123434 58459 123437
rect 101817 123434 101883 123437
rect 103982 123434 104042 123608
rect 145014 123472 145074 123918
rect 174822 123976 177691 123978
rect 174822 123920 177630 123976
rect 177686 123920 177691 123976
rect 174822 123918 177691 123920
rect 58393 123432 60956 123434
rect 58393 123376 58398 123432
rect 58454 123376 60956 123432
rect 58393 123374 60956 123376
rect 101817 123432 104042 123434
rect 101817 123376 101822 123432
rect 101878 123376 104042 123432
rect 174822 123404 174882 123918
rect 177625 123915 177691 123918
rect 185905 123842 185971 123845
rect 187886 123842 187946 124220
rect 185905 123840 187946 123842
rect 185905 123784 185910 123840
rect 185966 123784 187946 123840
rect 185905 123782 187946 123784
rect 185905 123779 185971 123782
rect 185721 123434 185787 123437
rect 187886 123434 187946 123676
rect 185721 123432 187946 123434
rect 101817 123374 104042 123376
rect 185721 123376 185726 123432
rect 185782 123376 187946 123432
rect 185721 123374 187946 123376
rect 58393 123371 58459 123374
rect 101817 123371 101883 123374
rect 185721 123371 185787 123374
rect 143585 123298 143651 123301
rect 143585 123296 145074 123298
rect 143585 123240 143590 123296
rect 143646 123240 145074 123296
rect 143585 123238 145074 123240
rect 143585 123235 143651 123238
rect 92709 123162 92775 123165
rect 90734 123160 92775 123162
rect 90734 123104 92714 123160
rect 92770 123104 92775 123160
rect 90734 123102 92775 123104
rect 47862 122618 47922 122996
rect 90734 122928 90794 123102
rect 92709 123099 92775 123102
rect 134477 123026 134543 123029
rect 131796 123024 134543 123026
rect 131796 122968 134482 123024
rect 134538 122968 134543 123024
rect 131796 122966 134543 122968
rect 134477 122963 134543 122966
rect 145014 122928 145074 123238
rect 177717 123026 177783 123029
rect 174822 123024 177783 123026
rect 174822 122968 177722 123024
rect 177778 122968 177783 123024
rect 174822 122966 177783 122968
rect 58209 122890 58275 122893
rect 58209 122888 60956 122890
rect 58209 122832 58214 122888
rect 58270 122832 60956 122888
rect 58209 122830 60956 122832
rect 58209 122827 58275 122830
rect 92801 122754 92867 122757
rect 90734 122752 92867 122754
rect 90734 122696 92806 122752
rect 92862 122696 92867 122752
rect 90734 122694 92867 122696
rect 50849 122618 50915 122621
rect 47862 122616 50915 122618
rect 47862 122560 50854 122616
rect 50910 122560 50915 122616
rect 47862 122558 50915 122560
rect 50849 122555 50915 122558
rect 47862 122346 47922 122452
rect 50205 122346 50271 122349
rect 47862 122344 50271 122346
rect 47862 122288 50210 122344
rect 50266 122288 50271 122344
rect 47862 122286 50271 122288
rect 50205 122283 50271 122286
rect 90734 122248 90794 122694
rect 92801 122691 92867 122694
rect 101633 122618 101699 122621
rect 103982 122618 104042 122928
rect 174822 122860 174882 122966
rect 177717 122963 177783 122966
rect 142849 122754 142915 122757
rect 177625 122754 177691 122757
rect 142849 122752 145074 122754
rect 142849 122696 142854 122752
rect 142910 122696 145074 122752
rect 142849 122694 145074 122696
rect 142849 122691 142915 122694
rect 101633 122616 104042 122618
rect 101633 122560 101638 122616
rect 101694 122560 104042 122616
rect 101633 122558 104042 122560
rect 101633 122555 101699 122558
rect 134937 122482 135003 122485
rect 131796 122480 135003 122482
rect 131796 122424 134942 122480
rect 134998 122424 135003 122480
rect 131796 122422 135003 122424
rect 134937 122419 135003 122422
rect 58301 122210 58367 122213
rect 58301 122208 60956 122210
rect 58301 122152 58306 122208
rect 58362 122152 60956 122208
rect 58301 122150 60956 122152
rect 58301 122147 58367 122150
rect 101449 122074 101515 122077
rect 103982 122074 104042 122384
rect 145014 122248 145074 122694
rect 174822 122752 177691 122754
rect 174822 122696 177630 122752
rect 177686 122696 177691 122752
rect 174822 122694 177691 122696
rect 174822 122180 174882 122694
rect 177625 122691 177691 122694
rect 185813 122618 185879 122621
rect 187886 122618 187946 122996
rect 185813 122616 187946 122618
rect 185813 122560 185818 122616
rect 185874 122560 187946 122616
rect 185813 122558 187946 122560
rect 185813 122555 185879 122558
rect 185537 122210 185603 122213
rect 187886 122210 187946 122452
rect 185537 122208 187946 122210
rect 185537 122152 185542 122208
rect 185598 122152 187946 122208
rect 185537 122150 187946 122152
rect 185537 122147 185603 122150
rect 101449 122072 104042 122074
rect 101449 122016 101454 122072
rect 101510 122016 104042 122072
rect 101449 122014 104042 122016
rect 101449 122011 101515 122014
rect 134477 121938 134543 121941
rect 131796 121936 134543 121938
rect 47862 121530 47922 121908
rect 131796 121880 134482 121936
rect 134538 121880 134543 121936
rect 131796 121878 134543 121880
rect 134477 121875 134543 121878
rect 92709 121802 92775 121805
rect 90734 121800 92775 121802
rect 90734 121744 92714 121800
rect 92770 121744 92775 121800
rect 90734 121742 92775 121744
rect 90734 121704 90794 121742
rect 92709 121739 92775 121742
rect 58209 121666 58275 121669
rect 58209 121664 60956 121666
rect 58209 121608 58214 121664
rect 58270 121608 60956 121664
rect 58209 121606 60956 121608
rect 58209 121603 58275 121606
rect 50205 121530 50271 121533
rect 92801 121530 92867 121533
rect 47862 121528 50271 121530
rect 47862 121472 50210 121528
rect 50266 121472 50271 121528
rect 47862 121470 50271 121472
rect 50205 121467 50271 121470
rect 90734 121528 92867 121530
rect 90734 121472 92806 121528
rect 92862 121472 92867 121528
rect 90734 121470 92867 121472
rect 47862 120986 47922 121364
rect 90734 121160 90794 121470
rect 92801 121467 92867 121470
rect 101725 121530 101791 121533
rect 103982 121530 104042 121840
rect 143033 121802 143099 121805
rect 177717 121802 177783 121805
rect 143033 121800 145074 121802
rect 143033 121744 143038 121800
rect 143094 121744 145074 121800
rect 143033 121742 145074 121744
rect 143033 121739 143099 121742
rect 145014 121704 145074 121742
rect 174822 121800 177783 121802
rect 174822 121744 177722 121800
rect 177778 121744 177783 121800
rect 174822 121742 177783 121744
rect 174822 121636 174882 121742
rect 177717 121739 177783 121742
rect 101725 121528 104042 121530
rect 101725 121472 101730 121528
rect 101786 121472 104042 121528
rect 101725 121470 104042 121472
rect 142757 121530 142823 121533
rect 177625 121530 177691 121533
rect 142757 121528 145074 121530
rect 142757 121472 142762 121528
rect 142818 121472 145074 121528
rect 142757 121470 145074 121472
rect 101725 121467 101791 121470
rect 142757 121467 142823 121470
rect 134661 121394 134727 121397
rect 131796 121392 134727 121394
rect 131796 121336 134666 121392
rect 134722 121336 134727 121392
rect 131796 121334 134727 121336
rect 134661 121331 134727 121334
rect 58301 121122 58367 121125
rect 101081 121122 101147 121125
rect 103982 121122 104042 121296
rect 145014 121160 145074 121470
rect 174822 121528 177691 121530
rect 174822 121472 177630 121528
rect 177686 121472 177691 121528
rect 174822 121470 177691 121472
rect 58301 121120 60956 121122
rect 58301 121064 58306 121120
rect 58362 121064 60956 121120
rect 58301 121062 60956 121064
rect 101081 121120 104042 121122
rect 101081 121064 101086 121120
rect 101142 121064 104042 121120
rect 174822 121092 174882 121470
rect 177625 121467 177691 121470
rect 185353 121530 185419 121533
rect 187886 121530 187946 121908
rect 185353 121528 187946 121530
rect 185353 121472 185358 121528
rect 185414 121472 187946 121528
rect 185353 121470 187946 121472
rect 185353 121467 185419 121470
rect 101081 121062 104042 121064
rect 58301 121059 58367 121062
rect 101081 121059 101147 121062
rect 51217 120986 51283 120989
rect 47862 120984 51283 120986
rect 47862 120928 51222 120984
rect 51278 120928 51283 120984
rect 47862 120926 51283 120928
rect 51217 120923 51283 120926
rect 51217 120850 51283 120853
rect 47678 120848 51283 120850
rect 47678 120792 51222 120848
rect 51278 120792 51283 120848
rect 47678 120790 51283 120792
rect 47678 120684 47738 120790
rect 51217 120787 51283 120790
rect 185169 120850 185235 120853
rect 187886 120850 187946 121364
rect 185169 120848 187946 120850
rect 185169 120792 185174 120848
rect 185230 120792 187946 120848
rect 185169 120790 187946 120792
rect 185169 120787 185235 120790
rect 101541 120714 101607 120717
rect 135397 120714 135463 120717
rect 101541 120712 104012 120714
rect 101541 120656 101546 120712
rect 101602 120656 104012 120712
rect 101541 120654 104012 120656
rect 131796 120712 135463 120714
rect 131796 120656 135402 120712
rect 135458 120656 135463 120712
rect 131796 120654 135463 120656
rect 101541 120651 101607 120654
rect 135397 120651 135463 120654
rect 185261 120714 185327 120717
rect 185261 120712 187762 120714
rect 185261 120656 185266 120712
rect 185322 120656 187762 120712
rect 185261 120654 187762 120656
rect 185261 120651 185327 120654
rect 92709 120578 92775 120581
rect 90734 120576 92775 120578
rect 90734 120520 92714 120576
rect 92770 120520 92775 120576
rect 90734 120518 92775 120520
rect 90734 120480 90794 120518
rect 92709 120515 92775 120518
rect 142941 120578 143007 120581
rect 177717 120578 177783 120581
rect 142941 120576 145074 120578
rect 142941 120520 142946 120576
rect 143002 120520 145074 120576
rect 142941 120518 145074 120520
rect 142941 120515 143007 120518
rect 145014 120480 145074 120518
rect 174822 120576 177783 120578
rect 174822 120520 177722 120576
rect 177778 120520 177783 120576
rect 174822 120518 177783 120520
rect 187702 120578 187762 120654
rect 187886 120578 187946 120684
rect 187702 120518 187946 120578
rect 58209 120442 58275 120445
rect 58209 120440 60956 120442
rect 58209 120384 58214 120440
rect 58270 120384 60956 120440
rect 174822 120412 174882 120518
rect 177717 120515 177783 120518
rect 58209 120382 60956 120384
rect 58209 120379 58275 120382
rect 143585 120306 143651 120309
rect 143585 120304 145074 120306
rect 143585 120248 143590 120304
rect 143646 120248 145074 120304
rect 143585 120246 145074 120248
rect 143585 120243 143651 120246
rect 92801 120170 92867 120173
rect 134477 120170 134543 120173
rect 90734 120168 92867 120170
rect 47862 119762 47922 120140
rect 90734 120112 92806 120168
rect 92862 120112 92867 120168
rect 90734 120110 92867 120112
rect 131796 120168 134543 120170
rect 131796 120112 134482 120168
rect 134538 120112 134543 120168
rect 131796 120110 134543 120112
rect 90734 119936 90794 120110
rect 92801 120107 92867 120110
rect 134477 120107 134543 120110
rect 58301 119898 58367 119901
rect 58301 119896 60956 119898
rect 58301 119840 58306 119896
rect 58362 119840 60956 119896
rect 58301 119838 60956 119840
rect 58301 119835 58367 119838
rect 51217 119762 51283 119765
rect 47862 119760 51283 119762
rect 47862 119704 51222 119760
rect 51278 119704 51283 119760
rect 47862 119702 51283 119704
rect 51217 119699 51283 119702
rect 101265 119762 101331 119765
rect 103982 119762 104042 120072
rect 145014 119936 145074 120246
rect 177625 120170 177691 120173
rect 174822 120168 177691 120170
rect 174822 120112 177630 120168
rect 177686 120112 177691 120168
rect 174822 120110 177691 120112
rect 174822 119868 174882 120110
rect 177625 120107 177691 120110
rect 101265 119760 104042 119762
rect 101265 119704 101270 119760
rect 101326 119704 104042 119760
rect 101265 119702 104042 119704
rect 185261 119762 185327 119765
rect 187886 119762 187946 120140
rect 185261 119760 187946 119762
rect 185261 119704 185266 119760
rect 185322 119704 187946 119760
rect 185261 119702 187946 119704
rect 101265 119699 101331 119702
rect 185261 119699 185327 119702
rect 135397 119626 135463 119629
rect 131796 119624 135463 119626
rect 47862 119354 47922 119596
rect 131796 119568 135402 119624
rect 135458 119568 135463 119624
rect 131796 119566 135463 119568
rect 135397 119563 135463 119566
rect 51217 119354 51283 119357
rect 47862 119352 51283 119354
rect 47862 119296 51222 119352
rect 51278 119296 51283 119352
rect 47862 119294 51283 119296
rect 51217 119291 51283 119294
rect 101357 119354 101423 119357
rect 103982 119354 104042 119528
rect 101357 119352 104042 119354
rect 101357 119296 101362 119352
rect 101418 119296 104042 119352
rect 101357 119294 104042 119296
rect 185169 119354 185235 119357
rect 187886 119354 187946 119596
rect 185169 119352 187946 119354
rect 185169 119296 185174 119352
rect 185230 119296 187946 119352
rect 185169 119294 187946 119296
rect 101357 119291 101423 119294
rect 185169 119291 185235 119294
rect 58209 119218 58275 119221
rect 92709 119218 92775 119221
rect 58209 119216 60956 119218
rect 58209 119160 58214 119216
rect 58270 119160 60956 119216
rect 58209 119158 60956 119160
rect 90764 119216 92775 119218
rect 90764 119160 92714 119216
rect 92770 119160 92775 119216
rect 90764 119158 92775 119160
rect 58209 119155 58275 119158
rect 92709 119155 92775 119158
rect 143585 119218 143651 119221
rect 143585 119216 145044 119218
rect 143585 119160 143590 119216
rect 143646 119160 145044 119216
rect 143585 119158 145044 119160
rect 143585 119155 143651 119158
rect 143585 119082 143651 119085
rect 174822 119082 174882 119188
rect 177717 119082 177783 119085
rect 143585 119080 145074 119082
rect 143585 119024 143590 119080
rect 143646 119024 145074 119080
rect 143585 119022 145074 119024
rect 174822 119080 177783 119082
rect 174822 119024 177722 119080
rect 177778 119024 177783 119080
rect 174822 119022 177783 119024
rect 143585 119019 143651 119022
rect 92801 118946 92867 118949
rect 134661 118946 134727 118949
rect 90734 118944 92867 118946
rect 47862 118538 47922 118916
rect 90734 118888 92806 118944
rect 92862 118888 92867 118944
rect 90734 118886 92867 118888
rect 131796 118944 134727 118946
rect 131796 118888 134666 118944
rect 134722 118888 134727 118944
rect 131796 118886 134727 118888
rect 90734 118712 90794 118886
rect 92801 118883 92867 118886
rect 134661 118883 134727 118886
rect 58301 118674 58367 118677
rect 58301 118672 60956 118674
rect 58301 118616 58306 118672
rect 58362 118616 60956 118672
rect 58301 118614 60956 118616
rect 58301 118611 58367 118614
rect 51217 118538 51283 118541
rect 92893 118538 92959 118541
rect 47862 118536 51283 118538
rect 47862 118480 51222 118536
rect 51278 118480 51283 118536
rect 47862 118478 51283 118480
rect 51217 118475 51283 118478
rect 90734 118536 92959 118538
rect 90734 118480 92898 118536
rect 92954 118480 92959 118536
rect 90734 118478 92959 118480
rect 47862 117994 47922 118372
rect 90734 118168 90794 118478
rect 92893 118475 92959 118478
rect 101357 118538 101423 118541
rect 103982 118538 104042 118848
rect 145014 118712 145074 119022
rect 177717 119019 177783 119022
rect 177717 118810 177783 118813
rect 174822 118808 177783 118810
rect 174822 118752 177722 118808
rect 177778 118752 177783 118808
rect 174822 118750 177783 118752
rect 174822 118644 174882 118750
rect 177717 118747 177783 118750
rect 101357 118536 104042 118538
rect 101357 118480 101362 118536
rect 101418 118480 104042 118536
rect 101357 118478 104042 118480
rect 142573 118538 142639 118541
rect 177625 118538 177691 118541
rect 142573 118536 145074 118538
rect 142573 118480 142578 118536
rect 142634 118480 145074 118536
rect 142573 118478 145074 118480
rect 101357 118475 101423 118478
rect 142573 118475 142639 118478
rect 134661 118402 134727 118405
rect 131796 118400 134727 118402
rect 131796 118344 134666 118400
rect 134722 118344 134727 118400
rect 131796 118342 134727 118344
rect 134661 118339 134727 118342
rect 58393 118130 58459 118133
rect 101725 118130 101791 118133
rect 103982 118130 104042 118304
rect 145014 118168 145074 118478
rect 174822 118536 177691 118538
rect 174822 118480 177630 118536
rect 177686 118480 177691 118536
rect 174822 118478 177691 118480
rect 58393 118128 60956 118130
rect 58393 118072 58398 118128
rect 58454 118072 60956 118128
rect 58393 118070 60956 118072
rect 101725 118128 104042 118130
rect 101725 118072 101730 118128
rect 101786 118072 104042 118128
rect 174822 118100 174882 118478
rect 177625 118475 177691 118478
rect 185261 118538 185327 118541
rect 187886 118538 187946 118916
rect 185261 118536 187946 118538
rect 185261 118480 185266 118536
rect 185322 118480 187946 118536
rect 185261 118478 187946 118480
rect 185261 118475 185327 118478
rect 101725 118070 104042 118072
rect 58393 118067 58459 118070
rect 101725 118067 101791 118070
rect 51217 117994 51283 117997
rect 47862 117992 51283 117994
rect 47862 117936 51222 117992
rect 51278 117936 51283 117992
rect 47862 117934 51283 117936
rect 51217 117931 51283 117934
rect 185169 117994 185235 117997
rect 187886 117994 187946 118372
rect 185169 117992 187946 117994
rect 185169 117936 185174 117992
rect 185230 117936 187946 117992
rect 185169 117934 187946 117936
rect 185169 117931 185235 117934
rect 134845 117858 134911 117861
rect 131796 117856 134911 117858
rect 18005 117042 18071 117045
rect 19894 117042 19954 117556
rect 47862 117450 47922 117828
rect 131796 117800 134850 117856
rect 134906 117800 134911 117856
rect 131796 117798 134911 117800
rect 134845 117795 134911 117798
rect 92709 117586 92775 117589
rect 90734 117584 92775 117586
rect 90734 117528 92714 117584
rect 92770 117528 92775 117584
rect 90734 117526 92775 117528
rect 90734 117488 90794 117526
rect 92709 117523 92775 117526
rect 51217 117450 51283 117453
rect 47862 117448 51283 117450
rect 47862 117392 51222 117448
rect 51278 117392 51283 117448
rect 47862 117390 51283 117392
rect 51217 117387 51283 117390
rect 58209 117450 58275 117453
rect 101173 117450 101239 117453
rect 103982 117450 104042 117760
rect 142573 117722 142639 117725
rect 142573 117720 145074 117722
rect 142573 117664 142578 117720
rect 142634 117664 145074 117720
rect 142573 117662 145074 117664
rect 142573 117659 142639 117662
rect 145014 117488 145074 117662
rect 177717 117586 177783 117589
rect 174822 117584 177783 117586
rect 174822 117528 177722 117584
rect 177778 117528 177783 117584
rect 174822 117526 177783 117528
rect 58209 117448 60956 117450
rect 58209 117392 58214 117448
rect 58270 117392 60956 117448
rect 58209 117390 60956 117392
rect 101173 117448 104042 117450
rect 101173 117392 101178 117448
rect 101234 117392 104042 117448
rect 174822 117420 174882 117526
rect 177717 117523 177783 117526
rect 185353 117450 185419 117453
rect 187886 117450 187946 117828
rect 185353 117448 187946 117450
rect 101173 117390 104042 117392
rect 185353 117392 185358 117448
rect 185414 117392 187946 117448
rect 185353 117390 187946 117392
rect 58209 117387 58275 117390
rect 101173 117387 101239 117390
rect 185353 117387 185419 117390
rect 92801 117314 92867 117317
rect 134937 117314 135003 117317
rect 90734 117312 92867 117314
rect 18005 117040 19954 117042
rect 18005 116984 18010 117040
rect 18066 116984 19954 117040
rect 18005 116982 19954 116984
rect 18005 116979 18071 116982
rect 47862 116770 47922 117284
rect 90734 117256 92806 117312
rect 92862 117256 92867 117312
rect 90734 117254 92867 117256
rect 131796 117312 135003 117314
rect 131796 117256 134942 117312
rect 134998 117256 135003 117312
rect 131796 117254 135003 117256
rect 90734 116944 90794 117254
rect 92801 117251 92867 117254
rect 134937 117251 135003 117254
rect 143217 117314 143283 117317
rect 177625 117314 177691 117317
rect 143217 117312 145074 117314
rect 143217 117256 143222 117312
rect 143278 117256 145074 117312
rect 143217 117254 145074 117256
rect 143217 117251 143283 117254
rect 58301 116906 58367 116909
rect 58301 116904 60956 116906
rect 58301 116848 58306 116904
rect 58362 116848 60956 116904
rect 58301 116846 60956 116848
rect 58301 116843 58367 116846
rect 50573 116770 50639 116773
rect 47862 116768 50639 116770
rect 47862 116712 50578 116768
rect 50634 116712 50639 116768
rect 47862 116710 50639 116712
rect 50573 116707 50639 116710
rect 101081 116770 101147 116773
rect 103982 116770 104042 117216
rect 145014 116944 145074 117254
rect 174822 117312 177691 117314
rect 174822 117256 177630 117312
rect 177686 117256 177691 117312
rect 215854 117314 215914 117556
rect 216909 117314 216975 117317
rect 217553 117314 217619 117317
rect 215854 117312 217619 117314
rect 174822 117254 177691 117256
rect 174822 116876 174882 117254
rect 177625 117251 177691 117254
rect 101081 116768 104042 116770
rect 101081 116712 101086 116768
rect 101142 116712 104042 116768
rect 101081 116710 104042 116712
rect 185261 116770 185327 116773
rect 187886 116770 187946 117284
rect 215854 117256 216914 117312
rect 216970 117256 217558 117312
rect 217614 117256 217619 117312
rect 215854 117254 217619 117256
rect 216909 117251 216975 117254
rect 217553 117251 217619 117254
rect 185261 116768 187946 116770
rect 185261 116712 185266 116768
rect 185322 116712 187946 116768
rect 185261 116710 187946 116712
rect 101081 116707 101147 116710
rect 185261 116707 185327 116710
rect 100989 116634 101055 116637
rect 134753 116634 134819 116637
rect 100989 116632 104012 116634
rect 47862 116498 47922 116604
rect 100989 116576 100994 116632
rect 101050 116576 104012 116632
rect 100989 116574 104012 116576
rect 131796 116632 134819 116634
rect 131796 116576 134758 116632
rect 134814 116576 134819 116632
rect 131796 116574 134819 116576
rect 100989 116571 101055 116574
rect 134753 116571 134819 116574
rect 50757 116498 50823 116501
rect 47862 116496 50823 116498
rect 47862 116440 50762 116496
rect 50818 116440 50823 116496
rect 47862 116438 50823 116440
rect 50757 116435 50823 116438
rect 185169 116498 185235 116501
rect 187886 116498 187946 116604
rect 185169 116496 187946 116498
rect 185169 116440 185174 116496
rect 185230 116440 187946 116496
rect 185169 116438 187946 116440
rect 185169 116435 185235 116438
rect 92709 116362 92775 116365
rect 90734 116360 92775 116362
rect 90734 116304 92714 116360
rect 92770 116304 92775 116360
rect 90734 116302 92775 116304
rect 90734 116264 90794 116302
rect 92709 116299 92775 116302
rect 142941 116362 143007 116365
rect 177717 116362 177783 116365
rect 142941 116360 145074 116362
rect 142941 116304 142946 116360
rect 143002 116304 145074 116360
rect 142941 116302 145074 116304
rect 142941 116299 143007 116302
rect 145014 116264 145074 116302
rect 174822 116360 177783 116362
rect 174822 116304 177722 116360
rect 177778 116304 177783 116360
rect 174822 116302 177783 116304
rect 58209 116226 58275 116229
rect 58209 116224 60956 116226
rect 58209 116168 58214 116224
rect 58270 116168 60956 116224
rect 174822 116196 174882 116302
rect 177717 116299 177783 116302
rect 58209 116166 60956 116168
rect 58209 116163 58275 116166
rect 135029 116090 135095 116093
rect 131796 116088 135095 116090
rect 47862 115682 47922 116060
rect 131796 116032 135034 116088
rect 135090 116032 135095 116088
rect 131796 116030 135095 116032
rect 135029 116027 135095 116030
rect 143585 116090 143651 116093
rect 143585 116088 145074 116090
rect 143585 116032 143590 116088
rect 143646 116032 145074 116088
rect 143585 116030 145074 116032
rect 143585 116027 143651 116030
rect 92801 115954 92867 115957
rect 90734 115952 92867 115954
rect 90734 115896 92806 115952
rect 92862 115896 92867 115952
rect 90734 115894 92867 115896
rect 90734 115720 90794 115894
rect 92801 115891 92867 115894
rect 50849 115682 50915 115685
rect 47862 115680 50915 115682
rect 47862 115624 50854 115680
rect 50910 115624 50915 115680
rect 47862 115622 50915 115624
rect 50849 115619 50915 115622
rect 58301 115682 58367 115685
rect 101081 115682 101147 115685
rect 103982 115682 104042 115992
rect 145014 115720 145074 116030
rect 177717 115954 177783 115957
rect 174822 115952 177783 115954
rect 174822 115896 177722 115952
rect 177778 115896 177783 115952
rect 174822 115894 177783 115896
rect 58301 115680 60956 115682
rect 58301 115624 58306 115680
rect 58362 115624 60956 115680
rect 58301 115622 60956 115624
rect 101081 115680 104042 115682
rect 101081 115624 101086 115680
rect 101142 115624 104042 115680
rect 174822 115652 174882 115894
rect 177717 115891 177783 115894
rect 185261 115682 185327 115685
rect 187886 115682 187946 116060
rect 185261 115680 187946 115682
rect 101081 115622 104042 115624
rect 185261 115624 185266 115680
rect 185322 115624 187946 115680
rect 185261 115622 187946 115624
rect 58301 115619 58367 115622
rect 101081 115619 101147 115622
rect 185261 115619 185327 115622
rect 92893 115546 92959 115549
rect 134845 115546 134911 115549
rect 90734 115544 92959 115546
rect 47862 115138 47922 115516
rect 90734 115488 92898 115544
rect 92954 115488 92959 115544
rect 90734 115486 92959 115488
rect 131796 115544 134911 115546
rect 131796 115488 134850 115544
rect 134906 115488 134911 115544
rect 131796 115486 134911 115488
rect 90734 115176 90794 115486
rect 92893 115483 92959 115486
rect 134845 115483 134911 115486
rect 142757 115546 142823 115549
rect 177073 115546 177139 115549
rect 142757 115544 145074 115546
rect 142757 115488 142762 115544
rect 142818 115488 145074 115544
rect 142757 115486 145074 115488
rect 142757 115483 142823 115486
rect 100989 115274 101055 115277
rect 103982 115274 104042 115448
rect 100989 115272 104042 115274
rect 100989 115216 100994 115272
rect 101050 115216 104042 115272
rect 100989 115214 104042 115216
rect 100989 115211 101055 115214
rect 145014 115176 145074 115486
rect 174822 115544 177139 115546
rect 174822 115488 177078 115544
rect 177134 115488 177139 115544
rect 174822 115486 177139 115488
rect 50665 115138 50731 115141
rect 47862 115136 50731 115138
rect 47862 115080 50670 115136
rect 50726 115080 50731 115136
rect 47862 115078 50731 115080
rect 50665 115075 50731 115078
rect 58393 115138 58459 115141
rect 58393 115136 60956 115138
rect 58393 115080 58398 115136
rect 58454 115080 60956 115136
rect 174822 115108 174882 115486
rect 177073 115483 177139 115486
rect 185169 115274 185235 115277
rect 187886 115274 187946 115516
rect 185169 115272 187946 115274
rect 185169 115216 185174 115272
rect 185230 115216 187946 115272
rect 185169 115214 187946 115216
rect 185169 115211 185235 115214
rect 58393 115078 60956 115080
rect 58393 115075 58459 115078
rect 9896 115002 10376 115032
rect 13313 115002 13379 115005
rect 9896 115000 13379 115002
rect 9896 114944 13318 115000
rect 13374 114944 13379 115000
rect 9896 114942 13379 114944
rect 9896 114912 10376 114942
rect 13313 114939 13379 114942
rect 135121 114866 135187 114869
rect 131796 114864 135187 114866
rect 47862 114458 47922 114836
rect 131796 114808 135126 114864
rect 135182 114808 135187 114864
rect 131796 114806 135187 114808
rect 135121 114803 135187 114806
rect 50941 114458 51007 114461
rect 47862 114456 51007 114458
rect 47862 114400 50946 114456
rect 51002 114400 51007 114456
rect 47862 114398 51007 114400
rect 50941 114395 51007 114398
rect 101817 114458 101883 114461
rect 103982 114458 104042 114768
rect 101817 114456 104042 114458
rect 101817 114400 101822 114456
rect 101878 114400 104042 114456
rect 101817 114398 104042 114400
rect 185813 114458 185879 114461
rect 187886 114458 187946 114836
rect 185813 114456 187946 114458
rect 185813 114400 185818 114456
rect 185874 114400 187946 114456
rect 185813 114398 187946 114400
rect 101817 114395 101883 114398
rect 185813 114395 185879 114398
rect 135305 114322 135371 114325
rect 131796 114320 135371 114322
rect 47862 114050 47922 114292
rect 131796 114264 135310 114320
rect 135366 114264 135371 114320
rect 131796 114262 135371 114264
rect 135305 114259 135371 114262
rect 51125 114050 51191 114053
rect 47862 114048 51191 114050
rect 47862 113992 51130 114048
rect 51186 113992 51191 114048
rect 47862 113990 51191 113992
rect 51125 113987 51191 113990
rect 51217 113914 51283 113917
rect 47678 113912 51283 113914
rect 47678 113856 51222 113912
rect 51278 113856 51283 113912
rect 47678 113854 51283 113856
rect 47678 113748 47738 113854
rect 51217 113851 51283 113854
rect 102001 113914 102067 113917
rect 103982 113914 104042 114224
rect 102001 113912 104042 113914
rect 102001 113856 102006 113912
rect 102062 113856 104042 113912
rect 102001 113854 104042 113856
rect 185997 113914 186063 113917
rect 187886 113914 187946 114292
rect 185997 113912 187946 113914
rect 185997 113856 186002 113912
rect 186058 113856 187946 113912
rect 185997 113854 187946 113856
rect 102001 113851 102067 113854
rect 185997 113851 186063 113854
rect 101633 113778 101699 113781
rect 135397 113778 135463 113781
rect 101633 113776 104012 113778
rect 101633 113720 101638 113776
rect 101694 113720 104012 113776
rect 101633 113718 104012 113720
rect 131796 113776 135463 113778
rect 131796 113720 135402 113776
rect 135458 113720 135463 113776
rect 131796 113718 135463 113720
rect 101633 113715 101699 113718
rect 135397 113715 135463 113718
rect 186181 113778 186247 113781
rect 186181 113776 187762 113778
rect 186181 113720 186186 113776
rect 186242 113720 187762 113776
rect 186181 113718 187762 113720
rect 186181 113715 186247 113718
rect 187702 113642 187762 113718
rect 187886 113642 187946 113748
rect 187702 113582 187946 113642
rect 135213 113234 135279 113237
rect 131796 113232 135279 113234
rect 47862 112826 47922 113204
rect 131796 113176 135218 113232
rect 135274 113176 135279 113232
rect 131796 113174 135279 113176
rect 135213 113171 135279 113174
rect 51033 112826 51099 112829
rect 47862 112824 51099 112826
rect 47862 112768 51038 112824
rect 51094 112768 51099 112824
rect 47862 112766 51099 112768
rect 51033 112763 51099 112766
rect 100989 112554 101055 112557
rect 103982 112554 104042 113136
rect 185169 112690 185235 112693
rect 187886 112690 187946 113204
rect 185169 112688 187946 112690
rect 185169 112632 185174 112688
rect 185230 112632 187946 112688
rect 185169 112630 187946 112632
rect 185169 112627 185235 112630
rect 100989 112552 104042 112554
rect 100989 112496 100994 112552
rect 101050 112496 104042 112552
rect 100989 112494 104042 112496
rect 100989 112491 101055 112494
rect 61889 111194 61955 111197
rect 108441 111196 108507 111197
rect 134017 111196 134083 111197
rect 62022 111194 62028 111196
rect 61889 111192 62028 111194
rect 61889 111136 61894 111192
rect 61950 111136 62028 111192
rect 61889 111134 62028 111136
rect 61889 111131 61955 111134
rect 62022 111132 62028 111134
rect 62092 111132 62098 111196
rect 108390 111132 108396 111196
rect 108460 111194 108507 111196
rect 133966 111194 133972 111196
rect 108460 111192 108552 111194
rect 108502 111136 108552 111192
rect 108460 111134 108552 111136
rect 133926 111134 133972 111194
rect 134036 111192 134083 111196
rect 134078 111136 134083 111192
rect 108460 111132 108507 111134
rect 133966 111132 133972 111134
rect 134036 111132 134083 111136
rect 108441 111131 108507 111132
rect 134017 111131 134083 111132
rect 222337 100586 222403 100589
rect 225416 100586 225896 100616
rect 222337 100584 225896 100586
rect 222337 100528 222342 100584
rect 222398 100528 225896 100584
rect 222337 100526 225896 100528
rect 222337 100523 222403 100526
rect 225416 100496 225896 100526
rect 98781 99770 98847 99773
rect 95702 99768 98847 99770
rect 95702 99712 98786 99768
rect 98842 99712 98847 99768
rect 95702 99710 98847 99712
rect 95702 99224 95762 99710
rect 98781 99707 98847 99710
rect 183697 99226 183763 99229
rect 179820 99224 183763 99226
rect 179820 99168 183702 99224
rect 183758 99168 183763 99224
rect 179820 99166 183763 99168
rect 183697 99163 183763 99166
rect 191977 98818 192043 98821
rect 191977 98816 193988 98818
rect 191977 98760 191982 98816
rect 192038 98760 193988 98816
rect 191977 98758 193988 98760
rect 191977 98755 192043 98758
rect 99517 98546 99583 98549
rect 95702 98544 99583 98546
rect 95702 98488 99522 98544
rect 99578 98488 99583 98544
rect 95702 98486 99583 98488
rect 95702 98000 95762 98486
rect 99517 98483 99583 98486
rect 106785 98546 106851 98549
rect 106785 98544 109900 98546
rect 106785 98488 106790 98544
rect 106846 98488 109900 98544
rect 106785 98486 109900 98488
rect 106785 98483 106851 98486
rect 183605 98002 183671 98005
rect 179820 98000 183671 98002
rect 179820 97944 183610 98000
rect 183666 97944 183671 98000
rect 179820 97942 183671 97944
rect 183605 97939 183671 97942
rect 99425 97050 99491 97053
rect 95702 97048 99491 97050
rect 95702 96992 99430 97048
rect 99486 96992 99491 97048
rect 95702 96990 99491 96992
rect 95702 96776 95762 96990
rect 99425 96987 99491 96990
rect 193766 96852 193772 96916
rect 193836 96852 193842 96916
rect 209825 96914 209891 96917
rect 209782 96912 209891 96914
rect 209782 96856 209830 96912
rect 209886 96856 209891 96912
rect 183513 96778 183579 96781
rect 179820 96776 183579 96778
rect 179820 96720 183518 96776
rect 183574 96720 183579 96776
rect 179820 96718 183579 96720
rect 193774 96778 193834 96852
rect 209782 96851 209891 96856
rect 209782 96780 209842 96851
rect 193774 96718 193988 96778
rect 183513 96715 183579 96718
rect 209774 96716 209780 96780
rect 209844 96716 209850 96780
rect 22329 96506 22395 96509
rect 211757 96506 211823 96509
rect 22329 96504 25996 96506
rect 22329 96448 22334 96504
rect 22390 96448 25996 96504
rect 22329 96446 25996 96448
rect 209812 96504 211823 96506
rect 209812 96448 211762 96504
rect 211818 96448 211823 96504
rect 209812 96446 211823 96448
rect 22329 96443 22395 96446
rect 211757 96443 211823 96446
rect 106785 96234 106851 96237
rect 106785 96232 109900 96234
rect 106785 96176 106790 96232
rect 106846 96176 109900 96232
rect 106785 96174 109900 96176
rect 106785 96171 106851 96174
rect 99241 95554 99307 95557
rect 183329 95554 183395 95557
rect 95732 95552 99307 95554
rect 95732 95496 99246 95552
rect 99302 95496 99307 95552
rect 95732 95494 99307 95496
rect 179820 95552 183395 95554
rect 179820 95496 183334 95552
rect 183390 95496 183395 95552
rect 179820 95494 183395 95496
rect 99241 95491 99307 95494
rect 183329 95491 183395 95494
rect 41833 95282 41899 95285
rect 41790 95280 41899 95282
rect 41790 95224 41838 95280
rect 41894 95224 41899 95280
rect 41790 95219 41899 95224
rect 41790 94708 41850 95219
rect 191977 94738 192043 94741
rect 191977 94736 193988 94738
rect 191977 94680 191982 94736
rect 192038 94680 193988 94736
rect 191977 94678 193988 94680
rect 191977 94675 192043 94678
rect 99333 94330 99399 94333
rect 183421 94330 183487 94333
rect 95732 94328 99399 94330
rect 95732 94272 99338 94328
rect 99394 94272 99399 94328
rect 95732 94270 99399 94272
rect 179820 94328 183487 94330
rect 179820 94272 183426 94328
rect 183482 94272 183487 94328
rect 179820 94270 183487 94272
rect 99333 94267 99399 94270
rect 183421 94267 183487 94270
rect 106509 93922 106575 93925
rect 106509 93920 109900 93922
rect 106509 93864 106514 93920
rect 106570 93864 109900 93920
rect 106509 93862 109900 93864
rect 106509 93859 106575 93862
rect 99149 93650 99215 93653
rect 95702 93648 99215 93650
rect 95702 93592 99154 93648
rect 99210 93592 99215 93648
rect 95702 93590 99215 93592
rect 95702 93104 95762 93590
rect 99149 93587 99215 93590
rect 183237 93106 183303 93109
rect 179820 93104 183303 93106
rect 179820 93048 183242 93104
rect 183298 93048 183303 93104
rect 179820 93046 183303 93048
rect 183237 93043 183303 93046
rect 191149 92834 191215 92837
rect 191149 92832 193988 92834
rect 191149 92776 191154 92832
rect 191210 92776 193988 92832
rect 191149 92774 193988 92776
rect 191149 92771 191215 92774
rect 99057 92426 99123 92429
rect 95702 92424 99123 92426
rect 95702 92368 99062 92424
rect 99118 92368 99123 92424
rect 95702 92366 99123 92368
rect 95702 91880 95762 92366
rect 99057 92363 99123 92366
rect 183145 91882 183211 91885
rect 179820 91880 183211 91882
rect 179820 91824 183150 91880
rect 183206 91824 183211 91880
rect 179820 91822 183211 91824
rect 183145 91819 183211 91822
rect 106785 91474 106851 91477
rect 106785 91472 109900 91474
rect 106785 91416 106790 91472
rect 106846 91416 109900 91472
rect 106785 91414 109900 91416
rect 106785 91411 106851 91414
rect 9896 91338 10376 91368
rect 13313 91338 13379 91341
rect 9896 91336 13379 91338
rect 9896 91280 13318 91336
rect 13374 91280 13379 91336
rect 9896 91278 13379 91280
rect 9896 91248 10376 91278
rect 13313 91275 13379 91278
rect 98965 91202 99031 91205
rect 95702 91200 99031 91202
rect 95702 91144 98970 91200
rect 99026 91144 99031 91200
rect 95702 91142 99031 91144
rect 95702 90656 95762 91142
rect 98965 91139 99031 91142
rect 190781 90794 190847 90797
rect 190781 90792 193988 90794
rect 190781 90736 190786 90792
rect 190842 90736 193988 90792
rect 190781 90734 193988 90736
rect 190781 90731 190847 90734
rect 183053 90658 183119 90661
rect 179820 90656 183119 90658
rect 179820 90600 183058 90656
rect 183114 90600 183119 90656
rect 179820 90598 183119 90600
rect 183053 90595 183119 90598
rect 98781 89978 98847 89981
rect 95702 89976 98847 89978
rect 95702 89920 98786 89976
rect 98842 89920 98847 89976
rect 95702 89918 98847 89920
rect 22329 89842 22395 89845
rect 22329 89840 25996 89842
rect 22329 89784 22334 89840
rect 22390 89784 25996 89840
rect 22329 89782 25996 89784
rect 22329 89779 22395 89782
rect 95702 89432 95762 89918
rect 98781 89915 98847 89918
rect 128497 89842 128563 89845
rect 211849 89842 211915 89845
rect 125724 89840 128563 89842
rect 125724 89784 128502 89840
rect 128558 89784 128563 89840
rect 125724 89782 128563 89784
rect 209812 89840 211915 89842
rect 209812 89784 211854 89840
rect 211910 89784 211915 89840
rect 209812 89782 211915 89784
rect 128497 89779 128563 89782
rect 211849 89779 211915 89782
rect 182869 89434 182935 89437
rect 179820 89432 182935 89434
rect 179820 89376 182874 89432
rect 182930 89376 182935 89432
rect 179820 89374 182935 89376
rect 182869 89371 182935 89374
rect 106785 89162 106851 89165
rect 106785 89160 109900 89162
rect 106785 89104 106790 89160
rect 106846 89104 109900 89160
rect 106785 89102 109900 89104
rect 106785 89099 106851 89102
rect 99517 88754 99583 88757
rect 95702 88752 99583 88754
rect 95702 88696 99522 88752
rect 99578 88696 99583 88752
rect 95702 88694 99583 88696
rect 95702 88208 95762 88694
rect 99517 88691 99583 88694
rect 191701 88754 191767 88757
rect 191701 88752 193988 88754
rect 191701 88696 191706 88752
rect 191762 88696 193988 88752
rect 191701 88694 193988 88696
rect 191701 88691 191767 88694
rect 183513 88210 183579 88213
rect 179820 88208 183579 88210
rect 179820 88152 183518 88208
rect 183574 88152 183579 88208
rect 179820 88150 183579 88152
rect 183513 88147 183579 88150
rect 98689 87394 98755 87397
rect 95702 87392 98755 87394
rect 95702 87336 98694 87392
rect 98750 87336 98755 87392
rect 95702 87334 98755 87336
rect 95702 87120 95762 87334
rect 98689 87331 98755 87334
rect 183697 87122 183763 87125
rect 179820 87120 183763 87122
rect 179820 87064 183702 87120
rect 183758 87064 183763 87120
rect 179820 87062 183763 87064
rect 183697 87059 183763 87062
rect 106785 86850 106851 86853
rect 191609 86850 191675 86853
rect 106785 86848 109900 86850
rect 106785 86792 106790 86848
rect 106846 86792 109900 86848
rect 106785 86790 109900 86792
rect 191609 86848 193988 86850
rect 191609 86792 191614 86848
rect 191670 86792 193988 86848
rect 191609 86790 193988 86792
rect 106785 86787 106851 86790
rect 191609 86787 191675 86790
rect 183697 85898 183763 85901
rect 179820 85896 183763 85898
rect 179820 85840 183702 85896
rect 183758 85840 183763 85896
rect 95702 85354 95762 85840
rect 179820 85838 183763 85840
rect 183697 85835 183763 85838
rect 99517 85354 99583 85357
rect 95702 85352 99583 85354
rect 95702 85296 99522 85352
rect 99578 85296 99583 85352
rect 95702 85294 99583 85296
rect 99517 85291 99583 85294
rect 44409 84810 44475 84813
rect 41820 84808 44475 84810
rect 41820 84752 44414 84808
rect 44470 84752 44475 84808
rect 41820 84750 44475 84752
rect 44409 84747 44475 84750
rect 191977 84810 192043 84813
rect 191977 84808 193988 84810
rect 191977 84752 191982 84808
rect 192038 84752 193988 84808
rect 191977 84750 193988 84752
rect 191977 84747 192043 84750
rect 99517 84674 99583 84677
rect 183697 84674 183763 84677
rect 95732 84672 99583 84674
rect 95732 84616 99522 84672
rect 99578 84616 99583 84672
rect 95732 84614 99583 84616
rect 179820 84672 183763 84674
rect 179820 84616 183702 84672
rect 183758 84616 183763 84672
rect 179820 84614 183763 84616
rect 99517 84611 99583 84614
rect 183697 84611 183763 84614
rect 107797 84402 107863 84405
rect 107797 84400 109900 84402
rect 107797 84344 107802 84400
rect 107858 84344 109900 84400
rect 107797 84342 109900 84344
rect 107797 84339 107863 84342
rect 99425 83994 99491 83997
rect 95702 83992 99491 83994
rect 95702 83936 99430 83992
rect 99486 83936 99491 83992
rect 95702 83934 99491 83936
rect 95702 83448 95762 83934
rect 99425 83931 99491 83934
rect 182501 83450 182567 83453
rect 179820 83448 182567 83450
rect 179820 83392 182506 83448
rect 182562 83392 182567 83448
rect 179820 83390 182567 83392
rect 182501 83387 182567 83390
rect 22329 83178 22395 83181
rect 212033 83178 212099 83181
rect 22329 83176 25996 83178
rect 22329 83120 22334 83176
rect 22390 83120 25996 83176
rect 22329 83118 25996 83120
rect 209812 83176 212099 83178
rect 209812 83120 212038 83176
rect 212094 83120 212099 83176
rect 209812 83118 212099 83120
rect 22329 83115 22395 83118
rect 212033 83115 212099 83118
rect 99517 82770 99583 82773
rect 95702 82768 99583 82770
rect 95702 82712 99522 82768
rect 99578 82712 99583 82768
rect 95702 82710 99583 82712
rect 95702 82224 95762 82710
rect 99517 82707 99583 82710
rect 191977 82770 192043 82773
rect 191977 82768 193988 82770
rect 191977 82712 191982 82768
rect 192038 82712 193988 82768
rect 191977 82710 193988 82712
rect 191977 82707 192043 82710
rect 183697 82226 183763 82229
rect 179820 82224 183763 82226
rect 179820 82168 183702 82224
rect 183758 82168 183763 82224
rect 179820 82166 183763 82168
rect 183697 82163 183763 82166
rect 106785 82090 106851 82093
rect 106785 82088 109900 82090
rect 106785 82032 106790 82088
rect 106846 82032 109900 82088
rect 106785 82030 109900 82032
rect 106785 82027 106851 82030
rect 99517 81546 99583 81549
rect 95702 81544 99583 81546
rect 95702 81488 99522 81544
rect 99578 81488 99583 81544
rect 95702 81486 99583 81488
rect 95702 81000 95762 81486
rect 99517 81483 99583 81486
rect 183237 81002 183303 81005
rect 179820 81000 183303 81002
rect 179820 80944 183242 81000
rect 183298 80944 183303 81000
rect 179820 80942 183303 80944
rect 183237 80939 183303 80942
rect 191885 80866 191951 80869
rect 191885 80864 193988 80866
rect 191885 80808 191890 80864
rect 191946 80808 193988 80864
rect 191885 80806 193988 80808
rect 191885 80803 191951 80806
rect 136869 80458 136935 80461
rect 136869 80456 140106 80458
rect 136869 80400 136874 80456
rect 136930 80400 140106 80456
rect 136869 80398 140106 80400
rect 136869 80395 136935 80398
rect 53333 79914 53399 79917
rect 53333 79912 55988 79914
rect 140046 79912 140106 80398
rect 53333 79856 53338 79912
rect 53394 79856 55988 79912
rect 53333 79854 55988 79856
rect 53333 79851 53399 79854
rect 99517 79778 99583 79781
rect 95732 79776 99583 79778
rect 95732 79720 99522 79776
rect 99578 79720 99583 79776
rect 95732 79718 99583 79720
rect 99517 79715 99583 79718
rect 106785 79778 106851 79781
rect 183697 79778 183763 79781
rect 106785 79776 109900 79778
rect 106785 79720 106790 79776
rect 106846 79720 109900 79776
rect 106785 79718 109900 79720
rect 179820 79776 183763 79778
rect 179820 79720 183702 79776
rect 183758 79720 183763 79776
rect 179820 79718 183763 79720
rect 106785 79715 106851 79718
rect 183697 79715 183763 79718
rect 191977 78826 192043 78829
rect 191977 78824 193988 78826
rect 191977 78768 191982 78824
rect 192038 78768 193988 78824
rect 191977 78766 193988 78768
rect 191977 78763 192043 78766
rect 183513 78554 183579 78557
rect 179820 78552 183579 78554
rect 179820 78496 183518 78552
rect 183574 78496 183579 78552
rect 95702 78010 95762 78496
rect 179820 78494 183579 78496
rect 183513 78491 183579 78494
rect 99517 78010 99583 78013
rect 95702 78008 99583 78010
rect 95702 77952 99522 78008
rect 99578 77952 99583 78008
rect 95702 77950 99583 77952
rect 99517 77947 99583 77950
rect 106509 77466 106575 77469
rect 106509 77464 109900 77466
rect 106509 77408 106514 77464
rect 106570 77408 109900 77464
rect 106509 77406 109900 77408
rect 106509 77403 106575 77406
rect 183053 77330 183119 77333
rect 179820 77328 183119 77330
rect 179820 77272 183058 77328
rect 183114 77272 183119 77328
rect 95702 76786 95762 77272
rect 179820 77270 183119 77272
rect 183053 77267 183119 77270
rect 209825 76922 209891 76925
rect 209782 76920 209891 76922
rect 209782 76864 209830 76920
rect 209886 76864 209891 76920
rect 209782 76859 209891 76864
rect 99517 76786 99583 76789
rect 95702 76784 99583 76786
rect 95702 76728 99522 76784
rect 99578 76728 99583 76784
rect 95702 76726 99583 76728
rect 99517 76723 99583 76726
rect 191977 76786 192043 76789
rect 191977 76784 193988 76786
rect 191977 76728 191982 76784
rect 192038 76728 193988 76784
rect 191977 76726 193988 76728
rect 191977 76723 192043 76726
rect 25590 76452 25596 76516
rect 25660 76514 25666 76516
rect 25660 76454 25996 76514
rect 25660 76452 25666 76454
rect 41782 76452 41788 76516
rect 41852 76514 41858 76516
rect 44409 76514 44475 76517
rect 41852 76512 44475 76514
rect 41852 76456 44414 76512
rect 44470 76456 44475 76512
rect 209782 76484 209842 76859
rect 41852 76454 44475 76456
rect 41852 76452 41858 76454
rect 44409 76451 44475 76454
rect 183237 76106 183303 76109
rect 179820 76104 183303 76106
rect 179820 76048 183242 76104
rect 183298 76048 183303 76104
rect 95702 75562 95762 76048
rect 179820 76046 183303 76048
rect 183237 76043 183303 76046
rect 98229 75562 98295 75565
rect 95702 75560 98295 75562
rect 95702 75504 98234 75560
rect 98290 75504 98295 75560
rect 95702 75502 98295 75504
rect 98229 75499 98295 75502
rect 106785 75018 106851 75021
rect 106785 75016 109900 75018
rect 106785 74960 106790 75016
rect 106846 74960 109900 75016
rect 106785 74958 109900 74960
rect 106785 74955 106851 74958
rect 183697 74882 183763 74885
rect 179820 74880 183763 74882
rect 179820 74824 183702 74880
rect 183758 74824 183763 74880
rect 44409 74746 44475 74749
rect 41820 74744 44475 74746
rect 41820 74688 44414 74744
rect 44470 74688 44475 74744
rect 41820 74686 44475 74688
rect 44409 74683 44475 74686
rect 95702 74338 95762 74824
rect 179820 74822 183763 74824
rect 183697 74819 183763 74822
rect 191517 74746 191583 74749
rect 191517 74744 193988 74746
rect 191517 74688 191522 74744
rect 191578 74688 193988 74744
rect 191517 74686 193988 74688
rect 191517 74683 191583 74686
rect 99425 74338 99491 74341
rect 95702 74336 99491 74338
rect 95702 74280 99430 74336
rect 99486 74280 99491 74336
rect 95702 74278 99491 74280
rect 99425 74275 99491 74278
rect 222337 74338 222403 74341
rect 225416 74338 225896 74368
rect 222337 74336 225896 74338
rect 222337 74280 222342 74336
rect 222398 74280 225896 74336
rect 222337 74278 225896 74280
rect 222337 74275 222403 74278
rect 225416 74248 225896 74278
rect 99517 73794 99583 73797
rect 183697 73794 183763 73797
rect 95732 73792 99583 73794
rect 95732 73736 99522 73792
rect 99578 73736 99583 73792
rect 95732 73734 99583 73736
rect 179820 73792 183763 73794
rect 179820 73736 183702 73792
rect 183758 73736 183763 73792
rect 179820 73734 183763 73736
rect 99517 73731 99583 73734
rect 183697 73731 183763 73734
rect 191977 72842 192043 72845
rect 191977 72840 193988 72842
rect 191977 72784 191982 72840
rect 192038 72784 193988 72840
rect 191977 72782 193988 72784
rect 191977 72779 192043 72782
rect 106785 72706 106851 72709
rect 106785 72704 109900 72706
rect 106785 72648 106790 72704
rect 106846 72648 109900 72704
rect 106785 72646 109900 72648
rect 106785 72643 106851 72646
rect 99517 72570 99583 72573
rect 183697 72570 183763 72573
rect 95732 72568 99583 72570
rect 95732 72512 99522 72568
rect 99578 72512 99583 72568
rect 95732 72510 99583 72512
rect 179820 72568 183763 72570
rect 179820 72512 183702 72568
rect 183758 72512 183763 72568
rect 179820 72510 183763 72512
rect 99517 72507 99583 72510
rect 183697 72507 183763 72510
rect 183697 71346 183763 71349
rect 179820 71344 183763 71346
rect 179820 71288 183702 71344
rect 183758 71288 183763 71344
rect 95702 71074 95762 71288
rect 179820 71286 183763 71288
rect 183697 71283 183763 71286
rect 99517 71074 99583 71077
rect 95702 71072 99583 71074
rect 95702 71016 99522 71072
rect 99578 71016 99583 71072
rect 95702 71014 99583 71016
rect 99517 71011 99583 71014
rect 190781 70802 190847 70805
rect 190781 70800 193988 70802
rect 190781 70744 190786 70800
rect 190842 70744 193988 70800
rect 190781 70742 193988 70744
rect 190781 70739 190847 70742
rect 106693 70394 106759 70397
rect 106693 70392 109900 70394
rect 106693 70336 106698 70392
rect 106754 70336 109900 70392
rect 106693 70334 109900 70336
rect 106693 70331 106759 70334
rect 182869 70122 182935 70125
rect 179820 70120 182935 70122
rect 179820 70064 182874 70120
rect 182930 70064 182935 70120
rect 25774 69516 25780 69580
rect 25844 69578 25850 69580
rect 25966 69578 26026 69820
rect 41782 69788 41788 69852
rect 41852 69850 41858 69852
rect 53333 69850 53399 69853
rect 41852 69848 53399 69850
rect 41852 69792 53338 69848
rect 53394 69792 53399 69848
rect 41852 69790 53399 69792
rect 95702 69850 95762 70064
rect 179820 70062 182935 70064
rect 182869 70059 182935 70062
rect 99517 69850 99583 69853
rect 128497 69850 128563 69853
rect 211430 69850 211436 69852
rect 95702 69848 99583 69850
rect 95702 69792 99522 69848
rect 99578 69792 99583 69848
rect 95702 69790 99583 69792
rect 125724 69848 128563 69850
rect 125724 69792 128502 69848
rect 128558 69792 128563 69848
rect 125724 69790 128563 69792
rect 209812 69790 211436 69850
rect 41852 69788 41858 69790
rect 53333 69787 53399 69790
rect 99517 69787 99583 69790
rect 128497 69787 128563 69790
rect 211430 69788 211436 69790
rect 211500 69788 211506 69852
rect 25844 69518 26026 69578
rect 25844 69516 25850 69518
rect 183053 68898 183119 68901
rect 179820 68896 183119 68898
rect 179820 68840 183058 68896
rect 183114 68840 183119 68896
rect 95702 68354 95762 68840
rect 179820 68838 183119 68840
rect 183053 68835 183119 68838
rect 190965 68762 191031 68765
rect 190965 68760 193988 68762
rect 190965 68704 190970 68760
rect 191026 68704 193988 68760
rect 190965 68702 193988 68704
rect 190965 68699 191031 68702
rect 98965 68354 99031 68357
rect 95702 68352 99031 68354
rect 95702 68296 98970 68352
rect 99026 68296 99031 68352
rect 95702 68294 99031 68296
rect 98965 68291 99031 68294
rect 106601 67946 106667 67949
rect 106601 67944 109900 67946
rect 106601 67888 106606 67944
rect 106662 67888 109900 67944
rect 106601 67886 109900 67888
rect 106601 67883 106667 67886
rect 9896 67810 10376 67840
rect 13313 67810 13379 67813
rect 9896 67808 13379 67810
rect 9896 67752 13318 67808
rect 13374 67752 13379 67808
rect 9896 67750 13379 67752
rect 9896 67720 10376 67750
rect 13313 67747 13379 67750
rect 183145 67674 183211 67677
rect 179820 67672 183211 67674
rect 179820 67616 183150 67672
rect 183206 67616 183211 67672
rect 95702 67130 95762 67616
rect 179820 67614 183211 67616
rect 183145 67611 183211 67614
rect 99057 67130 99123 67133
rect 95702 67128 99123 67130
rect 95702 67072 99062 67128
rect 99118 67072 99123 67128
rect 95702 67070 99123 67072
rect 99057 67067 99123 67070
rect 191333 66858 191399 66861
rect 191333 66856 193988 66858
rect 191333 66800 191338 66856
rect 191394 66800 193988 66856
rect 191333 66798 193988 66800
rect 191333 66795 191399 66798
rect 53425 66586 53491 66589
rect 53977 66586 54043 66589
rect 136869 66586 136935 66589
rect 53425 66584 55988 66586
rect 53425 66528 53430 66584
rect 53486 66528 53982 66584
rect 54038 66528 55988 66584
rect 53425 66526 55988 66528
rect 136869 66584 140076 66586
rect 136869 66528 136874 66584
rect 136930 66528 140076 66584
rect 136869 66526 140076 66528
rect 53425 66523 53491 66526
rect 53977 66523 54043 66526
rect 136869 66523 136935 66526
rect 183237 66450 183303 66453
rect 179820 66448 183303 66450
rect 179820 66392 183242 66448
rect 183298 66392 183303 66448
rect 95702 65906 95762 66392
rect 179820 66390 183303 66392
rect 183237 66387 183303 66390
rect 99149 65906 99215 65909
rect 95702 65904 99215 65906
rect 95702 65848 99154 65904
rect 99210 65848 99215 65904
rect 95702 65846 99215 65848
rect 99149 65843 99215 65846
rect 106509 65634 106575 65637
rect 106509 65632 109900 65634
rect 106509 65576 106514 65632
rect 106570 65576 109900 65632
rect 106509 65574 109900 65576
rect 106509 65571 106575 65574
rect 183329 65226 183395 65229
rect 179820 65224 183395 65226
rect 179820 65168 183334 65224
rect 183390 65168 183395 65224
rect 44501 64818 44567 64821
rect 41820 64816 44567 64818
rect 41820 64760 44506 64816
rect 44562 64760 44567 64816
rect 41820 64758 44567 64760
rect 44501 64755 44567 64758
rect 95702 64682 95762 65168
rect 179820 65166 183395 65168
rect 183329 65163 183395 65166
rect 191517 64818 191583 64821
rect 191517 64816 193988 64818
rect 191517 64760 191522 64816
rect 191578 64760 193988 64816
rect 191517 64758 193988 64760
rect 191517 64755 191583 64758
rect 99241 64682 99307 64685
rect 95702 64680 99307 64682
rect 95702 64624 99246 64680
rect 99302 64624 99307 64680
rect 95702 64622 99307 64624
rect 99241 64619 99307 64622
rect 183421 64002 183487 64005
rect 179820 64000 183487 64002
rect 179820 63944 183426 64000
rect 183482 63944 183487 64000
rect 95702 63458 95762 63944
rect 179820 63942 183487 63944
rect 183421 63939 183487 63942
rect 99333 63458 99399 63461
rect 95702 63456 99399 63458
rect 95702 63400 99338 63456
rect 99394 63400 99399 63456
rect 95702 63398 99399 63400
rect 99333 63395 99399 63398
rect 106601 63322 106667 63325
rect 106601 63320 109900 63322
rect 106601 63264 106606 63320
rect 106662 63264 109900 63320
rect 106601 63262 109900 63264
rect 106601 63259 106667 63262
rect 22329 63186 22395 63189
rect 211614 63186 211620 63188
rect 22329 63184 25996 63186
rect 22329 63128 22334 63184
rect 22390 63128 25996 63184
rect 22329 63126 25996 63128
rect 209812 63126 211620 63186
rect 22329 63123 22395 63126
rect 211614 63124 211620 63126
rect 211684 63186 211690 63188
rect 212677 63186 212743 63189
rect 211684 63184 212743 63186
rect 211684 63128 212682 63184
rect 212738 63128 212743 63184
rect 211684 63126 212743 63128
rect 211684 63124 211690 63126
rect 212677 63123 212743 63126
rect 98781 62778 98847 62781
rect 183605 62778 183671 62781
rect 95732 62776 98847 62778
rect 95732 62720 98786 62776
rect 98842 62720 98847 62776
rect 95732 62718 98847 62720
rect 179820 62776 183671 62778
rect 179820 62720 183610 62776
rect 183666 62720 183671 62776
rect 179820 62718 183671 62720
rect 98781 62715 98847 62718
rect 183605 62715 183671 62718
rect 189953 62778 190019 62781
rect 189953 62776 193988 62778
rect 189953 62720 189958 62776
rect 190014 62720 193988 62776
rect 189953 62718 193988 62720
rect 189953 62715 190019 62718
rect 99517 61554 99583 61557
rect 183697 61554 183763 61557
rect 95732 61552 99583 61554
rect 95732 61496 99522 61552
rect 99578 61496 99583 61552
rect 95732 61494 99583 61496
rect 179820 61552 183763 61554
rect 179820 61496 183702 61552
rect 183758 61496 183763 61552
rect 179820 61494 183763 61496
rect 99517 61491 99583 61494
rect 183697 61491 183763 61494
rect 107153 61010 107219 61013
rect 107153 61008 109900 61010
rect 107153 60952 107158 61008
rect 107214 60952 109900 61008
rect 107153 60950 109900 60952
rect 107153 60947 107219 60950
rect 191977 60874 192043 60877
rect 191977 60872 193988 60874
rect 191977 60816 191982 60872
rect 192038 60816 193988 60872
rect 191977 60814 193988 60816
rect 191977 60811 192043 60814
rect 182685 60466 182751 60469
rect 179820 60464 182751 60466
rect 179820 60408 182690 60464
rect 182746 60408 182751 60464
rect 95702 60058 95762 60408
rect 179820 60406 182751 60408
rect 182685 60403 182751 60406
rect 99517 60058 99583 60061
rect 95702 60056 99583 60058
rect 95702 60000 99522 60056
rect 99578 60000 99583 60056
rect 95702 59998 99583 60000
rect 99517 59995 99583 59998
rect 59221 58426 59287 58429
rect 140222 58426 140228 58428
rect 59221 58424 140228 58426
rect 59221 58368 59226 58424
rect 59282 58368 140228 58424
rect 59221 58366 140228 58368
rect 59221 58363 59287 58366
rect 140222 58364 140228 58366
rect 140292 58364 140298 58428
rect 222245 48090 222311 48093
rect 225416 48090 225896 48120
rect 222245 48088 225896 48090
rect 222245 48032 222250 48088
rect 222306 48032 225896 48088
rect 222245 48030 225896 48032
rect 222245 48027 222311 48030
rect 225416 48000 225896 48030
rect 152734 46940 152740 47004
rect 152804 47002 152810 47004
rect 164745 47002 164811 47005
rect 152804 47000 164811 47002
rect 152804 46944 164750 47000
rect 164806 46944 164811 47000
rect 152804 46942 164811 46944
rect 152804 46940 152810 46942
rect 164745 46939 164811 46942
rect 68830 46804 68836 46868
rect 68900 46866 68906 46868
rect 80749 46866 80815 46869
rect 68900 46864 80815 46866
rect 68900 46808 80754 46864
rect 80810 46808 80815 46864
rect 68900 46806 80815 46808
rect 68900 46804 68906 46806
rect 80749 46803 80815 46806
rect 149054 46804 149060 46868
rect 149124 46866 149130 46868
rect 161893 46866 161959 46869
rect 149124 46864 161959 46866
rect 149124 46808 161898 46864
rect 161954 46808 161959 46864
rect 149124 46806 161959 46808
rect 149124 46804 149130 46806
rect 161893 46803 161959 46806
rect 64966 46668 64972 46732
rect 65036 46730 65042 46732
rect 77805 46730 77871 46733
rect 65036 46728 77871 46730
rect 65036 46672 77810 46728
rect 77866 46672 77871 46728
rect 65036 46670 77871 46672
rect 65036 46668 65042 46670
rect 77805 46667 77871 46670
rect 146294 46668 146300 46732
rect 146364 46730 146370 46732
rect 158949 46730 159015 46733
rect 146364 46728 159015 46730
rect 146364 46672 158954 46728
rect 159010 46672 159015 46728
rect 146364 46670 159015 46672
rect 146364 46668 146370 46670
rect 158949 46667 159015 46670
rect 68462 46532 68468 46596
rect 68532 46594 68538 46596
rect 79277 46594 79343 46597
rect 68532 46592 79343 46594
rect 68532 46536 79282 46592
rect 79338 46536 79343 46592
rect 68532 46534 79343 46536
rect 68532 46532 68538 46534
rect 79277 46531 79343 46534
rect 101357 46594 101423 46597
rect 101357 46592 104042 46594
rect 101357 46536 101362 46592
rect 101418 46536 104042 46592
rect 101357 46534 104042 46536
rect 101357 46531 101423 46534
rect 103982 46500 104042 46534
rect 152550 46532 152556 46596
rect 152620 46594 152626 46596
rect 163273 46594 163339 46597
rect 152620 46592 163339 46594
rect 152620 46536 163278 46592
rect 163334 46536 163339 46592
rect 152620 46534 163339 46536
rect 152620 46532 152626 46534
rect 163273 46531 163339 46534
rect 63494 46396 63500 46460
rect 63564 46458 63570 46460
rect 74861 46458 74927 46461
rect 63564 46456 74927 46458
rect 63564 46400 74866 46456
rect 74922 46400 74927 46456
rect 63564 46398 74927 46400
rect 63564 46396 63570 46398
rect 74861 46395 74927 46398
rect 49929 46322 49995 46325
rect 47862 46320 49995 46322
rect 47862 46264 49934 46320
rect 49990 46264 49995 46320
rect 47862 46262 49995 46264
rect 47862 46224 47922 46262
rect 49929 46259 49995 46262
rect 62206 46260 62212 46324
rect 62276 46322 62282 46324
rect 73389 46322 73455 46325
rect 62276 46320 73455 46322
rect 62276 46264 73394 46320
rect 73450 46264 73455 46320
rect 62276 46262 73455 46264
rect 62276 46260 62282 46262
rect 73389 46259 73455 46262
rect 85717 46322 85783 46325
rect 89806 46322 89812 46324
rect 85717 46320 89812 46322
rect 85717 46264 85722 46320
rect 85778 46264 89812 46320
rect 85717 46262 89812 46264
rect 85717 46259 85783 46262
rect 89806 46260 89812 46262
rect 89876 46260 89882 46324
rect 131766 46322 131826 46496
rect 147766 46396 147772 46460
rect 147836 46458 147842 46460
rect 160329 46458 160395 46461
rect 147836 46456 160395 46458
rect 147836 46400 160334 46456
rect 160390 46400 160395 46456
rect 147836 46398 160395 46400
rect 147836 46396 147842 46398
rect 160329 46395 160395 46398
rect 135397 46322 135463 46325
rect 131766 46320 135463 46322
rect 131766 46264 135402 46320
rect 135458 46264 135463 46320
rect 131766 46262 135463 46264
rect 135397 46259 135463 46262
rect 146110 46260 146116 46324
rect 146180 46322 146186 46324
rect 157569 46322 157635 46325
rect 146180 46320 157635 46322
rect 146180 46264 157574 46320
rect 157630 46264 157635 46320
rect 146180 46262 157635 46264
rect 146180 46260 146186 46262
rect 157569 46259 157635 46262
rect 63310 46124 63316 46188
rect 63380 46186 63386 46188
rect 76333 46186 76399 46189
rect 63380 46184 76399 46186
rect 63380 46128 76338 46184
rect 76394 46128 76399 46184
rect 63380 46126 76399 46128
rect 63380 46124 63386 46126
rect 76333 46123 76399 46126
rect 87097 46186 87163 46189
rect 89070 46186 89076 46188
rect 87097 46184 89076 46186
rect 87097 46128 87102 46184
rect 87158 46128 89076 46184
rect 87097 46126 89076 46128
rect 87097 46123 87163 46126
rect 89070 46124 89076 46126
rect 89140 46124 89146 46188
rect 147030 46124 147036 46188
rect 147100 46186 147106 46188
rect 154257 46186 154323 46189
rect 147100 46184 154323 46186
rect 147100 46128 154262 46184
rect 154318 46128 154323 46184
rect 147100 46126 154323 46128
rect 147100 46124 147106 46126
rect 154257 46123 154323 46126
rect 169897 46186 169963 46189
rect 172974 46186 172980 46188
rect 169897 46184 172980 46186
rect 169897 46128 169902 46184
rect 169958 46128 172980 46184
rect 169897 46126 172980 46128
rect 169897 46123 169963 46126
rect 172974 46124 172980 46126
rect 173044 46124 173050 46188
rect 185905 46186 185971 46189
rect 187886 46186 187946 46496
rect 185905 46184 187946 46186
rect 185905 46128 185910 46184
rect 185966 46128 187946 46184
rect 185905 46126 187946 46128
rect 185905 46123 185971 46126
rect 103430 45922 104012 45982
rect 101725 45914 101791 45917
rect 103430 45914 103490 45922
rect 101725 45912 103490 45914
rect 101725 45856 101730 45912
rect 101786 45856 103490 45912
rect 101725 45854 103490 45856
rect 101725 45851 101791 45854
rect 47862 45234 47922 45680
rect 131766 45506 131826 45952
rect 135397 45506 135463 45509
rect 131766 45504 135463 45506
rect 131766 45448 135402 45504
rect 135458 45448 135463 45504
rect 131766 45446 135463 45448
rect 135397 45443 135463 45446
rect 185169 45506 185235 45509
rect 187886 45506 187946 45952
rect 185169 45504 187946 45506
rect 185169 45448 185174 45504
rect 185230 45448 187946 45504
rect 185169 45446 187946 45448
rect 185169 45443 185235 45446
rect 103430 45242 104012 45302
rect 53333 45234 53399 45237
rect 47862 45232 53399 45234
rect 47862 45176 53338 45232
rect 53394 45176 53399 45232
rect 47862 45174 53399 45176
rect 53333 45171 53399 45174
rect 101817 45234 101883 45237
rect 103430 45234 103490 45242
rect 101817 45232 103490 45234
rect 101817 45176 101822 45232
rect 101878 45176 103490 45232
rect 101817 45174 103490 45176
rect 101817 45171 101883 45174
rect 131766 45098 131826 45272
rect 135397 45098 135463 45101
rect 131766 45096 135463 45098
rect 131766 45040 135402 45096
rect 135458 45040 135463 45096
rect 131766 45038 135463 45040
rect 135397 45035 135463 45038
rect 47862 44962 47922 45000
rect 53241 44962 53307 44965
rect 47862 44960 53307 44962
rect 47862 44904 53246 44960
rect 53302 44904 53307 44960
rect 47862 44902 53307 44904
rect 53241 44899 53307 44902
rect 185813 44962 185879 44965
rect 187886 44962 187946 45272
rect 185813 44960 187946 44962
rect 185813 44904 185818 44960
rect 185874 44904 187946 44960
rect 185813 44902 187946 44904
rect 185813 44899 185879 44902
rect 101265 44826 101331 44829
rect 135397 44826 135463 44829
rect 101265 44824 103490 44826
rect 101265 44768 101270 44824
rect 101326 44768 103490 44824
rect 101265 44766 103490 44768
rect 101265 44763 101331 44766
rect 103430 44762 103490 44766
rect 131766 44824 135463 44826
rect 131766 44768 135402 44824
rect 135458 44768 135463 44824
rect 131766 44766 135463 44768
rect 103430 44702 104012 44762
rect 131766 44728 131826 44766
rect 135397 44763 135463 44766
rect 171369 44826 171435 44829
rect 173342 44826 173348 44828
rect 171369 44824 173348 44826
rect 171369 44768 171374 44824
rect 171430 44768 173348 44824
rect 171369 44766 173348 44768
rect 171369 44763 171435 44766
rect 173342 44764 173348 44766
rect 173412 44764 173418 44828
rect 185445 44826 185511 44829
rect 185445 44824 187946 44826
rect 185445 44768 185450 44824
rect 185506 44768 187946 44824
rect 185445 44766 187946 44768
rect 185445 44763 185511 44766
rect 187886 44728 187946 44766
rect 143677 44690 143743 44693
rect 172933 44690 172999 44693
rect 173894 44690 173900 44692
rect 143677 44688 145074 44690
rect 143677 44632 143682 44688
rect 143738 44632 145074 44688
rect 143677 44630 145074 44632
rect 143677 44627 143743 44630
rect 145014 44456 145074 44630
rect 172933 44688 173900 44690
rect 172933 44632 172938 44688
rect 172994 44632 173900 44688
rect 172933 44630 173900 44632
rect 172933 44627 172999 44630
rect 173894 44628 173900 44630
rect 173964 44628 173970 44692
rect 9896 44146 10376 44176
rect 13405 44146 13471 44149
rect 9896 44144 13471 44146
rect 9896 44088 13410 44144
rect 13466 44088 13471 44144
rect 9896 44086 13471 44088
rect 9896 44056 10376 44086
rect 13405 44083 13471 44086
rect 47862 44010 47922 44456
rect 58945 44418 59011 44421
rect 92709 44418 92775 44421
rect 177717 44418 177783 44421
rect 58945 44416 60956 44418
rect 58945 44360 58950 44416
rect 59006 44360 60956 44416
rect 58945 44358 60956 44360
rect 90764 44416 92775 44418
rect 90764 44360 92714 44416
rect 92770 44360 92775 44416
rect 90764 44358 92775 44360
rect 174852 44416 177783 44418
rect 174852 44360 177722 44416
rect 177778 44360 177783 44416
rect 174852 44358 177783 44360
rect 58945 44355 59011 44358
rect 92709 44355 92775 44358
rect 177717 44355 177783 44358
rect 92801 44282 92867 44285
rect 90734 44280 92867 44282
rect 90734 44224 92806 44280
rect 92862 44224 92867 44280
rect 90734 44222 92867 44224
rect 50021 44010 50087 44013
rect 47862 44008 50087 44010
rect 47862 43952 50026 44008
rect 50082 43952 50087 44008
rect 47862 43950 50087 43952
rect 50021 43947 50087 43950
rect 90734 43912 90794 44222
rect 92801 44219 92867 44222
rect 143493 44146 143559 44149
rect 143493 44144 145074 44146
rect 143493 44088 143498 44144
rect 143554 44088 145074 44144
rect 143493 44086 145074 44088
rect 143493 44083 143559 44086
rect 103430 44018 104012 44078
rect 101633 44010 101699 44013
rect 103430 44010 103490 44018
rect 101633 44008 103490 44010
rect 101633 43952 101638 44008
rect 101694 43952 103490 44008
rect 101633 43950 103490 43952
rect 101633 43947 101699 43950
rect 58209 43874 58275 43877
rect 58209 43872 60956 43874
rect 58209 43816 58214 43872
rect 58270 43816 60956 43872
rect 58209 43814 60956 43816
rect 58209 43811 58275 43814
rect 47862 43602 47922 43776
rect 131766 43738 131826 44048
rect 145014 43912 145074 44086
rect 177717 43874 177783 43877
rect 174852 43872 177783 43874
rect 174852 43816 177722 43872
rect 177778 43816 177783 43872
rect 174852 43814 177783 43816
rect 177717 43811 177783 43814
rect 135397 43738 135463 43741
rect 131766 43736 135463 43738
rect 131766 43680 135402 43736
rect 135458 43680 135463 43736
rect 131766 43678 135463 43680
rect 135397 43675 135463 43678
rect 185169 43738 185235 43741
rect 187886 43738 187946 44048
rect 185169 43736 187946 43738
rect 185169 43680 185174 43736
rect 185230 43680 187946 43736
rect 185169 43678 187946 43680
rect 185169 43675 185235 43678
rect 49929 43602 49995 43605
rect 47862 43600 49995 43602
rect 47862 43544 49934 43600
rect 49990 43544 49995 43600
rect 47862 43542 49995 43544
rect 49929 43539 49995 43542
rect 103430 43474 104012 43534
rect 100805 43466 100871 43469
rect 103430 43466 103490 43474
rect 100805 43464 103490 43466
rect 100805 43408 100810 43464
rect 100866 43408 103490 43464
rect 100805 43406 103490 43408
rect 131766 43466 131826 43504
rect 135213 43466 135279 43469
rect 131766 43464 135279 43466
rect 131766 43408 135218 43464
rect 135274 43408 135279 43464
rect 131766 43406 135279 43408
rect 100805 43403 100871 43406
rect 135213 43403 135279 43406
rect 184985 43466 185051 43469
rect 187886 43466 187946 43504
rect 184985 43464 187946 43466
rect 184985 43408 184990 43464
rect 185046 43408 187946 43464
rect 184985 43406 187946 43408
rect 184985 43403 185051 43406
rect 142297 43330 142363 43333
rect 142297 43328 144522 43330
rect 142297 43272 142302 43328
rect 142358 43272 144522 43328
rect 142297 43270 144522 43272
rect 142297 43267 142363 43270
rect 144462 43262 144522 43270
rect 47862 42786 47922 43232
rect 144462 43202 145044 43262
rect 59037 43194 59103 43197
rect 92709 43194 92775 43197
rect 177717 43194 177783 43197
rect 59037 43192 60956 43194
rect 59037 43136 59042 43192
rect 59098 43136 60956 43192
rect 59037 43134 60956 43136
rect 90764 43192 92775 43194
rect 90764 43136 92714 43192
rect 92770 43136 92775 43192
rect 90764 43134 92775 43136
rect 174852 43192 177783 43194
rect 174852 43136 177722 43192
rect 177778 43136 177783 43192
rect 174852 43134 177783 43136
rect 59037 43131 59103 43134
rect 92709 43131 92775 43134
rect 177717 43131 177783 43134
rect 142205 43058 142271 43061
rect 142205 43056 145074 43058
rect 142205 43000 142210 43056
rect 142266 43000 145074 43056
rect 142205 42998 145074 43000
rect 142205 42995 142271 42998
rect 92893 42922 92959 42925
rect 90734 42920 92959 42922
rect 90734 42864 92898 42920
rect 92954 42864 92959 42920
rect 90734 42862 92959 42864
rect 50021 42786 50087 42789
rect 47862 42784 50087 42786
rect 47862 42728 50026 42784
rect 50082 42728 50087 42784
rect 47862 42726 50087 42728
rect 50021 42723 50087 42726
rect 90734 42688 90794 42862
rect 92893 42859 92959 42862
rect 103430 42794 104012 42854
rect 101725 42786 101791 42789
rect 103430 42786 103490 42794
rect 101725 42784 103490 42786
rect 101725 42728 101730 42784
rect 101786 42728 103490 42784
rect 101725 42726 103490 42728
rect 101725 42723 101791 42726
rect 58209 42650 58275 42653
rect 58209 42648 60956 42650
rect 58209 42592 58214 42648
rect 58270 42592 60956 42648
rect 58209 42590 60956 42592
rect 58209 42587 58275 42590
rect 47862 42514 47922 42552
rect 49929 42514 49995 42517
rect 92801 42514 92867 42517
rect 47862 42512 49995 42514
rect 47862 42456 49934 42512
rect 49990 42456 49995 42512
rect 47862 42454 49995 42456
rect 49929 42451 49995 42454
rect 90734 42512 92867 42514
rect 90734 42456 92806 42512
rect 92862 42456 92867 42512
rect 90734 42454 92867 42456
rect 131766 42514 131826 42824
rect 145014 42688 145074 42998
rect 177809 42650 177875 42653
rect 174852 42648 177875 42650
rect 174852 42592 177814 42648
rect 177870 42592 177875 42648
rect 174852 42590 177875 42592
rect 177809 42587 177875 42590
rect 135397 42514 135463 42517
rect 131766 42512 135463 42514
rect 131766 42456 135402 42512
rect 135458 42456 135463 42512
rect 131766 42454 135463 42456
rect 90734 42144 90794 42454
rect 92801 42451 92867 42454
rect 135397 42451 135463 42454
rect 142757 42514 142823 42517
rect 185169 42514 185235 42517
rect 187886 42514 187946 42824
rect 142757 42512 145074 42514
rect 142757 42456 142762 42512
rect 142818 42456 145074 42512
rect 142757 42454 145074 42456
rect 142757 42451 142823 42454
rect 103430 42250 104012 42310
rect 100897 42242 100963 42245
rect 103430 42242 103490 42250
rect 100897 42240 103490 42242
rect 100897 42184 100902 42240
rect 100958 42184 103490 42240
rect 100897 42182 103490 42184
rect 131766 42242 131826 42280
rect 135213 42242 135279 42245
rect 131766 42240 135279 42242
rect 131766 42184 135218 42240
rect 135274 42184 135279 42240
rect 131766 42182 135279 42184
rect 100897 42179 100963 42182
rect 135213 42179 135279 42182
rect 145014 42144 145074 42454
rect 185169 42512 187946 42514
rect 185169 42456 185174 42512
rect 185230 42456 187946 42512
rect 185169 42454 187946 42456
rect 185169 42451 185235 42454
rect 49929 42106 49995 42109
rect 47862 42104 49995 42106
rect 47862 42048 49934 42104
rect 49990 42048 49995 42104
rect 47862 42046 49995 42048
rect 47862 42008 47922 42046
rect 49929 42043 49995 42046
rect 58301 42106 58367 42109
rect 177717 42106 177783 42109
rect 58301 42104 60956 42106
rect 58301 42048 58306 42104
rect 58362 42048 60956 42104
rect 58301 42046 60956 42048
rect 174852 42104 177783 42106
rect 174852 42048 177722 42104
rect 177778 42048 177783 42104
rect 174852 42046 177783 42048
rect 58301 42043 58367 42046
rect 177717 42043 177783 42046
rect 185077 42106 185143 42109
rect 187886 42106 187946 42280
rect 185077 42104 187946 42106
rect 185077 42048 185082 42104
rect 185138 42048 187946 42104
rect 185077 42046 187946 42048
rect 185077 42043 185143 42046
rect 18097 41970 18163 41973
rect 18097 41968 19402 41970
rect 18097 41912 18102 41968
rect 18158 41912 19402 41968
rect 18097 41910 19402 41912
rect 18097 41907 18163 41910
rect 19342 41902 19402 41910
rect 19342 41842 19924 41902
rect 143401 41834 143467 41837
rect 143401 41832 145074 41834
rect 143401 41776 143406 41832
rect 143462 41776 145074 41832
rect 143401 41774 145074 41776
rect 143401 41771 143467 41774
rect 92709 41698 92775 41701
rect 90734 41696 92775 41698
rect 90734 41640 92714 41696
rect 92770 41640 92775 41696
rect 90734 41638 92775 41640
rect 90734 41464 90794 41638
rect 92709 41635 92775 41638
rect 103430 41570 104012 41630
rect 100989 41562 101055 41565
rect 103430 41562 103490 41570
rect 100989 41560 103490 41562
rect 100989 41504 100994 41560
rect 101050 41504 103490 41560
rect 100989 41502 103490 41504
rect 100989 41499 101055 41502
rect 58209 41426 58275 41429
rect 58209 41424 60956 41426
rect 58209 41368 58214 41424
rect 58270 41368 60956 41424
rect 58209 41366 60956 41368
rect 58209 41363 58275 41366
rect 47862 41018 47922 41328
rect 131766 41290 131826 41600
rect 145014 41464 145074 41774
rect 177717 41426 177783 41429
rect 174852 41424 177783 41426
rect 174852 41368 177722 41424
rect 177778 41368 177783 41424
rect 174852 41366 177783 41368
rect 177717 41363 177783 41366
rect 135397 41290 135463 41293
rect 131766 41288 135463 41290
rect 131766 41232 135402 41288
rect 135458 41232 135463 41288
rect 131766 41230 135463 41232
rect 135397 41227 135463 41230
rect 143309 41290 143375 41293
rect 185169 41290 185235 41293
rect 187886 41290 187946 41600
rect 143309 41288 145074 41290
rect 143309 41232 143314 41288
rect 143370 41232 145074 41288
rect 143309 41230 145074 41232
rect 143309 41227 143375 41230
rect 92801 41154 92867 41157
rect 90734 41152 92867 41154
rect 90734 41096 92806 41152
rect 92862 41096 92867 41152
rect 90734 41094 92867 41096
rect 50021 41018 50087 41021
rect 47862 41016 50087 41018
rect 47862 40960 50026 41016
rect 50082 40960 50087 41016
rect 47862 40958 50087 40960
rect 50021 40955 50087 40958
rect 90734 40920 90794 41094
rect 92801 41091 92867 41094
rect 103430 41026 104012 41086
rect 100805 41018 100871 41021
rect 103430 41018 103490 41026
rect 100805 41016 103490 41018
rect 100805 40960 100810 41016
rect 100866 40960 103490 41016
rect 100805 40958 103490 40960
rect 100805 40955 100871 40958
rect 58301 40882 58367 40885
rect 131766 40882 131826 41056
rect 145014 40920 145074 41230
rect 185169 41288 187946 41290
rect 185169 41232 185174 41288
rect 185230 41232 187946 41288
rect 185169 41230 187946 41232
rect 185169 41227 185235 41230
rect 135213 40882 135279 40885
rect 177625 40882 177691 40885
rect 58301 40880 60956 40882
rect 58301 40824 58306 40880
rect 58362 40824 60956 40880
rect 58301 40822 60956 40824
rect 131766 40880 135279 40882
rect 131766 40824 135218 40880
rect 135274 40824 135279 40880
rect 131766 40822 135279 40824
rect 174852 40880 177691 40882
rect 174852 40824 177630 40880
rect 177686 40824 177691 40880
rect 174852 40822 177691 40824
rect 58301 40819 58367 40822
rect 135213 40819 135279 40822
rect 177625 40819 177691 40822
rect 47862 40746 47922 40784
rect 49929 40746 49995 40749
rect 47862 40744 49995 40746
rect 47862 40688 49934 40744
rect 49990 40688 49995 40744
rect 47862 40686 49995 40688
rect 49929 40683 49995 40686
rect 184985 40610 185051 40613
rect 187886 40610 187946 41056
rect 184985 40608 187946 40610
rect 184985 40552 184990 40608
rect 185046 40552 187946 40608
rect 184985 40550 187946 40552
rect 184985 40547 185051 40550
rect 143677 40474 143743 40477
rect 143677 40472 145074 40474
rect 143677 40416 143682 40472
rect 143738 40416 145074 40472
rect 143677 40414 145074 40416
rect 143677 40411 143743 40414
rect 103430 40346 104012 40406
rect 101081 40338 101147 40341
rect 103430 40338 103490 40346
rect 101081 40336 103490 40338
rect 101081 40280 101086 40336
rect 101142 40280 103490 40336
rect 101081 40278 103490 40280
rect 101081 40275 101147 40278
rect 58393 40202 58459 40205
rect 92709 40202 92775 40205
rect 58393 40200 60956 40202
rect 58393 40144 58398 40200
rect 58454 40144 60956 40200
rect 58393 40142 60956 40144
rect 90764 40200 92775 40202
rect 90764 40144 92714 40200
rect 92770 40144 92775 40200
rect 90764 40142 92775 40144
rect 58393 40139 58459 40142
rect 92709 40139 92775 40142
rect 47862 39794 47922 40104
rect 92801 40066 92867 40069
rect 90734 40064 92867 40066
rect 90734 40008 92806 40064
rect 92862 40008 92867 40064
rect 90734 40006 92867 40008
rect 131766 40066 131826 40376
rect 145014 40240 145074 40414
rect 177717 40202 177783 40205
rect 174852 40200 177783 40202
rect 174852 40144 177722 40200
rect 177778 40144 177783 40200
rect 174852 40142 177783 40144
rect 177717 40139 177783 40142
rect 135213 40066 135279 40069
rect 131766 40064 135279 40066
rect 131766 40008 135218 40064
rect 135274 40008 135279 40064
rect 131766 40006 135279 40008
rect 51125 39794 51191 39797
rect 47862 39792 51191 39794
rect 47862 39736 51130 39792
rect 51186 39736 51191 39792
rect 47862 39734 51191 39736
rect 51125 39731 51191 39734
rect 90734 39696 90794 40006
rect 92801 40003 92867 40006
rect 135213 40003 135279 40006
rect 142481 40066 142547 40069
rect 185261 40066 185327 40069
rect 187886 40066 187946 40376
rect 142481 40064 145074 40066
rect 142481 40008 142486 40064
rect 142542 40008 145074 40064
rect 142481 40006 145074 40008
rect 142481 40003 142547 40006
rect 103430 39802 104012 39862
rect 100989 39794 101055 39797
rect 103430 39794 103490 39802
rect 100989 39792 103490 39794
rect 100989 39736 100994 39792
rect 101050 39736 103490 39792
rect 100989 39734 103490 39736
rect 100989 39731 101055 39734
rect 58209 39658 58275 39661
rect 58209 39656 60956 39658
rect 58209 39600 58214 39656
rect 58270 39600 60956 39656
rect 58209 39598 60956 39600
rect 58209 39595 58275 39598
rect 47862 39386 47922 39560
rect 131766 39522 131826 39832
rect 145014 39696 145074 40006
rect 185261 40064 187946 40066
rect 185261 40008 185266 40064
rect 185322 40008 187946 40064
rect 185261 40006 187946 40008
rect 185261 40003 185327 40006
rect 177257 39658 177323 39661
rect 174852 39656 177323 39658
rect 174852 39600 177262 39656
rect 177318 39600 177323 39656
rect 174852 39598 177323 39600
rect 177257 39595 177323 39598
rect 135397 39522 135463 39525
rect 131766 39520 135463 39522
rect 131766 39464 135402 39520
rect 135458 39464 135463 39520
rect 131766 39462 135463 39464
rect 135397 39459 135463 39462
rect 51217 39386 51283 39389
rect 47862 39384 51283 39386
rect 47862 39328 51222 39384
rect 51278 39328 51283 39384
rect 47862 39326 51283 39328
rect 51217 39323 51283 39326
rect 185169 39386 185235 39389
rect 187886 39386 187946 39832
rect 185169 39384 187946 39386
rect 185169 39328 185174 39384
rect 185230 39328 187946 39384
rect 185169 39326 187946 39328
rect 185169 39323 185235 39326
rect 103430 39122 104012 39182
rect 58301 39114 58367 39117
rect 92709 39114 92775 39117
rect 58301 39112 60956 39114
rect 58301 39056 58306 39112
rect 58362 39056 60956 39112
rect 58301 39054 60956 39056
rect 90764 39112 92775 39114
rect 90764 39056 92714 39112
rect 92770 39056 92775 39112
rect 90764 39054 92775 39056
rect 58301 39051 58367 39054
rect 92709 39051 92775 39054
rect 101173 39114 101239 39117
rect 103430 39114 103490 39122
rect 101173 39112 103490 39114
rect 101173 39056 101178 39112
rect 101234 39056 103490 39112
rect 101173 39054 103490 39056
rect 101173 39051 101239 39054
rect 47862 38570 47922 38880
rect 131766 38842 131826 39152
rect 143677 39114 143743 39117
rect 177257 39114 177323 39117
rect 143677 39112 145044 39114
rect 143677 39056 143682 39112
rect 143738 39056 145044 39112
rect 143677 39054 145044 39056
rect 174852 39112 177323 39114
rect 174852 39056 177262 39112
rect 177318 39056 177323 39112
rect 174852 39054 177323 39056
rect 143677 39051 143743 39054
rect 177257 39051 177323 39054
rect 142849 38978 142915 38981
rect 142849 38976 145074 38978
rect 142849 38920 142854 38976
rect 142910 38920 145074 38976
rect 142849 38918 145074 38920
rect 142849 38915 142915 38918
rect 135213 38842 135279 38845
rect 131766 38840 135279 38842
rect 131766 38784 135218 38840
rect 135274 38784 135279 38840
rect 131766 38782 135279 38784
rect 135213 38779 135279 38782
rect 92801 38706 92867 38709
rect 90734 38704 92867 38706
rect 90734 38648 92806 38704
rect 92862 38648 92867 38704
rect 90734 38646 92867 38648
rect 51125 38570 51191 38573
rect 47862 38568 51191 38570
rect 47862 38512 51130 38568
rect 51186 38512 51191 38568
rect 47862 38510 51191 38512
rect 51125 38507 51191 38510
rect 90734 38472 90794 38646
rect 92801 38643 92867 38646
rect 103430 38578 104012 38638
rect 100989 38570 101055 38573
rect 103430 38570 103490 38578
rect 100989 38568 103490 38570
rect 100989 38512 100994 38568
rect 101050 38512 103490 38568
rect 100989 38510 103490 38512
rect 100989 38507 101055 38510
rect 58209 38434 58275 38437
rect 58209 38432 60956 38434
rect 58209 38376 58214 38432
rect 58270 38376 60956 38432
rect 58209 38374 60956 38376
rect 58209 38371 58275 38374
rect 47862 38162 47922 38336
rect 92893 38298 92959 38301
rect 90734 38296 92959 38298
rect 90734 38240 92898 38296
rect 92954 38240 92959 38296
rect 90734 38238 92959 38240
rect 131766 38298 131826 38608
rect 145014 38472 145074 38918
rect 185261 38842 185327 38845
rect 187886 38842 187946 39152
rect 185261 38840 187946 38842
rect 185261 38784 185266 38840
rect 185322 38784 187946 38840
rect 185261 38782 187946 38784
rect 185261 38779 185327 38782
rect 177349 38434 177415 38437
rect 174852 38432 177415 38434
rect 174852 38376 177354 38432
rect 177410 38376 177415 38432
rect 174852 38374 177415 38376
rect 177349 38371 177415 38374
rect 135397 38298 135463 38301
rect 131766 38296 135463 38298
rect 131766 38240 135402 38296
rect 135458 38240 135463 38296
rect 131766 38238 135463 38240
rect 51217 38162 51283 38165
rect 47862 38160 51283 38162
rect 47862 38104 51222 38160
rect 51278 38104 51283 38160
rect 47862 38102 51283 38104
rect 51217 38099 51283 38102
rect 90734 37928 90794 38238
rect 92893 38235 92959 38238
rect 135397 38235 135463 38238
rect 143401 38298 143467 38301
rect 143401 38296 145074 38298
rect 143401 38240 143406 38296
rect 143462 38240 145074 38296
rect 143401 38238 145074 38240
rect 143401 38235 143467 38238
rect 103430 37898 104012 37958
rect 145014 37928 145074 38238
rect 185169 38162 185235 38165
rect 187886 38162 187946 38608
rect 185169 38160 187946 38162
rect 185169 38104 185174 38160
rect 185230 38104 187946 38160
rect 185169 38102 187946 38104
rect 185169 38099 185235 38102
rect 58393 37890 58459 37893
rect 100529 37890 100595 37893
rect 103430 37890 103490 37898
rect 58393 37888 60956 37890
rect 58393 37832 58398 37888
rect 58454 37832 60956 37888
rect 58393 37830 60956 37832
rect 100529 37888 103490 37890
rect 100529 37832 100534 37888
rect 100590 37832 103490 37888
rect 100529 37830 103490 37832
rect 131766 37890 131826 37928
rect 135397 37890 135463 37893
rect 177717 37890 177783 37893
rect 131766 37888 135463 37890
rect 131766 37832 135402 37888
rect 135458 37832 135463 37888
rect 131766 37830 135463 37832
rect 174852 37888 177783 37890
rect 174852 37832 177722 37888
rect 177778 37832 177783 37888
rect 174852 37830 177783 37832
rect 58393 37827 58459 37830
rect 100529 37827 100595 37830
rect 135397 37827 135463 37830
rect 177717 37827 177783 37830
rect 184985 37890 185051 37893
rect 187886 37890 187946 37928
rect 184985 37888 187946 37890
rect 184985 37832 184990 37888
rect 185046 37832 187946 37888
rect 184985 37830 187946 37832
rect 184985 37827 185051 37830
rect 47862 37346 47922 37656
rect 92709 37482 92775 37485
rect 90734 37480 92775 37482
rect 90734 37424 92714 37480
rect 92770 37424 92775 37480
rect 90734 37422 92775 37424
rect 50205 37346 50271 37349
rect 47862 37344 50271 37346
rect 47862 37288 50210 37344
rect 50266 37288 50271 37344
rect 47862 37286 50271 37288
rect 50205 37283 50271 37286
rect 90734 37248 90794 37422
rect 92709 37419 92775 37422
rect 143677 37482 143743 37485
rect 143677 37480 145074 37482
rect 143677 37424 143682 37480
rect 143738 37424 145074 37480
rect 143677 37422 145074 37424
rect 143677 37419 143743 37422
rect 103430 37354 104012 37414
rect 100989 37346 101055 37349
rect 103430 37346 103490 37354
rect 100989 37344 103490 37346
rect 100989 37288 100994 37344
rect 101050 37288 103490 37344
rect 100989 37286 103490 37288
rect 100989 37283 101055 37286
rect 58209 37210 58275 37213
rect 58209 37208 60956 37210
rect 58209 37152 58214 37208
rect 58270 37152 60956 37208
rect 58209 37150 60956 37152
rect 58209 37147 58275 37150
rect 47862 36802 47922 37112
rect 92801 37074 92867 37077
rect 90734 37072 92867 37074
rect 90734 37016 92806 37072
rect 92862 37016 92867 37072
rect 90734 37014 92867 37016
rect 51217 36802 51283 36805
rect 47862 36800 51283 36802
rect 47862 36744 51222 36800
rect 51278 36744 51283 36800
rect 47862 36742 51283 36744
rect 51217 36739 51283 36742
rect 90734 36704 90794 37014
rect 92801 37011 92867 37014
rect 131766 36938 131826 37384
rect 145014 37248 145074 37422
rect 177717 37210 177783 37213
rect 174852 37208 177783 37210
rect 174852 37152 177722 37208
rect 177778 37152 177783 37208
rect 174852 37150 177783 37152
rect 177717 37147 177783 37150
rect 135397 36938 135463 36941
rect 131766 36936 135463 36938
rect 131766 36880 135402 36936
rect 135458 36880 135463 36936
rect 131766 36878 135463 36880
rect 135397 36875 135463 36878
rect 143493 36938 143559 36941
rect 185169 36938 185235 36941
rect 187886 36938 187946 37384
rect 143493 36936 145074 36938
rect 143493 36880 143498 36936
rect 143554 36880 145074 36936
rect 143493 36878 145074 36880
rect 143493 36875 143559 36878
rect 103430 36674 104012 36734
rect 145014 36704 145074 36878
rect 185169 36936 187946 36938
rect 185169 36880 185174 36936
rect 185230 36880 187946 36936
rect 185169 36878 187946 36880
rect 185169 36875 185235 36878
rect 58301 36666 58367 36669
rect 100897 36666 100963 36669
rect 103430 36666 103490 36674
rect 58301 36664 60956 36666
rect 58301 36608 58306 36664
rect 58362 36608 60956 36664
rect 58301 36606 60956 36608
rect 100897 36664 103490 36666
rect 100897 36608 100902 36664
rect 100958 36608 103490 36664
rect 100897 36606 103490 36608
rect 131766 36666 131826 36704
rect 134661 36666 134727 36669
rect 177441 36666 177507 36669
rect 131766 36664 134727 36666
rect 131766 36608 134666 36664
rect 134722 36608 134727 36664
rect 131766 36606 134727 36608
rect 174852 36664 177507 36666
rect 174852 36608 177446 36664
rect 177502 36608 177507 36664
rect 174852 36606 177507 36608
rect 58301 36603 58367 36606
rect 100897 36603 100963 36606
rect 134661 36603 134727 36606
rect 177441 36603 177507 36606
rect 51125 36530 51191 36533
rect 47862 36528 51191 36530
rect 47862 36472 51130 36528
rect 51186 36472 51191 36528
rect 47862 36470 51191 36472
rect 47862 36432 47922 36470
rect 51125 36467 51191 36470
rect 185077 36530 185143 36533
rect 187886 36530 187946 36704
rect 185077 36528 187946 36530
rect 185077 36472 185082 36528
rect 185138 36472 187946 36528
rect 185077 36470 187946 36472
rect 185077 36467 185143 36470
rect 103430 36130 104012 36190
rect 58209 36122 58275 36125
rect 92709 36122 92775 36125
rect 58209 36120 60956 36122
rect 58209 36064 58214 36120
rect 58270 36064 60956 36120
rect 58209 36062 60956 36064
rect 90764 36120 92775 36122
rect 90764 36064 92714 36120
rect 92770 36064 92775 36120
rect 90764 36062 92775 36064
rect 58209 36059 58275 36062
rect 92709 36059 92775 36062
rect 100989 36122 101055 36125
rect 103430 36122 103490 36130
rect 100989 36120 103490 36122
rect 100989 36064 100994 36120
rect 101050 36064 103490 36120
rect 100989 36062 103490 36064
rect 100989 36059 101055 36062
rect 92801 35986 92867 35989
rect 90734 35984 92867 35986
rect 90734 35928 92806 35984
rect 92862 35928 92867 35984
rect 90734 35926 92867 35928
rect 47862 35714 47922 35888
rect 51217 35714 51283 35717
rect 47862 35712 51283 35714
rect 47862 35656 51222 35712
rect 51278 35656 51283 35712
rect 47862 35654 51283 35656
rect 51217 35651 51283 35654
rect 90734 35480 90794 35926
rect 92801 35923 92867 35926
rect 131766 35714 131826 36160
rect 143677 36122 143743 36125
rect 177441 36122 177507 36125
rect 143677 36120 145044 36122
rect 143677 36064 143682 36120
rect 143738 36064 145044 36120
rect 143677 36062 145044 36064
rect 174852 36120 177507 36122
rect 174852 36064 177446 36120
rect 177502 36064 177507 36120
rect 174852 36062 177507 36064
rect 143677 36059 143743 36062
rect 177441 36059 177507 36062
rect 143033 35986 143099 35989
rect 143033 35984 145074 35986
rect 143033 35928 143038 35984
rect 143094 35928 145074 35984
rect 143033 35926 145074 35928
rect 143033 35923 143099 35926
rect 135397 35714 135463 35717
rect 131766 35712 135463 35714
rect 131766 35656 135402 35712
rect 135458 35656 135463 35712
rect 131766 35654 135463 35656
rect 135397 35651 135463 35654
rect 103430 35450 104012 35510
rect 145014 35480 145074 35926
rect 185445 35714 185511 35717
rect 187886 35714 187946 36160
rect 185445 35712 187946 35714
rect 185445 35656 185450 35712
rect 185506 35656 187946 35712
rect 185445 35654 187946 35656
rect 185445 35651 185511 35654
rect 58301 35442 58367 35445
rect 100713 35442 100779 35445
rect 103430 35442 103490 35450
rect 58301 35440 60956 35442
rect 58301 35384 58306 35440
rect 58362 35384 60956 35440
rect 58301 35382 60956 35384
rect 100713 35440 103490 35442
rect 100713 35384 100718 35440
rect 100774 35384 103490 35440
rect 100713 35382 103490 35384
rect 58301 35379 58367 35382
rect 100713 35379 100779 35382
rect 131766 35306 131826 35480
rect 177349 35442 177415 35445
rect 174852 35440 177415 35442
rect 174852 35384 177354 35440
rect 177410 35384 177415 35440
rect 174852 35382 177415 35384
rect 177349 35379 177415 35382
rect 135213 35306 135279 35309
rect 131766 35304 135279 35306
rect 131766 35248 135218 35304
rect 135274 35248 135279 35304
rect 131766 35246 135279 35248
rect 135213 35243 135279 35246
rect 184893 35306 184959 35309
rect 187886 35306 187946 35480
rect 184893 35304 187946 35306
rect 184893 35248 184898 35304
rect 184954 35248 187946 35304
rect 184893 35246 187946 35248
rect 184893 35243 184959 35246
rect 47862 35170 47922 35208
rect 51217 35170 51283 35173
rect 47862 35168 51283 35170
rect 47862 35112 51222 35168
rect 51278 35112 51283 35168
rect 47862 35110 51283 35112
rect 51217 35107 51283 35110
rect 103430 34906 104012 34966
rect 58301 34898 58367 34901
rect 92709 34898 92775 34901
rect 58301 34896 60956 34898
rect 58301 34840 58306 34896
rect 58362 34840 60956 34896
rect 58301 34838 60956 34840
rect 90764 34896 92775 34898
rect 90764 34840 92714 34896
rect 92770 34840 92775 34896
rect 90764 34838 92775 34840
rect 58301 34835 58367 34838
rect 92709 34835 92775 34838
rect 101081 34898 101147 34901
rect 103430 34898 103490 34906
rect 101081 34896 103490 34898
rect 101081 34840 101086 34896
rect 101142 34840 103490 34896
rect 101081 34838 103490 34840
rect 101081 34835 101147 34838
rect 47862 34218 47922 34664
rect 92801 34626 92867 34629
rect 90734 34624 92867 34626
rect 90734 34568 92806 34624
rect 92862 34568 92867 34624
rect 90734 34566 92867 34568
rect 90734 34256 90794 34566
rect 92801 34563 92867 34566
rect 131766 34490 131826 34936
rect 143677 34898 143743 34901
rect 177257 34898 177323 34901
rect 143677 34896 145044 34898
rect 143677 34840 143682 34896
rect 143738 34840 145044 34896
rect 143677 34838 145044 34840
rect 174852 34896 177323 34898
rect 174852 34840 177262 34896
rect 177318 34840 177323 34896
rect 174852 34838 177323 34840
rect 143677 34835 143743 34838
rect 177257 34835 177323 34838
rect 142389 34626 142455 34629
rect 142389 34624 145074 34626
rect 142389 34568 142394 34624
rect 142450 34568 145074 34624
rect 142389 34566 145074 34568
rect 142389 34563 142455 34566
rect 135213 34490 135279 34493
rect 131766 34488 135279 34490
rect 131766 34432 135218 34488
rect 135274 34432 135279 34488
rect 131766 34430 135279 34432
rect 135213 34427 135279 34430
rect 103430 34226 104012 34286
rect 145014 34256 145074 34566
rect 185261 34490 185327 34493
rect 187886 34490 187946 34936
rect 185261 34488 187946 34490
rect 185261 34432 185266 34488
rect 185322 34432 187946 34488
rect 185261 34430 187946 34432
rect 185261 34427 185327 34430
rect 51125 34218 51191 34221
rect 47862 34216 51191 34218
rect 47862 34160 51130 34216
rect 51186 34160 51191 34216
rect 47862 34158 51191 34160
rect 51125 34155 51191 34158
rect 58209 34218 58275 34221
rect 100989 34218 101055 34221
rect 103430 34218 103490 34226
rect 58209 34216 60956 34218
rect 58209 34160 58214 34216
rect 58270 34160 60956 34216
rect 58209 34158 60956 34160
rect 100989 34216 103490 34218
rect 100989 34160 100994 34216
rect 101050 34160 103490 34216
rect 100989 34158 103490 34160
rect 58209 34155 58275 34158
rect 100989 34155 101055 34158
rect 47862 33946 47922 33984
rect 51217 33946 51283 33949
rect 47862 33944 51283 33946
rect 47862 33888 51222 33944
rect 51278 33888 51283 33944
rect 47862 33886 51283 33888
rect 131766 33946 131826 34256
rect 177717 34218 177783 34221
rect 174852 34216 177783 34218
rect 174852 34160 177722 34216
rect 177778 34160 177783 34216
rect 174852 34158 177783 34160
rect 177717 34155 177783 34158
rect 135397 33946 135463 33949
rect 131766 33944 135463 33946
rect 131766 33888 135402 33944
rect 135458 33888 135463 33944
rect 131766 33886 135463 33888
rect 51217 33883 51283 33886
rect 135397 33883 135463 33886
rect 185169 33946 185235 33949
rect 187886 33946 187946 34256
rect 185169 33944 187946 33946
rect 185169 33888 185174 33944
rect 185230 33888 187946 33944
rect 185169 33886 187946 33888
rect 185169 33883 185235 33886
rect 100805 33810 100871 33813
rect 134661 33810 134727 33813
rect 100805 33808 103490 33810
rect 100805 33752 100810 33808
rect 100866 33752 103490 33808
rect 100805 33750 103490 33752
rect 100805 33747 100871 33750
rect 103430 33746 103490 33750
rect 131766 33808 134727 33810
rect 131766 33752 134666 33808
rect 134722 33752 134727 33808
rect 131766 33750 134727 33752
rect 103430 33686 104012 33746
rect 131766 33712 131826 33750
rect 134661 33747 134727 33750
rect 184985 33810 185051 33813
rect 184985 33808 187946 33810
rect 184985 33752 184990 33808
rect 185046 33752 187946 33808
rect 184985 33750 187946 33752
rect 184985 33747 185051 33750
rect 187886 33712 187946 33750
rect 59221 33674 59287 33677
rect 92709 33674 92775 33677
rect 59221 33672 60956 33674
rect 59221 33616 59226 33672
rect 59282 33616 60956 33672
rect 59221 33614 60956 33616
rect 90764 33672 92775 33674
rect 90764 33616 92714 33672
rect 92770 33616 92775 33672
rect 90764 33614 92775 33616
rect 59221 33611 59287 33614
rect 92709 33611 92775 33614
rect 143677 33674 143743 33677
rect 177625 33674 177691 33677
rect 143677 33672 145044 33674
rect 143677 33616 143682 33672
rect 143738 33616 145044 33672
rect 143677 33614 145044 33616
rect 174852 33672 177691 33674
rect 174852 33616 177630 33672
rect 177686 33616 177691 33672
rect 174852 33614 177691 33616
rect 143677 33611 143743 33614
rect 177625 33611 177691 33614
rect 47862 33130 47922 33440
rect 92801 33402 92867 33405
rect 90734 33400 92867 33402
rect 90734 33344 92806 33400
rect 92862 33344 92867 33400
rect 90734 33342 92867 33344
rect 90734 33168 90794 33342
rect 92801 33339 92867 33342
rect 143309 33402 143375 33405
rect 143309 33400 145074 33402
rect 143309 33344 143314 33400
rect 143370 33344 145074 33400
rect 143309 33342 145074 33344
rect 143309 33339 143375 33342
rect 103430 33138 104012 33198
rect 145014 33168 145074 33342
rect 50021 33130 50087 33133
rect 47862 33128 50087 33130
rect 47862 33072 50026 33128
rect 50082 33072 50087 33128
rect 47862 33070 50087 33072
rect 50021 33067 50087 33070
rect 58209 33130 58275 33133
rect 100989 33130 101055 33133
rect 103430 33130 103490 33138
rect 58209 33128 60956 33130
rect 58209 33072 58214 33128
rect 58270 33072 60956 33128
rect 58209 33070 60956 33072
rect 100989 33128 103490 33130
rect 100989 33072 100994 33128
rect 101050 33072 103490 33128
rect 100989 33070 103490 33072
rect 58209 33067 58275 33070
rect 100989 33067 101055 33070
rect 92893 32994 92959 32997
rect 90734 32992 92959 32994
rect 90734 32936 92898 32992
rect 92954 32936 92959 32992
rect 90734 32934 92959 32936
rect 47862 32586 47922 32896
rect 51217 32586 51283 32589
rect 47862 32584 51283 32586
rect 47862 32528 51222 32584
rect 51278 32528 51283 32584
rect 47862 32526 51283 32528
rect 51217 32523 51283 32526
rect 19342 32458 19924 32518
rect 90734 32488 90794 32934
rect 92893 32931 92959 32934
rect 131766 32722 131826 33168
rect 177717 33130 177783 33133
rect 174852 33128 177783 33130
rect 174852 33072 177722 33128
rect 177778 33072 177783 33128
rect 174852 33070 177783 33072
rect 177717 33067 177783 33070
rect 142757 32994 142823 32997
rect 142757 32992 145074 32994
rect 142757 32936 142762 32992
rect 142818 32936 145074 32992
rect 142757 32934 145074 32936
rect 142757 32931 142823 32934
rect 135397 32722 135463 32725
rect 131766 32720 135463 32722
rect 131766 32664 135402 32720
rect 135458 32664 135463 32720
rect 131766 32662 135463 32664
rect 135397 32659 135463 32662
rect 103430 32458 104012 32518
rect 145014 32488 145074 32934
rect 185169 32722 185235 32725
rect 187886 32722 187946 33168
rect 185169 32720 187946 32722
rect 185169 32664 185174 32720
rect 185230 32664 187946 32720
rect 185169 32662 187946 32664
rect 185169 32659 185235 32662
rect 18097 32450 18163 32453
rect 19342 32450 19402 32458
rect 18097 32448 19402 32450
rect 18097 32392 18102 32448
rect 18158 32392 19402 32448
rect 18097 32390 19402 32392
rect 58301 32450 58367 32453
rect 100897 32450 100963 32453
rect 103430 32450 103490 32458
rect 58301 32448 60956 32450
rect 58301 32392 58306 32448
rect 58362 32392 60956 32448
rect 58301 32390 60956 32392
rect 100897 32448 103490 32450
rect 100897 32392 100902 32448
rect 100958 32392 103490 32448
rect 100897 32390 103490 32392
rect 131766 32450 131826 32488
rect 135213 32450 135279 32453
rect 177809 32450 177875 32453
rect 131766 32448 135279 32450
rect 131766 32392 135218 32448
rect 135274 32392 135279 32448
rect 131766 32390 135279 32392
rect 174852 32448 177875 32450
rect 174852 32392 177814 32448
rect 177870 32392 177875 32448
rect 174852 32390 177875 32392
rect 18097 32387 18163 32390
rect 58301 32387 58367 32390
rect 100897 32387 100963 32390
rect 135213 32387 135279 32390
rect 177809 32387 177875 32390
rect 185077 32314 185143 32317
rect 187886 32314 187946 32488
rect 185077 32312 187946 32314
rect 185077 32256 185082 32312
rect 185138 32256 187946 32312
rect 185077 32254 187946 32256
rect 185077 32251 185143 32254
rect 47862 31906 47922 32216
rect 143677 32178 143743 32181
rect 143677 32176 145074 32178
rect 143677 32120 143682 32176
rect 143738 32120 145074 32176
rect 143677 32118 145074 32120
rect 143677 32115 143743 32118
rect 103430 31914 104012 31974
rect 145014 31944 145074 32118
rect 50021 31906 50087 31909
rect 47862 31904 50087 31906
rect 47862 31848 50026 31904
rect 50082 31848 50087 31904
rect 47862 31846 50087 31848
rect 50021 31843 50087 31846
rect 58209 31906 58275 31909
rect 92709 31906 92775 31909
rect 58209 31904 60956 31906
rect 58209 31848 58214 31904
rect 58270 31848 60956 31904
rect 58209 31846 60956 31848
rect 90764 31904 92775 31906
rect 90764 31848 92714 31904
rect 92770 31848 92775 31904
rect 90764 31846 92775 31848
rect 58209 31843 58275 31846
rect 92709 31843 92775 31846
rect 100989 31906 101055 31909
rect 103430 31906 103490 31914
rect 100989 31904 103490 31906
rect 100989 31848 100994 31904
rect 101050 31848 103490 31904
rect 100989 31846 103490 31848
rect 100989 31843 101055 31846
rect 92801 31770 92867 31773
rect 90734 31768 92867 31770
rect 90734 31712 92806 31768
rect 92862 31712 92867 31768
rect 90734 31710 92867 31712
rect 47862 31498 47922 31672
rect 51217 31498 51283 31501
rect 47862 31496 51283 31498
rect 47862 31440 51222 31496
rect 51278 31440 51283 31496
rect 47862 31438 51283 31440
rect 51217 31435 51283 31438
rect 90734 31264 90794 31710
rect 92801 31707 92867 31710
rect 131766 31498 131826 31944
rect 177717 31906 177783 31909
rect 174852 31904 177783 31906
rect 174852 31848 177722 31904
rect 177778 31848 177783 31904
rect 174852 31846 177783 31848
rect 177717 31843 177783 31846
rect 142573 31770 142639 31773
rect 142573 31768 145074 31770
rect 142573 31712 142578 31768
rect 142634 31712 145074 31768
rect 142573 31710 145074 31712
rect 142573 31707 142639 31710
rect 135397 31498 135463 31501
rect 131766 31496 135463 31498
rect 131766 31440 135402 31496
rect 135458 31440 135463 31496
rect 131766 31438 135463 31440
rect 135397 31435 135463 31438
rect 103430 31234 104012 31294
rect 145014 31264 145074 31710
rect 185169 31498 185235 31501
rect 187886 31498 187946 31944
rect 185169 31496 187946 31498
rect 185169 31440 185174 31496
rect 185230 31440 187946 31496
rect 185169 31438 187946 31440
rect 185169 31435 185235 31438
rect 58301 31226 58367 31229
rect 100805 31226 100871 31229
rect 103430 31226 103490 31234
rect 58301 31224 60956 31226
rect 58301 31168 58306 31224
rect 58362 31168 60956 31224
rect 58301 31166 60956 31168
rect 100805 31224 103490 31226
rect 100805 31168 100810 31224
rect 100866 31168 103490 31224
rect 100805 31166 103490 31168
rect 131766 31226 131826 31264
rect 135213 31226 135279 31229
rect 177625 31226 177691 31229
rect 131766 31224 135279 31226
rect 131766 31168 135218 31224
rect 135274 31168 135279 31224
rect 131766 31166 135279 31168
rect 174852 31224 177691 31226
rect 174852 31168 177630 31224
rect 177686 31168 177691 31224
rect 174852 31166 177691 31168
rect 58301 31163 58367 31166
rect 100805 31163 100871 31166
rect 135213 31163 135279 31166
rect 177625 31163 177691 31166
rect 47862 30954 47922 30992
rect 51217 30954 51283 30957
rect 47862 30952 51283 30954
rect 47862 30896 51222 30952
rect 51278 30896 51283 30952
rect 47862 30894 51283 30896
rect 51217 30891 51283 30894
rect 184985 30954 185051 30957
rect 187886 30954 187946 31264
rect 184985 30952 187946 30954
rect 184985 30896 184990 30952
rect 185046 30896 187946 30952
rect 184985 30894 187946 30896
rect 184985 30891 185051 30894
rect 103430 30690 104012 30750
rect 58301 30682 58367 30685
rect 92709 30682 92775 30685
rect 58301 30680 60956 30682
rect 58301 30624 58306 30680
rect 58362 30624 60956 30680
rect 58301 30622 60956 30624
rect 90764 30680 92775 30682
rect 90764 30624 92714 30680
rect 92770 30624 92775 30680
rect 90764 30622 92775 30624
rect 58301 30619 58367 30622
rect 92709 30619 92775 30622
rect 101081 30682 101147 30685
rect 103430 30682 103490 30690
rect 101081 30680 103490 30682
rect 101081 30624 101086 30680
rect 101142 30624 103490 30680
rect 101081 30622 103490 30624
rect 131766 30682 131826 30720
rect 135213 30682 135279 30685
rect 131766 30680 135279 30682
rect 131766 30624 135218 30680
rect 135274 30624 135279 30680
rect 131766 30622 135279 30624
rect 101081 30619 101147 30622
rect 135213 30619 135279 30622
rect 143677 30682 143743 30685
rect 177441 30682 177507 30685
rect 143677 30680 145044 30682
rect 143677 30624 143682 30680
rect 143738 30624 145044 30680
rect 143677 30622 145044 30624
rect 174852 30680 177507 30682
rect 174852 30624 177446 30680
rect 177502 30624 177507 30680
rect 174852 30622 177507 30624
rect 143677 30619 143743 30622
rect 177441 30619 177507 30622
rect 92801 30546 92867 30549
rect 90734 30544 92867 30546
rect 90734 30488 92806 30544
rect 92862 30488 92867 30544
rect 90734 30486 92867 30488
rect 47862 30002 47922 30448
rect 90734 30176 90794 30486
rect 92801 30483 92867 30486
rect 142757 30546 142823 30549
rect 142757 30544 145074 30546
rect 142757 30488 142762 30544
rect 142818 30488 145074 30544
rect 142757 30486 145074 30488
rect 142757 30483 142823 30486
rect 145014 30176 145074 30486
rect 185261 30274 185327 30277
rect 187886 30274 187946 30720
rect 185261 30272 187946 30274
rect 185261 30216 185266 30272
rect 185322 30216 187946 30272
rect 185261 30214 187946 30216
rect 185261 30211 185327 30214
rect 58209 30138 58275 30141
rect 177717 30138 177783 30141
rect 58209 30136 60956 30138
rect 58209 30080 58214 30136
rect 58270 30080 60956 30136
rect 58209 30078 60956 30080
rect 174852 30136 177783 30138
rect 174852 30080 177722 30136
rect 177778 30080 177783 30136
rect 174852 30078 177783 30080
rect 58209 30075 58275 30078
rect 177717 30075 177783 30078
rect 103430 30010 104012 30070
rect 51125 30002 51191 30005
rect 47862 30000 51191 30002
rect 47862 29944 51130 30000
rect 51186 29944 51191 30000
rect 47862 29942 51191 29944
rect 51125 29939 51191 29942
rect 100989 30002 101055 30005
rect 103430 30002 103490 30010
rect 100989 30000 103490 30002
rect 100989 29944 100994 30000
rect 101050 29944 103490 30000
rect 100989 29942 103490 29944
rect 100989 29939 101055 29942
rect 131766 29866 131826 30040
rect 135397 29866 135463 29869
rect 131766 29864 135463 29866
rect 131766 29808 135402 29864
rect 135458 29808 135463 29864
rect 131766 29806 135463 29808
rect 135397 29803 135463 29806
rect 47862 29730 47922 29768
rect 51217 29730 51283 29733
rect 47862 29728 51283 29730
rect 47862 29672 51222 29728
rect 51278 29672 51283 29728
rect 47862 29670 51283 29672
rect 51217 29667 51283 29670
rect 185169 29730 185235 29733
rect 187886 29730 187946 30040
rect 185169 29728 187946 29730
rect 185169 29672 185174 29728
rect 185230 29672 187946 29728
rect 185169 29670 187946 29672
rect 185169 29667 185235 29670
rect 103430 29466 104012 29526
rect 58393 29458 58459 29461
rect 92709 29458 92775 29461
rect 58393 29456 60956 29458
rect 58393 29400 58398 29456
rect 58454 29400 60956 29456
rect 58393 29398 60956 29400
rect 90764 29456 92775 29458
rect 90764 29400 92714 29456
rect 92770 29400 92775 29456
rect 90764 29398 92775 29400
rect 58393 29395 58459 29398
rect 92709 29395 92775 29398
rect 101725 29458 101791 29461
rect 103430 29458 103490 29466
rect 101725 29456 103490 29458
rect 101725 29400 101730 29456
rect 101786 29400 103490 29456
rect 101725 29398 103490 29400
rect 101725 29395 101791 29398
rect 131766 29322 131826 29496
rect 143677 29458 143743 29461
rect 177257 29458 177323 29461
rect 143677 29456 145044 29458
rect 143677 29400 143682 29456
rect 143738 29400 145044 29456
rect 143677 29398 145044 29400
rect 174852 29456 177323 29458
rect 174852 29400 177262 29456
rect 177318 29400 177323 29456
rect 174852 29398 177323 29400
rect 143677 29395 143743 29398
rect 177257 29395 177323 29398
rect 135213 29322 135279 29325
rect 131766 29320 135279 29322
rect 131766 29264 135218 29320
rect 135274 29264 135279 29320
rect 131766 29262 135279 29264
rect 135213 29259 135279 29262
rect 47862 28778 47922 29224
rect 92893 29186 92959 29189
rect 90734 29184 92959 29186
rect 90734 29128 92898 29184
rect 92954 29128 92959 29184
rect 90734 29126 92959 29128
rect 90734 28952 90794 29126
rect 92893 29123 92959 29126
rect 143585 29186 143651 29189
rect 143585 29184 145074 29186
rect 143585 29128 143590 29184
rect 143646 29128 145074 29184
rect 143585 29126 145074 29128
rect 143585 29123 143651 29126
rect 145014 28952 145074 29126
rect 185353 29050 185419 29053
rect 187886 29050 187946 29496
rect 185353 29048 187946 29050
rect 185353 28992 185358 29048
rect 185414 28992 187946 29048
rect 185353 28990 187946 28992
rect 185353 28987 185419 28990
rect 58209 28914 58275 28917
rect 177717 28914 177783 28917
rect 58209 28912 60956 28914
rect 58209 28856 58214 28912
rect 58270 28856 60956 28912
rect 58209 28854 60956 28856
rect 174852 28912 177783 28914
rect 174852 28856 177722 28912
rect 177778 28856 177783 28912
rect 174852 28854 177783 28856
rect 58209 28851 58275 28854
rect 177717 28851 177783 28854
rect 103430 28786 104012 28846
rect 51125 28778 51191 28781
rect 92801 28778 92867 28781
rect 47862 28776 51191 28778
rect 47862 28720 51130 28776
rect 51186 28720 51191 28776
rect 47862 28718 51191 28720
rect 51125 28715 51191 28718
rect 90734 28776 92867 28778
rect 90734 28720 92806 28776
rect 92862 28720 92867 28776
rect 90734 28718 92867 28720
rect 47862 28370 47922 28544
rect 51217 28370 51283 28373
rect 47862 28368 51283 28370
rect 47862 28312 51222 28368
rect 51278 28312 51283 28368
rect 47862 28310 51283 28312
rect 51217 28307 51283 28310
rect 90734 28272 90794 28718
rect 92801 28715 92867 28718
rect 101909 28778 101975 28781
rect 103430 28778 103490 28786
rect 101909 28776 103490 28778
rect 101909 28720 101914 28776
rect 101970 28720 103490 28776
rect 101909 28718 103490 28720
rect 101909 28715 101975 28718
rect 131766 28506 131826 28816
rect 142757 28778 142823 28781
rect 142757 28776 145074 28778
rect 142757 28720 142762 28776
rect 142818 28720 145074 28776
rect 142757 28718 145074 28720
rect 142757 28715 142823 28718
rect 135397 28506 135463 28509
rect 131766 28504 135463 28506
rect 131766 28448 135402 28504
rect 135458 28448 135463 28504
rect 131766 28446 135463 28448
rect 135397 28443 135463 28446
rect 135397 28370 135463 28373
rect 131766 28368 135463 28370
rect 131766 28312 135402 28368
rect 135458 28312 135463 28368
rect 131766 28310 135463 28312
rect 103430 28242 104012 28302
rect 131766 28272 131826 28310
rect 135397 28307 135463 28310
rect 145014 28272 145074 28718
rect 185261 28506 185327 28509
rect 187886 28506 187946 28816
rect 185261 28504 187946 28506
rect 185261 28448 185266 28504
rect 185322 28448 187946 28504
rect 185261 28446 187946 28448
rect 185261 28443 185327 28446
rect 58301 28234 58367 28237
rect 100989 28234 101055 28237
rect 103430 28234 103490 28242
rect 177441 28234 177507 28237
rect 58301 28232 60956 28234
rect 58301 28176 58306 28232
rect 58362 28176 60956 28232
rect 58301 28174 60956 28176
rect 100989 28232 103490 28234
rect 100989 28176 100994 28232
rect 101050 28176 103490 28232
rect 100989 28174 103490 28176
rect 174852 28232 177507 28234
rect 174852 28176 177446 28232
rect 177502 28176 177507 28232
rect 174852 28174 177507 28176
rect 58301 28171 58367 28174
rect 100989 28171 101055 28174
rect 177441 28171 177507 28174
rect 185169 28234 185235 28237
rect 187886 28234 187946 28272
rect 185169 28232 187946 28234
rect 185169 28176 185174 28232
rect 185230 28176 187946 28232
rect 185169 28174 187946 28176
rect 185169 28171 185235 28174
rect 47862 27554 47922 28000
rect 143677 27962 143743 27965
rect 143677 27960 145074 27962
rect 143677 27904 143682 27960
rect 143738 27904 145074 27960
rect 143677 27902 145074 27904
rect 143677 27899 143743 27902
rect 145014 27728 145074 27902
rect 58301 27690 58367 27693
rect 92709 27690 92775 27693
rect 177717 27690 177783 27693
rect 58301 27688 60956 27690
rect 58301 27632 58306 27688
rect 58362 27632 60956 27688
rect 58301 27630 60956 27632
rect 90764 27688 92775 27690
rect 90764 27632 92714 27688
rect 92770 27632 92775 27688
rect 90764 27630 92775 27632
rect 174852 27688 177783 27690
rect 174852 27632 177722 27688
rect 177778 27632 177783 27688
rect 174852 27630 177783 27632
rect 58301 27627 58367 27630
rect 92709 27627 92775 27630
rect 177717 27627 177783 27630
rect 103430 27562 104012 27622
rect 50021 27554 50087 27557
rect 47862 27552 50087 27554
rect 47862 27496 50026 27552
rect 50082 27496 50087 27552
rect 47862 27494 50087 27496
rect 50021 27491 50087 27494
rect 100989 27554 101055 27557
rect 103430 27554 103490 27562
rect 100989 27552 103490 27554
rect 100989 27496 100994 27552
rect 101050 27496 103490 27552
rect 100989 27494 103490 27496
rect 100989 27491 101055 27494
rect 92801 27418 92867 27421
rect 90734 27416 92867 27418
rect 90734 27360 92806 27416
rect 92862 27360 92867 27416
rect 90734 27358 92867 27360
rect 47862 27146 47922 27320
rect 90734 27184 90794 27358
rect 92801 27355 92867 27358
rect 131766 27282 131826 27592
rect 143401 27554 143467 27557
rect 143401 27552 145074 27554
rect 143401 27496 143406 27552
rect 143462 27496 145074 27552
rect 143401 27494 145074 27496
rect 143401 27491 143467 27494
rect 135397 27282 135463 27285
rect 131766 27280 135463 27282
rect 131766 27224 135402 27280
rect 135458 27224 135463 27280
rect 131766 27222 135463 27224
rect 135397 27219 135463 27222
rect 145014 27184 145074 27494
rect 185169 27282 185235 27285
rect 187886 27282 187946 27592
rect 185169 27280 187946 27282
rect 185169 27224 185174 27280
rect 185230 27224 187946 27280
rect 185169 27222 187946 27224
rect 185169 27219 185235 27222
rect 51217 27146 51283 27149
rect 47862 27144 51283 27146
rect 47862 27088 51222 27144
rect 51278 27088 51283 27144
rect 47862 27086 51283 27088
rect 51217 27083 51283 27086
rect 58209 27146 58275 27149
rect 177349 27146 177415 27149
rect 58209 27144 60956 27146
rect 58209 27088 58214 27144
rect 58270 27088 60956 27144
rect 58209 27086 60956 27088
rect 174852 27144 177415 27146
rect 174852 27088 177354 27144
rect 177410 27088 177415 27144
rect 174852 27086 177415 27088
rect 58209 27083 58275 27086
rect 177349 27083 177415 27086
rect 103430 27018 104012 27078
rect 101173 27010 101239 27013
rect 103430 27010 103490 27018
rect 101173 27008 103490 27010
rect 101173 26952 101178 27008
rect 101234 26952 103490 27008
rect 101173 26950 103490 26952
rect 131766 27010 131826 27048
rect 135213 27010 135279 27013
rect 131766 27008 135279 27010
rect 131766 26952 135218 27008
rect 135274 26952 135279 27008
rect 131766 26950 135279 26952
rect 101173 26947 101239 26950
rect 135213 26947 135279 26950
rect 51125 26874 51191 26877
rect 47862 26872 51191 26874
rect 47862 26816 51130 26872
rect 51186 26816 51191 26872
rect 47862 26814 51191 26816
rect 47862 26776 47922 26814
rect 51125 26811 51191 26814
rect 185813 26874 185879 26877
rect 187886 26874 187946 27048
rect 185813 26872 187946 26874
rect 185813 26816 185818 26872
rect 185874 26816 187946 26872
rect 185813 26814 187946 26816
rect 185813 26811 185879 26814
rect 92893 26738 92959 26741
rect 90734 26736 92959 26738
rect 90734 26680 92898 26736
rect 92954 26680 92959 26736
rect 90734 26678 92959 26680
rect 90734 26504 90794 26678
rect 92893 26675 92959 26678
rect 58209 26466 58275 26469
rect 143677 26466 143743 26469
rect 177625 26466 177691 26469
rect 58209 26464 60956 26466
rect 58209 26408 58214 26464
rect 58270 26408 60956 26464
rect 58209 26406 60956 26408
rect 143677 26464 145044 26466
rect 143677 26408 143682 26464
rect 143738 26408 145044 26464
rect 143677 26406 145044 26408
rect 174852 26464 177691 26466
rect 174852 26408 177630 26464
rect 177686 26408 177691 26464
rect 174852 26406 177691 26408
rect 58209 26403 58275 26406
rect 143677 26403 143743 26406
rect 177625 26403 177691 26406
rect 103430 26338 104012 26398
rect 92709 26330 92775 26333
rect 90734 26328 92775 26330
rect 90734 26272 92714 26328
rect 92770 26272 92775 26328
rect 90734 26270 92775 26272
rect 47862 25786 47922 26096
rect 90734 25960 90794 26270
rect 92709 26267 92775 26270
rect 101081 26330 101147 26333
rect 103430 26330 103490 26338
rect 101081 26328 103490 26330
rect 101081 26272 101086 26328
rect 101142 26272 103490 26328
rect 101081 26270 103490 26272
rect 101081 26267 101147 26270
rect 131766 26058 131826 26368
rect 143585 26330 143651 26333
rect 143585 26328 145074 26330
rect 143585 26272 143590 26328
rect 143646 26272 145074 26328
rect 143585 26270 145074 26272
rect 143585 26267 143651 26270
rect 135213 26058 135279 26061
rect 131766 26056 135279 26058
rect 131766 26000 135218 26056
rect 135274 26000 135279 26056
rect 131766 25998 135279 26000
rect 135213 25995 135279 25998
rect 145014 25960 145074 26270
rect 185261 26058 185327 26061
rect 187886 26058 187946 26368
rect 185261 26056 187946 26058
rect 185261 26000 185266 26056
rect 185322 26000 187946 26056
rect 185261 25998 187946 26000
rect 185261 25995 185327 25998
rect 58301 25922 58367 25925
rect 177717 25922 177783 25925
rect 58301 25920 60956 25922
rect 58301 25864 58306 25920
rect 58362 25864 60956 25920
rect 58301 25862 60956 25864
rect 174852 25920 177783 25922
rect 174852 25864 177722 25920
rect 177778 25864 177783 25920
rect 174852 25862 177783 25864
rect 58301 25859 58367 25862
rect 177717 25859 177783 25862
rect 103430 25794 104012 25854
rect 51125 25786 51191 25789
rect 47862 25784 51191 25786
rect 47862 25728 51130 25784
rect 51186 25728 51191 25784
rect 47862 25726 51191 25728
rect 51125 25723 51191 25726
rect 100989 25786 101055 25789
rect 103430 25786 103490 25794
rect 100989 25784 103490 25786
rect 100989 25728 100994 25784
rect 101050 25728 103490 25784
rect 100989 25726 103490 25728
rect 100989 25723 101055 25726
rect 131766 25650 131826 25824
rect 135397 25650 135463 25653
rect 131766 25648 135463 25650
rect 131766 25592 135402 25648
rect 135458 25592 135463 25648
rect 131766 25590 135463 25592
rect 135397 25587 135463 25590
rect 185721 25650 185787 25653
rect 187886 25650 187946 25824
rect 185721 25648 187946 25650
rect 185721 25592 185726 25648
rect 185782 25592 187946 25648
rect 185721 25590 187946 25592
rect 185721 25587 185787 25590
rect 47862 25514 47922 25552
rect 51217 25514 51283 25517
rect 47862 25512 51283 25514
rect 47862 25456 51222 25512
rect 51278 25456 51283 25512
rect 47862 25454 51283 25456
rect 51217 25451 51283 25454
rect 59037 25242 59103 25245
rect 92893 25242 92959 25245
rect 59037 25240 60956 25242
rect 59037 25184 59042 25240
rect 59098 25184 60956 25240
rect 59037 25182 60956 25184
rect 90764 25240 92959 25242
rect 90764 25184 92898 25240
rect 92954 25184 92959 25240
rect 90764 25182 92959 25184
rect 59037 25179 59103 25182
rect 92893 25179 92959 25182
rect 143125 25242 143191 25245
rect 177717 25242 177783 25245
rect 143125 25240 145044 25242
rect 143125 25184 143130 25240
rect 143186 25184 145044 25240
rect 143125 25182 145044 25184
rect 174852 25240 177783 25242
rect 174852 25184 177722 25240
rect 177778 25184 177783 25240
rect 174852 25182 177783 25184
rect 143125 25179 143191 25182
rect 177717 25179 177783 25182
rect 103430 25114 104012 25174
rect 101081 25106 101147 25109
rect 103430 25106 103490 25114
rect 101081 25104 103490 25106
rect 101081 25048 101086 25104
rect 101142 25048 103490 25104
rect 101081 25046 103490 25048
rect 101081 25043 101147 25046
rect 92801 24970 92867 24973
rect 90734 24968 92867 24970
rect 90734 24912 92806 24968
rect 92862 24912 92867 24968
rect 90734 24910 92867 24912
rect 47862 24562 47922 24872
rect 90734 24736 90794 24910
rect 92801 24907 92867 24910
rect 131766 24834 131826 25144
rect 143677 25106 143743 25109
rect 143677 25104 145074 25106
rect 143677 25048 143682 25104
rect 143738 25048 145074 25104
rect 143677 25046 145074 25048
rect 143677 25043 143743 25046
rect 135029 24834 135095 24837
rect 131766 24832 135095 24834
rect 131766 24776 135034 24832
rect 135090 24776 135095 24832
rect 131766 24774 135095 24776
rect 135029 24771 135095 24774
rect 145014 24736 145074 25046
rect 185169 24834 185235 24837
rect 187886 24834 187946 25144
rect 185169 24832 187946 24834
rect 185169 24776 185174 24832
rect 185230 24776 187946 24832
rect 185169 24774 187946 24776
rect 185169 24771 185235 24774
rect 59497 24698 59563 24701
rect 177809 24698 177875 24701
rect 59497 24696 60956 24698
rect 59497 24640 59502 24696
rect 59558 24640 60956 24696
rect 59497 24638 60956 24640
rect 174852 24696 177875 24698
rect 174852 24640 177814 24696
rect 177870 24640 177875 24696
rect 174852 24638 177875 24640
rect 59497 24635 59563 24638
rect 177809 24635 177875 24638
rect 103430 24570 104012 24630
rect 51125 24562 51191 24565
rect 92709 24562 92775 24565
rect 47862 24560 51191 24562
rect 47862 24504 51130 24560
rect 51186 24504 51191 24560
rect 47862 24502 51191 24504
rect 51125 24499 51191 24502
rect 90734 24560 92775 24562
rect 90734 24504 92714 24560
rect 92770 24504 92775 24560
rect 90734 24502 92775 24504
rect 47862 24290 47922 24328
rect 51217 24290 51283 24293
rect 47862 24288 51283 24290
rect 47862 24232 51222 24288
rect 51278 24232 51283 24288
rect 47862 24230 51283 24232
rect 51217 24227 51283 24230
rect 90734 24192 90794 24502
rect 92709 24499 92775 24502
rect 100989 24562 101055 24565
rect 103430 24562 103490 24570
rect 100989 24560 103490 24562
rect 100989 24504 100994 24560
rect 101050 24504 103490 24560
rect 100989 24502 103490 24504
rect 100989 24499 101055 24502
rect 131766 24426 131826 24600
rect 143493 24562 143559 24565
rect 143493 24560 145074 24562
rect 143493 24504 143498 24560
rect 143554 24504 145074 24560
rect 143493 24502 145074 24504
rect 143493 24499 143559 24502
rect 135397 24426 135463 24429
rect 131766 24424 135463 24426
rect 131766 24368 135402 24424
rect 135458 24368 135463 24424
rect 131766 24366 135463 24368
rect 135397 24363 135463 24366
rect 145014 24192 145074 24502
rect 59405 24154 59471 24157
rect 177349 24154 177415 24157
rect 59405 24152 60956 24154
rect 59405 24096 59410 24152
rect 59466 24096 60956 24152
rect 59405 24094 60956 24096
rect 174852 24152 177415 24154
rect 174852 24096 177354 24152
rect 177410 24096 177415 24152
rect 174852 24094 177415 24096
rect 59405 24091 59471 24094
rect 177349 24091 177415 24094
rect 185261 24154 185327 24157
rect 187886 24154 187946 24600
rect 185261 24152 187946 24154
rect 185261 24096 185266 24152
rect 185322 24096 187946 24152
rect 185261 24094 187946 24096
rect 185261 24091 185327 24094
rect 143677 24018 143743 24021
rect 143677 24016 145074 24018
rect 143677 23960 143682 24016
rect 143738 23960 145074 24016
rect 143677 23958 145074 23960
rect 143677 23955 143743 23958
rect 103430 23890 104012 23950
rect 100989 23882 101055 23885
rect 103430 23882 103490 23890
rect 100989 23880 103490 23882
rect 100989 23824 100994 23880
rect 101050 23824 103490 23880
rect 100989 23822 103490 23824
rect 100989 23819 101055 23822
rect 92709 23746 92775 23749
rect 90734 23744 92775 23746
rect 90734 23688 92714 23744
rect 92770 23688 92775 23744
rect 90734 23686 92775 23688
rect 131766 23746 131826 23920
rect 134477 23746 134543 23749
rect 131766 23744 134543 23746
rect 131766 23688 134482 23744
rect 134538 23688 134543 23744
rect 131766 23686 134543 23688
rect 47862 23338 47922 23648
rect 90734 23512 90794 23686
rect 92709 23683 92775 23686
rect 134477 23683 134543 23686
rect 145014 23512 145074 23958
rect 185261 23610 185327 23613
rect 187886 23610 187946 23920
rect 185261 23608 187946 23610
rect 185261 23552 185266 23608
rect 185322 23552 187946 23608
rect 185261 23550 187946 23552
rect 185261 23547 185327 23550
rect 58209 23474 58275 23477
rect 177625 23474 177691 23477
rect 58209 23472 60956 23474
rect 58209 23416 58214 23472
rect 58270 23416 60956 23472
rect 58209 23414 60956 23416
rect 174852 23472 177691 23474
rect 174852 23416 177630 23472
rect 177686 23416 177691 23472
rect 174852 23414 177691 23416
rect 58209 23411 58275 23414
rect 177625 23411 177691 23414
rect 103430 23346 104012 23406
rect 50389 23338 50455 23341
rect 92801 23338 92867 23341
rect 47862 23336 50455 23338
rect 47862 23280 50394 23336
rect 50450 23280 50455 23336
rect 47862 23278 50455 23280
rect 50389 23275 50455 23278
rect 90734 23336 92867 23338
rect 90734 23280 92806 23336
rect 92862 23280 92867 23336
rect 90734 23278 92867 23280
rect 19702 23208 19708 23272
rect 19772 23270 19778 23272
rect 19772 23210 19924 23270
rect 19772 23208 19778 23210
rect 47862 22930 47922 23104
rect 90734 22968 90794 23278
rect 92801 23275 92867 23278
rect 101081 23338 101147 23341
rect 103430 23338 103490 23346
rect 101081 23336 103490 23338
rect 101081 23280 101086 23336
rect 101142 23280 103490 23336
rect 101081 23278 103490 23280
rect 101081 23275 101147 23278
rect 131766 23066 131826 23376
rect 143585 23338 143651 23341
rect 143585 23336 145074 23338
rect 143585 23280 143590 23336
rect 143646 23280 145074 23336
rect 143585 23278 145074 23280
rect 143585 23275 143651 23278
rect 135397 23066 135463 23069
rect 131766 23064 135463 23066
rect 131766 23008 135402 23064
rect 135458 23008 135463 23064
rect 131766 23006 135463 23008
rect 135397 23003 135463 23006
rect 145014 22968 145074 23278
rect 51217 22930 51283 22933
rect 47862 22928 51283 22930
rect 47862 22872 51222 22928
rect 51278 22872 51283 22928
rect 47862 22870 51283 22872
rect 51217 22867 51283 22870
rect 58301 22930 58367 22933
rect 177349 22930 177415 22933
rect 58301 22928 60956 22930
rect 58301 22872 58306 22928
rect 58362 22872 60956 22928
rect 58301 22870 60956 22872
rect 174852 22928 177415 22930
rect 174852 22872 177354 22928
rect 177410 22872 177415 22928
rect 174852 22870 177415 22872
rect 58301 22867 58367 22870
rect 177349 22867 177415 22870
rect 185169 22930 185235 22933
rect 187886 22930 187946 23376
rect 185169 22928 187946 22930
rect 185169 22872 185174 22928
rect 185230 22872 187946 22928
rect 185169 22870 187946 22872
rect 185169 22867 185235 22870
rect 53977 22796 54043 22797
rect 53926 22732 53932 22796
rect 53996 22794 54043 22796
rect 53996 22792 54088 22794
rect 54038 22736 54088 22792
rect 53996 22734 54088 22736
rect 53996 22732 54043 22734
rect 53977 22731 54043 22732
rect 103430 22666 104012 22726
rect 101173 22658 101239 22661
rect 103430 22658 103490 22666
rect 101173 22656 103490 22658
rect 101173 22600 101178 22656
rect 101234 22600 103490 22656
rect 101173 22598 103490 22600
rect 131766 22658 131826 22696
rect 135305 22658 135371 22661
rect 131766 22656 135371 22658
rect 131766 22600 135310 22656
rect 135366 22600 135371 22656
rect 131766 22598 135371 22600
rect 101173 22595 101239 22598
rect 135305 22595 135371 22598
rect 185261 22658 185327 22661
rect 187886 22658 187946 22696
rect 185261 22656 187946 22658
rect 185261 22600 185266 22656
rect 185322 22600 187946 22656
rect 185261 22598 187946 22600
rect 185261 22595 185327 22598
rect 135029 22522 135095 22525
rect 131766 22520 135095 22522
rect 131766 22464 135034 22520
rect 135090 22464 135095 22520
rect 131766 22462 135095 22464
rect 47862 22114 47922 22424
rect 58209 22250 58275 22253
rect 92709 22250 92775 22253
rect 58209 22248 60956 22250
rect 58209 22192 58214 22248
rect 58270 22192 60956 22248
rect 58209 22190 60956 22192
rect 90764 22248 92775 22250
rect 90764 22192 92714 22248
rect 92770 22192 92775 22248
rect 90764 22190 92775 22192
rect 58209 22187 58275 22190
rect 92709 22187 92775 22190
rect 100989 22250 101055 22253
rect 100989 22248 103490 22250
rect 100989 22192 100994 22248
rect 101050 22192 103490 22248
rect 100989 22190 103490 22192
rect 100989 22187 101055 22190
rect 103430 22186 103490 22190
rect 103430 22126 104012 22186
rect 131766 22152 131826 22462
rect 135029 22459 135095 22462
rect 142757 22522 142823 22525
rect 142757 22520 145074 22522
rect 142757 22464 142762 22520
rect 142818 22464 145074 22520
rect 142757 22462 145074 22464
rect 142757 22459 142823 22462
rect 145014 22288 145074 22462
rect 185169 22386 185235 22389
rect 185169 22384 187946 22386
rect 185169 22328 185174 22384
rect 185230 22328 187946 22384
rect 185169 22326 187946 22328
rect 185169 22323 185235 22326
rect 177625 22250 177691 22253
rect 174852 22248 177691 22250
rect 174852 22192 177630 22248
rect 177686 22192 177691 22248
rect 174852 22190 177691 22192
rect 177625 22187 177691 22190
rect 187886 22152 187946 22326
rect 50573 22114 50639 22117
rect 92801 22114 92867 22117
rect 47862 22112 50639 22114
rect 47862 22056 50578 22112
rect 50634 22056 50639 22112
rect 47862 22054 50639 22056
rect 50573 22051 50639 22054
rect 90734 22112 92867 22114
rect 90734 22056 92806 22112
rect 92862 22056 92867 22112
rect 90734 22054 92867 22056
rect 50941 21978 51007 21981
rect 47862 21976 51007 21978
rect 47862 21920 50946 21976
rect 51002 21920 51007 21976
rect 47862 21918 51007 21920
rect 47862 21880 47922 21918
rect 50941 21915 51007 21918
rect 90734 21744 90794 22054
rect 92801 22051 92867 22054
rect 143309 22114 143375 22117
rect 143309 22112 145074 22114
rect 143309 22056 143314 22112
rect 143370 22056 145074 22112
rect 143309 22054 145074 22056
rect 143309 22051 143375 22054
rect 135121 21978 135187 21981
rect 131766 21976 135187 21978
rect 131766 21920 135126 21976
rect 135182 21920 135187 21976
rect 131766 21918 135187 21920
rect 58301 21706 58367 21709
rect 58301 21704 60956 21706
rect 58301 21648 58306 21704
rect 58362 21648 60956 21704
rect 58301 21646 60956 21648
rect 58301 21643 58367 21646
rect 101081 21570 101147 21573
rect 101081 21568 103490 21570
rect 101081 21512 101086 21568
rect 101142 21512 103490 21568
rect 101081 21510 103490 21512
rect 101081 21507 101147 21510
rect 103430 21506 103490 21510
rect 103430 21446 104012 21506
rect 131766 21472 131826 21918
rect 135121 21915 135187 21918
rect 145014 21744 145074 22054
rect 185118 21916 185124 21980
rect 185188 21978 185194 21980
rect 220313 21978 220379 21981
rect 225416 21978 225896 22008
rect 185188 21918 187946 21978
rect 185188 21916 185194 21918
rect 177717 21706 177783 21709
rect 174852 21704 177783 21706
rect 174852 21648 177722 21704
rect 177778 21648 177783 21704
rect 174852 21646 177783 21648
rect 177717 21643 177783 21646
rect 187886 21472 187946 21918
rect 220313 21976 225896 21978
rect 220313 21920 220318 21976
rect 220374 21920 225896 21976
rect 220313 21918 225896 21920
rect 220313 21915 220379 21918
rect 225416 21888 225896 21918
rect 47862 21162 47922 21200
rect 50297 21162 50363 21165
rect 47862 21160 50363 21162
rect 47862 21104 50302 21160
rect 50358 21104 50363 21160
rect 47862 21102 50363 21104
rect 50297 21099 50363 21102
rect 58209 21162 58275 21165
rect 92709 21162 92775 21165
rect 134937 21162 135003 21165
rect 58209 21160 60956 21162
rect 58209 21104 58214 21160
rect 58270 21104 60956 21160
rect 58209 21102 60956 21104
rect 90764 21160 92775 21162
rect 90764 21104 92714 21160
rect 92770 21104 92775 21160
rect 90764 21102 92775 21104
rect 58209 21099 58275 21102
rect 92709 21099 92775 21102
rect 131766 21160 135003 21162
rect 131766 21104 134942 21160
rect 134998 21104 135003 21160
rect 131766 21102 135003 21104
rect 50849 21026 50915 21029
rect 47862 21024 50915 21026
rect 47862 20968 50854 21024
rect 50910 20968 50915 21024
rect 47862 20966 50915 20968
rect 47862 20656 47922 20966
rect 50849 20963 50915 20966
rect 61705 21026 61771 21029
rect 63269 21028 63335 21029
rect 62206 21026 62212 21028
rect 61705 21024 62212 21026
rect 61705 20968 61710 21024
rect 61766 20968 62212 21024
rect 61705 20966 62212 20968
rect 61705 20963 61771 20966
rect 62206 20964 62212 20966
rect 62276 20964 62282 21028
rect 63269 21026 63316 21028
rect 63224 21024 63316 21026
rect 63224 20968 63274 21024
rect 63224 20966 63316 20968
rect 63269 20964 63316 20966
rect 63380 20964 63386 21028
rect 64741 21026 64807 21029
rect 64966 21026 64972 21028
rect 64741 21024 64972 21026
rect 64741 20968 64746 21024
rect 64802 20968 64972 21024
rect 64741 20966 64972 20968
rect 63269 20963 63335 20964
rect 64741 20963 64807 20966
rect 64966 20964 64972 20966
rect 65036 20964 65042 21028
rect 65753 21026 65819 21029
rect 68462 21026 68468 21028
rect 65753 21024 68468 21026
rect 65753 20968 65758 21024
rect 65814 20968 68468 21024
rect 65753 20966 68468 20968
rect 65753 20963 65819 20966
rect 68462 20964 68468 20966
rect 68532 20964 68538 21028
rect 103430 20898 104012 20958
rect 131766 20928 131826 21102
rect 134937 21099 135003 21102
rect 143677 21162 143743 21165
rect 177717 21162 177783 21165
rect 143677 21160 145044 21162
rect 143677 21104 143682 21160
rect 143738 21104 145044 21160
rect 143677 21102 145044 21104
rect 174852 21160 177783 21162
rect 174852 21104 177722 21160
rect 177778 21104 177783 21160
rect 174852 21102 177783 21104
rect 143677 21099 143743 21102
rect 177717 21099 177783 21102
rect 146253 21028 146319 21029
rect 147725 21028 147791 21029
rect 146253 21026 146300 21028
rect 146208 21024 146300 21026
rect 146208 20968 146258 21024
rect 146208 20966 146300 20968
rect 146253 20964 146300 20966
rect 146364 20964 146370 21028
rect 147725 21026 147772 21028
rect 147680 21024 147772 21026
rect 147680 20968 147730 21024
rect 147680 20966 147772 20968
rect 147725 20964 147772 20966
rect 147836 20964 147842 21028
rect 148737 21026 148803 21029
rect 149054 21026 149060 21028
rect 148737 21024 149060 21026
rect 148737 20968 148742 21024
rect 148798 20968 149060 21024
rect 148737 20966 149060 20968
rect 146253 20963 146319 20964
rect 147725 20963 147791 20964
rect 148737 20963 148803 20966
rect 149054 20964 149060 20966
rect 149124 20964 149130 21028
rect 62717 20890 62783 20893
rect 63494 20890 63500 20892
rect 62717 20888 63500 20890
rect 62717 20832 62722 20888
rect 62778 20832 63500 20888
rect 62717 20830 63500 20832
rect 62717 20827 62783 20830
rect 63494 20828 63500 20830
rect 63564 20828 63570 20892
rect 66857 20890 66923 20893
rect 68830 20890 68836 20892
rect 66857 20888 68836 20890
rect 66857 20832 66862 20888
rect 66918 20832 68836 20888
rect 66857 20830 68836 20832
rect 66857 20827 66923 20830
rect 68830 20828 68836 20830
rect 68900 20828 68906 20892
rect 101030 20828 101036 20892
rect 101100 20890 101106 20892
rect 103430 20890 103490 20898
rect 101100 20830 103490 20890
rect 145701 20890 145767 20893
rect 146110 20890 146116 20892
rect 145701 20888 146116 20890
rect 145701 20832 145706 20888
rect 145762 20832 146116 20888
rect 145701 20830 146116 20832
rect 101100 20828 101106 20830
rect 145701 20827 145767 20830
rect 146110 20828 146116 20830
rect 146180 20828 146186 20892
rect 185486 20828 185492 20892
rect 185556 20890 185562 20892
rect 187886 20890 187946 20928
rect 185556 20830 187946 20890
rect 185556 20828 185562 20830
rect 134845 20754 134911 20757
rect 131766 20752 134911 20754
rect 131766 20696 134850 20752
rect 134906 20696 134911 20752
rect 131766 20694 134911 20696
rect 9896 20618 10376 20648
rect 13313 20618 13379 20621
rect 9896 20616 13379 20618
rect 9896 20560 13318 20616
rect 13374 20560 13379 20616
rect 9896 20558 13379 20560
rect 9896 20528 10376 20558
rect 13313 20555 13379 20558
rect 51033 20482 51099 20485
rect 47862 20480 51099 20482
rect 47862 20424 51038 20480
rect 51094 20424 51099 20480
rect 47862 20422 51099 20424
rect 47862 19976 47922 20422
rect 51033 20419 51099 20422
rect 103430 20218 104012 20278
rect 131766 20248 131826 20694
rect 134845 20691 134911 20694
rect 150531 20754 150597 20757
rect 152734 20754 152740 20756
rect 150531 20752 152740 20754
rect 150531 20696 150536 20752
rect 150592 20696 152740 20752
rect 150531 20694 152740 20696
rect 150531 20691 150597 20694
rect 152734 20692 152740 20694
rect 152804 20692 152810 20756
rect 185118 20692 185124 20756
rect 185188 20754 185194 20756
rect 185188 20694 187946 20754
rect 185188 20692 185194 20694
rect 187886 20248 187946 20694
rect 101030 20148 101036 20212
rect 101100 20210 101106 20212
rect 103430 20210 103490 20218
rect 101100 20150 103490 20210
rect 101100 20148 101106 20150
rect 50481 19802 50547 19805
rect 47862 19800 50547 19802
rect 47862 19744 50486 19800
rect 50542 19744 50547 19800
rect 47862 19742 50547 19744
rect 47862 19432 47922 19742
rect 50481 19739 50547 19742
rect 100989 19802 101055 19805
rect 134661 19802 134727 19805
rect 100989 19800 103490 19802
rect 100989 19744 100994 19800
rect 101050 19744 103490 19800
rect 100989 19742 103490 19744
rect 100989 19739 101055 19742
rect 103430 19738 103490 19742
rect 131766 19800 134727 19802
rect 131766 19744 134666 19800
rect 134722 19744 134727 19800
rect 131766 19742 134727 19744
rect 103430 19678 104012 19738
rect 131766 19704 131826 19742
rect 134661 19739 134727 19742
rect 185169 19802 185235 19805
rect 185169 19800 187946 19802
rect 185169 19744 185174 19800
rect 185230 19744 187946 19800
rect 185169 19742 187946 19744
rect 185169 19739 185235 19742
rect 187886 19704 187946 19742
rect 134753 19530 134819 19533
rect 131766 19528 134819 19530
rect 131766 19472 134758 19528
rect 134814 19472 134819 19528
rect 131766 19470 134819 19472
rect 50757 19258 50823 19261
rect 47862 19256 50823 19258
rect 47862 19200 50762 19256
rect 50818 19200 50823 19256
rect 47862 19198 50823 19200
rect 47862 18888 47922 19198
rect 50757 19195 50823 19198
rect 101081 19258 101147 19261
rect 101081 19256 103490 19258
rect 101081 19200 101086 19256
rect 101142 19200 103490 19256
rect 101081 19198 103490 19200
rect 101081 19195 101147 19198
rect 103430 19194 103490 19198
rect 103430 19134 104012 19194
rect 131766 19160 131826 19470
rect 134753 19467 134819 19470
rect 185261 19530 185327 19533
rect 185261 19528 187946 19530
rect 185261 19472 185266 19528
rect 185322 19472 187946 19528
rect 185261 19470 187946 19472
rect 185261 19467 185327 19470
rect 187886 19160 187946 19470
rect 151822 18518 152250 18578
rect 149749 18306 149815 18309
rect 151822 18306 151882 18518
rect 152190 18442 152250 18518
rect 152550 18442 152556 18444
rect 152190 18382 152556 18442
rect 152550 18380 152556 18382
rect 152620 18380 152626 18444
rect 211389 18442 211455 18445
rect 213454 18442 213460 18444
rect 211389 18440 213460 18442
rect 211389 18384 211394 18440
rect 211450 18384 213460 18440
rect 211389 18382 213460 18384
rect 211389 18379 211455 18382
rect 213454 18380 213460 18382
rect 213524 18380 213530 18444
rect 149749 18304 151882 18306
rect 149749 18248 149754 18304
rect 149810 18248 151882 18304
rect 149749 18246 151882 18248
rect 149749 18243 149815 18246
rect 129049 17082 129115 17085
rect 147030 17082 147036 17084
rect 129049 17080 147036 17082
rect 129049 17024 129054 17080
rect 129110 17024 147036 17080
rect 129049 17022 147036 17024
rect 129049 17019 129115 17022
rect 147030 17020 147036 17022
rect 147100 17020 147106 17084
rect 201821 17082 201887 17085
rect 212534 17082 212540 17084
rect 201821 17080 212540 17082
rect 201821 17024 201826 17080
rect 201882 17024 212540 17080
rect 201821 17022 212540 17024
rect 201821 17019 201887 17022
rect 212534 17020 212540 17022
rect 212604 17020 212610 17084
<< via3 >>
rect 23572 236524 23636 236588
rect 88524 235164 88588 235228
rect 139492 235224 139556 235228
rect 139492 235168 139506 235224
rect 139506 235168 139556 235224
rect 139492 235164 139556 235168
rect 171324 235164 171388 235228
rect 88524 208916 88588 208980
rect 171324 208916 171388 208980
rect 140228 195180 140292 195244
rect 209964 190752 210028 190756
rect 209964 190696 209978 190752
rect 209978 190696 210028 190752
rect 209964 190692 210028 190696
rect 193956 190556 194020 190620
rect 25780 178724 25844 178788
rect 41972 178588 42036 178652
rect 212540 164852 212604 164916
rect 139492 164716 139556 164780
rect 25780 163628 25844 163692
rect 41788 163764 41852 163828
rect 23572 157100 23636 157164
rect 62028 111132 62092 111196
rect 108396 111192 108460 111196
rect 108396 111136 108446 111192
rect 108446 111136 108460 111192
rect 108396 111132 108460 111136
rect 133972 111192 134036 111196
rect 133972 111136 134022 111192
rect 134022 111136 134036 111192
rect 133972 111132 134036 111136
rect 193772 96852 193836 96916
rect 209780 96716 209844 96780
rect 25596 76452 25660 76516
rect 41788 76452 41852 76516
rect 25780 69516 25844 69580
rect 41788 69788 41852 69852
rect 211436 69788 211500 69852
rect 211620 63124 211684 63188
rect 140228 58364 140292 58428
rect 152740 46940 152804 47004
rect 68836 46804 68900 46868
rect 149060 46804 149124 46868
rect 64972 46668 65036 46732
rect 146300 46668 146364 46732
rect 68468 46532 68532 46596
rect 152556 46532 152620 46596
rect 63500 46396 63564 46460
rect 62212 46260 62276 46324
rect 89812 46260 89876 46324
rect 147772 46396 147836 46460
rect 146116 46260 146180 46324
rect 63316 46124 63380 46188
rect 89076 46124 89140 46188
rect 147036 46124 147100 46188
rect 172980 46124 173044 46188
rect 173348 44764 173412 44828
rect 173900 44628 173964 44692
rect 19708 23208 19772 23272
rect 53932 22792 53996 22796
rect 53932 22736 53982 22792
rect 53982 22736 53996 22792
rect 53932 22732 53996 22736
rect 185124 21916 185188 21980
rect 62212 20964 62276 21028
rect 63316 21024 63380 21028
rect 63316 20968 63330 21024
rect 63330 20968 63380 21024
rect 63316 20964 63380 20968
rect 64972 20964 65036 21028
rect 68468 20964 68532 21028
rect 146300 21024 146364 21028
rect 146300 20968 146314 21024
rect 146314 20968 146364 21024
rect 146300 20964 146364 20968
rect 147772 21024 147836 21028
rect 147772 20968 147786 21024
rect 147786 20968 147836 21024
rect 147772 20964 147836 20968
rect 149060 20964 149124 21028
rect 63500 20828 63564 20892
rect 68836 20828 68900 20892
rect 101036 20828 101100 20892
rect 146116 20828 146180 20892
rect 185492 20828 185556 20892
rect 152740 20692 152804 20756
rect 185124 20692 185188 20756
rect 101036 20148 101100 20212
rect 152556 18380 152620 18444
rect 213460 18380 213524 18444
rect 147036 17020 147100 17084
rect 212540 17020 212604 17084
<< metal4 >>
rect 0 253078 4000 253200
rect 0 252842 122 253078
rect 358 252842 442 253078
rect 678 252842 762 253078
rect 998 252842 1082 253078
rect 1318 252842 1402 253078
rect 1638 252842 1722 253078
rect 1958 252842 2042 253078
rect 2278 252842 2362 253078
rect 2598 252842 2682 253078
rect 2918 252842 3002 253078
rect 3238 252842 3322 253078
rect 3558 252842 3642 253078
rect 3878 252842 4000 253078
rect 0 252758 4000 252842
rect 0 252522 122 252758
rect 358 252522 442 252758
rect 678 252522 762 252758
rect 998 252522 1082 252758
rect 1318 252522 1402 252758
rect 1638 252522 1722 252758
rect 1958 252522 2042 252758
rect 2278 252522 2362 252758
rect 2598 252522 2682 252758
rect 2918 252522 3002 252758
rect 3238 252522 3322 252758
rect 3558 252522 3642 252758
rect 3878 252522 4000 252758
rect 0 252438 4000 252522
rect 0 252202 122 252438
rect 358 252202 442 252438
rect 678 252202 762 252438
rect 998 252202 1082 252438
rect 1318 252202 1402 252438
rect 1638 252202 1722 252438
rect 1958 252202 2042 252438
rect 2278 252202 2362 252438
rect 2598 252202 2682 252438
rect 2918 252202 3002 252438
rect 3238 252202 3322 252438
rect 3558 252202 3642 252438
rect 3878 252202 4000 252438
rect 0 252118 4000 252202
rect 0 251882 122 252118
rect 358 251882 442 252118
rect 678 251882 762 252118
rect 998 251882 1082 252118
rect 1318 251882 1402 252118
rect 1638 251882 1722 252118
rect 1958 251882 2042 252118
rect 2278 251882 2362 252118
rect 2598 251882 2682 252118
rect 2918 251882 3002 252118
rect 3238 251882 3322 252118
rect 3558 251882 3642 252118
rect 3878 251882 4000 252118
rect 0 251798 4000 251882
rect 0 251562 122 251798
rect 358 251562 442 251798
rect 678 251562 762 251798
rect 998 251562 1082 251798
rect 1318 251562 1402 251798
rect 1638 251562 1722 251798
rect 1958 251562 2042 251798
rect 2278 251562 2362 251798
rect 2598 251562 2682 251798
rect 2918 251562 3002 251798
rect 3238 251562 3322 251798
rect 3558 251562 3642 251798
rect 3878 251562 4000 251798
rect 0 251478 4000 251562
rect 0 251242 122 251478
rect 358 251242 442 251478
rect 678 251242 762 251478
rect 998 251242 1082 251478
rect 1318 251242 1402 251478
rect 1638 251242 1722 251478
rect 1958 251242 2042 251478
rect 2278 251242 2362 251478
rect 2598 251242 2682 251478
rect 2918 251242 3002 251478
rect 3238 251242 3322 251478
rect 3558 251242 3642 251478
rect 3878 251242 4000 251478
rect 0 251158 4000 251242
rect 0 250922 122 251158
rect 358 250922 442 251158
rect 678 250922 762 251158
rect 998 250922 1082 251158
rect 1318 250922 1402 251158
rect 1638 250922 1722 251158
rect 1958 250922 2042 251158
rect 2278 250922 2362 251158
rect 2598 250922 2682 251158
rect 2918 250922 3002 251158
rect 3238 250922 3322 251158
rect 3558 250922 3642 251158
rect 3878 250922 4000 251158
rect 0 250838 4000 250922
rect 0 250602 122 250838
rect 358 250602 442 250838
rect 678 250602 762 250838
rect 998 250602 1082 250838
rect 1318 250602 1402 250838
rect 1638 250602 1722 250838
rect 1958 250602 2042 250838
rect 2278 250602 2362 250838
rect 2598 250602 2682 250838
rect 2918 250602 3002 250838
rect 3238 250602 3322 250838
rect 3558 250602 3642 250838
rect 3878 250602 4000 250838
rect 0 250518 4000 250602
rect 0 250282 122 250518
rect 358 250282 442 250518
rect 678 250282 762 250518
rect 998 250282 1082 250518
rect 1318 250282 1402 250518
rect 1638 250282 1722 250518
rect 1958 250282 2042 250518
rect 2278 250282 2362 250518
rect 2598 250282 2682 250518
rect 2918 250282 3002 250518
rect 3238 250282 3322 250518
rect 3558 250282 3642 250518
rect 3878 250282 4000 250518
rect 0 250198 4000 250282
rect 0 249962 122 250198
rect 358 249962 442 250198
rect 678 249962 762 250198
rect 998 249962 1082 250198
rect 1318 249962 1402 250198
rect 1638 249962 1722 250198
rect 1958 249962 2042 250198
rect 2278 249962 2362 250198
rect 2598 249962 2682 250198
rect 2918 249962 3002 250198
rect 3238 249962 3322 250198
rect 3558 249962 3642 250198
rect 3878 249962 4000 250198
rect 0 249878 4000 249962
rect 0 249642 122 249878
rect 358 249642 442 249878
rect 678 249642 762 249878
rect 998 249642 1082 249878
rect 1318 249642 1402 249878
rect 1638 249642 1722 249878
rect 1958 249642 2042 249878
rect 2278 249642 2362 249878
rect 2598 249642 2682 249878
rect 2918 249642 3002 249878
rect 3238 249642 3322 249878
rect 3558 249642 3642 249878
rect 3878 249642 4000 249878
rect 0 249558 4000 249642
rect 0 249322 122 249558
rect 358 249322 442 249558
rect 678 249322 762 249558
rect 998 249322 1082 249558
rect 1318 249322 1402 249558
rect 1638 249322 1722 249558
rect 1958 249322 2042 249558
rect 2278 249322 2362 249558
rect 2598 249322 2682 249558
rect 2918 249322 3002 249558
rect 3238 249322 3322 249558
rect 3558 249322 3642 249558
rect 3878 249322 4000 249558
rect 0 228918 4000 249322
rect 231716 253078 235716 253200
rect 231716 252842 231838 253078
rect 232074 252842 232158 253078
rect 232394 252842 232478 253078
rect 232714 252842 232798 253078
rect 233034 252842 233118 253078
rect 233354 252842 233438 253078
rect 233674 252842 233758 253078
rect 233994 252842 234078 253078
rect 234314 252842 234398 253078
rect 234634 252842 234718 253078
rect 234954 252842 235038 253078
rect 235274 252842 235358 253078
rect 235594 252842 235716 253078
rect 231716 252758 235716 252842
rect 231716 252522 231838 252758
rect 232074 252522 232158 252758
rect 232394 252522 232478 252758
rect 232714 252522 232798 252758
rect 233034 252522 233118 252758
rect 233354 252522 233438 252758
rect 233674 252522 233758 252758
rect 233994 252522 234078 252758
rect 234314 252522 234398 252758
rect 234634 252522 234718 252758
rect 234954 252522 235038 252758
rect 235274 252522 235358 252758
rect 235594 252522 235716 252758
rect 231716 252438 235716 252522
rect 231716 252202 231838 252438
rect 232074 252202 232158 252438
rect 232394 252202 232478 252438
rect 232714 252202 232798 252438
rect 233034 252202 233118 252438
rect 233354 252202 233438 252438
rect 233674 252202 233758 252438
rect 233994 252202 234078 252438
rect 234314 252202 234398 252438
rect 234634 252202 234718 252438
rect 234954 252202 235038 252438
rect 235274 252202 235358 252438
rect 235594 252202 235716 252438
rect 231716 252118 235716 252202
rect 231716 251882 231838 252118
rect 232074 251882 232158 252118
rect 232394 251882 232478 252118
rect 232714 251882 232798 252118
rect 233034 251882 233118 252118
rect 233354 251882 233438 252118
rect 233674 251882 233758 252118
rect 233994 251882 234078 252118
rect 234314 251882 234398 252118
rect 234634 251882 234718 252118
rect 234954 251882 235038 252118
rect 235274 251882 235358 252118
rect 235594 251882 235716 252118
rect 231716 251798 235716 251882
rect 231716 251562 231838 251798
rect 232074 251562 232158 251798
rect 232394 251562 232478 251798
rect 232714 251562 232798 251798
rect 233034 251562 233118 251798
rect 233354 251562 233438 251798
rect 233674 251562 233758 251798
rect 233994 251562 234078 251798
rect 234314 251562 234398 251798
rect 234634 251562 234718 251798
rect 234954 251562 235038 251798
rect 235274 251562 235358 251798
rect 235594 251562 235716 251798
rect 231716 251478 235716 251562
rect 231716 251242 231838 251478
rect 232074 251242 232158 251478
rect 232394 251242 232478 251478
rect 232714 251242 232798 251478
rect 233034 251242 233118 251478
rect 233354 251242 233438 251478
rect 233674 251242 233758 251478
rect 233994 251242 234078 251478
rect 234314 251242 234398 251478
rect 234634 251242 234718 251478
rect 234954 251242 235038 251478
rect 235274 251242 235358 251478
rect 235594 251242 235716 251478
rect 231716 251158 235716 251242
rect 231716 250922 231838 251158
rect 232074 250922 232158 251158
rect 232394 250922 232478 251158
rect 232714 250922 232798 251158
rect 233034 250922 233118 251158
rect 233354 250922 233438 251158
rect 233674 250922 233758 251158
rect 233994 250922 234078 251158
rect 234314 250922 234398 251158
rect 234634 250922 234718 251158
rect 234954 250922 235038 251158
rect 235274 250922 235358 251158
rect 235594 250922 235716 251158
rect 231716 250838 235716 250922
rect 231716 250602 231838 250838
rect 232074 250602 232158 250838
rect 232394 250602 232478 250838
rect 232714 250602 232798 250838
rect 233034 250602 233118 250838
rect 233354 250602 233438 250838
rect 233674 250602 233758 250838
rect 233994 250602 234078 250838
rect 234314 250602 234398 250838
rect 234634 250602 234718 250838
rect 234954 250602 235038 250838
rect 235274 250602 235358 250838
rect 235594 250602 235716 250838
rect 231716 250518 235716 250602
rect 231716 250282 231838 250518
rect 232074 250282 232158 250518
rect 232394 250282 232478 250518
rect 232714 250282 232798 250518
rect 233034 250282 233118 250518
rect 233354 250282 233438 250518
rect 233674 250282 233758 250518
rect 233994 250282 234078 250518
rect 234314 250282 234398 250518
rect 234634 250282 234718 250518
rect 234954 250282 235038 250518
rect 235274 250282 235358 250518
rect 235594 250282 235716 250518
rect 231716 250198 235716 250282
rect 231716 249962 231838 250198
rect 232074 249962 232158 250198
rect 232394 249962 232478 250198
rect 232714 249962 232798 250198
rect 233034 249962 233118 250198
rect 233354 249962 233438 250198
rect 233674 249962 233758 250198
rect 233994 249962 234078 250198
rect 234314 249962 234398 250198
rect 234634 249962 234718 250198
rect 234954 249962 235038 250198
rect 235274 249962 235358 250198
rect 235594 249962 235716 250198
rect 231716 249878 235716 249962
rect 231716 249642 231838 249878
rect 232074 249642 232158 249878
rect 232394 249642 232478 249878
rect 232714 249642 232798 249878
rect 233034 249642 233118 249878
rect 233354 249642 233438 249878
rect 233674 249642 233758 249878
rect 233994 249642 234078 249878
rect 234314 249642 234398 249878
rect 234634 249642 234718 249878
rect 234954 249642 235038 249878
rect 235274 249642 235358 249878
rect 235594 249642 235716 249878
rect 231716 249558 235716 249642
rect 231716 249322 231838 249558
rect 232074 249322 232158 249558
rect 232394 249322 232478 249558
rect 232714 249322 232798 249558
rect 233034 249322 233118 249558
rect 233354 249322 233438 249558
rect 233674 249322 233758 249558
rect 233994 249322 234078 249558
rect 234314 249322 234398 249558
rect 234634 249322 234718 249558
rect 234954 249322 235038 249558
rect 235274 249322 235358 249558
rect 235594 249322 235716 249558
rect 0 228682 122 228918
rect 358 228682 442 228918
rect 678 228682 762 228918
rect 998 228682 1082 228918
rect 1318 228682 1402 228918
rect 1638 228682 1722 228918
rect 1958 228682 2042 228918
rect 2278 228682 2362 228918
rect 2598 228682 2682 228918
rect 2918 228682 3002 228918
rect 3238 228682 3322 228918
rect 3558 228682 3642 228918
rect 3878 228682 4000 228918
rect 0 206518 4000 228682
rect 0 206282 122 206518
rect 358 206282 442 206518
rect 678 206282 762 206518
rect 998 206282 1082 206518
rect 1318 206282 1402 206518
rect 1638 206282 1722 206518
rect 1958 206282 2042 206518
rect 2278 206282 2362 206518
rect 2598 206282 2682 206518
rect 2918 206282 3002 206518
rect 3238 206282 3322 206518
rect 3558 206282 3642 206518
rect 3878 206282 4000 206518
rect 0 184118 4000 206282
rect 0 183882 122 184118
rect 358 183882 442 184118
rect 678 183882 762 184118
rect 998 183882 1082 184118
rect 1318 183882 1402 184118
rect 1638 183882 1722 184118
rect 1958 183882 2042 184118
rect 2278 183882 2362 184118
rect 2598 183882 2682 184118
rect 2918 183882 3002 184118
rect 3238 183882 3322 184118
rect 3558 183882 3642 184118
rect 3878 183882 4000 184118
rect 0 161718 4000 183882
rect 0 161482 122 161718
rect 358 161482 442 161718
rect 678 161482 762 161718
rect 998 161482 1082 161718
rect 1318 161482 1402 161718
rect 1638 161482 1722 161718
rect 1958 161482 2042 161718
rect 2278 161482 2362 161718
rect 2598 161482 2682 161718
rect 2918 161482 3002 161718
rect 3238 161482 3322 161718
rect 3558 161482 3642 161718
rect 3878 161482 4000 161718
rect 0 139318 4000 161482
rect 0 139082 122 139318
rect 358 139082 442 139318
rect 678 139082 762 139318
rect 998 139082 1082 139318
rect 1318 139082 1402 139318
rect 1638 139082 1722 139318
rect 1958 139082 2042 139318
rect 2278 139082 2362 139318
rect 2598 139082 2682 139318
rect 2918 139082 3002 139318
rect 3238 139082 3322 139318
rect 3558 139082 3642 139318
rect 3878 139082 4000 139318
rect 0 116918 4000 139082
rect 0 116682 122 116918
rect 358 116682 442 116918
rect 678 116682 762 116918
rect 998 116682 1082 116918
rect 1318 116682 1402 116918
rect 1638 116682 1722 116918
rect 1958 116682 2042 116918
rect 2278 116682 2362 116918
rect 2598 116682 2682 116918
rect 2918 116682 3002 116918
rect 3238 116682 3322 116918
rect 3558 116682 3642 116918
rect 3878 116682 4000 116918
rect 0 94518 4000 116682
rect 0 94282 122 94518
rect 358 94282 442 94518
rect 678 94282 762 94518
rect 998 94282 1082 94518
rect 1318 94282 1402 94518
rect 1638 94282 1722 94518
rect 1958 94282 2042 94518
rect 2278 94282 2362 94518
rect 2598 94282 2682 94518
rect 2918 94282 3002 94518
rect 3238 94282 3322 94518
rect 3558 94282 3642 94518
rect 3878 94282 4000 94518
rect 0 72118 4000 94282
rect 0 71882 122 72118
rect 358 71882 442 72118
rect 678 71882 762 72118
rect 998 71882 1082 72118
rect 1318 71882 1402 72118
rect 1638 71882 1722 72118
rect 1958 71882 2042 72118
rect 2278 71882 2362 72118
rect 2598 71882 2682 72118
rect 2918 71882 3002 72118
rect 3238 71882 3322 72118
rect 3558 71882 3642 72118
rect 3878 71882 4000 72118
rect 0 49718 4000 71882
rect 0 49482 122 49718
rect 358 49482 442 49718
rect 678 49482 762 49718
rect 998 49482 1082 49718
rect 1318 49482 1402 49718
rect 1638 49482 1722 49718
rect 1958 49482 2042 49718
rect 2278 49482 2362 49718
rect 2598 49482 2682 49718
rect 2918 49482 3002 49718
rect 3238 49482 3322 49718
rect 3558 49482 3642 49718
rect 3878 49482 4000 49718
rect 0 27318 4000 49482
rect 0 27082 122 27318
rect 358 27082 442 27318
rect 678 27082 762 27318
rect 998 27082 1082 27318
rect 1318 27082 1402 27318
rect 1638 27082 1722 27318
rect 1958 27082 2042 27318
rect 2278 27082 2362 27318
rect 2598 27082 2682 27318
rect 2918 27082 3002 27318
rect 3238 27082 3322 27318
rect 3558 27082 3642 27318
rect 3878 27082 4000 27318
rect 0 3878 4000 27082
rect 5000 248078 9000 248200
rect 5000 247842 5122 248078
rect 5358 247842 5442 248078
rect 5678 247842 5762 248078
rect 5998 247842 6082 248078
rect 6318 247842 6402 248078
rect 6638 247842 6722 248078
rect 6958 247842 7042 248078
rect 7278 247842 7362 248078
rect 7598 247842 7682 248078
rect 7918 247842 8002 248078
rect 8238 247842 8322 248078
rect 8558 247842 8642 248078
rect 8878 247842 9000 248078
rect 5000 247758 9000 247842
rect 5000 247522 5122 247758
rect 5358 247522 5442 247758
rect 5678 247522 5762 247758
rect 5998 247522 6082 247758
rect 6318 247522 6402 247758
rect 6638 247522 6722 247758
rect 6958 247522 7042 247758
rect 7278 247522 7362 247758
rect 7598 247522 7682 247758
rect 7918 247522 8002 247758
rect 8238 247522 8322 247758
rect 8558 247522 8642 247758
rect 8878 247522 9000 247758
rect 5000 247438 9000 247522
rect 5000 247202 5122 247438
rect 5358 247202 5442 247438
rect 5678 247202 5762 247438
rect 5998 247202 6082 247438
rect 6318 247202 6402 247438
rect 6638 247202 6722 247438
rect 6958 247202 7042 247438
rect 7278 247202 7362 247438
rect 7598 247202 7682 247438
rect 7918 247202 8002 247438
rect 8238 247202 8322 247438
rect 8558 247202 8642 247438
rect 8878 247202 9000 247438
rect 5000 247118 9000 247202
rect 5000 246882 5122 247118
rect 5358 246882 5442 247118
rect 5678 246882 5762 247118
rect 5998 246882 6082 247118
rect 6318 246882 6402 247118
rect 6638 246882 6722 247118
rect 6958 246882 7042 247118
rect 7278 246882 7362 247118
rect 7598 246882 7682 247118
rect 7918 246882 8002 247118
rect 8238 246882 8322 247118
rect 8558 246882 8642 247118
rect 8878 246882 9000 247118
rect 5000 246798 9000 246882
rect 5000 246562 5122 246798
rect 5358 246562 5442 246798
rect 5678 246562 5762 246798
rect 5998 246562 6082 246798
rect 6318 246562 6402 246798
rect 6638 246562 6722 246798
rect 6958 246562 7042 246798
rect 7278 246562 7362 246798
rect 7598 246562 7682 246798
rect 7918 246562 8002 246798
rect 8238 246562 8322 246798
rect 8558 246562 8642 246798
rect 8878 246562 9000 246798
rect 5000 246478 9000 246562
rect 5000 246242 5122 246478
rect 5358 246242 5442 246478
rect 5678 246242 5762 246478
rect 5998 246242 6082 246478
rect 6318 246242 6402 246478
rect 6638 246242 6722 246478
rect 6958 246242 7042 246478
rect 7278 246242 7362 246478
rect 7598 246242 7682 246478
rect 7918 246242 8002 246478
rect 8238 246242 8322 246478
rect 8558 246242 8642 246478
rect 8878 246242 9000 246478
rect 5000 246158 9000 246242
rect 5000 245922 5122 246158
rect 5358 245922 5442 246158
rect 5678 245922 5762 246158
rect 5998 245922 6082 246158
rect 6318 245922 6402 246158
rect 6638 245922 6722 246158
rect 6958 245922 7042 246158
rect 7278 245922 7362 246158
rect 7598 245922 7682 246158
rect 7918 245922 8002 246158
rect 8238 245922 8322 246158
rect 8558 245922 8642 246158
rect 8878 245922 9000 246158
rect 5000 245838 9000 245922
rect 5000 245602 5122 245838
rect 5358 245602 5442 245838
rect 5678 245602 5762 245838
rect 5998 245602 6082 245838
rect 6318 245602 6402 245838
rect 6638 245602 6722 245838
rect 6958 245602 7042 245838
rect 7278 245602 7362 245838
rect 7598 245602 7682 245838
rect 7918 245602 8002 245838
rect 8238 245602 8322 245838
rect 8558 245602 8642 245838
rect 8878 245602 9000 245838
rect 5000 245518 9000 245602
rect 5000 245282 5122 245518
rect 5358 245282 5442 245518
rect 5678 245282 5762 245518
rect 5998 245282 6082 245518
rect 6318 245282 6402 245518
rect 6638 245282 6722 245518
rect 6958 245282 7042 245518
rect 7278 245282 7362 245518
rect 7598 245282 7682 245518
rect 7918 245282 8002 245518
rect 8238 245282 8322 245518
rect 8558 245282 8642 245518
rect 8878 245282 9000 245518
rect 5000 245198 9000 245282
rect 5000 244962 5122 245198
rect 5358 244962 5442 245198
rect 5678 244962 5762 245198
rect 5998 244962 6082 245198
rect 6318 244962 6402 245198
rect 6638 244962 6722 245198
rect 6958 244962 7042 245198
rect 7278 244962 7362 245198
rect 7598 244962 7682 245198
rect 7918 244962 8002 245198
rect 8238 244962 8322 245198
rect 8558 244962 8642 245198
rect 8878 244962 9000 245198
rect 5000 244878 9000 244962
rect 5000 244642 5122 244878
rect 5358 244642 5442 244878
rect 5678 244642 5762 244878
rect 5998 244642 6082 244878
rect 6318 244642 6402 244878
rect 6638 244642 6722 244878
rect 6958 244642 7042 244878
rect 7278 244642 7362 244878
rect 7598 244642 7682 244878
rect 7918 244642 8002 244878
rect 8238 244642 8322 244878
rect 8558 244642 8642 244878
rect 8878 244642 9000 244878
rect 5000 244558 9000 244642
rect 5000 244322 5122 244558
rect 5358 244322 5442 244558
rect 5678 244322 5762 244558
rect 5998 244322 6082 244558
rect 6318 244322 6402 244558
rect 6638 244322 6722 244558
rect 6958 244322 7042 244558
rect 7278 244322 7362 244558
rect 7598 244322 7682 244558
rect 7918 244322 8002 244558
rect 8238 244322 8322 244558
rect 8558 244322 8642 244558
rect 8878 244322 9000 244558
rect 5000 240118 9000 244322
rect 5000 239882 5122 240118
rect 5358 239882 5442 240118
rect 5678 239882 5762 240118
rect 5998 239882 6082 240118
rect 6318 239882 6402 240118
rect 6638 239882 6722 240118
rect 6958 239882 7042 240118
rect 7278 239882 7362 240118
rect 7598 239882 7682 240118
rect 7918 239882 8002 240118
rect 8238 239882 8322 240118
rect 8558 239882 8642 240118
rect 8878 239882 9000 240118
rect 5000 217718 9000 239882
rect 226716 248078 230716 248200
rect 226716 247842 226838 248078
rect 227074 247842 227158 248078
rect 227394 247842 227478 248078
rect 227714 247842 227798 248078
rect 228034 247842 228118 248078
rect 228354 247842 228438 248078
rect 228674 247842 228758 248078
rect 228994 247842 229078 248078
rect 229314 247842 229398 248078
rect 229634 247842 229718 248078
rect 229954 247842 230038 248078
rect 230274 247842 230358 248078
rect 230594 247842 230716 248078
rect 226716 247758 230716 247842
rect 226716 247522 226838 247758
rect 227074 247522 227158 247758
rect 227394 247522 227478 247758
rect 227714 247522 227798 247758
rect 228034 247522 228118 247758
rect 228354 247522 228438 247758
rect 228674 247522 228758 247758
rect 228994 247522 229078 247758
rect 229314 247522 229398 247758
rect 229634 247522 229718 247758
rect 229954 247522 230038 247758
rect 230274 247522 230358 247758
rect 230594 247522 230716 247758
rect 226716 247438 230716 247522
rect 226716 247202 226838 247438
rect 227074 247202 227158 247438
rect 227394 247202 227478 247438
rect 227714 247202 227798 247438
rect 228034 247202 228118 247438
rect 228354 247202 228438 247438
rect 228674 247202 228758 247438
rect 228994 247202 229078 247438
rect 229314 247202 229398 247438
rect 229634 247202 229718 247438
rect 229954 247202 230038 247438
rect 230274 247202 230358 247438
rect 230594 247202 230716 247438
rect 226716 247118 230716 247202
rect 226716 246882 226838 247118
rect 227074 246882 227158 247118
rect 227394 246882 227478 247118
rect 227714 246882 227798 247118
rect 228034 246882 228118 247118
rect 228354 246882 228438 247118
rect 228674 246882 228758 247118
rect 228994 246882 229078 247118
rect 229314 246882 229398 247118
rect 229634 246882 229718 247118
rect 229954 246882 230038 247118
rect 230274 246882 230358 247118
rect 230594 246882 230716 247118
rect 226716 246798 230716 246882
rect 226716 246562 226838 246798
rect 227074 246562 227158 246798
rect 227394 246562 227478 246798
rect 227714 246562 227798 246798
rect 228034 246562 228118 246798
rect 228354 246562 228438 246798
rect 228674 246562 228758 246798
rect 228994 246562 229078 246798
rect 229314 246562 229398 246798
rect 229634 246562 229718 246798
rect 229954 246562 230038 246798
rect 230274 246562 230358 246798
rect 230594 246562 230716 246798
rect 226716 246478 230716 246562
rect 226716 246242 226838 246478
rect 227074 246242 227158 246478
rect 227394 246242 227478 246478
rect 227714 246242 227798 246478
rect 228034 246242 228118 246478
rect 228354 246242 228438 246478
rect 228674 246242 228758 246478
rect 228994 246242 229078 246478
rect 229314 246242 229398 246478
rect 229634 246242 229718 246478
rect 229954 246242 230038 246478
rect 230274 246242 230358 246478
rect 230594 246242 230716 246478
rect 226716 246158 230716 246242
rect 226716 245922 226838 246158
rect 227074 245922 227158 246158
rect 227394 245922 227478 246158
rect 227714 245922 227798 246158
rect 228034 245922 228118 246158
rect 228354 245922 228438 246158
rect 228674 245922 228758 246158
rect 228994 245922 229078 246158
rect 229314 245922 229398 246158
rect 229634 245922 229718 246158
rect 229954 245922 230038 246158
rect 230274 245922 230358 246158
rect 230594 245922 230716 246158
rect 226716 245838 230716 245922
rect 226716 245602 226838 245838
rect 227074 245602 227158 245838
rect 227394 245602 227478 245838
rect 227714 245602 227798 245838
rect 228034 245602 228118 245838
rect 228354 245602 228438 245838
rect 228674 245602 228758 245838
rect 228994 245602 229078 245838
rect 229314 245602 229398 245838
rect 229634 245602 229718 245838
rect 229954 245602 230038 245838
rect 230274 245602 230358 245838
rect 230594 245602 230716 245838
rect 226716 245518 230716 245602
rect 226716 245282 226838 245518
rect 227074 245282 227158 245518
rect 227394 245282 227478 245518
rect 227714 245282 227798 245518
rect 228034 245282 228118 245518
rect 228354 245282 228438 245518
rect 228674 245282 228758 245518
rect 228994 245282 229078 245518
rect 229314 245282 229398 245518
rect 229634 245282 229718 245518
rect 229954 245282 230038 245518
rect 230274 245282 230358 245518
rect 230594 245282 230716 245518
rect 226716 245198 230716 245282
rect 226716 244962 226838 245198
rect 227074 244962 227158 245198
rect 227394 244962 227478 245198
rect 227714 244962 227798 245198
rect 228034 244962 228118 245198
rect 228354 244962 228438 245198
rect 228674 244962 228758 245198
rect 228994 244962 229078 245198
rect 229314 244962 229398 245198
rect 229634 244962 229718 245198
rect 229954 244962 230038 245198
rect 230274 244962 230358 245198
rect 230594 244962 230716 245198
rect 226716 244878 230716 244962
rect 226716 244642 226838 244878
rect 227074 244642 227158 244878
rect 227394 244642 227478 244878
rect 227714 244642 227798 244878
rect 228034 244642 228118 244878
rect 228354 244642 228438 244878
rect 228674 244642 228758 244878
rect 228994 244642 229078 244878
rect 229314 244642 229398 244878
rect 229634 244642 229718 244878
rect 229954 244642 230038 244878
rect 230274 244642 230358 244878
rect 230594 244642 230716 244878
rect 226716 244558 230716 244642
rect 226716 244322 226838 244558
rect 227074 244322 227158 244558
rect 227394 244322 227478 244558
rect 227714 244322 227798 244558
rect 228034 244322 228118 244558
rect 228354 244322 228438 244558
rect 228674 244322 228758 244558
rect 228994 244322 229078 244558
rect 229314 244322 229398 244558
rect 229634 244322 229718 244558
rect 229954 244322 230038 244558
rect 230274 244322 230358 244558
rect 230594 244322 230716 244558
rect 226716 240118 230716 244322
rect 226716 239882 226838 240118
rect 227074 239882 227158 240118
rect 227394 239882 227478 240118
rect 227714 239882 227798 240118
rect 228034 239882 228118 240118
rect 228354 239882 228438 240118
rect 228674 239882 228758 240118
rect 228994 239882 229078 240118
rect 229314 239882 229398 240118
rect 229634 239882 229718 240118
rect 229954 239882 230038 240118
rect 230274 239882 230358 240118
rect 230594 239882 230716 240118
rect 23571 236588 23637 236589
rect 23571 236524 23572 236588
rect 23636 236524 23637 236588
rect 23571 236523 23637 236524
rect 5000 217482 5122 217718
rect 5358 217482 5442 217718
rect 5678 217482 5762 217718
rect 5998 217482 6082 217718
rect 6318 217482 6402 217718
rect 6638 217482 6722 217718
rect 6958 217482 7042 217718
rect 7278 217482 7362 217718
rect 7598 217482 7682 217718
rect 7918 217482 8002 217718
rect 8238 217482 8322 217718
rect 8558 217482 8642 217718
rect 8878 217482 9000 217718
rect 5000 195318 9000 217482
rect 5000 195082 5122 195318
rect 5358 195082 5442 195318
rect 5678 195082 5762 195318
rect 5998 195082 6082 195318
rect 6318 195082 6402 195318
rect 6638 195082 6722 195318
rect 6958 195082 7042 195318
rect 7278 195082 7362 195318
rect 7598 195082 7682 195318
rect 7918 195082 8002 195318
rect 8238 195082 8322 195318
rect 8558 195082 8642 195318
rect 8878 195082 9000 195318
rect 5000 172918 9000 195082
rect 5000 172682 5122 172918
rect 5358 172682 5442 172918
rect 5678 172682 5762 172918
rect 5998 172682 6082 172918
rect 6318 172682 6402 172918
rect 6638 172682 6722 172918
rect 6958 172682 7042 172918
rect 7278 172682 7362 172918
rect 7598 172682 7682 172918
rect 7918 172682 8002 172918
rect 8238 172682 8322 172918
rect 8558 172682 8642 172918
rect 8878 172682 9000 172918
rect 5000 150518 9000 172682
rect 23574 157165 23634 236523
rect 88523 235228 88589 235229
rect 88523 235164 88524 235228
rect 88588 235164 88589 235228
rect 88523 235163 88589 235164
rect 139491 235228 139557 235229
rect 139491 235164 139492 235228
rect 139556 235164 139557 235228
rect 139491 235163 139557 235164
rect 171323 235228 171389 235229
rect 171323 235164 171324 235228
rect 171388 235164 171389 235228
rect 171323 235163 171389 235164
rect 29885 228918 30205 228960
rect 29885 228682 29927 228918
rect 30163 228682 30205 228918
rect 29885 228640 30205 228682
rect 71840 228918 72160 228960
rect 71840 228682 71882 228918
rect 72118 228682 72160 228918
rect 71840 228640 72160 228682
rect 25219 217718 25539 217760
rect 25219 217482 25261 217718
rect 25497 217482 25539 217718
rect 25219 217440 25539 217482
rect 66840 217718 67160 217760
rect 66840 217482 66882 217718
rect 67118 217482 67160 217718
rect 66840 217440 67160 217482
rect 88526 208981 88586 235163
rect 114173 228918 114493 228960
rect 114173 228682 114215 228918
rect 114451 228682 114493 228918
rect 114173 228640 114493 228682
rect 109507 217718 109827 217760
rect 109507 217482 109549 217718
rect 109785 217482 109827 217718
rect 109507 217440 109827 217482
rect 88523 208980 88589 208981
rect 88523 208916 88524 208980
rect 88588 208916 88589 208980
rect 88523 208915 88589 208916
rect 32173 184118 32493 184160
rect 32173 183882 32215 184118
rect 32451 183882 32493 184118
rect 32173 183840 32493 183882
rect 75464 184118 75784 184160
rect 75464 183882 75506 184118
rect 75742 183882 75784 184118
rect 75464 183840 75784 183882
rect 116173 184118 116493 184160
rect 116173 183882 116215 184118
rect 116451 183882 116493 184118
rect 116173 183840 116493 183882
rect 25779 178788 25845 178789
rect 25779 178724 25780 178788
rect 25844 178786 25845 178788
rect 25844 178726 26578 178786
rect 25844 178724 25845 178726
rect 25779 178723 25845 178724
rect 26518 178602 26578 178726
rect 41971 178652 42037 178653
rect 41971 178602 41972 178652
rect 42036 178602 42037 178652
rect 29507 172918 29827 172960
rect 29507 172682 29549 172918
rect 29785 172682 29827 172918
rect 29507 172640 29827 172682
rect 60104 172918 60424 172960
rect 60104 172682 60146 172918
rect 60382 172682 60424 172918
rect 60104 172640 60424 172682
rect 113507 172918 113827 172960
rect 113507 172682 113549 172918
rect 113785 172682 113827 172918
rect 113507 172640 113827 172682
rect 139494 165002 139554 235163
rect 155840 228918 156160 228960
rect 155840 228682 155882 228918
rect 156118 228682 156160 228918
rect 155840 228640 156160 228682
rect 150840 217718 151160 217760
rect 150840 217482 150882 217718
rect 151118 217482 151160 217718
rect 150840 217440 151160 217482
rect 171326 208981 171386 235163
rect 198173 228918 198493 228960
rect 198173 228682 198215 228918
rect 198451 228682 198493 228918
rect 198173 228640 198493 228682
rect 193507 217718 193827 217760
rect 193507 217482 193549 217718
rect 193785 217482 193827 217718
rect 193507 217440 193827 217482
rect 226716 217718 230716 239882
rect 226716 217482 226838 217718
rect 227074 217482 227158 217718
rect 227394 217482 227478 217718
rect 227714 217482 227798 217718
rect 228034 217482 228118 217718
rect 228354 217482 228438 217718
rect 228674 217482 228758 217718
rect 228994 217482 229078 217718
rect 229314 217482 229398 217718
rect 229634 217482 229718 217718
rect 229954 217482 230038 217718
rect 230274 217482 230358 217718
rect 230594 217482 230716 217718
rect 171323 208980 171389 208981
rect 171323 208916 171324 208980
rect 171388 208916 171389 208980
rect 171323 208915 171389 208916
rect 226716 195318 230716 217482
rect 140227 195244 140293 195245
rect 140227 195180 140228 195244
rect 140292 195180 140293 195244
rect 140227 195179 140293 195180
rect 139491 164716 139492 164766
rect 139556 164716 139557 164766
rect 139491 164715 139557 164716
rect 41787 163828 41853 163829
rect 25782 163766 26578 163826
rect 25782 163693 25842 163766
rect 25779 163692 25845 163693
rect 25779 163628 25780 163692
rect 25844 163628 25845 163692
rect 26518 163642 26578 163766
rect 41787 163764 41788 163828
rect 41852 163764 41853 163828
rect 41787 163763 41853 163764
rect 41790 163642 41850 163763
rect 25779 163627 25845 163628
rect 32173 161718 32493 161760
rect 32173 161482 32215 161718
rect 32451 161482 32493 161718
rect 32173 161440 32493 161482
rect 75464 161718 75784 161760
rect 75464 161482 75506 161718
rect 75742 161482 75784 161718
rect 75464 161440 75784 161482
rect 116173 161718 116493 161760
rect 116173 161482 116215 161718
rect 116451 161482 116493 161718
rect 116173 161440 116493 161482
rect 23571 157164 23637 157165
rect 23571 157100 23572 157164
rect 23636 157100 23637 157164
rect 23571 157099 23637 157100
rect 5000 150282 5122 150518
rect 5358 150282 5442 150518
rect 5678 150282 5762 150518
rect 5998 150282 6082 150518
rect 6318 150282 6402 150518
rect 6638 150282 6722 150518
rect 6958 150282 7042 150518
rect 7278 150282 7362 150518
rect 7598 150282 7682 150518
rect 7918 150282 8002 150518
rect 8238 150282 8322 150518
rect 8558 150282 8642 150518
rect 8878 150282 9000 150518
rect 5000 128118 9000 150282
rect 5000 127882 5122 128118
rect 5358 127882 5442 128118
rect 5678 127882 5762 128118
rect 5998 127882 6082 128118
rect 6318 127882 6402 128118
rect 6638 127882 6722 128118
rect 6958 127882 7042 128118
rect 7278 127882 7362 128118
rect 7598 127882 7682 128118
rect 7918 127882 8002 128118
rect 8238 127882 8322 128118
rect 8558 127882 8642 128118
rect 8878 127882 9000 128118
rect 5000 105718 9000 127882
rect 25507 128118 25827 128160
rect 25507 127882 25549 128118
rect 25785 127882 25827 128118
rect 25507 127840 25827 127882
rect 66840 128118 67160 128160
rect 66840 127882 66882 128118
rect 67118 127882 67160 128118
rect 66840 127840 67160 127882
rect 109507 128118 109827 128160
rect 109507 127882 109549 128118
rect 109785 127882 109827 128118
rect 109507 127840 109827 127882
rect 30173 116918 30493 116960
rect 30173 116682 30215 116918
rect 30451 116682 30493 116918
rect 30173 116640 30493 116682
rect 114173 116918 114493 116960
rect 114173 116682 114215 116918
rect 114451 116682 114493 116918
rect 114173 116640 114493 116682
rect 5000 105482 5122 105718
rect 5358 105482 5442 105718
rect 5678 105482 5762 105718
rect 5998 105482 6082 105718
rect 6318 105482 6402 105718
rect 6638 105482 6722 105718
rect 6958 105482 7042 105718
rect 7278 105482 7362 105718
rect 7598 105482 7682 105718
rect 7918 105482 8002 105718
rect 8238 105482 8322 105718
rect 8558 105482 8642 105718
rect 8878 105482 9000 105718
rect 5000 83318 9000 105482
rect 32173 94518 32493 94560
rect 32173 94282 32215 94518
rect 32451 94282 32493 94518
rect 32173 94240 32493 94282
rect 75464 94518 75784 94560
rect 75464 94282 75506 94518
rect 75742 94282 75784 94518
rect 75464 94240 75784 94282
rect 116173 94518 116493 94560
rect 116173 94282 116215 94518
rect 116451 94282 116493 94518
rect 116173 94240 116493 94282
rect 5000 83082 5122 83318
rect 5358 83082 5442 83318
rect 5678 83082 5762 83318
rect 5998 83082 6082 83318
rect 6318 83082 6402 83318
rect 6638 83082 6722 83318
rect 6958 83082 7042 83318
rect 7278 83082 7362 83318
rect 7598 83082 7682 83318
rect 7918 83082 8002 83318
rect 8238 83082 8322 83318
rect 8558 83082 8642 83318
rect 8878 83082 9000 83318
rect 5000 60918 9000 83082
rect 29507 83318 29827 83360
rect 29507 83082 29549 83318
rect 29785 83082 29827 83318
rect 29507 83040 29827 83082
rect 60104 83318 60424 83360
rect 60104 83082 60146 83318
rect 60382 83082 60424 83318
rect 60104 83040 60424 83082
rect 113507 83318 113827 83360
rect 113507 83082 113549 83318
rect 113785 83082 113827 83318
rect 113507 83040 113827 83082
rect 32173 72118 32493 72160
rect 32173 71882 32215 72118
rect 32451 71882 32493 72118
rect 32173 71840 32493 71882
rect 75464 72118 75784 72160
rect 75464 71882 75506 72118
rect 75742 71882 75784 72118
rect 75464 71840 75784 71882
rect 116173 72118 116493 72160
rect 116173 71882 116215 72118
rect 116451 71882 116493 72118
rect 116173 71840 116493 71882
rect 41787 69852 41853 69853
rect 41787 69802 41788 69852
rect 41852 69802 41853 69852
rect 25779 69516 25780 69566
rect 25844 69516 25845 69566
rect 25779 69515 25845 69516
rect 5000 60682 5122 60918
rect 5358 60682 5442 60918
rect 5678 60682 5762 60918
rect 5998 60682 6082 60918
rect 6318 60682 6402 60918
rect 6638 60682 6722 60918
rect 6958 60682 7042 60918
rect 7278 60682 7362 60918
rect 7598 60682 7682 60918
rect 7918 60682 8002 60918
rect 8238 60682 8322 60918
rect 8558 60682 8642 60918
rect 8878 60682 9000 60918
rect 5000 38518 9000 60682
rect 140230 58429 140290 195179
rect 226716 195082 226838 195318
rect 227074 195082 227158 195318
rect 227394 195082 227478 195318
rect 227714 195082 227798 195318
rect 228034 195082 228118 195318
rect 228354 195082 228438 195318
rect 228674 195082 228758 195318
rect 228994 195082 229078 195318
rect 229314 195082 229398 195318
rect 229634 195082 229718 195318
rect 229954 195082 230038 195318
rect 230274 195082 230358 195318
rect 230594 195082 230716 195318
rect 193955 190556 193956 190606
rect 194020 190556 194021 190606
rect 193955 190555 194021 190556
rect 159464 184118 159784 184160
rect 159464 183882 159506 184118
rect 159742 183882 159784 184118
rect 159464 183840 159784 183882
rect 200173 184118 200493 184160
rect 200173 183882 200215 184118
rect 200451 183882 200493 184118
rect 200173 183840 200493 183882
rect 144104 172918 144424 172960
rect 144104 172682 144146 172918
rect 144382 172682 144424 172918
rect 144104 172640 144424 172682
rect 197507 172918 197827 172960
rect 197507 172682 197549 172918
rect 197785 172682 197827 172918
rect 197507 172640 197827 172682
rect 226716 172918 230716 195082
rect 226716 172682 226838 172918
rect 227074 172682 227158 172918
rect 227394 172682 227478 172918
rect 227714 172682 227798 172918
rect 228034 172682 228118 172918
rect 228354 172682 228438 172918
rect 228674 172682 228758 172918
rect 228994 172682 229078 172918
rect 229314 172682 229398 172918
rect 229634 172682 229718 172918
rect 229954 172682 230038 172918
rect 230274 172682 230358 172918
rect 230594 172682 230716 172918
rect 159464 161718 159784 161760
rect 159464 161482 159506 161718
rect 159742 161482 159784 161718
rect 159464 161440 159784 161482
rect 200173 161718 200493 161760
rect 200173 161482 200215 161718
rect 200451 161482 200493 161718
rect 200173 161440 200493 161482
rect 226716 150518 230716 172682
rect 226716 150282 226838 150518
rect 227074 150282 227158 150518
rect 227394 150282 227478 150518
rect 227714 150282 227798 150518
rect 228034 150282 228118 150518
rect 228354 150282 228438 150518
rect 228674 150282 228758 150518
rect 228994 150282 229078 150518
rect 229314 150282 229398 150518
rect 229634 150282 229718 150518
rect 229954 150282 230038 150518
rect 230274 150282 230358 150518
rect 230594 150282 230716 150518
rect 150840 128118 151160 128160
rect 150840 127882 150882 128118
rect 151118 127882 151160 128118
rect 150840 127840 151160 127882
rect 193507 128118 193827 128160
rect 193507 127882 193549 128118
rect 193785 127882 193827 128118
rect 193507 127840 193827 127882
rect 226716 128118 230716 150282
rect 226716 127882 226838 128118
rect 227074 127882 227158 128118
rect 227394 127882 227478 128118
rect 227714 127882 227798 128118
rect 228034 127882 228118 128118
rect 228354 127882 228438 128118
rect 228674 127882 228758 128118
rect 228994 127882 229078 128118
rect 229314 127882 229398 128118
rect 229634 127882 229718 128118
rect 229954 127882 230038 128118
rect 230274 127882 230358 128118
rect 230594 127882 230716 128118
rect 198173 116918 198493 116960
rect 198173 116682 198215 116918
rect 198451 116682 198493 116918
rect 198173 116640 198493 116682
rect 226716 105718 230716 127882
rect 226716 105482 226838 105718
rect 227074 105482 227158 105718
rect 227394 105482 227478 105718
rect 227714 105482 227798 105718
rect 228034 105482 228118 105718
rect 228354 105482 228438 105718
rect 228674 105482 228758 105718
rect 228994 105482 229078 105718
rect 229314 105482 229398 105718
rect 229634 105482 229718 105718
rect 229954 105482 230038 105718
rect 230274 105482 230358 105718
rect 230594 105482 230716 105718
rect 209779 96716 209780 96766
rect 209844 96716 209845 96766
rect 209779 96715 209845 96716
rect 159464 94518 159784 94560
rect 159464 94282 159506 94518
rect 159742 94282 159784 94518
rect 159464 94240 159784 94282
rect 200173 94518 200493 94560
rect 200173 94282 200215 94518
rect 200451 94282 200493 94518
rect 200173 94240 200493 94282
rect 144104 83318 144424 83360
rect 144104 83082 144146 83318
rect 144382 83082 144424 83318
rect 144104 83040 144424 83082
rect 197507 83318 197827 83360
rect 197507 83082 197549 83318
rect 197785 83082 197827 83318
rect 197507 83040 197827 83082
rect 226716 83318 230716 105482
rect 226716 83082 226838 83318
rect 227074 83082 227158 83318
rect 227394 83082 227478 83318
rect 227714 83082 227798 83318
rect 228034 83082 228118 83318
rect 228354 83082 228438 83318
rect 228674 83082 228758 83318
rect 228994 83082 229078 83318
rect 229314 83082 229398 83318
rect 229634 83082 229718 83318
rect 229954 83082 230038 83318
rect 230274 83082 230358 83318
rect 230594 83082 230716 83318
rect 159464 72118 159784 72160
rect 159464 71882 159506 72118
rect 159742 71882 159784 72118
rect 159464 71840 159784 71882
rect 200173 72118 200493 72160
rect 200173 71882 200215 72118
rect 200451 71882 200493 72118
rect 200173 71840 200493 71882
rect 211435 69852 211501 69853
rect 211435 69788 211436 69852
rect 211500 69788 211501 69852
rect 211435 69787 211501 69788
rect 140227 58428 140293 58429
rect 140227 58364 140228 58428
rect 140292 58364 140293 58428
rect 140227 58363 140293 58364
rect 152739 47004 152805 47005
rect 152739 46940 152740 47004
rect 152804 46940 152805 47004
rect 152739 46939 152805 46940
rect 68835 46868 68901 46869
rect 68835 46804 68836 46868
rect 68900 46804 68901 46868
rect 68835 46803 68901 46804
rect 149059 46868 149125 46869
rect 149059 46804 149060 46868
rect 149124 46804 149125 46868
rect 149059 46803 149125 46804
rect 64971 46732 65037 46733
rect 64971 46668 64972 46732
rect 65036 46668 65037 46732
rect 64971 46667 65037 46668
rect 63499 46460 63565 46461
rect 63499 46396 63500 46460
rect 63564 46396 63565 46460
rect 63499 46395 63565 46396
rect 62211 46324 62277 46325
rect 62211 46260 62212 46324
rect 62276 46260 62277 46324
rect 62211 46259 62277 46260
rect 5000 38282 5122 38518
rect 5358 38282 5442 38518
rect 5678 38282 5762 38518
rect 5998 38282 6082 38518
rect 6318 38282 6402 38518
rect 6638 38282 6722 38518
rect 6958 38282 7042 38518
rect 7278 38282 7362 38518
rect 7598 38282 7682 38518
rect 7918 38282 8002 38518
rect 8238 38282 8322 38518
rect 8558 38282 8642 38518
rect 8878 38282 9000 38518
rect 5000 16118 9000 38282
rect 25507 38518 25827 38560
rect 25507 38282 25549 38518
rect 25785 38282 25827 38518
rect 25507 38240 25827 38282
rect 30173 27318 30493 27360
rect 30173 27082 30215 27318
rect 30451 27082 30493 27318
rect 30173 27040 30493 27082
rect 19707 23272 19773 23273
rect 19707 23208 19708 23272
rect 19772 23208 19773 23272
rect 19707 23207 19773 23208
rect 19710 22882 19770 23207
rect 62214 21029 62274 46259
rect 63315 46188 63381 46189
rect 63315 46124 63316 46188
rect 63380 46124 63381 46188
rect 63315 46123 63381 46124
rect 63318 21029 63378 46123
rect 62211 21028 62277 21029
rect 62211 20964 62212 21028
rect 62276 20964 62277 21028
rect 62211 20963 62277 20964
rect 63315 21028 63381 21029
rect 63315 20964 63316 21028
rect 63380 20964 63381 21028
rect 63315 20963 63381 20964
rect 63502 20893 63562 46395
rect 64974 21029 65034 46667
rect 68467 46596 68533 46597
rect 68467 46532 68468 46596
rect 68532 46532 68533 46596
rect 68467 46531 68533 46532
rect 66840 38518 67160 38560
rect 66840 38282 66882 38518
rect 67118 38282 67160 38518
rect 66840 38240 67160 38282
rect 68470 21029 68530 46531
rect 64971 21028 65037 21029
rect 64971 20964 64972 21028
rect 65036 20964 65037 21028
rect 64971 20963 65037 20964
rect 68467 21028 68533 21029
rect 68467 20964 68468 21028
rect 68532 20964 68533 21028
rect 68467 20963 68533 20964
rect 68838 20893 68898 46803
rect 146299 46732 146365 46733
rect 146299 46668 146300 46732
rect 146364 46668 146365 46732
rect 146299 46667 146365 46668
rect 89811 46324 89877 46325
rect 89811 46260 89812 46324
rect 89876 46260 89877 46324
rect 89811 46259 89877 46260
rect 146115 46324 146181 46325
rect 146115 46260 146116 46324
rect 146180 46260 146181 46324
rect 146115 46259 146181 46260
rect 89075 46188 89141 46189
rect 89075 46124 89076 46188
rect 89140 46124 89141 46188
rect 89075 46123 89141 46124
rect 71840 27318 72160 27360
rect 71840 27082 71882 27318
rect 72118 27082 72160 27318
rect 71840 27040 72160 27082
rect 63499 20892 63565 20893
rect 63499 20828 63500 20892
rect 63564 20828 63565 20892
rect 63499 20827 63565 20828
rect 68835 20892 68901 20893
rect 68835 20828 68836 20892
rect 68900 20828 68901 20892
rect 89078 20842 89138 46123
rect 68835 20827 68901 20828
rect 89814 20162 89874 46259
rect 109507 38518 109827 38560
rect 109507 38282 109549 38518
rect 109785 38282 109827 38518
rect 109507 38240 109827 38282
rect 114173 27318 114493 27360
rect 114173 27082 114215 27318
rect 114451 27082 114493 27318
rect 114173 27040 114493 27082
rect 146118 20893 146178 46259
rect 146302 21029 146362 46667
rect 147771 46460 147837 46461
rect 147771 46396 147772 46460
rect 147836 46396 147837 46460
rect 147771 46395 147837 46396
rect 147035 46188 147101 46189
rect 147035 46124 147036 46188
rect 147100 46124 147101 46188
rect 147035 46123 147101 46124
rect 146299 21028 146365 21029
rect 146299 20964 146300 21028
rect 146364 20964 146365 21028
rect 146299 20963 146365 20964
rect 101035 20892 101101 20893
rect 101035 20842 101036 20892
rect 101100 20842 101101 20892
rect 146115 20892 146181 20893
rect 146115 20828 146116 20892
rect 146180 20828 146181 20892
rect 146115 20827 146181 20828
rect 101035 20212 101101 20213
rect 101035 20162 101036 20212
rect 101100 20162 101101 20212
rect 147038 17085 147098 46123
rect 147774 21029 147834 46395
rect 149062 21029 149122 46803
rect 152555 46596 152621 46597
rect 152555 46532 152556 46596
rect 152620 46532 152621 46596
rect 152555 46531 152621 46532
rect 150840 38518 151160 38560
rect 150840 38282 150882 38518
rect 151118 38282 151160 38518
rect 150840 38240 151160 38282
rect 147771 21028 147837 21029
rect 147771 20964 147772 21028
rect 147836 20964 147837 21028
rect 147771 20963 147837 20964
rect 149059 21028 149125 21029
rect 149059 20964 149060 21028
rect 149124 20964 149125 21028
rect 149059 20963 149125 20964
rect 152558 18445 152618 46531
rect 152742 20757 152802 46939
rect 172979 46188 173045 46189
rect 172979 46124 172980 46188
rect 173044 46124 173045 46188
rect 172979 46123 173045 46124
rect 155840 27318 156160 27360
rect 155840 27082 155882 27318
rect 156118 27082 156160 27318
rect 155840 27040 156160 27082
rect 172982 20842 173042 46123
rect 211438 45322 211498 69787
rect 211619 63188 211685 63189
rect 211619 63124 211620 63188
rect 211684 63124 211685 63188
rect 211619 63123 211685 63124
rect 211622 49994 211682 63123
rect 226716 60918 230716 83082
rect 226716 60682 226838 60918
rect 227074 60682 227158 60918
rect 227394 60682 227478 60918
rect 227714 60682 227798 60918
rect 228034 60682 228118 60918
rect 228354 60682 228438 60918
rect 228674 60682 228758 60918
rect 228994 60682 229078 60918
rect 229314 60682 229398 60918
rect 229634 60682 229718 60918
rect 229954 60682 230038 60918
rect 230274 60682 230358 60918
rect 230594 60682 230716 60918
rect 211622 49934 212602 49994
rect 212542 45234 212602 49934
rect 212542 45174 213338 45234
rect 173347 44828 173413 44829
rect 173347 44764 173348 44828
rect 173412 44764 173413 44828
rect 173347 44763 173413 44764
rect 152739 20756 152805 20757
rect 152739 20692 152740 20756
rect 152804 20692 152805 20756
rect 152739 20691 152805 20692
rect 173350 20162 173410 44763
rect 173899 44692 173965 44693
rect 173899 44628 173900 44692
rect 173964 44628 173965 44692
rect 173899 44627 173965 44628
rect 173902 22202 173962 44627
rect 193507 38518 193827 38560
rect 193507 38282 193549 38518
rect 193785 38282 193827 38518
rect 193507 38240 193827 38282
rect 213278 37754 213338 45174
rect 213278 37694 213522 37754
rect 213462 35034 213522 37694
rect 213830 37074 213890 45086
rect 226716 38518 230716 60682
rect 226716 38282 226838 38518
rect 227074 38282 227158 38518
rect 227394 38282 227478 38518
rect 227714 38282 227798 38518
rect 228034 38282 228118 38518
rect 228354 38282 228438 38518
rect 228674 38282 228758 38518
rect 228994 38282 229078 38518
rect 229314 38282 229398 38518
rect 229634 38282 229718 38518
rect 229954 38282 230038 38518
rect 230274 38282 230358 38518
rect 230594 38282 230716 38518
rect 213830 37014 214258 37074
rect 214198 35714 214258 37014
rect 213830 35654 214258 35714
rect 213830 35122 213890 35654
rect 213278 34974 213522 35034
rect 212726 27554 212786 34886
rect 213278 30274 213338 34974
rect 213278 30214 213522 30274
rect 212726 27494 213338 27554
rect 198173 27318 198493 27360
rect 198173 27082 198215 27318
rect 198451 27082 198493 27318
rect 198173 27040 198493 27082
rect 213278 24154 213338 27494
rect 212726 24094 213338 24154
rect 185123 21916 185124 21966
rect 185188 21916 185189 21966
rect 185123 21915 185189 21916
rect 185491 20892 185557 20893
rect 185491 20828 185492 20892
rect 185556 20828 185557 20892
rect 185491 20827 185557 20828
rect 185494 20162 185554 20827
rect 212726 20074 212786 24094
rect 212542 20014 212786 20074
rect 152555 18444 152621 18445
rect 152555 18380 152556 18444
rect 152620 18380 152621 18444
rect 152555 18379 152621 18380
rect 212542 17085 212602 20014
rect 213462 18445 213522 30214
rect 213459 18444 213525 18445
rect 213459 18380 213460 18444
rect 213524 18380 213525 18444
rect 213459 18379 213525 18380
rect 147035 17084 147101 17085
rect 147035 17020 147036 17084
rect 147100 17020 147101 17084
rect 147035 17019 147101 17020
rect 212539 17084 212605 17085
rect 212539 17020 212540 17084
rect 212604 17020 212605 17084
rect 212539 17019 212605 17020
rect 5000 15882 5122 16118
rect 5358 15882 5442 16118
rect 5678 15882 5762 16118
rect 5998 15882 6082 16118
rect 6318 15882 6402 16118
rect 6638 15882 6722 16118
rect 6958 15882 7042 16118
rect 7278 15882 7362 16118
rect 7598 15882 7682 16118
rect 7918 15882 8002 16118
rect 8238 15882 8322 16118
rect 8558 15882 8642 16118
rect 8878 15882 9000 16118
rect 5000 8878 9000 15882
rect 5000 8642 5122 8878
rect 5358 8642 5442 8878
rect 5678 8642 5762 8878
rect 5998 8642 6082 8878
rect 6318 8642 6402 8878
rect 6638 8642 6722 8878
rect 6958 8642 7042 8878
rect 7278 8642 7362 8878
rect 7598 8642 7682 8878
rect 7918 8642 8002 8878
rect 8238 8642 8322 8878
rect 8558 8642 8642 8878
rect 8878 8642 9000 8878
rect 5000 8558 9000 8642
rect 5000 8322 5122 8558
rect 5358 8322 5442 8558
rect 5678 8322 5762 8558
rect 5998 8322 6082 8558
rect 6318 8322 6402 8558
rect 6638 8322 6722 8558
rect 6958 8322 7042 8558
rect 7278 8322 7362 8558
rect 7598 8322 7682 8558
rect 7918 8322 8002 8558
rect 8238 8322 8322 8558
rect 8558 8322 8642 8558
rect 8878 8322 9000 8558
rect 5000 8238 9000 8322
rect 5000 8002 5122 8238
rect 5358 8002 5442 8238
rect 5678 8002 5762 8238
rect 5998 8002 6082 8238
rect 6318 8002 6402 8238
rect 6638 8002 6722 8238
rect 6958 8002 7042 8238
rect 7278 8002 7362 8238
rect 7598 8002 7682 8238
rect 7918 8002 8002 8238
rect 8238 8002 8322 8238
rect 8558 8002 8642 8238
rect 8878 8002 9000 8238
rect 5000 7918 9000 8002
rect 5000 7682 5122 7918
rect 5358 7682 5442 7918
rect 5678 7682 5762 7918
rect 5998 7682 6082 7918
rect 6318 7682 6402 7918
rect 6638 7682 6722 7918
rect 6958 7682 7042 7918
rect 7278 7682 7362 7918
rect 7598 7682 7682 7918
rect 7918 7682 8002 7918
rect 8238 7682 8322 7918
rect 8558 7682 8642 7918
rect 8878 7682 9000 7918
rect 5000 7598 9000 7682
rect 5000 7362 5122 7598
rect 5358 7362 5442 7598
rect 5678 7362 5762 7598
rect 5998 7362 6082 7598
rect 6318 7362 6402 7598
rect 6638 7362 6722 7598
rect 6958 7362 7042 7598
rect 7278 7362 7362 7598
rect 7598 7362 7682 7598
rect 7918 7362 8002 7598
rect 8238 7362 8322 7598
rect 8558 7362 8642 7598
rect 8878 7362 9000 7598
rect 5000 7278 9000 7362
rect 5000 7042 5122 7278
rect 5358 7042 5442 7278
rect 5678 7042 5762 7278
rect 5998 7042 6082 7278
rect 6318 7042 6402 7278
rect 6638 7042 6722 7278
rect 6958 7042 7042 7278
rect 7278 7042 7362 7278
rect 7598 7042 7682 7278
rect 7918 7042 8002 7278
rect 8238 7042 8322 7278
rect 8558 7042 8642 7278
rect 8878 7042 9000 7278
rect 5000 6958 9000 7042
rect 5000 6722 5122 6958
rect 5358 6722 5442 6958
rect 5678 6722 5762 6958
rect 5998 6722 6082 6958
rect 6318 6722 6402 6958
rect 6638 6722 6722 6958
rect 6958 6722 7042 6958
rect 7278 6722 7362 6958
rect 7598 6722 7682 6958
rect 7918 6722 8002 6958
rect 8238 6722 8322 6958
rect 8558 6722 8642 6958
rect 8878 6722 9000 6958
rect 5000 6638 9000 6722
rect 5000 6402 5122 6638
rect 5358 6402 5442 6638
rect 5678 6402 5762 6638
rect 5998 6402 6082 6638
rect 6318 6402 6402 6638
rect 6638 6402 6722 6638
rect 6958 6402 7042 6638
rect 7278 6402 7362 6638
rect 7598 6402 7682 6638
rect 7918 6402 8002 6638
rect 8238 6402 8322 6638
rect 8558 6402 8642 6638
rect 8878 6402 9000 6638
rect 5000 6318 9000 6402
rect 5000 6082 5122 6318
rect 5358 6082 5442 6318
rect 5678 6082 5762 6318
rect 5998 6082 6082 6318
rect 6318 6082 6402 6318
rect 6638 6082 6722 6318
rect 6958 6082 7042 6318
rect 7278 6082 7362 6318
rect 7598 6082 7682 6318
rect 7918 6082 8002 6318
rect 8238 6082 8322 6318
rect 8558 6082 8642 6318
rect 8878 6082 9000 6318
rect 5000 5998 9000 6082
rect 5000 5762 5122 5998
rect 5358 5762 5442 5998
rect 5678 5762 5762 5998
rect 5998 5762 6082 5998
rect 6318 5762 6402 5998
rect 6638 5762 6722 5998
rect 6958 5762 7042 5998
rect 7278 5762 7362 5998
rect 7598 5762 7682 5998
rect 7918 5762 8002 5998
rect 8238 5762 8322 5998
rect 8558 5762 8642 5998
rect 8878 5762 9000 5998
rect 5000 5678 9000 5762
rect 5000 5442 5122 5678
rect 5358 5442 5442 5678
rect 5678 5442 5762 5678
rect 5998 5442 6082 5678
rect 6318 5442 6402 5678
rect 6638 5442 6722 5678
rect 6958 5442 7042 5678
rect 7278 5442 7362 5678
rect 7598 5442 7682 5678
rect 7918 5442 8002 5678
rect 8238 5442 8322 5678
rect 8558 5442 8642 5678
rect 8878 5442 9000 5678
rect 5000 5358 9000 5442
rect 5000 5122 5122 5358
rect 5358 5122 5442 5358
rect 5678 5122 5762 5358
rect 5998 5122 6082 5358
rect 6318 5122 6402 5358
rect 6638 5122 6722 5358
rect 6958 5122 7042 5358
rect 7278 5122 7362 5358
rect 7598 5122 7682 5358
rect 7918 5122 8002 5358
rect 8238 5122 8322 5358
rect 8558 5122 8642 5358
rect 8878 5122 9000 5358
rect 5000 5000 9000 5122
rect 226716 16118 230716 38282
rect 226716 15882 226838 16118
rect 227074 15882 227158 16118
rect 227394 15882 227478 16118
rect 227714 15882 227798 16118
rect 228034 15882 228118 16118
rect 228354 15882 228438 16118
rect 228674 15882 228758 16118
rect 228994 15882 229078 16118
rect 229314 15882 229398 16118
rect 229634 15882 229718 16118
rect 229954 15882 230038 16118
rect 230274 15882 230358 16118
rect 230594 15882 230716 16118
rect 226716 8878 230716 15882
rect 226716 8642 226838 8878
rect 227074 8642 227158 8878
rect 227394 8642 227478 8878
rect 227714 8642 227798 8878
rect 228034 8642 228118 8878
rect 228354 8642 228438 8878
rect 228674 8642 228758 8878
rect 228994 8642 229078 8878
rect 229314 8642 229398 8878
rect 229634 8642 229718 8878
rect 229954 8642 230038 8878
rect 230274 8642 230358 8878
rect 230594 8642 230716 8878
rect 226716 8558 230716 8642
rect 226716 8322 226838 8558
rect 227074 8322 227158 8558
rect 227394 8322 227478 8558
rect 227714 8322 227798 8558
rect 228034 8322 228118 8558
rect 228354 8322 228438 8558
rect 228674 8322 228758 8558
rect 228994 8322 229078 8558
rect 229314 8322 229398 8558
rect 229634 8322 229718 8558
rect 229954 8322 230038 8558
rect 230274 8322 230358 8558
rect 230594 8322 230716 8558
rect 226716 8238 230716 8322
rect 226716 8002 226838 8238
rect 227074 8002 227158 8238
rect 227394 8002 227478 8238
rect 227714 8002 227798 8238
rect 228034 8002 228118 8238
rect 228354 8002 228438 8238
rect 228674 8002 228758 8238
rect 228994 8002 229078 8238
rect 229314 8002 229398 8238
rect 229634 8002 229718 8238
rect 229954 8002 230038 8238
rect 230274 8002 230358 8238
rect 230594 8002 230716 8238
rect 226716 7918 230716 8002
rect 226716 7682 226838 7918
rect 227074 7682 227158 7918
rect 227394 7682 227478 7918
rect 227714 7682 227798 7918
rect 228034 7682 228118 7918
rect 228354 7682 228438 7918
rect 228674 7682 228758 7918
rect 228994 7682 229078 7918
rect 229314 7682 229398 7918
rect 229634 7682 229718 7918
rect 229954 7682 230038 7918
rect 230274 7682 230358 7918
rect 230594 7682 230716 7918
rect 226716 7598 230716 7682
rect 226716 7362 226838 7598
rect 227074 7362 227158 7598
rect 227394 7362 227478 7598
rect 227714 7362 227798 7598
rect 228034 7362 228118 7598
rect 228354 7362 228438 7598
rect 228674 7362 228758 7598
rect 228994 7362 229078 7598
rect 229314 7362 229398 7598
rect 229634 7362 229718 7598
rect 229954 7362 230038 7598
rect 230274 7362 230358 7598
rect 230594 7362 230716 7598
rect 226716 7278 230716 7362
rect 226716 7042 226838 7278
rect 227074 7042 227158 7278
rect 227394 7042 227478 7278
rect 227714 7042 227798 7278
rect 228034 7042 228118 7278
rect 228354 7042 228438 7278
rect 228674 7042 228758 7278
rect 228994 7042 229078 7278
rect 229314 7042 229398 7278
rect 229634 7042 229718 7278
rect 229954 7042 230038 7278
rect 230274 7042 230358 7278
rect 230594 7042 230716 7278
rect 226716 6958 230716 7042
rect 226716 6722 226838 6958
rect 227074 6722 227158 6958
rect 227394 6722 227478 6958
rect 227714 6722 227798 6958
rect 228034 6722 228118 6958
rect 228354 6722 228438 6958
rect 228674 6722 228758 6958
rect 228994 6722 229078 6958
rect 229314 6722 229398 6958
rect 229634 6722 229718 6958
rect 229954 6722 230038 6958
rect 230274 6722 230358 6958
rect 230594 6722 230716 6958
rect 226716 6638 230716 6722
rect 226716 6402 226838 6638
rect 227074 6402 227158 6638
rect 227394 6402 227478 6638
rect 227714 6402 227798 6638
rect 228034 6402 228118 6638
rect 228354 6402 228438 6638
rect 228674 6402 228758 6638
rect 228994 6402 229078 6638
rect 229314 6402 229398 6638
rect 229634 6402 229718 6638
rect 229954 6402 230038 6638
rect 230274 6402 230358 6638
rect 230594 6402 230716 6638
rect 226716 6318 230716 6402
rect 226716 6082 226838 6318
rect 227074 6082 227158 6318
rect 227394 6082 227478 6318
rect 227714 6082 227798 6318
rect 228034 6082 228118 6318
rect 228354 6082 228438 6318
rect 228674 6082 228758 6318
rect 228994 6082 229078 6318
rect 229314 6082 229398 6318
rect 229634 6082 229718 6318
rect 229954 6082 230038 6318
rect 230274 6082 230358 6318
rect 230594 6082 230716 6318
rect 226716 5998 230716 6082
rect 226716 5762 226838 5998
rect 227074 5762 227158 5998
rect 227394 5762 227478 5998
rect 227714 5762 227798 5998
rect 228034 5762 228118 5998
rect 228354 5762 228438 5998
rect 228674 5762 228758 5998
rect 228994 5762 229078 5998
rect 229314 5762 229398 5998
rect 229634 5762 229718 5998
rect 229954 5762 230038 5998
rect 230274 5762 230358 5998
rect 230594 5762 230716 5998
rect 226716 5678 230716 5762
rect 226716 5442 226838 5678
rect 227074 5442 227158 5678
rect 227394 5442 227478 5678
rect 227714 5442 227798 5678
rect 228034 5442 228118 5678
rect 228354 5442 228438 5678
rect 228674 5442 228758 5678
rect 228994 5442 229078 5678
rect 229314 5442 229398 5678
rect 229634 5442 229718 5678
rect 229954 5442 230038 5678
rect 230274 5442 230358 5678
rect 230594 5442 230716 5678
rect 226716 5358 230716 5442
rect 226716 5122 226838 5358
rect 227074 5122 227158 5358
rect 227394 5122 227478 5358
rect 227714 5122 227798 5358
rect 228034 5122 228118 5358
rect 228354 5122 228438 5358
rect 228674 5122 228758 5358
rect 228994 5122 229078 5358
rect 229314 5122 229398 5358
rect 229634 5122 229718 5358
rect 229954 5122 230038 5358
rect 230274 5122 230358 5358
rect 230594 5122 230716 5358
rect 226716 5000 230716 5122
rect 231716 228918 235716 249322
rect 231716 228682 231838 228918
rect 232074 228682 232158 228918
rect 232394 228682 232478 228918
rect 232714 228682 232798 228918
rect 233034 228682 233118 228918
rect 233354 228682 233438 228918
rect 233674 228682 233758 228918
rect 233994 228682 234078 228918
rect 234314 228682 234398 228918
rect 234634 228682 234718 228918
rect 234954 228682 235038 228918
rect 235274 228682 235358 228918
rect 235594 228682 235716 228918
rect 231716 206518 235716 228682
rect 231716 206282 231838 206518
rect 232074 206282 232158 206518
rect 232394 206282 232478 206518
rect 232714 206282 232798 206518
rect 233034 206282 233118 206518
rect 233354 206282 233438 206518
rect 233674 206282 233758 206518
rect 233994 206282 234078 206518
rect 234314 206282 234398 206518
rect 234634 206282 234718 206518
rect 234954 206282 235038 206518
rect 235274 206282 235358 206518
rect 235594 206282 235716 206518
rect 231716 184118 235716 206282
rect 231716 183882 231838 184118
rect 232074 183882 232158 184118
rect 232394 183882 232478 184118
rect 232714 183882 232798 184118
rect 233034 183882 233118 184118
rect 233354 183882 233438 184118
rect 233674 183882 233758 184118
rect 233994 183882 234078 184118
rect 234314 183882 234398 184118
rect 234634 183882 234718 184118
rect 234954 183882 235038 184118
rect 235274 183882 235358 184118
rect 235594 183882 235716 184118
rect 231716 161718 235716 183882
rect 231716 161482 231838 161718
rect 232074 161482 232158 161718
rect 232394 161482 232478 161718
rect 232714 161482 232798 161718
rect 233034 161482 233118 161718
rect 233354 161482 233438 161718
rect 233674 161482 233758 161718
rect 233994 161482 234078 161718
rect 234314 161482 234398 161718
rect 234634 161482 234718 161718
rect 234954 161482 235038 161718
rect 235274 161482 235358 161718
rect 235594 161482 235716 161718
rect 231716 139318 235716 161482
rect 231716 139082 231838 139318
rect 232074 139082 232158 139318
rect 232394 139082 232478 139318
rect 232714 139082 232798 139318
rect 233034 139082 233118 139318
rect 233354 139082 233438 139318
rect 233674 139082 233758 139318
rect 233994 139082 234078 139318
rect 234314 139082 234398 139318
rect 234634 139082 234718 139318
rect 234954 139082 235038 139318
rect 235274 139082 235358 139318
rect 235594 139082 235716 139318
rect 231716 116918 235716 139082
rect 231716 116682 231838 116918
rect 232074 116682 232158 116918
rect 232394 116682 232478 116918
rect 232714 116682 232798 116918
rect 233034 116682 233118 116918
rect 233354 116682 233438 116918
rect 233674 116682 233758 116918
rect 233994 116682 234078 116918
rect 234314 116682 234398 116918
rect 234634 116682 234718 116918
rect 234954 116682 235038 116918
rect 235274 116682 235358 116918
rect 235594 116682 235716 116918
rect 231716 94518 235716 116682
rect 231716 94282 231838 94518
rect 232074 94282 232158 94518
rect 232394 94282 232478 94518
rect 232714 94282 232798 94518
rect 233034 94282 233118 94518
rect 233354 94282 233438 94518
rect 233674 94282 233758 94518
rect 233994 94282 234078 94518
rect 234314 94282 234398 94518
rect 234634 94282 234718 94518
rect 234954 94282 235038 94518
rect 235274 94282 235358 94518
rect 235594 94282 235716 94518
rect 231716 72118 235716 94282
rect 231716 71882 231838 72118
rect 232074 71882 232158 72118
rect 232394 71882 232478 72118
rect 232714 71882 232798 72118
rect 233034 71882 233118 72118
rect 233354 71882 233438 72118
rect 233674 71882 233758 72118
rect 233994 71882 234078 72118
rect 234314 71882 234398 72118
rect 234634 71882 234718 72118
rect 234954 71882 235038 72118
rect 235274 71882 235358 72118
rect 235594 71882 235716 72118
rect 231716 49718 235716 71882
rect 231716 49482 231838 49718
rect 232074 49482 232158 49718
rect 232394 49482 232478 49718
rect 232714 49482 232798 49718
rect 233034 49482 233118 49718
rect 233354 49482 233438 49718
rect 233674 49482 233758 49718
rect 233994 49482 234078 49718
rect 234314 49482 234398 49718
rect 234634 49482 234718 49718
rect 234954 49482 235038 49718
rect 235274 49482 235358 49718
rect 235594 49482 235716 49718
rect 231716 27318 235716 49482
rect 231716 27082 231838 27318
rect 232074 27082 232158 27318
rect 232394 27082 232478 27318
rect 232714 27082 232798 27318
rect 233034 27082 233118 27318
rect 233354 27082 233438 27318
rect 233674 27082 233758 27318
rect 233994 27082 234078 27318
rect 234314 27082 234398 27318
rect 234634 27082 234718 27318
rect 234954 27082 235038 27318
rect 235274 27082 235358 27318
rect 235594 27082 235716 27318
rect 0 3642 122 3878
rect 358 3642 442 3878
rect 678 3642 762 3878
rect 998 3642 1082 3878
rect 1318 3642 1402 3878
rect 1638 3642 1722 3878
rect 1958 3642 2042 3878
rect 2278 3642 2362 3878
rect 2598 3642 2682 3878
rect 2918 3642 3002 3878
rect 3238 3642 3322 3878
rect 3558 3642 3642 3878
rect 3878 3642 4000 3878
rect 0 3558 4000 3642
rect 0 3322 122 3558
rect 358 3322 442 3558
rect 678 3322 762 3558
rect 998 3322 1082 3558
rect 1318 3322 1402 3558
rect 1638 3322 1722 3558
rect 1958 3322 2042 3558
rect 2278 3322 2362 3558
rect 2598 3322 2682 3558
rect 2918 3322 3002 3558
rect 3238 3322 3322 3558
rect 3558 3322 3642 3558
rect 3878 3322 4000 3558
rect 0 3238 4000 3322
rect 0 3002 122 3238
rect 358 3002 442 3238
rect 678 3002 762 3238
rect 998 3002 1082 3238
rect 1318 3002 1402 3238
rect 1638 3002 1722 3238
rect 1958 3002 2042 3238
rect 2278 3002 2362 3238
rect 2598 3002 2682 3238
rect 2918 3002 3002 3238
rect 3238 3002 3322 3238
rect 3558 3002 3642 3238
rect 3878 3002 4000 3238
rect 0 2918 4000 3002
rect 0 2682 122 2918
rect 358 2682 442 2918
rect 678 2682 762 2918
rect 998 2682 1082 2918
rect 1318 2682 1402 2918
rect 1638 2682 1722 2918
rect 1958 2682 2042 2918
rect 2278 2682 2362 2918
rect 2598 2682 2682 2918
rect 2918 2682 3002 2918
rect 3238 2682 3322 2918
rect 3558 2682 3642 2918
rect 3878 2682 4000 2918
rect 0 2598 4000 2682
rect 0 2362 122 2598
rect 358 2362 442 2598
rect 678 2362 762 2598
rect 998 2362 1082 2598
rect 1318 2362 1402 2598
rect 1638 2362 1722 2598
rect 1958 2362 2042 2598
rect 2278 2362 2362 2598
rect 2598 2362 2682 2598
rect 2918 2362 3002 2598
rect 3238 2362 3322 2598
rect 3558 2362 3642 2598
rect 3878 2362 4000 2598
rect 0 2278 4000 2362
rect 0 2042 122 2278
rect 358 2042 442 2278
rect 678 2042 762 2278
rect 998 2042 1082 2278
rect 1318 2042 1402 2278
rect 1638 2042 1722 2278
rect 1958 2042 2042 2278
rect 2278 2042 2362 2278
rect 2598 2042 2682 2278
rect 2918 2042 3002 2278
rect 3238 2042 3322 2278
rect 3558 2042 3642 2278
rect 3878 2042 4000 2278
rect 0 1958 4000 2042
rect 0 1722 122 1958
rect 358 1722 442 1958
rect 678 1722 762 1958
rect 998 1722 1082 1958
rect 1318 1722 1402 1958
rect 1638 1722 1722 1958
rect 1958 1722 2042 1958
rect 2278 1722 2362 1958
rect 2598 1722 2682 1958
rect 2918 1722 3002 1958
rect 3238 1722 3322 1958
rect 3558 1722 3642 1958
rect 3878 1722 4000 1958
rect 0 1638 4000 1722
rect 0 1402 122 1638
rect 358 1402 442 1638
rect 678 1402 762 1638
rect 998 1402 1082 1638
rect 1318 1402 1402 1638
rect 1638 1402 1722 1638
rect 1958 1402 2042 1638
rect 2278 1402 2362 1638
rect 2598 1402 2682 1638
rect 2918 1402 3002 1638
rect 3238 1402 3322 1638
rect 3558 1402 3642 1638
rect 3878 1402 4000 1638
rect 0 1318 4000 1402
rect 0 1082 122 1318
rect 358 1082 442 1318
rect 678 1082 762 1318
rect 998 1082 1082 1318
rect 1318 1082 1402 1318
rect 1638 1082 1722 1318
rect 1958 1082 2042 1318
rect 2278 1082 2362 1318
rect 2598 1082 2682 1318
rect 2918 1082 3002 1318
rect 3238 1082 3322 1318
rect 3558 1082 3642 1318
rect 3878 1082 4000 1318
rect 0 998 4000 1082
rect 0 762 122 998
rect 358 762 442 998
rect 678 762 762 998
rect 998 762 1082 998
rect 1318 762 1402 998
rect 1638 762 1722 998
rect 1958 762 2042 998
rect 2278 762 2362 998
rect 2598 762 2682 998
rect 2918 762 3002 998
rect 3238 762 3322 998
rect 3558 762 3642 998
rect 3878 762 4000 998
rect 0 678 4000 762
rect 0 442 122 678
rect 358 442 442 678
rect 678 442 762 678
rect 998 442 1082 678
rect 1318 442 1402 678
rect 1638 442 1722 678
rect 1958 442 2042 678
rect 2278 442 2362 678
rect 2598 442 2682 678
rect 2918 442 3002 678
rect 3238 442 3322 678
rect 3558 442 3642 678
rect 3878 442 4000 678
rect 0 358 4000 442
rect 0 122 122 358
rect 358 122 442 358
rect 678 122 762 358
rect 998 122 1082 358
rect 1318 122 1402 358
rect 1638 122 1722 358
rect 1958 122 2042 358
rect 2278 122 2362 358
rect 2598 122 2682 358
rect 2918 122 3002 358
rect 3238 122 3322 358
rect 3558 122 3642 358
rect 3878 122 4000 358
rect 0 0 4000 122
rect 231716 3878 235716 27082
rect 231716 3642 231838 3878
rect 232074 3642 232158 3878
rect 232394 3642 232478 3878
rect 232714 3642 232798 3878
rect 233034 3642 233118 3878
rect 233354 3642 233438 3878
rect 233674 3642 233758 3878
rect 233994 3642 234078 3878
rect 234314 3642 234398 3878
rect 234634 3642 234718 3878
rect 234954 3642 235038 3878
rect 235274 3642 235358 3878
rect 235594 3642 235716 3878
rect 231716 3558 235716 3642
rect 231716 3322 231838 3558
rect 232074 3322 232158 3558
rect 232394 3322 232478 3558
rect 232714 3322 232798 3558
rect 233034 3322 233118 3558
rect 233354 3322 233438 3558
rect 233674 3322 233758 3558
rect 233994 3322 234078 3558
rect 234314 3322 234398 3558
rect 234634 3322 234718 3558
rect 234954 3322 235038 3558
rect 235274 3322 235358 3558
rect 235594 3322 235716 3558
rect 231716 3238 235716 3322
rect 231716 3002 231838 3238
rect 232074 3002 232158 3238
rect 232394 3002 232478 3238
rect 232714 3002 232798 3238
rect 233034 3002 233118 3238
rect 233354 3002 233438 3238
rect 233674 3002 233758 3238
rect 233994 3002 234078 3238
rect 234314 3002 234398 3238
rect 234634 3002 234718 3238
rect 234954 3002 235038 3238
rect 235274 3002 235358 3238
rect 235594 3002 235716 3238
rect 231716 2918 235716 3002
rect 231716 2682 231838 2918
rect 232074 2682 232158 2918
rect 232394 2682 232478 2918
rect 232714 2682 232798 2918
rect 233034 2682 233118 2918
rect 233354 2682 233438 2918
rect 233674 2682 233758 2918
rect 233994 2682 234078 2918
rect 234314 2682 234398 2918
rect 234634 2682 234718 2918
rect 234954 2682 235038 2918
rect 235274 2682 235358 2918
rect 235594 2682 235716 2918
rect 231716 2598 235716 2682
rect 231716 2362 231838 2598
rect 232074 2362 232158 2598
rect 232394 2362 232478 2598
rect 232714 2362 232798 2598
rect 233034 2362 233118 2598
rect 233354 2362 233438 2598
rect 233674 2362 233758 2598
rect 233994 2362 234078 2598
rect 234314 2362 234398 2598
rect 234634 2362 234718 2598
rect 234954 2362 235038 2598
rect 235274 2362 235358 2598
rect 235594 2362 235716 2598
rect 231716 2278 235716 2362
rect 231716 2042 231838 2278
rect 232074 2042 232158 2278
rect 232394 2042 232478 2278
rect 232714 2042 232798 2278
rect 233034 2042 233118 2278
rect 233354 2042 233438 2278
rect 233674 2042 233758 2278
rect 233994 2042 234078 2278
rect 234314 2042 234398 2278
rect 234634 2042 234718 2278
rect 234954 2042 235038 2278
rect 235274 2042 235358 2278
rect 235594 2042 235716 2278
rect 231716 1958 235716 2042
rect 231716 1722 231838 1958
rect 232074 1722 232158 1958
rect 232394 1722 232478 1958
rect 232714 1722 232798 1958
rect 233034 1722 233118 1958
rect 233354 1722 233438 1958
rect 233674 1722 233758 1958
rect 233994 1722 234078 1958
rect 234314 1722 234398 1958
rect 234634 1722 234718 1958
rect 234954 1722 235038 1958
rect 235274 1722 235358 1958
rect 235594 1722 235716 1958
rect 231716 1638 235716 1722
rect 231716 1402 231838 1638
rect 232074 1402 232158 1638
rect 232394 1402 232478 1638
rect 232714 1402 232798 1638
rect 233034 1402 233118 1638
rect 233354 1402 233438 1638
rect 233674 1402 233758 1638
rect 233994 1402 234078 1638
rect 234314 1402 234398 1638
rect 234634 1402 234718 1638
rect 234954 1402 235038 1638
rect 235274 1402 235358 1638
rect 235594 1402 235716 1638
rect 231716 1318 235716 1402
rect 231716 1082 231838 1318
rect 232074 1082 232158 1318
rect 232394 1082 232478 1318
rect 232714 1082 232798 1318
rect 233034 1082 233118 1318
rect 233354 1082 233438 1318
rect 233674 1082 233758 1318
rect 233994 1082 234078 1318
rect 234314 1082 234398 1318
rect 234634 1082 234718 1318
rect 234954 1082 235038 1318
rect 235274 1082 235358 1318
rect 235594 1082 235716 1318
rect 231716 998 235716 1082
rect 231716 762 231838 998
rect 232074 762 232158 998
rect 232394 762 232478 998
rect 232714 762 232798 998
rect 233034 762 233118 998
rect 233354 762 233438 998
rect 233674 762 233758 998
rect 233994 762 234078 998
rect 234314 762 234398 998
rect 234634 762 234718 998
rect 234954 762 235038 998
rect 235274 762 235358 998
rect 235594 762 235716 998
rect 231716 678 235716 762
rect 231716 442 231838 678
rect 232074 442 232158 678
rect 232394 442 232478 678
rect 232714 442 232798 678
rect 233034 442 233118 678
rect 233354 442 233438 678
rect 233674 442 233758 678
rect 233994 442 234078 678
rect 234314 442 234398 678
rect 234634 442 234718 678
rect 234954 442 235038 678
rect 235274 442 235358 678
rect 235594 442 235716 678
rect 231716 358 235716 442
rect 231716 122 231838 358
rect 232074 122 232158 358
rect 232394 122 232478 358
rect 232714 122 232798 358
rect 233034 122 233118 358
rect 233354 122 233438 358
rect 233674 122 233758 358
rect 233994 122 234078 358
rect 234314 122 234398 358
rect 234634 122 234718 358
rect 234954 122 235038 358
rect 235274 122 235358 358
rect 235594 122 235716 358
rect 231716 0 235716 122
<< via4 >>
rect 122 252842 358 253078
rect 442 252842 678 253078
rect 762 252842 998 253078
rect 1082 252842 1318 253078
rect 1402 252842 1638 253078
rect 1722 252842 1958 253078
rect 2042 252842 2278 253078
rect 2362 252842 2598 253078
rect 2682 252842 2918 253078
rect 3002 252842 3238 253078
rect 3322 252842 3558 253078
rect 3642 252842 3878 253078
rect 122 252522 358 252758
rect 442 252522 678 252758
rect 762 252522 998 252758
rect 1082 252522 1318 252758
rect 1402 252522 1638 252758
rect 1722 252522 1958 252758
rect 2042 252522 2278 252758
rect 2362 252522 2598 252758
rect 2682 252522 2918 252758
rect 3002 252522 3238 252758
rect 3322 252522 3558 252758
rect 3642 252522 3878 252758
rect 122 252202 358 252438
rect 442 252202 678 252438
rect 762 252202 998 252438
rect 1082 252202 1318 252438
rect 1402 252202 1638 252438
rect 1722 252202 1958 252438
rect 2042 252202 2278 252438
rect 2362 252202 2598 252438
rect 2682 252202 2918 252438
rect 3002 252202 3238 252438
rect 3322 252202 3558 252438
rect 3642 252202 3878 252438
rect 122 251882 358 252118
rect 442 251882 678 252118
rect 762 251882 998 252118
rect 1082 251882 1318 252118
rect 1402 251882 1638 252118
rect 1722 251882 1958 252118
rect 2042 251882 2278 252118
rect 2362 251882 2598 252118
rect 2682 251882 2918 252118
rect 3002 251882 3238 252118
rect 3322 251882 3558 252118
rect 3642 251882 3878 252118
rect 122 251562 358 251798
rect 442 251562 678 251798
rect 762 251562 998 251798
rect 1082 251562 1318 251798
rect 1402 251562 1638 251798
rect 1722 251562 1958 251798
rect 2042 251562 2278 251798
rect 2362 251562 2598 251798
rect 2682 251562 2918 251798
rect 3002 251562 3238 251798
rect 3322 251562 3558 251798
rect 3642 251562 3878 251798
rect 122 251242 358 251478
rect 442 251242 678 251478
rect 762 251242 998 251478
rect 1082 251242 1318 251478
rect 1402 251242 1638 251478
rect 1722 251242 1958 251478
rect 2042 251242 2278 251478
rect 2362 251242 2598 251478
rect 2682 251242 2918 251478
rect 3002 251242 3238 251478
rect 3322 251242 3558 251478
rect 3642 251242 3878 251478
rect 122 250922 358 251158
rect 442 250922 678 251158
rect 762 250922 998 251158
rect 1082 250922 1318 251158
rect 1402 250922 1638 251158
rect 1722 250922 1958 251158
rect 2042 250922 2278 251158
rect 2362 250922 2598 251158
rect 2682 250922 2918 251158
rect 3002 250922 3238 251158
rect 3322 250922 3558 251158
rect 3642 250922 3878 251158
rect 122 250602 358 250838
rect 442 250602 678 250838
rect 762 250602 998 250838
rect 1082 250602 1318 250838
rect 1402 250602 1638 250838
rect 1722 250602 1958 250838
rect 2042 250602 2278 250838
rect 2362 250602 2598 250838
rect 2682 250602 2918 250838
rect 3002 250602 3238 250838
rect 3322 250602 3558 250838
rect 3642 250602 3878 250838
rect 122 250282 358 250518
rect 442 250282 678 250518
rect 762 250282 998 250518
rect 1082 250282 1318 250518
rect 1402 250282 1638 250518
rect 1722 250282 1958 250518
rect 2042 250282 2278 250518
rect 2362 250282 2598 250518
rect 2682 250282 2918 250518
rect 3002 250282 3238 250518
rect 3322 250282 3558 250518
rect 3642 250282 3878 250518
rect 122 249962 358 250198
rect 442 249962 678 250198
rect 762 249962 998 250198
rect 1082 249962 1318 250198
rect 1402 249962 1638 250198
rect 1722 249962 1958 250198
rect 2042 249962 2278 250198
rect 2362 249962 2598 250198
rect 2682 249962 2918 250198
rect 3002 249962 3238 250198
rect 3322 249962 3558 250198
rect 3642 249962 3878 250198
rect 122 249642 358 249878
rect 442 249642 678 249878
rect 762 249642 998 249878
rect 1082 249642 1318 249878
rect 1402 249642 1638 249878
rect 1722 249642 1958 249878
rect 2042 249642 2278 249878
rect 2362 249642 2598 249878
rect 2682 249642 2918 249878
rect 3002 249642 3238 249878
rect 3322 249642 3558 249878
rect 3642 249642 3878 249878
rect 122 249322 358 249558
rect 442 249322 678 249558
rect 762 249322 998 249558
rect 1082 249322 1318 249558
rect 1402 249322 1638 249558
rect 1722 249322 1958 249558
rect 2042 249322 2278 249558
rect 2362 249322 2598 249558
rect 2682 249322 2918 249558
rect 3002 249322 3238 249558
rect 3322 249322 3558 249558
rect 3642 249322 3878 249558
rect 231838 252842 232074 253078
rect 232158 252842 232394 253078
rect 232478 252842 232714 253078
rect 232798 252842 233034 253078
rect 233118 252842 233354 253078
rect 233438 252842 233674 253078
rect 233758 252842 233994 253078
rect 234078 252842 234314 253078
rect 234398 252842 234634 253078
rect 234718 252842 234954 253078
rect 235038 252842 235274 253078
rect 235358 252842 235594 253078
rect 231838 252522 232074 252758
rect 232158 252522 232394 252758
rect 232478 252522 232714 252758
rect 232798 252522 233034 252758
rect 233118 252522 233354 252758
rect 233438 252522 233674 252758
rect 233758 252522 233994 252758
rect 234078 252522 234314 252758
rect 234398 252522 234634 252758
rect 234718 252522 234954 252758
rect 235038 252522 235274 252758
rect 235358 252522 235594 252758
rect 231838 252202 232074 252438
rect 232158 252202 232394 252438
rect 232478 252202 232714 252438
rect 232798 252202 233034 252438
rect 233118 252202 233354 252438
rect 233438 252202 233674 252438
rect 233758 252202 233994 252438
rect 234078 252202 234314 252438
rect 234398 252202 234634 252438
rect 234718 252202 234954 252438
rect 235038 252202 235274 252438
rect 235358 252202 235594 252438
rect 231838 251882 232074 252118
rect 232158 251882 232394 252118
rect 232478 251882 232714 252118
rect 232798 251882 233034 252118
rect 233118 251882 233354 252118
rect 233438 251882 233674 252118
rect 233758 251882 233994 252118
rect 234078 251882 234314 252118
rect 234398 251882 234634 252118
rect 234718 251882 234954 252118
rect 235038 251882 235274 252118
rect 235358 251882 235594 252118
rect 231838 251562 232074 251798
rect 232158 251562 232394 251798
rect 232478 251562 232714 251798
rect 232798 251562 233034 251798
rect 233118 251562 233354 251798
rect 233438 251562 233674 251798
rect 233758 251562 233994 251798
rect 234078 251562 234314 251798
rect 234398 251562 234634 251798
rect 234718 251562 234954 251798
rect 235038 251562 235274 251798
rect 235358 251562 235594 251798
rect 231838 251242 232074 251478
rect 232158 251242 232394 251478
rect 232478 251242 232714 251478
rect 232798 251242 233034 251478
rect 233118 251242 233354 251478
rect 233438 251242 233674 251478
rect 233758 251242 233994 251478
rect 234078 251242 234314 251478
rect 234398 251242 234634 251478
rect 234718 251242 234954 251478
rect 235038 251242 235274 251478
rect 235358 251242 235594 251478
rect 231838 250922 232074 251158
rect 232158 250922 232394 251158
rect 232478 250922 232714 251158
rect 232798 250922 233034 251158
rect 233118 250922 233354 251158
rect 233438 250922 233674 251158
rect 233758 250922 233994 251158
rect 234078 250922 234314 251158
rect 234398 250922 234634 251158
rect 234718 250922 234954 251158
rect 235038 250922 235274 251158
rect 235358 250922 235594 251158
rect 231838 250602 232074 250838
rect 232158 250602 232394 250838
rect 232478 250602 232714 250838
rect 232798 250602 233034 250838
rect 233118 250602 233354 250838
rect 233438 250602 233674 250838
rect 233758 250602 233994 250838
rect 234078 250602 234314 250838
rect 234398 250602 234634 250838
rect 234718 250602 234954 250838
rect 235038 250602 235274 250838
rect 235358 250602 235594 250838
rect 231838 250282 232074 250518
rect 232158 250282 232394 250518
rect 232478 250282 232714 250518
rect 232798 250282 233034 250518
rect 233118 250282 233354 250518
rect 233438 250282 233674 250518
rect 233758 250282 233994 250518
rect 234078 250282 234314 250518
rect 234398 250282 234634 250518
rect 234718 250282 234954 250518
rect 235038 250282 235274 250518
rect 235358 250282 235594 250518
rect 231838 249962 232074 250198
rect 232158 249962 232394 250198
rect 232478 249962 232714 250198
rect 232798 249962 233034 250198
rect 233118 249962 233354 250198
rect 233438 249962 233674 250198
rect 233758 249962 233994 250198
rect 234078 249962 234314 250198
rect 234398 249962 234634 250198
rect 234718 249962 234954 250198
rect 235038 249962 235274 250198
rect 235358 249962 235594 250198
rect 231838 249642 232074 249878
rect 232158 249642 232394 249878
rect 232478 249642 232714 249878
rect 232798 249642 233034 249878
rect 233118 249642 233354 249878
rect 233438 249642 233674 249878
rect 233758 249642 233994 249878
rect 234078 249642 234314 249878
rect 234398 249642 234634 249878
rect 234718 249642 234954 249878
rect 235038 249642 235274 249878
rect 235358 249642 235594 249878
rect 231838 249322 232074 249558
rect 232158 249322 232394 249558
rect 232478 249322 232714 249558
rect 232798 249322 233034 249558
rect 233118 249322 233354 249558
rect 233438 249322 233674 249558
rect 233758 249322 233994 249558
rect 234078 249322 234314 249558
rect 234398 249322 234634 249558
rect 234718 249322 234954 249558
rect 235038 249322 235274 249558
rect 235358 249322 235594 249558
rect 122 228682 358 228918
rect 442 228682 678 228918
rect 762 228682 998 228918
rect 1082 228682 1318 228918
rect 1402 228682 1638 228918
rect 1722 228682 1958 228918
rect 2042 228682 2278 228918
rect 2362 228682 2598 228918
rect 2682 228682 2918 228918
rect 3002 228682 3238 228918
rect 3322 228682 3558 228918
rect 3642 228682 3878 228918
rect 122 206282 358 206518
rect 442 206282 678 206518
rect 762 206282 998 206518
rect 1082 206282 1318 206518
rect 1402 206282 1638 206518
rect 1722 206282 1958 206518
rect 2042 206282 2278 206518
rect 2362 206282 2598 206518
rect 2682 206282 2918 206518
rect 3002 206282 3238 206518
rect 3322 206282 3558 206518
rect 3642 206282 3878 206518
rect 122 183882 358 184118
rect 442 183882 678 184118
rect 762 183882 998 184118
rect 1082 183882 1318 184118
rect 1402 183882 1638 184118
rect 1722 183882 1958 184118
rect 2042 183882 2278 184118
rect 2362 183882 2598 184118
rect 2682 183882 2918 184118
rect 3002 183882 3238 184118
rect 3322 183882 3558 184118
rect 3642 183882 3878 184118
rect 122 161482 358 161718
rect 442 161482 678 161718
rect 762 161482 998 161718
rect 1082 161482 1318 161718
rect 1402 161482 1638 161718
rect 1722 161482 1958 161718
rect 2042 161482 2278 161718
rect 2362 161482 2598 161718
rect 2682 161482 2918 161718
rect 3002 161482 3238 161718
rect 3322 161482 3558 161718
rect 3642 161482 3878 161718
rect 122 139082 358 139318
rect 442 139082 678 139318
rect 762 139082 998 139318
rect 1082 139082 1318 139318
rect 1402 139082 1638 139318
rect 1722 139082 1958 139318
rect 2042 139082 2278 139318
rect 2362 139082 2598 139318
rect 2682 139082 2918 139318
rect 3002 139082 3238 139318
rect 3322 139082 3558 139318
rect 3642 139082 3878 139318
rect 122 116682 358 116918
rect 442 116682 678 116918
rect 762 116682 998 116918
rect 1082 116682 1318 116918
rect 1402 116682 1638 116918
rect 1722 116682 1958 116918
rect 2042 116682 2278 116918
rect 2362 116682 2598 116918
rect 2682 116682 2918 116918
rect 3002 116682 3238 116918
rect 3322 116682 3558 116918
rect 3642 116682 3878 116918
rect 122 94282 358 94518
rect 442 94282 678 94518
rect 762 94282 998 94518
rect 1082 94282 1318 94518
rect 1402 94282 1638 94518
rect 1722 94282 1958 94518
rect 2042 94282 2278 94518
rect 2362 94282 2598 94518
rect 2682 94282 2918 94518
rect 3002 94282 3238 94518
rect 3322 94282 3558 94518
rect 3642 94282 3878 94518
rect 122 71882 358 72118
rect 442 71882 678 72118
rect 762 71882 998 72118
rect 1082 71882 1318 72118
rect 1402 71882 1638 72118
rect 1722 71882 1958 72118
rect 2042 71882 2278 72118
rect 2362 71882 2598 72118
rect 2682 71882 2918 72118
rect 3002 71882 3238 72118
rect 3322 71882 3558 72118
rect 3642 71882 3878 72118
rect 122 49482 358 49718
rect 442 49482 678 49718
rect 762 49482 998 49718
rect 1082 49482 1318 49718
rect 1402 49482 1638 49718
rect 1722 49482 1958 49718
rect 2042 49482 2278 49718
rect 2362 49482 2598 49718
rect 2682 49482 2918 49718
rect 3002 49482 3238 49718
rect 3322 49482 3558 49718
rect 3642 49482 3878 49718
rect 122 27082 358 27318
rect 442 27082 678 27318
rect 762 27082 998 27318
rect 1082 27082 1318 27318
rect 1402 27082 1638 27318
rect 1722 27082 1958 27318
rect 2042 27082 2278 27318
rect 2362 27082 2598 27318
rect 2682 27082 2918 27318
rect 3002 27082 3238 27318
rect 3322 27082 3558 27318
rect 3642 27082 3878 27318
rect 5122 247842 5358 248078
rect 5442 247842 5678 248078
rect 5762 247842 5998 248078
rect 6082 247842 6318 248078
rect 6402 247842 6638 248078
rect 6722 247842 6958 248078
rect 7042 247842 7278 248078
rect 7362 247842 7598 248078
rect 7682 247842 7918 248078
rect 8002 247842 8238 248078
rect 8322 247842 8558 248078
rect 8642 247842 8878 248078
rect 5122 247522 5358 247758
rect 5442 247522 5678 247758
rect 5762 247522 5998 247758
rect 6082 247522 6318 247758
rect 6402 247522 6638 247758
rect 6722 247522 6958 247758
rect 7042 247522 7278 247758
rect 7362 247522 7598 247758
rect 7682 247522 7918 247758
rect 8002 247522 8238 247758
rect 8322 247522 8558 247758
rect 8642 247522 8878 247758
rect 5122 247202 5358 247438
rect 5442 247202 5678 247438
rect 5762 247202 5998 247438
rect 6082 247202 6318 247438
rect 6402 247202 6638 247438
rect 6722 247202 6958 247438
rect 7042 247202 7278 247438
rect 7362 247202 7598 247438
rect 7682 247202 7918 247438
rect 8002 247202 8238 247438
rect 8322 247202 8558 247438
rect 8642 247202 8878 247438
rect 5122 246882 5358 247118
rect 5442 246882 5678 247118
rect 5762 246882 5998 247118
rect 6082 246882 6318 247118
rect 6402 246882 6638 247118
rect 6722 246882 6958 247118
rect 7042 246882 7278 247118
rect 7362 246882 7598 247118
rect 7682 246882 7918 247118
rect 8002 246882 8238 247118
rect 8322 246882 8558 247118
rect 8642 246882 8878 247118
rect 5122 246562 5358 246798
rect 5442 246562 5678 246798
rect 5762 246562 5998 246798
rect 6082 246562 6318 246798
rect 6402 246562 6638 246798
rect 6722 246562 6958 246798
rect 7042 246562 7278 246798
rect 7362 246562 7598 246798
rect 7682 246562 7918 246798
rect 8002 246562 8238 246798
rect 8322 246562 8558 246798
rect 8642 246562 8878 246798
rect 5122 246242 5358 246478
rect 5442 246242 5678 246478
rect 5762 246242 5998 246478
rect 6082 246242 6318 246478
rect 6402 246242 6638 246478
rect 6722 246242 6958 246478
rect 7042 246242 7278 246478
rect 7362 246242 7598 246478
rect 7682 246242 7918 246478
rect 8002 246242 8238 246478
rect 8322 246242 8558 246478
rect 8642 246242 8878 246478
rect 5122 245922 5358 246158
rect 5442 245922 5678 246158
rect 5762 245922 5998 246158
rect 6082 245922 6318 246158
rect 6402 245922 6638 246158
rect 6722 245922 6958 246158
rect 7042 245922 7278 246158
rect 7362 245922 7598 246158
rect 7682 245922 7918 246158
rect 8002 245922 8238 246158
rect 8322 245922 8558 246158
rect 8642 245922 8878 246158
rect 5122 245602 5358 245838
rect 5442 245602 5678 245838
rect 5762 245602 5998 245838
rect 6082 245602 6318 245838
rect 6402 245602 6638 245838
rect 6722 245602 6958 245838
rect 7042 245602 7278 245838
rect 7362 245602 7598 245838
rect 7682 245602 7918 245838
rect 8002 245602 8238 245838
rect 8322 245602 8558 245838
rect 8642 245602 8878 245838
rect 5122 245282 5358 245518
rect 5442 245282 5678 245518
rect 5762 245282 5998 245518
rect 6082 245282 6318 245518
rect 6402 245282 6638 245518
rect 6722 245282 6958 245518
rect 7042 245282 7278 245518
rect 7362 245282 7598 245518
rect 7682 245282 7918 245518
rect 8002 245282 8238 245518
rect 8322 245282 8558 245518
rect 8642 245282 8878 245518
rect 5122 244962 5358 245198
rect 5442 244962 5678 245198
rect 5762 244962 5998 245198
rect 6082 244962 6318 245198
rect 6402 244962 6638 245198
rect 6722 244962 6958 245198
rect 7042 244962 7278 245198
rect 7362 244962 7598 245198
rect 7682 244962 7918 245198
rect 8002 244962 8238 245198
rect 8322 244962 8558 245198
rect 8642 244962 8878 245198
rect 5122 244642 5358 244878
rect 5442 244642 5678 244878
rect 5762 244642 5998 244878
rect 6082 244642 6318 244878
rect 6402 244642 6638 244878
rect 6722 244642 6958 244878
rect 7042 244642 7278 244878
rect 7362 244642 7598 244878
rect 7682 244642 7918 244878
rect 8002 244642 8238 244878
rect 8322 244642 8558 244878
rect 8642 244642 8878 244878
rect 5122 244322 5358 244558
rect 5442 244322 5678 244558
rect 5762 244322 5998 244558
rect 6082 244322 6318 244558
rect 6402 244322 6638 244558
rect 6722 244322 6958 244558
rect 7042 244322 7278 244558
rect 7362 244322 7598 244558
rect 7682 244322 7918 244558
rect 8002 244322 8238 244558
rect 8322 244322 8558 244558
rect 8642 244322 8878 244558
rect 5122 239882 5358 240118
rect 5442 239882 5678 240118
rect 5762 239882 5998 240118
rect 6082 239882 6318 240118
rect 6402 239882 6638 240118
rect 6722 239882 6958 240118
rect 7042 239882 7278 240118
rect 7362 239882 7598 240118
rect 7682 239882 7918 240118
rect 8002 239882 8238 240118
rect 8322 239882 8558 240118
rect 8642 239882 8878 240118
rect 226838 247842 227074 248078
rect 227158 247842 227394 248078
rect 227478 247842 227714 248078
rect 227798 247842 228034 248078
rect 228118 247842 228354 248078
rect 228438 247842 228674 248078
rect 228758 247842 228994 248078
rect 229078 247842 229314 248078
rect 229398 247842 229634 248078
rect 229718 247842 229954 248078
rect 230038 247842 230274 248078
rect 230358 247842 230594 248078
rect 226838 247522 227074 247758
rect 227158 247522 227394 247758
rect 227478 247522 227714 247758
rect 227798 247522 228034 247758
rect 228118 247522 228354 247758
rect 228438 247522 228674 247758
rect 228758 247522 228994 247758
rect 229078 247522 229314 247758
rect 229398 247522 229634 247758
rect 229718 247522 229954 247758
rect 230038 247522 230274 247758
rect 230358 247522 230594 247758
rect 226838 247202 227074 247438
rect 227158 247202 227394 247438
rect 227478 247202 227714 247438
rect 227798 247202 228034 247438
rect 228118 247202 228354 247438
rect 228438 247202 228674 247438
rect 228758 247202 228994 247438
rect 229078 247202 229314 247438
rect 229398 247202 229634 247438
rect 229718 247202 229954 247438
rect 230038 247202 230274 247438
rect 230358 247202 230594 247438
rect 226838 246882 227074 247118
rect 227158 246882 227394 247118
rect 227478 246882 227714 247118
rect 227798 246882 228034 247118
rect 228118 246882 228354 247118
rect 228438 246882 228674 247118
rect 228758 246882 228994 247118
rect 229078 246882 229314 247118
rect 229398 246882 229634 247118
rect 229718 246882 229954 247118
rect 230038 246882 230274 247118
rect 230358 246882 230594 247118
rect 226838 246562 227074 246798
rect 227158 246562 227394 246798
rect 227478 246562 227714 246798
rect 227798 246562 228034 246798
rect 228118 246562 228354 246798
rect 228438 246562 228674 246798
rect 228758 246562 228994 246798
rect 229078 246562 229314 246798
rect 229398 246562 229634 246798
rect 229718 246562 229954 246798
rect 230038 246562 230274 246798
rect 230358 246562 230594 246798
rect 226838 246242 227074 246478
rect 227158 246242 227394 246478
rect 227478 246242 227714 246478
rect 227798 246242 228034 246478
rect 228118 246242 228354 246478
rect 228438 246242 228674 246478
rect 228758 246242 228994 246478
rect 229078 246242 229314 246478
rect 229398 246242 229634 246478
rect 229718 246242 229954 246478
rect 230038 246242 230274 246478
rect 230358 246242 230594 246478
rect 226838 245922 227074 246158
rect 227158 245922 227394 246158
rect 227478 245922 227714 246158
rect 227798 245922 228034 246158
rect 228118 245922 228354 246158
rect 228438 245922 228674 246158
rect 228758 245922 228994 246158
rect 229078 245922 229314 246158
rect 229398 245922 229634 246158
rect 229718 245922 229954 246158
rect 230038 245922 230274 246158
rect 230358 245922 230594 246158
rect 226838 245602 227074 245838
rect 227158 245602 227394 245838
rect 227478 245602 227714 245838
rect 227798 245602 228034 245838
rect 228118 245602 228354 245838
rect 228438 245602 228674 245838
rect 228758 245602 228994 245838
rect 229078 245602 229314 245838
rect 229398 245602 229634 245838
rect 229718 245602 229954 245838
rect 230038 245602 230274 245838
rect 230358 245602 230594 245838
rect 226838 245282 227074 245518
rect 227158 245282 227394 245518
rect 227478 245282 227714 245518
rect 227798 245282 228034 245518
rect 228118 245282 228354 245518
rect 228438 245282 228674 245518
rect 228758 245282 228994 245518
rect 229078 245282 229314 245518
rect 229398 245282 229634 245518
rect 229718 245282 229954 245518
rect 230038 245282 230274 245518
rect 230358 245282 230594 245518
rect 226838 244962 227074 245198
rect 227158 244962 227394 245198
rect 227478 244962 227714 245198
rect 227798 244962 228034 245198
rect 228118 244962 228354 245198
rect 228438 244962 228674 245198
rect 228758 244962 228994 245198
rect 229078 244962 229314 245198
rect 229398 244962 229634 245198
rect 229718 244962 229954 245198
rect 230038 244962 230274 245198
rect 230358 244962 230594 245198
rect 226838 244642 227074 244878
rect 227158 244642 227394 244878
rect 227478 244642 227714 244878
rect 227798 244642 228034 244878
rect 228118 244642 228354 244878
rect 228438 244642 228674 244878
rect 228758 244642 228994 244878
rect 229078 244642 229314 244878
rect 229398 244642 229634 244878
rect 229718 244642 229954 244878
rect 230038 244642 230274 244878
rect 230358 244642 230594 244878
rect 226838 244322 227074 244558
rect 227158 244322 227394 244558
rect 227478 244322 227714 244558
rect 227798 244322 228034 244558
rect 228118 244322 228354 244558
rect 228438 244322 228674 244558
rect 228758 244322 228994 244558
rect 229078 244322 229314 244558
rect 229398 244322 229634 244558
rect 229718 244322 229954 244558
rect 230038 244322 230274 244558
rect 230358 244322 230594 244558
rect 226838 239882 227074 240118
rect 227158 239882 227394 240118
rect 227478 239882 227714 240118
rect 227798 239882 228034 240118
rect 228118 239882 228354 240118
rect 228438 239882 228674 240118
rect 228758 239882 228994 240118
rect 229078 239882 229314 240118
rect 229398 239882 229634 240118
rect 229718 239882 229954 240118
rect 230038 239882 230274 240118
rect 230358 239882 230594 240118
rect 5122 217482 5358 217718
rect 5442 217482 5678 217718
rect 5762 217482 5998 217718
rect 6082 217482 6318 217718
rect 6402 217482 6638 217718
rect 6722 217482 6958 217718
rect 7042 217482 7278 217718
rect 7362 217482 7598 217718
rect 7682 217482 7918 217718
rect 8002 217482 8238 217718
rect 8322 217482 8558 217718
rect 8642 217482 8878 217718
rect 5122 195082 5358 195318
rect 5442 195082 5678 195318
rect 5762 195082 5998 195318
rect 6082 195082 6318 195318
rect 6402 195082 6638 195318
rect 6722 195082 6958 195318
rect 7042 195082 7278 195318
rect 7362 195082 7598 195318
rect 7682 195082 7918 195318
rect 8002 195082 8238 195318
rect 8322 195082 8558 195318
rect 8642 195082 8878 195318
rect 5122 172682 5358 172918
rect 5442 172682 5678 172918
rect 5762 172682 5998 172918
rect 6082 172682 6318 172918
rect 6402 172682 6638 172918
rect 6722 172682 6958 172918
rect 7042 172682 7278 172918
rect 7362 172682 7598 172918
rect 7682 172682 7918 172918
rect 8002 172682 8238 172918
rect 8322 172682 8558 172918
rect 8642 172682 8878 172918
rect 29927 228682 30163 228918
rect 71882 228682 72118 228918
rect 25261 217482 25497 217718
rect 66882 217482 67118 217718
rect 114215 228682 114451 228918
rect 109549 217482 109785 217718
rect 32215 183882 32451 184118
rect 75506 183882 75742 184118
rect 116215 183882 116451 184118
rect 26430 178366 26666 178602
rect 41886 178588 41972 178602
rect 41972 178588 42036 178602
rect 42036 178588 42122 178602
rect 41886 178366 42122 178588
rect 29549 172682 29785 172918
rect 60146 172682 60382 172918
rect 113549 172682 113785 172918
rect 155882 228682 156118 228918
rect 150882 217482 151118 217718
rect 198215 228682 198451 228918
rect 193549 217482 193785 217718
rect 226838 217482 227074 217718
rect 227158 217482 227394 217718
rect 227478 217482 227714 217718
rect 227798 217482 228034 217718
rect 228118 217482 228354 217718
rect 228438 217482 228674 217718
rect 228758 217482 228994 217718
rect 229078 217482 229314 217718
rect 229398 217482 229634 217718
rect 229718 217482 229954 217718
rect 230038 217482 230274 217718
rect 230358 217482 230594 217718
rect 139406 164780 139642 165002
rect 139406 164766 139492 164780
rect 139492 164766 139556 164780
rect 139556 164766 139642 164780
rect 26430 163406 26666 163642
rect 41702 163406 41938 163642
rect 32215 161482 32451 161718
rect 75506 161482 75742 161718
rect 116215 161482 116451 161718
rect 5122 150282 5358 150518
rect 5442 150282 5678 150518
rect 5762 150282 5998 150518
rect 6082 150282 6318 150518
rect 6402 150282 6638 150518
rect 6722 150282 6958 150518
rect 7042 150282 7278 150518
rect 7362 150282 7598 150518
rect 7682 150282 7918 150518
rect 8002 150282 8238 150518
rect 8322 150282 8558 150518
rect 8642 150282 8878 150518
rect 5122 127882 5358 128118
rect 5442 127882 5678 128118
rect 5762 127882 5998 128118
rect 6082 127882 6318 128118
rect 6402 127882 6638 128118
rect 6722 127882 6958 128118
rect 7042 127882 7278 128118
rect 7362 127882 7598 128118
rect 7682 127882 7918 128118
rect 8002 127882 8238 128118
rect 8322 127882 8558 128118
rect 8642 127882 8878 128118
rect 25549 127882 25785 128118
rect 66882 127882 67118 128118
rect 109549 127882 109785 128118
rect 30215 116682 30451 116918
rect 114215 116682 114451 116918
rect 61942 111196 62178 111282
rect 61942 111132 62028 111196
rect 62028 111132 62092 111196
rect 62092 111132 62178 111196
rect 61942 111046 62178 111132
rect 108310 111196 108546 111282
rect 108310 111132 108396 111196
rect 108396 111132 108460 111196
rect 108460 111132 108546 111196
rect 108310 111046 108546 111132
rect 133886 111196 134122 111282
rect 133886 111132 133972 111196
rect 133972 111132 134036 111196
rect 134036 111132 134122 111196
rect 133886 111046 134122 111132
rect 5122 105482 5358 105718
rect 5442 105482 5678 105718
rect 5762 105482 5998 105718
rect 6082 105482 6318 105718
rect 6402 105482 6638 105718
rect 6722 105482 6958 105718
rect 7042 105482 7278 105718
rect 7362 105482 7598 105718
rect 7682 105482 7918 105718
rect 8002 105482 8238 105718
rect 8322 105482 8558 105718
rect 8642 105482 8878 105718
rect 32215 94282 32451 94518
rect 75506 94282 75742 94518
rect 116215 94282 116451 94518
rect 5122 83082 5358 83318
rect 5442 83082 5678 83318
rect 5762 83082 5998 83318
rect 6082 83082 6318 83318
rect 6402 83082 6638 83318
rect 6722 83082 6958 83318
rect 7042 83082 7278 83318
rect 7362 83082 7598 83318
rect 7682 83082 7918 83318
rect 8002 83082 8238 83318
rect 8322 83082 8558 83318
rect 8642 83082 8878 83318
rect 29549 83082 29785 83318
rect 60146 83082 60382 83318
rect 113549 83082 113785 83318
rect 25510 76516 25746 76602
rect 25510 76452 25596 76516
rect 25596 76452 25660 76516
rect 25660 76452 25746 76516
rect 25510 76366 25746 76452
rect 41702 76516 41938 76602
rect 41702 76452 41788 76516
rect 41788 76452 41852 76516
rect 41852 76452 41938 76516
rect 41702 76366 41938 76452
rect 32215 71882 32451 72118
rect 75506 71882 75742 72118
rect 116215 71882 116451 72118
rect 25694 69580 25930 69802
rect 25694 69566 25780 69580
rect 25780 69566 25844 69580
rect 25844 69566 25930 69580
rect 41702 69788 41788 69802
rect 41788 69788 41852 69802
rect 41852 69788 41938 69802
rect 41702 69566 41938 69788
rect 5122 60682 5358 60918
rect 5442 60682 5678 60918
rect 5762 60682 5998 60918
rect 6082 60682 6318 60918
rect 6402 60682 6638 60918
rect 6722 60682 6958 60918
rect 7042 60682 7278 60918
rect 7362 60682 7598 60918
rect 7682 60682 7918 60918
rect 8002 60682 8238 60918
rect 8322 60682 8558 60918
rect 8642 60682 8878 60918
rect 226838 195082 227074 195318
rect 227158 195082 227394 195318
rect 227478 195082 227714 195318
rect 227798 195082 228034 195318
rect 228118 195082 228354 195318
rect 228438 195082 228674 195318
rect 228758 195082 228994 195318
rect 229078 195082 229314 195318
rect 229398 195082 229634 195318
rect 229718 195082 229954 195318
rect 230038 195082 230274 195318
rect 230358 195082 230594 195318
rect 193870 190620 194106 190842
rect 193870 190606 193956 190620
rect 193956 190606 194020 190620
rect 194020 190606 194106 190620
rect 209878 190756 210114 190842
rect 209878 190692 209964 190756
rect 209964 190692 210028 190756
rect 210028 190692 210114 190756
rect 209878 190606 210114 190692
rect 159506 183882 159742 184118
rect 200215 183882 200451 184118
rect 144146 172682 144382 172918
rect 197549 172682 197785 172918
rect 226838 172682 227074 172918
rect 227158 172682 227394 172918
rect 227478 172682 227714 172918
rect 227798 172682 228034 172918
rect 228118 172682 228354 172918
rect 228438 172682 228674 172918
rect 228758 172682 228994 172918
rect 229078 172682 229314 172918
rect 229398 172682 229634 172918
rect 229718 172682 229954 172918
rect 230038 172682 230274 172918
rect 230358 172682 230594 172918
rect 212454 164916 212690 165002
rect 212454 164852 212540 164916
rect 212540 164852 212604 164916
rect 212604 164852 212690 164916
rect 212454 164766 212690 164852
rect 159506 161482 159742 161718
rect 200215 161482 200451 161718
rect 226838 150282 227074 150518
rect 227158 150282 227394 150518
rect 227478 150282 227714 150518
rect 227798 150282 228034 150518
rect 228118 150282 228354 150518
rect 228438 150282 228674 150518
rect 228758 150282 228994 150518
rect 229078 150282 229314 150518
rect 229398 150282 229634 150518
rect 229718 150282 229954 150518
rect 230038 150282 230274 150518
rect 230358 150282 230594 150518
rect 150882 127882 151118 128118
rect 193549 127882 193785 128118
rect 226838 127882 227074 128118
rect 227158 127882 227394 128118
rect 227478 127882 227714 128118
rect 227798 127882 228034 128118
rect 228118 127882 228354 128118
rect 228438 127882 228674 128118
rect 228758 127882 228994 128118
rect 229078 127882 229314 128118
rect 229398 127882 229634 128118
rect 229718 127882 229954 128118
rect 230038 127882 230274 128118
rect 230358 127882 230594 128118
rect 198215 116682 198451 116918
rect 226838 105482 227074 105718
rect 227158 105482 227394 105718
rect 227478 105482 227714 105718
rect 227798 105482 228034 105718
rect 228118 105482 228354 105718
rect 228438 105482 228674 105718
rect 228758 105482 228994 105718
rect 229078 105482 229314 105718
rect 229398 105482 229634 105718
rect 229718 105482 229954 105718
rect 230038 105482 230274 105718
rect 230358 105482 230594 105718
rect 193686 96916 193922 97002
rect 193686 96852 193772 96916
rect 193772 96852 193836 96916
rect 193836 96852 193922 96916
rect 193686 96766 193922 96852
rect 209694 96780 209930 97002
rect 209694 96766 209780 96780
rect 209780 96766 209844 96780
rect 209844 96766 209930 96780
rect 159506 94282 159742 94518
rect 200215 94282 200451 94518
rect 144146 83082 144382 83318
rect 197549 83082 197785 83318
rect 226838 83082 227074 83318
rect 227158 83082 227394 83318
rect 227478 83082 227714 83318
rect 227798 83082 228034 83318
rect 228118 83082 228354 83318
rect 228438 83082 228674 83318
rect 228758 83082 228994 83318
rect 229078 83082 229314 83318
rect 229398 83082 229634 83318
rect 229718 83082 229954 83318
rect 230038 83082 230274 83318
rect 230358 83082 230594 83318
rect 159506 71882 159742 72118
rect 200215 71882 200451 72118
rect 5122 38282 5358 38518
rect 5442 38282 5678 38518
rect 5762 38282 5998 38518
rect 6082 38282 6318 38518
rect 6402 38282 6638 38518
rect 6722 38282 6958 38518
rect 7042 38282 7278 38518
rect 7362 38282 7598 38518
rect 7682 38282 7918 38518
rect 8002 38282 8238 38518
rect 8322 38282 8558 38518
rect 8642 38282 8878 38518
rect 25549 38282 25785 38518
rect 30215 27082 30451 27318
rect 19622 22646 19858 22882
rect 53846 22796 54082 22882
rect 53846 22732 53932 22796
rect 53932 22732 53996 22796
rect 53996 22732 54082 22796
rect 53846 22646 54082 22732
rect 66882 38282 67118 38518
rect 71882 27082 72118 27318
rect 88990 20606 89226 20842
rect 109549 38282 109785 38518
rect 114215 27082 114451 27318
rect 100950 20828 101036 20842
rect 101036 20828 101100 20842
rect 101100 20828 101186 20842
rect 100950 20606 101186 20828
rect 89726 19926 89962 20162
rect 100950 20148 101036 20162
rect 101036 20148 101100 20162
rect 101100 20148 101186 20162
rect 100950 19926 101186 20148
rect 150882 38282 151118 38518
rect 155882 27082 156118 27318
rect 226838 60682 227074 60918
rect 227158 60682 227394 60918
rect 227478 60682 227714 60918
rect 227798 60682 228034 60918
rect 228118 60682 228354 60918
rect 228438 60682 228674 60918
rect 228758 60682 228994 60918
rect 229078 60682 229314 60918
rect 229398 60682 229634 60918
rect 229718 60682 229954 60918
rect 230038 60682 230274 60918
rect 230358 60682 230594 60918
rect 211350 45086 211586 45322
rect 172894 20606 173130 20842
rect 193549 38282 193785 38518
rect 213742 45086 213978 45322
rect 212638 34886 212874 35122
rect 226838 38282 227074 38518
rect 227158 38282 227394 38518
rect 227478 38282 227714 38518
rect 227798 38282 228034 38518
rect 228118 38282 228354 38518
rect 228438 38282 228674 38518
rect 228758 38282 228994 38518
rect 229078 38282 229314 38518
rect 229398 38282 229634 38518
rect 229718 38282 229954 38518
rect 230038 38282 230274 38518
rect 230358 38282 230594 38518
rect 213742 34886 213978 35122
rect 198215 27082 198451 27318
rect 173814 21966 174050 22202
rect 185038 21980 185274 22202
rect 185038 21966 185124 21980
rect 185124 21966 185188 21980
rect 185188 21966 185274 21980
rect 185038 20756 185274 20842
rect 185038 20692 185124 20756
rect 185124 20692 185188 20756
rect 185188 20692 185274 20756
rect 185038 20606 185274 20692
rect 173262 19926 173498 20162
rect 185406 19926 185642 20162
rect 5122 15882 5358 16118
rect 5442 15882 5678 16118
rect 5762 15882 5998 16118
rect 6082 15882 6318 16118
rect 6402 15882 6638 16118
rect 6722 15882 6958 16118
rect 7042 15882 7278 16118
rect 7362 15882 7598 16118
rect 7682 15882 7918 16118
rect 8002 15882 8238 16118
rect 8322 15882 8558 16118
rect 8642 15882 8878 16118
rect 5122 8642 5358 8878
rect 5442 8642 5678 8878
rect 5762 8642 5998 8878
rect 6082 8642 6318 8878
rect 6402 8642 6638 8878
rect 6722 8642 6958 8878
rect 7042 8642 7278 8878
rect 7362 8642 7598 8878
rect 7682 8642 7918 8878
rect 8002 8642 8238 8878
rect 8322 8642 8558 8878
rect 8642 8642 8878 8878
rect 5122 8322 5358 8558
rect 5442 8322 5678 8558
rect 5762 8322 5998 8558
rect 6082 8322 6318 8558
rect 6402 8322 6638 8558
rect 6722 8322 6958 8558
rect 7042 8322 7278 8558
rect 7362 8322 7598 8558
rect 7682 8322 7918 8558
rect 8002 8322 8238 8558
rect 8322 8322 8558 8558
rect 8642 8322 8878 8558
rect 5122 8002 5358 8238
rect 5442 8002 5678 8238
rect 5762 8002 5998 8238
rect 6082 8002 6318 8238
rect 6402 8002 6638 8238
rect 6722 8002 6958 8238
rect 7042 8002 7278 8238
rect 7362 8002 7598 8238
rect 7682 8002 7918 8238
rect 8002 8002 8238 8238
rect 8322 8002 8558 8238
rect 8642 8002 8878 8238
rect 5122 7682 5358 7918
rect 5442 7682 5678 7918
rect 5762 7682 5998 7918
rect 6082 7682 6318 7918
rect 6402 7682 6638 7918
rect 6722 7682 6958 7918
rect 7042 7682 7278 7918
rect 7362 7682 7598 7918
rect 7682 7682 7918 7918
rect 8002 7682 8238 7918
rect 8322 7682 8558 7918
rect 8642 7682 8878 7918
rect 5122 7362 5358 7598
rect 5442 7362 5678 7598
rect 5762 7362 5998 7598
rect 6082 7362 6318 7598
rect 6402 7362 6638 7598
rect 6722 7362 6958 7598
rect 7042 7362 7278 7598
rect 7362 7362 7598 7598
rect 7682 7362 7918 7598
rect 8002 7362 8238 7598
rect 8322 7362 8558 7598
rect 8642 7362 8878 7598
rect 5122 7042 5358 7278
rect 5442 7042 5678 7278
rect 5762 7042 5998 7278
rect 6082 7042 6318 7278
rect 6402 7042 6638 7278
rect 6722 7042 6958 7278
rect 7042 7042 7278 7278
rect 7362 7042 7598 7278
rect 7682 7042 7918 7278
rect 8002 7042 8238 7278
rect 8322 7042 8558 7278
rect 8642 7042 8878 7278
rect 5122 6722 5358 6958
rect 5442 6722 5678 6958
rect 5762 6722 5998 6958
rect 6082 6722 6318 6958
rect 6402 6722 6638 6958
rect 6722 6722 6958 6958
rect 7042 6722 7278 6958
rect 7362 6722 7598 6958
rect 7682 6722 7918 6958
rect 8002 6722 8238 6958
rect 8322 6722 8558 6958
rect 8642 6722 8878 6958
rect 5122 6402 5358 6638
rect 5442 6402 5678 6638
rect 5762 6402 5998 6638
rect 6082 6402 6318 6638
rect 6402 6402 6638 6638
rect 6722 6402 6958 6638
rect 7042 6402 7278 6638
rect 7362 6402 7598 6638
rect 7682 6402 7918 6638
rect 8002 6402 8238 6638
rect 8322 6402 8558 6638
rect 8642 6402 8878 6638
rect 5122 6082 5358 6318
rect 5442 6082 5678 6318
rect 5762 6082 5998 6318
rect 6082 6082 6318 6318
rect 6402 6082 6638 6318
rect 6722 6082 6958 6318
rect 7042 6082 7278 6318
rect 7362 6082 7598 6318
rect 7682 6082 7918 6318
rect 8002 6082 8238 6318
rect 8322 6082 8558 6318
rect 8642 6082 8878 6318
rect 5122 5762 5358 5998
rect 5442 5762 5678 5998
rect 5762 5762 5998 5998
rect 6082 5762 6318 5998
rect 6402 5762 6638 5998
rect 6722 5762 6958 5998
rect 7042 5762 7278 5998
rect 7362 5762 7598 5998
rect 7682 5762 7918 5998
rect 8002 5762 8238 5998
rect 8322 5762 8558 5998
rect 8642 5762 8878 5998
rect 5122 5442 5358 5678
rect 5442 5442 5678 5678
rect 5762 5442 5998 5678
rect 6082 5442 6318 5678
rect 6402 5442 6638 5678
rect 6722 5442 6958 5678
rect 7042 5442 7278 5678
rect 7362 5442 7598 5678
rect 7682 5442 7918 5678
rect 8002 5442 8238 5678
rect 8322 5442 8558 5678
rect 8642 5442 8878 5678
rect 5122 5122 5358 5358
rect 5442 5122 5678 5358
rect 5762 5122 5998 5358
rect 6082 5122 6318 5358
rect 6402 5122 6638 5358
rect 6722 5122 6958 5358
rect 7042 5122 7278 5358
rect 7362 5122 7598 5358
rect 7682 5122 7918 5358
rect 8002 5122 8238 5358
rect 8322 5122 8558 5358
rect 8642 5122 8878 5358
rect 226838 15882 227074 16118
rect 227158 15882 227394 16118
rect 227478 15882 227714 16118
rect 227798 15882 228034 16118
rect 228118 15882 228354 16118
rect 228438 15882 228674 16118
rect 228758 15882 228994 16118
rect 229078 15882 229314 16118
rect 229398 15882 229634 16118
rect 229718 15882 229954 16118
rect 230038 15882 230274 16118
rect 230358 15882 230594 16118
rect 226838 8642 227074 8878
rect 227158 8642 227394 8878
rect 227478 8642 227714 8878
rect 227798 8642 228034 8878
rect 228118 8642 228354 8878
rect 228438 8642 228674 8878
rect 228758 8642 228994 8878
rect 229078 8642 229314 8878
rect 229398 8642 229634 8878
rect 229718 8642 229954 8878
rect 230038 8642 230274 8878
rect 230358 8642 230594 8878
rect 226838 8322 227074 8558
rect 227158 8322 227394 8558
rect 227478 8322 227714 8558
rect 227798 8322 228034 8558
rect 228118 8322 228354 8558
rect 228438 8322 228674 8558
rect 228758 8322 228994 8558
rect 229078 8322 229314 8558
rect 229398 8322 229634 8558
rect 229718 8322 229954 8558
rect 230038 8322 230274 8558
rect 230358 8322 230594 8558
rect 226838 8002 227074 8238
rect 227158 8002 227394 8238
rect 227478 8002 227714 8238
rect 227798 8002 228034 8238
rect 228118 8002 228354 8238
rect 228438 8002 228674 8238
rect 228758 8002 228994 8238
rect 229078 8002 229314 8238
rect 229398 8002 229634 8238
rect 229718 8002 229954 8238
rect 230038 8002 230274 8238
rect 230358 8002 230594 8238
rect 226838 7682 227074 7918
rect 227158 7682 227394 7918
rect 227478 7682 227714 7918
rect 227798 7682 228034 7918
rect 228118 7682 228354 7918
rect 228438 7682 228674 7918
rect 228758 7682 228994 7918
rect 229078 7682 229314 7918
rect 229398 7682 229634 7918
rect 229718 7682 229954 7918
rect 230038 7682 230274 7918
rect 230358 7682 230594 7918
rect 226838 7362 227074 7598
rect 227158 7362 227394 7598
rect 227478 7362 227714 7598
rect 227798 7362 228034 7598
rect 228118 7362 228354 7598
rect 228438 7362 228674 7598
rect 228758 7362 228994 7598
rect 229078 7362 229314 7598
rect 229398 7362 229634 7598
rect 229718 7362 229954 7598
rect 230038 7362 230274 7598
rect 230358 7362 230594 7598
rect 226838 7042 227074 7278
rect 227158 7042 227394 7278
rect 227478 7042 227714 7278
rect 227798 7042 228034 7278
rect 228118 7042 228354 7278
rect 228438 7042 228674 7278
rect 228758 7042 228994 7278
rect 229078 7042 229314 7278
rect 229398 7042 229634 7278
rect 229718 7042 229954 7278
rect 230038 7042 230274 7278
rect 230358 7042 230594 7278
rect 226838 6722 227074 6958
rect 227158 6722 227394 6958
rect 227478 6722 227714 6958
rect 227798 6722 228034 6958
rect 228118 6722 228354 6958
rect 228438 6722 228674 6958
rect 228758 6722 228994 6958
rect 229078 6722 229314 6958
rect 229398 6722 229634 6958
rect 229718 6722 229954 6958
rect 230038 6722 230274 6958
rect 230358 6722 230594 6958
rect 226838 6402 227074 6638
rect 227158 6402 227394 6638
rect 227478 6402 227714 6638
rect 227798 6402 228034 6638
rect 228118 6402 228354 6638
rect 228438 6402 228674 6638
rect 228758 6402 228994 6638
rect 229078 6402 229314 6638
rect 229398 6402 229634 6638
rect 229718 6402 229954 6638
rect 230038 6402 230274 6638
rect 230358 6402 230594 6638
rect 226838 6082 227074 6318
rect 227158 6082 227394 6318
rect 227478 6082 227714 6318
rect 227798 6082 228034 6318
rect 228118 6082 228354 6318
rect 228438 6082 228674 6318
rect 228758 6082 228994 6318
rect 229078 6082 229314 6318
rect 229398 6082 229634 6318
rect 229718 6082 229954 6318
rect 230038 6082 230274 6318
rect 230358 6082 230594 6318
rect 226838 5762 227074 5998
rect 227158 5762 227394 5998
rect 227478 5762 227714 5998
rect 227798 5762 228034 5998
rect 228118 5762 228354 5998
rect 228438 5762 228674 5998
rect 228758 5762 228994 5998
rect 229078 5762 229314 5998
rect 229398 5762 229634 5998
rect 229718 5762 229954 5998
rect 230038 5762 230274 5998
rect 230358 5762 230594 5998
rect 226838 5442 227074 5678
rect 227158 5442 227394 5678
rect 227478 5442 227714 5678
rect 227798 5442 228034 5678
rect 228118 5442 228354 5678
rect 228438 5442 228674 5678
rect 228758 5442 228994 5678
rect 229078 5442 229314 5678
rect 229398 5442 229634 5678
rect 229718 5442 229954 5678
rect 230038 5442 230274 5678
rect 230358 5442 230594 5678
rect 226838 5122 227074 5358
rect 227158 5122 227394 5358
rect 227478 5122 227714 5358
rect 227798 5122 228034 5358
rect 228118 5122 228354 5358
rect 228438 5122 228674 5358
rect 228758 5122 228994 5358
rect 229078 5122 229314 5358
rect 229398 5122 229634 5358
rect 229718 5122 229954 5358
rect 230038 5122 230274 5358
rect 230358 5122 230594 5358
rect 231838 228682 232074 228918
rect 232158 228682 232394 228918
rect 232478 228682 232714 228918
rect 232798 228682 233034 228918
rect 233118 228682 233354 228918
rect 233438 228682 233674 228918
rect 233758 228682 233994 228918
rect 234078 228682 234314 228918
rect 234398 228682 234634 228918
rect 234718 228682 234954 228918
rect 235038 228682 235274 228918
rect 235358 228682 235594 228918
rect 231838 206282 232074 206518
rect 232158 206282 232394 206518
rect 232478 206282 232714 206518
rect 232798 206282 233034 206518
rect 233118 206282 233354 206518
rect 233438 206282 233674 206518
rect 233758 206282 233994 206518
rect 234078 206282 234314 206518
rect 234398 206282 234634 206518
rect 234718 206282 234954 206518
rect 235038 206282 235274 206518
rect 235358 206282 235594 206518
rect 231838 183882 232074 184118
rect 232158 183882 232394 184118
rect 232478 183882 232714 184118
rect 232798 183882 233034 184118
rect 233118 183882 233354 184118
rect 233438 183882 233674 184118
rect 233758 183882 233994 184118
rect 234078 183882 234314 184118
rect 234398 183882 234634 184118
rect 234718 183882 234954 184118
rect 235038 183882 235274 184118
rect 235358 183882 235594 184118
rect 231838 161482 232074 161718
rect 232158 161482 232394 161718
rect 232478 161482 232714 161718
rect 232798 161482 233034 161718
rect 233118 161482 233354 161718
rect 233438 161482 233674 161718
rect 233758 161482 233994 161718
rect 234078 161482 234314 161718
rect 234398 161482 234634 161718
rect 234718 161482 234954 161718
rect 235038 161482 235274 161718
rect 235358 161482 235594 161718
rect 231838 139082 232074 139318
rect 232158 139082 232394 139318
rect 232478 139082 232714 139318
rect 232798 139082 233034 139318
rect 233118 139082 233354 139318
rect 233438 139082 233674 139318
rect 233758 139082 233994 139318
rect 234078 139082 234314 139318
rect 234398 139082 234634 139318
rect 234718 139082 234954 139318
rect 235038 139082 235274 139318
rect 235358 139082 235594 139318
rect 231838 116682 232074 116918
rect 232158 116682 232394 116918
rect 232478 116682 232714 116918
rect 232798 116682 233034 116918
rect 233118 116682 233354 116918
rect 233438 116682 233674 116918
rect 233758 116682 233994 116918
rect 234078 116682 234314 116918
rect 234398 116682 234634 116918
rect 234718 116682 234954 116918
rect 235038 116682 235274 116918
rect 235358 116682 235594 116918
rect 231838 94282 232074 94518
rect 232158 94282 232394 94518
rect 232478 94282 232714 94518
rect 232798 94282 233034 94518
rect 233118 94282 233354 94518
rect 233438 94282 233674 94518
rect 233758 94282 233994 94518
rect 234078 94282 234314 94518
rect 234398 94282 234634 94518
rect 234718 94282 234954 94518
rect 235038 94282 235274 94518
rect 235358 94282 235594 94518
rect 231838 71882 232074 72118
rect 232158 71882 232394 72118
rect 232478 71882 232714 72118
rect 232798 71882 233034 72118
rect 233118 71882 233354 72118
rect 233438 71882 233674 72118
rect 233758 71882 233994 72118
rect 234078 71882 234314 72118
rect 234398 71882 234634 72118
rect 234718 71882 234954 72118
rect 235038 71882 235274 72118
rect 235358 71882 235594 72118
rect 231838 49482 232074 49718
rect 232158 49482 232394 49718
rect 232478 49482 232714 49718
rect 232798 49482 233034 49718
rect 233118 49482 233354 49718
rect 233438 49482 233674 49718
rect 233758 49482 233994 49718
rect 234078 49482 234314 49718
rect 234398 49482 234634 49718
rect 234718 49482 234954 49718
rect 235038 49482 235274 49718
rect 235358 49482 235594 49718
rect 231838 27082 232074 27318
rect 232158 27082 232394 27318
rect 232478 27082 232714 27318
rect 232798 27082 233034 27318
rect 233118 27082 233354 27318
rect 233438 27082 233674 27318
rect 233758 27082 233994 27318
rect 234078 27082 234314 27318
rect 234398 27082 234634 27318
rect 234718 27082 234954 27318
rect 235038 27082 235274 27318
rect 235358 27082 235594 27318
rect 122 3642 358 3878
rect 442 3642 678 3878
rect 762 3642 998 3878
rect 1082 3642 1318 3878
rect 1402 3642 1638 3878
rect 1722 3642 1958 3878
rect 2042 3642 2278 3878
rect 2362 3642 2598 3878
rect 2682 3642 2918 3878
rect 3002 3642 3238 3878
rect 3322 3642 3558 3878
rect 3642 3642 3878 3878
rect 122 3322 358 3558
rect 442 3322 678 3558
rect 762 3322 998 3558
rect 1082 3322 1318 3558
rect 1402 3322 1638 3558
rect 1722 3322 1958 3558
rect 2042 3322 2278 3558
rect 2362 3322 2598 3558
rect 2682 3322 2918 3558
rect 3002 3322 3238 3558
rect 3322 3322 3558 3558
rect 3642 3322 3878 3558
rect 122 3002 358 3238
rect 442 3002 678 3238
rect 762 3002 998 3238
rect 1082 3002 1318 3238
rect 1402 3002 1638 3238
rect 1722 3002 1958 3238
rect 2042 3002 2278 3238
rect 2362 3002 2598 3238
rect 2682 3002 2918 3238
rect 3002 3002 3238 3238
rect 3322 3002 3558 3238
rect 3642 3002 3878 3238
rect 122 2682 358 2918
rect 442 2682 678 2918
rect 762 2682 998 2918
rect 1082 2682 1318 2918
rect 1402 2682 1638 2918
rect 1722 2682 1958 2918
rect 2042 2682 2278 2918
rect 2362 2682 2598 2918
rect 2682 2682 2918 2918
rect 3002 2682 3238 2918
rect 3322 2682 3558 2918
rect 3642 2682 3878 2918
rect 122 2362 358 2598
rect 442 2362 678 2598
rect 762 2362 998 2598
rect 1082 2362 1318 2598
rect 1402 2362 1638 2598
rect 1722 2362 1958 2598
rect 2042 2362 2278 2598
rect 2362 2362 2598 2598
rect 2682 2362 2918 2598
rect 3002 2362 3238 2598
rect 3322 2362 3558 2598
rect 3642 2362 3878 2598
rect 122 2042 358 2278
rect 442 2042 678 2278
rect 762 2042 998 2278
rect 1082 2042 1318 2278
rect 1402 2042 1638 2278
rect 1722 2042 1958 2278
rect 2042 2042 2278 2278
rect 2362 2042 2598 2278
rect 2682 2042 2918 2278
rect 3002 2042 3238 2278
rect 3322 2042 3558 2278
rect 3642 2042 3878 2278
rect 122 1722 358 1958
rect 442 1722 678 1958
rect 762 1722 998 1958
rect 1082 1722 1318 1958
rect 1402 1722 1638 1958
rect 1722 1722 1958 1958
rect 2042 1722 2278 1958
rect 2362 1722 2598 1958
rect 2682 1722 2918 1958
rect 3002 1722 3238 1958
rect 3322 1722 3558 1958
rect 3642 1722 3878 1958
rect 122 1402 358 1638
rect 442 1402 678 1638
rect 762 1402 998 1638
rect 1082 1402 1318 1638
rect 1402 1402 1638 1638
rect 1722 1402 1958 1638
rect 2042 1402 2278 1638
rect 2362 1402 2598 1638
rect 2682 1402 2918 1638
rect 3002 1402 3238 1638
rect 3322 1402 3558 1638
rect 3642 1402 3878 1638
rect 122 1082 358 1318
rect 442 1082 678 1318
rect 762 1082 998 1318
rect 1082 1082 1318 1318
rect 1402 1082 1638 1318
rect 1722 1082 1958 1318
rect 2042 1082 2278 1318
rect 2362 1082 2598 1318
rect 2682 1082 2918 1318
rect 3002 1082 3238 1318
rect 3322 1082 3558 1318
rect 3642 1082 3878 1318
rect 122 762 358 998
rect 442 762 678 998
rect 762 762 998 998
rect 1082 762 1318 998
rect 1402 762 1638 998
rect 1722 762 1958 998
rect 2042 762 2278 998
rect 2362 762 2598 998
rect 2682 762 2918 998
rect 3002 762 3238 998
rect 3322 762 3558 998
rect 3642 762 3878 998
rect 122 442 358 678
rect 442 442 678 678
rect 762 442 998 678
rect 1082 442 1318 678
rect 1402 442 1638 678
rect 1722 442 1958 678
rect 2042 442 2278 678
rect 2362 442 2598 678
rect 2682 442 2918 678
rect 3002 442 3238 678
rect 3322 442 3558 678
rect 3642 442 3878 678
rect 122 122 358 358
rect 442 122 678 358
rect 762 122 998 358
rect 1082 122 1318 358
rect 1402 122 1638 358
rect 1722 122 1958 358
rect 2042 122 2278 358
rect 2362 122 2598 358
rect 2682 122 2918 358
rect 3002 122 3238 358
rect 3322 122 3558 358
rect 3642 122 3878 358
rect 231838 3642 232074 3878
rect 232158 3642 232394 3878
rect 232478 3642 232714 3878
rect 232798 3642 233034 3878
rect 233118 3642 233354 3878
rect 233438 3642 233674 3878
rect 233758 3642 233994 3878
rect 234078 3642 234314 3878
rect 234398 3642 234634 3878
rect 234718 3642 234954 3878
rect 235038 3642 235274 3878
rect 235358 3642 235594 3878
rect 231838 3322 232074 3558
rect 232158 3322 232394 3558
rect 232478 3322 232714 3558
rect 232798 3322 233034 3558
rect 233118 3322 233354 3558
rect 233438 3322 233674 3558
rect 233758 3322 233994 3558
rect 234078 3322 234314 3558
rect 234398 3322 234634 3558
rect 234718 3322 234954 3558
rect 235038 3322 235274 3558
rect 235358 3322 235594 3558
rect 231838 3002 232074 3238
rect 232158 3002 232394 3238
rect 232478 3002 232714 3238
rect 232798 3002 233034 3238
rect 233118 3002 233354 3238
rect 233438 3002 233674 3238
rect 233758 3002 233994 3238
rect 234078 3002 234314 3238
rect 234398 3002 234634 3238
rect 234718 3002 234954 3238
rect 235038 3002 235274 3238
rect 235358 3002 235594 3238
rect 231838 2682 232074 2918
rect 232158 2682 232394 2918
rect 232478 2682 232714 2918
rect 232798 2682 233034 2918
rect 233118 2682 233354 2918
rect 233438 2682 233674 2918
rect 233758 2682 233994 2918
rect 234078 2682 234314 2918
rect 234398 2682 234634 2918
rect 234718 2682 234954 2918
rect 235038 2682 235274 2918
rect 235358 2682 235594 2918
rect 231838 2362 232074 2598
rect 232158 2362 232394 2598
rect 232478 2362 232714 2598
rect 232798 2362 233034 2598
rect 233118 2362 233354 2598
rect 233438 2362 233674 2598
rect 233758 2362 233994 2598
rect 234078 2362 234314 2598
rect 234398 2362 234634 2598
rect 234718 2362 234954 2598
rect 235038 2362 235274 2598
rect 235358 2362 235594 2598
rect 231838 2042 232074 2278
rect 232158 2042 232394 2278
rect 232478 2042 232714 2278
rect 232798 2042 233034 2278
rect 233118 2042 233354 2278
rect 233438 2042 233674 2278
rect 233758 2042 233994 2278
rect 234078 2042 234314 2278
rect 234398 2042 234634 2278
rect 234718 2042 234954 2278
rect 235038 2042 235274 2278
rect 235358 2042 235594 2278
rect 231838 1722 232074 1958
rect 232158 1722 232394 1958
rect 232478 1722 232714 1958
rect 232798 1722 233034 1958
rect 233118 1722 233354 1958
rect 233438 1722 233674 1958
rect 233758 1722 233994 1958
rect 234078 1722 234314 1958
rect 234398 1722 234634 1958
rect 234718 1722 234954 1958
rect 235038 1722 235274 1958
rect 235358 1722 235594 1958
rect 231838 1402 232074 1638
rect 232158 1402 232394 1638
rect 232478 1402 232714 1638
rect 232798 1402 233034 1638
rect 233118 1402 233354 1638
rect 233438 1402 233674 1638
rect 233758 1402 233994 1638
rect 234078 1402 234314 1638
rect 234398 1402 234634 1638
rect 234718 1402 234954 1638
rect 235038 1402 235274 1638
rect 235358 1402 235594 1638
rect 231838 1082 232074 1318
rect 232158 1082 232394 1318
rect 232478 1082 232714 1318
rect 232798 1082 233034 1318
rect 233118 1082 233354 1318
rect 233438 1082 233674 1318
rect 233758 1082 233994 1318
rect 234078 1082 234314 1318
rect 234398 1082 234634 1318
rect 234718 1082 234954 1318
rect 235038 1082 235274 1318
rect 235358 1082 235594 1318
rect 231838 762 232074 998
rect 232158 762 232394 998
rect 232478 762 232714 998
rect 232798 762 233034 998
rect 233118 762 233354 998
rect 233438 762 233674 998
rect 233758 762 233994 998
rect 234078 762 234314 998
rect 234398 762 234634 998
rect 234718 762 234954 998
rect 235038 762 235274 998
rect 235358 762 235594 998
rect 231838 442 232074 678
rect 232158 442 232394 678
rect 232478 442 232714 678
rect 232798 442 233034 678
rect 233118 442 233354 678
rect 233438 442 233674 678
rect 233758 442 233994 678
rect 234078 442 234314 678
rect 234398 442 234634 678
rect 234718 442 234954 678
rect 235038 442 235274 678
rect 235358 442 235594 678
rect 231838 122 232074 358
rect 232158 122 232394 358
rect 232478 122 232714 358
rect 232798 122 233034 358
rect 233118 122 233354 358
rect 233438 122 233674 358
rect 233758 122 233994 358
rect 234078 122 234314 358
rect 234398 122 234634 358
rect 234718 122 234954 358
rect 235038 122 235274 358
rect 235358 122 235594 358
<< metal5 >>
rect 0 253078 235716 253200
rect 0 252842 122 253078
rect 358 252842 442 253078
rect 678 252842 762 253078
rect 998 252842 1082 253078
rect 1318 252842 1402 253078
rect 1638 252842 1722 253078
rect 1958 252842 2042 253078
rect 2278 252842 2362 253078
rect 2598 252842 2682 253078
rect 2918 252842 3002 253078
rect 3238 252842 3322 253078
rect 3558 252842 3642 253078
rect 3878 252842 231838 253078
rect 232074 252842 232158 253078
rect 232394 252842 232478 253078
rect 232714 252842 232798 253078
rect 233034 252842 233118 253078
rect 233354 252842 233438 253078
rect 233674 252842 233758 253078
rect 233994 252842 234078 253078
rect 234314 252842 234398 253078
rect 234634 252842 234718 253078
rect 234954 252842 235038 253078
rect 235274 252842 235358 253078
rect 235594 252842 235716 253078
rect 0 252758 235716 252842
rect 0 252522 122 252758
rect 358 252522 442 252758
rect 678 252522 762 252758
rect 998 252522 1082 252758
rect 1318 252522 1402 252758
rect 1638 252522 1722 252758
rect 1958 252522 2042 252758
rect 2278 252522 2362 252758
rect 2598 252522 2682 252758
rect 2918 252522 3002 252758
rect 3238 252522 3322 252758
rect 3558 252522 3642 252758
rect 3878 252522 231838 252758
rect 232074 252522 232158 252758
rect 232394 252522 232478 252758
rect 232714 252522 232798 252758
rect 233034 252522 233118 252758
rect 233354 252522 233438 252758
rect 233674 252522 233758 252758
rect 233994 252522 234078 252758
rect 234314 252522 234398 252758
rect 234634 252522 234718 252758
rect 234954 252522 235038 252758
rect 235274 252522 235358 252758
rect 235594 252522 235716 252758
rect 0 252438 235716 252522
rect 0 252202 122 252438
rect 358 252202 442 252438
rect 678 252202 762 252438
rect 998 252202 1082 252438
rect 1318 252202 1402 252438
rect 1638 252202 1722 252438
rect 1958 252202 2042 252438
rect 2278 252202 2362 252438
rect 2598 252202 2682 252438
rect 2918 252202 3002 252438
rect 3238 252202 3322 252438
rect 3558 252202 3642 252438
rect 3878 252202 231838 252438
rect 232074 252202 232158 252438
rect 232394 252202 232478 252438
rect 232714 252202 232798 252438
rect 233034 252202 233118 252438
rect 233354 252202 233438 252438
rect 233674 252202 233758 252438
rect 233994 252202 234078 252438
rect 234314 252202 234398 252438
rect 234634 252202 234718 252438
rect 234954 252202 235038 252438
rect 235274 252202 235358 252438
rect 235594 252202 235716 252438
rect 0 252118 235716 252202
rect 0 251882 122 252118
rect 358 251882 442 252118
rect 678 251882 762 252118
rect 998 251882 1082 252118
rect 1318 251882 1402 252118
rect 1638 251882 1722 252118
rect 1958 251882 2042 252118
rect 2278 251882 2362 252118
rect 2598 251882 2682 252118
rect 2918 251882 3002 252118
rect 3238 251882 3322 252118
rect 3558 251882 3642 252118
rect 3878 251882 231838 252118
rect 232074 251882 232158 252118
rect 232394 251882 232478 252118
rect 232714 251882 232798 252118
rect 233034 251882 233118 252118
rect 233354 251882 233438 252118
rect 233674 251882 233758 252118
rect 233994 251882 234078 252118
rect 234314 251882 234398 252118
rect 234634 251882 234718 252118
rect 234954 251882 235038 252118
rect 235274 251882 235358 252118
rect 235594 251882 235716 252118
rect 0 251798 235716 251882
rect 0 251562 122 251798
rect 358 251562 442 251798
rect 678 251562 762 251798
rect 998 251562 1082 251798
rect 1318 251562 1402 251798
rect 1638 251562 1722 251798
rect 1958 251562 2042 251798
rect 2278 251562 2362 251798
rect 2598 251562 2682 251798
rect 2918 251562 3002 251798
rect 3238 251562 3322 251798
rect 3558 251562 3642 251798
rect 3878 251562 231838 251798
rect 232074 251562 232158 251798
rect 232394 251562 232478 251798
rect 232714 251562 232798 251798
rect 233034 251562 233118 251798
rect 233354 251562 233438 251798
rect 233674 251562 233758 251798
rect 233994 251562 234078 251798
rect 234314 251562 234398 251798
rect 234634 251562 234718 251798
rect 234954 251562 235038 251798
rect 235274 251562 235358 251798
rect 235594 251562 235716 251798
rect 0 251478 235716 251562
rect 0 251242 122 251478
rect 358 251242 442 251478
rect 678 251242 762 251478
rect 998 251242 1082 251478
rect 1318 251242 1402 251478
rect 1638 251242 1722 251478
rect 1958 251242 2042 251478
rect 2278 251242 2362 251478
rect 2598 251242 2682 251478
rect 2918 251242 3002 251478
rect 3238 251242 3322 251478
rect 3558 251242 3642 251478
rect 3878 251242 231838 251478
rect 232074 251242 232158 251478
rect 232394 251242 232478 251478
rect 232714 251242 232798 251478
rect 233034 251242 233118 251478
rect 233354 251242 233438 251478
rect 233674 251242 233758 251478
rect 233994 251242 234078 251478
rect 234314 251242 234398 251478
rect 234634 251242 234718 251478
rect 234954 251242 235038 251478
rect 235274 251242 235358 251478
rect 235594 251242 235716 251478
rect 0 251158 235716 251242
rect 0 250922 122 251158
rect 358 250922 442 251158
rect 678 250922 762 251158
rect 998 250922 1082 251158
rect 1318 250922 1402 251158
rect 1638 250922 1722 251158
rect 1958 250922 2042 251158
rect 2278 250922 2362 251158
rect 2598 250922 2682 251158
rect 2918 250922 3002 251158
rect 3238 250922 3322 251158
rect 3558 250922 3642 251158
rect 3878 250922 231838 251158
rect 232074 250922 232158 251158
rect 232394 250922 232478 251158
rect 232714 250922 232798 251158
rect 233034 250922 233118 251158
rect 233354 250922 233438 251158
rect 233674 250922 233758 251158
rect 233994 250922 234078 251158
rect 234314 250922 234398 251158
rect 234634 250922 234718 251158
rect 234954 250922 235038 251158
rect 235274 250922 235358 251158
rect 235594 250922 235716 251158
rect 0 250838 235716 250922
rect 0 250602 122 250838
rect 358 250602 442 250838
rect 678 250602 762 250838
rect 998 250602 1082 250838
rect 1318 250602 1402 250838
rect 1638 250602 1722 250838
rect 1958 250602 2042 250838
rect 2278 250602 2362 250838
rect 2598 250602 2682 250838
rect 2918 250602 3002 250838
rect 3238 250602 3322 250838
rect 3558 250602 3642 250838
rect 3878 250602 231838 250838
rect 232074 250602 232158 250838
rect 232394 250602 232478 250838
rect 232714 250602 232798 250838
rect 233034 250602 233118 250838
rect 233354 250602 233438 250838
rect 233674 250602 233758 250838
rect 233994 250602 234078 250838
rect 234314 250602 234398 250838
rect 234634 250602 234718 250838
rect 234954 250602 235038 250838
rect 235274 250602 235358 250838
rect 235594 250602 235716 250838
rect 0 250518 235716 250602
rect 0 250282 122 250518
rect 358 250282 442 250518
rect 678 250282 762 250518
rect 998 250282 1082 250518
rect 1318 250282 1402 250518
rect 1638 250282 1722 250518
rect 1958 250282 2042 250518
rect 2278 250282 2362 250518
rect 2598 250282 2682 250518
rect 2918 250282 3002 250518
rect 3238 250282 3322 250518
rect 3558 250282 3642 250518
rect 3878 250282 231838 250518
rect 232074 250282 232158 250518
rect 232394 250282 232478 250518
rect 232714 250282 232798 250518
rect 233034 250282 233118 250518
rect 233354 250282 233438 250518
rect 233674 250282 233758 250518
rect 233994 250282 234078 250518
rect 234314 250282 234398 250518
rect 234634 250282 234718 250518
rect 234954 250282 235038 250518
rect 235274 250282 235358 250518
rect 235594 250282 235716 250518
rect 0 250198 235716 250282
rect 0 249962 122 250198
rect 358 249962 442 250198
rect 678 249962 762 250198
rect 998 249962 1082 250198
rect 1318 249962 1402 250198
rect 1638 249962 1722 250198
rect 1958 249962 2042 250198
rect 2278 249962 2362 250198
rect 2598 249962 2682 250198
rect 2918 249962 3002 250198
rect 3238 249962 3322 250198
rect 3558 249962 3642 250198
rect 3878 249962 231838 250198
rect 232074 249962 232158 250198
rect 232394 249962 232478 250198
rect 232714 249962 232798 250198
rect 233034 249962 233118 250198
rect 233354 249962 233438 250198
rect 233674 249962 233758 250198
rect 233994 249962 234078 250198
rect 234314 249962 234398 250198
rect 234634 249962 234718 250198
rect 234954 249962 235038 250198
rect 235274 249962 235358 250198
rect 235594 249962 235716 250198
rect 0 249878 235716 249962
rect 0 249642 122 249878
rect 358 249642 442 249878
rect 678 249642 762 249878
rect 998 249642 1082 249878
rect 1318 249642 1402 249878
rect 1638 249642 1722 249878
rect 1958 249642 2042 249878
rect 2278 249642 2362 249878
rect 2598 249642 2682 249878
rect 2918 249642 3002 249878
rect 3238 249642 3322 249878
rect 3558 249642 3642 249878
rect 3878 249642 231838 249878
rect 232074 249642 232158 249878
rect 232394 249642 232478 249878
rect 232714 249642 232798 249878
rect 233034 249642 233118 249878
rect 233354 249642 233438 249878
rect 233674 249642 233758 249878
rect 233994 249642 234078 249878
rect 234314 249642 234398 249878
rect 234634 249642 234718 249878
rect 234954 249642 235038 249878
rect 235274 249642 235358 249878
rect 235594 249642 235716 249878
rect 0 249558 235716 249642
rect 0 249322 122 249558
rect 358 249322 442 249558
rect 678 249322 762 249558
rect 998 249322 1082 249558
rect 1318 249322 1402 249558
rect 1638 249322 1722 249558
rect 1958 249322 2042 249558
rect 2278 249322 2362 249558
rect 2598 249322 2682 249558
rect 2918 249322 3002 249558
rect 3238 249322 3322 249558
rect 3558 249322 3642 249558
rect 3878 249322 231838 249558
rect 232074 249322 232158 249558
rect 232394 249322 232478 249558
rect 232714 249322 232798 249558
rect 233034 249322 233118 249558
rect 233354 249322 233438 249558
rect 233674 249322 233758 249558
rect 233994 249322 234078 249558
rect 234314 249322 234398 249558
rect 234634 249322 234718 249558
rect 234954 249322 235038 249558
rect 235274 249322 235358 249558
rect 235594 249322 235716 249558
rect 0 249200 235716 249322
rect 5000 248078 230716 248200
rect 5000 247842 5122 248078
rect 5358 247842 5442 248078
rect 5678 247842 5762 248078
rect 5998 247842 6082 248078
rect 6318 247842 6402 248078
rect 6638 247842 6722 248078
rect 6958 247842 7042 248078
rect 7278 247842 7362 248078
rect 7598 247842 7682 248078
rect 7918 247842 8002 248078
rect 8238 247842 8322 248078
rect 8558 247842 8642 248078
rect 8878 247842 226838 248078
rect 227074 247842 227158 248078
rect 227394 247842 227478 248078
rect 227714 247842 227798 248078
rect 228034 247842 228118 248078
rect 228354 247842 228438 248078
rect 228674 247842 228758 248078
rect 228994 247842 229078 248078
rect 229314 247842 229398 248078
rect 229634 247842 229718 248078
rect 229954 247842 230038 248078
rect 230274 247842 230358 248078
rect 230594 247842 230716 248078
rect 5000 247758 230716 247842
rect 5000 247522 5122 247758
rect 5358 247522 5442 247758
rect 5678 247522 5762 247758
rect 5998 247522 6082 247758
rect 6318 247522 6402 247758
rect 6638 247522 6722 247758
rect 6958 247522 7042 247758
rect 7278 247522 7362 247758
rect 7598 247522 7682 247758
rect 7918 247522 8002 247758
rect 8238 247522 8322 247758
rect 8558 247522 8642 247758
rect 8878 247522 226838 247758
rect 227074 247522 227158 247758
rect 227394 247522 227478 247758
rect 227714 247522 227798 247758
rect 228034 247522 228118 247758
rect 228354 247522 228438 247758
rect 228674 247522 228758 247758
rect 228994 247522 229078 247758
rect 229314 247522 229398 247758
rect 229634 247522 229718 247758
rect 229954 247522 230038 247758
rect 230274 247522 230358 247758
rect 230594 247522 230716 247758
rect 5000 247438 230716 247522
rect 5000 247202 5122 247438
rect 5358 247202 5442 247438
rect 5678 247202 5762 247438
rect 5998 247202 6082 247438
rect 6318 247202 6402 247438
rect 6638 247202 6722 247438
rect 6958 247202 7042 247438
rect 7278 247202 7362 247438
rect 7598 247202 7682 247438
rect 7918 247202 8002 247438
rect 8238 247202 8322 247438
rect 8558 247202 8642 247438
rect 8878 247202 226838 247438
rect 227074 247202 227158 247438
rect 227394 247202 227478 247438
rect 227714 247202 227798 247438
rect 228034 247202 228118 247438
rect 228354 247202 228438 247438
rect 228674 247202 228758 247438
rect 228994 247202 229078 247438
rect 229314 247202 229398 247438
rect 229634 247202 229718 247438
rect 229954 247202 230038 247438
rect 230274 247202 230358 247438
rect 230594 247202 230716 247438
rect 5000 247118 230716 247202
rect 5000 246882 5122 247118
rect 5358 246882 5442 247118
rect 5678 246882 5762 247118
rect 5998 246882 6082 247118
rect 6318 246882 6402 247118
rect 6638 246882 6722 247118
rect 6958 246882 7042 247118
rect 7278 246882 7362 247118
rect 7598 246882 7682 247118
rect 7918 246882 8002 247118
rect 8238 246882 8322 247118
rect 8558 246882 8642 247118
rect 8878 246882 226838 247118
rect 227074 246882 227158 247118
rect 227394 246882 227478 247118
rect 227714 246882 227798 247118
rect 228034 246882 228118 247118
rect 228354 246882 228438 247118
rect 228674 246882 228758 247118
rect 228994 246882 229078 247118
rect 229314 246882 229398 247118
rect 229634 246882 229718 247118
rect 229954 246882 230038 247118
rect 230274 246882 230358 247118
rect 230594 246882 230716 247118
rect 5000 246798 230716 246882
rect 5000 246562 5122 246798
rect 5358 246562 5442 246798
rect 5678 246562 5762 246798
rect 5998 246562 6082 246798
rect 6318 246562 6402 246798
rect 6638 246562 6722 246798
rect 6958 246562 7042 246798
rect 7278 246562 7362 246798
rect 7598 246562 7682 246798
rect 7918 246562 8002 246798
rect 8238 246562 8322 246798
rect 8558 246562 8642 246798
rect 8878 246562 226838 246798
rect 227074 246562 227158 246798
rect 227394 246562 227478 246798
rect 227714 246562 227798 246798
rect 228034 246562 228118 246798
rect 228354 246562 228438 246798
rect 228674 246562 228758 246798
rect 228994 246562 229078 246798
rect 229314 246562 229398 246798
rect 229634 246562 229718 246798
rect 229954 246562 230038 246798
rect 230274 246562 230358 246798
rect 230594 246562 230716 246798
rect 5000 246478 230716 246562
rect 5000 246242 5122 246478
rect 5358 246242 5442 246478
rect 5678 246242 5762 246478
rect 5998 246242 6082 246478
rect 6318 246242 6402 246478
rect 6638 246242 6722 246478
rect 6958 246242 7042 246478
rect 7278 246242 7362 246478
rect 7598 246242 7682 246478
rect 7918 246242 8002 246478
rect 8238 246242 8322 246478
rect 8558 246242 8642 246478
rect 8878 246242 226838 246478
rect 227074 246242 227158 246478
rect 227394 246242 227478 246478
rect 227714 246242 227798 246478
rect 228034 246242 228118 246478
rect 228354 246242 228438 246478
rect 228674 246242 228758 246478
rect 228994 246242 229078 246478
rect 229314 246242 229398 246478
rect 229634 246242 229718 246478
rect 229954 246242 230038 246478
rect 230274 246242 230358 246478
rect 230594 246242 230716 246478
rect 5000 246158 230716 246242
rect 5000 245922 5122 246158
rect 5358 245922 5442 246158
rect 5678 245922 5762 246158
rect 5998 245922 6082 246158
rect 6318 245922 6402 246158
rect 6638 245922 6722 246158
rect 6958 245922 7042 246158
rect 7278 245922 7362 246158
rect 7598 245922 7682 246158
rect 7918 245922 8002 246158
rect 8238 245922 8322 246158
rect 8558 245922 8642 246158
rect 8878 245922 226838 246158
rect 227074 245922 227158 246158
rect 227394 245922 227478 246158
rect 227714 245922 227798 246158
rect 228034 245922 228118 246158
rect 228354 245922 228438 246158
rect 228674 245922 228758 246158
rect 228994 245922 229078 246158
rect 229314 245922 229398 246158
rect 229634 245922 229718 246158
rect 229954 245922 230038 246158
rect 230274 245922 230358 246158
rect 230594 245922 230716 246158
rect 5000 245838 230716 245922
rect 5000 245602 5122 245838
rect 5358 245602 5442 245838
rect 5678 245602 5762 245838
rect 5998 245602 6082 245838
rect 6318 245602 6402 245838
rect 6638 245602 6722 245838
rect 6958 245602 7042 245838
rect 7278 245602 7362 245838
rect 7598 245602 7682 245838
rect 7918 245602 8002 245838
rect 8238 245602 8322 245838
rect 8558 245602 8642 245838
rect 8878 245602 226838 245838
rect 227074 245602 227158 245838
rect 227394 245602 227478 245838
rect 227714 245602 227798 245838
rect 228034 245602 228118 245838
rect 228354 245602 228438 245838
rect 228674 245602 228758 245838
rect 228994 245602 229078 245838
rect 229314 245602 229398 245838
rect 229634 245602 229718 245838
rect 229954 245602 230038 245838
rect 230274 245602 230358 245838
rect 230594 245602 230716 245838
rect 5000 245518 230716 245602
rect 5000 245282 5122 245518
rect 5358 245282 5442 245518
rect 5678 245282 5762 245518
rect 5998 245282 6082 245518
rect 6318 245282 6402 245518
rect 6638 245282 6722 245518
rect 6958 245282 7042 245518
rect 7278 245282 7362 245518
rect 7598 245282 7682 245518
rect 7918 245282 8002 245518
rect 8238 245282 8322 245518
rect 8558 245282 8642 245518
rect 8878 245282 226838 245518
rect 227074 245282 227158 245518
rect 227394 245282 227478 245518
rect 227714 245282 227798 245518
rect 228034 245282 228118 245518
rect 228354 245282 228438 245518
rect 228674 245282 228758 245518
rect 228994 245282 229078 245518
rect 229314 245282 229398 245518
rect 229634 245282 229718 245518
rect 229954 245282 230038 245518
rect 230274 245282 230358 245518
rect 230594 245282 230716 245518
rect 5000 245198 230716 245282
rect 5000 244962 5122 245198
rect 5358 244962 5442 245198
rect 5678 244962 5762 245198
rect 5998 244962 6082 245198
rect 6318 244962 6402 245198
rect 6638 244962 6722 245198
rect 6958 244962 7042 245198
rect 7278 244962 7362 245198
rect 7598 244962 7682 245198
rect 7918 244962 8002 245198
rect 8238 244962 8322 245198
rect 8558 244962 8642 245198
rect 8878 244962 226838 245198
rect 227074 244962 227158 245198
rect 227394 244962 227478 245198
rect 227714 244962 227798 245198
rect 228034 244962 228118 245198
rect 228354 244962 228438 245198
rect 228674 244962 228758 245198
rect 228994 244962 229078 245198
rect 229314 244962 229398 245198
rect 229634 244962 229718 245198
rect 229954 244962 230038 245198
rect 230274 244962 230358 245198
rect 230594 244962 230716 245198
rect 5000 244878 230716 244962
rect 5000 244642 5122 244878
rect 5358 244642 5442 244878
rect 5678 244642 5762 244878
rect 5998 244642 6082 244878
rect 6318 244642 6402 244878
rect 6638 244642 6722 244878
rect 6958 244642 7042 244878
rect 7278 244642 7362 244878
rect 7598 244642 7682 244878
rect 7918 244642 8002 244878
rect 8238 244642 8322 244878
rect 8558 244642 8642 244878
rect 8878 244642 226838 244878
rect 227074 244642 227158 244878
rect 227394 244642 227478 244878
rect 227714 244642 227798 244878
rect 228034 244642 228118 244878
rect 228354 244642 228438 244878
rect 228674 244642 228758 244878
rect 228994 244642 229078 244878
rect 229314 244642 229398 244878
rect 229634 244642 229718 244878
rect 229954 244642 230038 244878
rect 230274 244642 230358 244878
rect 230594 244642 230716 244878
rect 5000 244558 230716 244642
rect 5000 244322 5122 244558
rect 5358 244322 5442 244558
rect 5678 244322 5762 244558
rect 5998 244322 6082 244558
rect 6318 244322 6402 244558
rect 6638 244322 6722 244558
rect 6958 244322 7042 244558
rect 7278 244322 7362 244558
rect 7598 244322 7682 244558
rect 7918 244322 8002 244558
rect 8238 244322 8322 244558
rect 8558 244322 8642 244558
rect 8878 244322 226838 244558
rect 227074 244322 227158 244558
rect 227394 244322 227478 244558
rect 227714 244322 227798 244558
rect 228034 244322 228118 244558
rect 228354 244322 228438 244558
rect 228674 244322 228758 244558
rect 228994 244322 229078 244558
rect 229314 244322 229398 244558
rect 229634 244322 229718 244558
rect 229954 244322 230038 244558
rect 230274 244322 230358 244558
rect 230594 244322 230716 244558
rect 5000 244200 230716 244322
rect 0 240118 235716 240160
rect 0 239882 5122 240118
rect 5358 239882 5442 240118
rect 5678 239882 5762 240118
rect 5998 239882 6082 240118
rect 6318 239882 6402 240118
rect 6638 239882 6722 240118
rect 6958 239882 7042 240118
rect 7278 239882 7362 240118
rect 7598 239882 7682 240118
rect 7918 239882 8002 240118
rect 8238 239882 8322 240118
rect 8558 239882 8642 240118
rect 8878 239882 226838 240118
rect 227074 239882 227158 240118
rect 227394 239882 227478 240118
rect 227714 239882 227798 240118
rect 228034 239882 228118 240118
rect 228354 239882 228438 240118
rect 228674 239882 228758 240118
rect 228994 239882 229078 240118
rect 229314 239882 229398 240118
rect 229634 239882 229718 240118
rect 229954 239882 230038 240118
rect 230274 239882 230358 240118
rect 230594 239882 235716 240118
rect 0 239840 235716 239882
rect 0 228918 235716 228960
rect 0 228682 122 228918
rect 358 228682 442 228918
rect 678 228682 762 228918
rect 998 228682 1082 228918
rect 1318 228682 1402 228918
rect 1638 228682 1722 228918
rect 1958 228682 2042 228918
rect 2278 228682 2362 228918
rect 2598 228682 2682 228918
rect 2918 228682 3002 228918
rect 3238 228682 3322 228918
rect 3558 228682 3642 228918
rect 3878 228682 29927 228918
rect 30163 228682 71882 228918
rect 72118 228682 114215 228918
rect 114451 228682 155882 228918
rect 156118 228682 198215 228918
rect 198451 228682 231838 228918
rect 232074 228682 232158 228918
rect 232394 228682 232478 228918
rect 232714 228682 232798 228918
rect 233034 228682 233118 228918
rect 233354 228682 233438 228918
rect 233674 228682 233758 228918
rect 233994 228682 234078 228918
rect 234314 228682 234398 228918
rect 234634 228682 234718 228918
rect 234954 228682 235038 228918
rect 235274 228682 235358 228918
rect 235594 228682 235716 228918
rect 0 228640 235716 228682
rect 0 217718 235716 217760
rect 0 217482 5122 217718
rect 5358 217482 5442 217718
rect 5678 217482 5762 217718
rect 5998 217482 6082 217718
rect 6318 217482 6402 217718
rect 6638 217482 6722 217718
rect 6958 217482 7042 217718
rect 7278 217482 7362 217718
rect 7598 217482 7682 217718
rect 7918 217482 8002 217718
rect 8238 217482 8322 217718
rect 8558 217482 8642 217718
rect 8878 217482 25261 217718
rect 25497 217482 66882 217718
rect 67118 217482 109549 217718
rect 109785 217482 150882 217718
rect 151118 217482 193549 217718
rect 193785 217482 226838 217718
rect 227074 217482 227158 217718
rect 227394 217482 227478 217718
rect 227714 217482 227798 217718
rect 228034 217482 228118 217718
rect 228354 217482 228438 217718
rect 228674 217482 228758 217718
rect 228994 217482 229078 217718
rect 229314 217482 229398 217718
rect 229634 217482 229718 217718
rect 229954 217482 230038 217718
rect 230274 217482 230358 217718
rect 230594 217482 235716 217718
rect 0 217440 235716 217482
rect 0 206518 235716 206560
rect 0 206282 122 206518
rect 358 206282 442 206518
rect 678 206282 762 206518
rect 998 206282 1082 206518
rect 1318 206282 1402 206518
rect 1638 206282 1722 206518
rect 1958 206282 2042 206518
rect 2278 206282 2362 206518
rect 2598 206282 2682 206518
rect 2918 206282 3002 206518
rect 3238 206282 3322 206518
rect 3558 206282 3642 206518
rect 3878 206282 231838 206518
rect 232074 206282 232158 206518
rect 232394 206282 232478 206518
rect 232714 206282 232798 206518
rect 233034 206282 233118 206518
rect 233354 206282 233438 206518
rect 233674 206282 233758 206518
rect 233994 206282 234078 206518
rect 234314 206282 234398 206518
rect 234634 206282 234718 206518
rect 234954 206282 235038 206518
rect 235274 206282 235358 206518
rect 235594 206282 235716 206518
rect 0 206240 235716 206282
rect 0 195318 235716 195360
rect 0 195082 5122 195318
rect 5358 195082 5442 195318
rect 5678 195082 5762 195318
rect 5998 195082 6082 195318
rect 6318 195082 6402 195318
rect 6638 195082 6722 195318
rect 6958 195082 7042 195318
rect 7278 195082 7362 195318
rect 7598 195082 7682 195318
rect 7918 195082 8002 195318
rect 8238 195082 8322 195318
rect 8558 195082 8642 195318
rect 8878 195082 226838 195318
rect 227074 195082 227158 195318
rect 227394 195082 227478 195318
rect 227714 195082 227798 195318
rect 228034 195082 228118 195318
rect 228354 195082 228438 195318
rect 228674 195082 228758 195318
rect 228994 195082 229078 195318
rect 229314 195082 229398 195318
rect 229634 195082 229718 195318
rect 229954 195082 230038 195318
rect 230274 195082 230358 195318
rect 230594 195082 235716 195318
rect 0 195040 235716 195082
rect 193828 190842 210156 190884
rect 193828 190606 193870 190842
rect 194106 190606 209878 190842
rect 210114 190606 210156 190842
rect 193828 190564 210156 190606
rect 0 184118 235716 184160
rect 0 183882 122 184118
rect 358 183882 442 184118
rect 678 183882 762 184118
rect 998 183882 1082 184118
rect 1318 183882 1402 184118
rect 1638 183882 1722 184118
rect 1958 183882 2042 184118
rect 2278 183882 2362 184118
rect 2598 183882 2682 184118
rect 2918 183882 3002 184118
rect 3238 183882 3322 184118
rect 3558 183882 3642 184118
rect 3878 183882 32215 184118
rect 32451 183882 75506 184118
rect 75742 183882 116215 184118
rect 116451 183882 159506 184118
rect 159742 183882 200215 184118
rect 200451 183882 231838 184118
rect 232074 183882 232158 184118
rect 232394 183882 232478 184118
rect 232714 183882 232798 184118
rect 233034 183882 233118 184118
rect 233354 183882 233438 184118
rect 233674 183882 233758 184118
rect 233994 183882 234078 184118
rect 234314 183882 234398 184118
rect 234634 183882 234718 184118
rect 234954 183882 235038 184118
rect 235274 183882 235358 184118
rect 235594 183882 235716 184118
rect 0 183840 235716 183882
rect 26388 178602 42164 178644
rect 26388 178366 26430 178602
rect 26666 178366 41886 178602
rect 42122 178366 42164 178602
rect 26388 178324 42164 178366
rect 0 172918 235716 172960
rect 0 172682 5122 172918
rect 5358 172682 5442 172918
rect 5678 172682 5762 172918
rect 5998 172682 6082 172918
rect 6318 172682 6402 172918
rect 6638 172682 6722 172918
rect 6958 172682 7042 172918
rect 7278 172682 7362 172918
rect 7598 172682 7682 172918
rect 7918 172682 8002 172918
rect 8238 172682 8322 172918
rect 8558 172682 8642 172918
rect 8878 172682 29549 172918
rect 29785 172682 60146 172918
rect 60382 172682 113549 172918
rect 113785 172682 144146 172918
rect 144382 172682 197549 172918
rect 197785 172682 226838 172918
rect 227074 172682 227158 172918
rect 227394 172682 227478 172918
rect 227714 172682 227798 172918
rect 228034 172682 228118 172918
rect 228354 172682 228438 172918
rect 228674 172682 228758 172918
rect 228994 172682 229078 172918
rect 229314 172682 229398 172918
rect 229634 172682 229718 172918
rect 229954 172682 230038 172918
rect 230274 172682 230358 172918
rect 230594 172682 235716 172918
rect 0 172640 235716 172682
rect 139364 165002 212732 165044
rect 139364 164766 139406 165002
rect 139642 164766 212454 165002
rect 212690 164766 212732 165002
rect 139364 164724 212732 164766
rect 26388 163642 41980 163684
rect 26388 163406 26430 163642
rect 26666 163406 41702 163642
rect 41938 163406 41980 163642
rect 26388 163364 41980 163406
rect 0 161718 235716 161760
rect 0 161482 122 161718
rect 358 161482 442 161718
rect 678 161482 762 161718
rect 998 161482 1082 161718
rect 1318 161482 1402 161718
rect 1638 161482 1722 161718
rect 1958 161482 2042 161718
rect 2278 161482 2362 161718
rect 2598 161482 2682 161718
rect 2918 161482 3002 161718
rect 3238 161482 3322 161718
rect 3558 161482 3642 161718
rect 3878 161482 32215 161718
rect 32451 161482 75506 161718
rect 75742 161482 116215 161718
rect 116451 161482 159506 161718
rect 159742 161482 200215 161718
rect 200451 161482 231838 161718
rect 232074 161482 232158 161718
rect 232394 161482 232478 161718
rect 232714 161482 232798 161718
rect 233034 161482 233118 161718
rect 233354 161482 233438 161718
rect 233674 161482 233758 161718
rect 233994 161482 234078 161718
rect 234314 161482 234398 161718
rect 234634 161482 234718 161718
rect 234954 161482 235038 161718
rect 235274 161482 235358 161718
rect 235594 161482 235716 161718
rect 0 161440 235716 161482
rect 0 150518 235716 150560
rect 0 150282 5122 150518
rect 5358 150282 5442 150518
rect 5678 150282 5762 150518
rect 5998 150282 6082 150518
rect 6318 150282 6402 150518
rect 6638 150282 6722 150518
rect 6958 150282 7042 150518
rect 7278 150282 7362 150518
rect 7598 150282 7682 150518
rect 7918 150282 8002 150518
rect 8238 150282 8322 150518
rect 8558 150282 8642 150518
rect 8878 150282 226838 150518
rect 227074 150282 227158 150518
rect 227394 150282 227478 150518
rect 227714 150282 227798 150518
rect 228034 150282 228118 150518
rect 228354 150282 228438 150518
rect 228674 150282 228758 150518
rect 228994 150282 229078 150518
rect 229314 150282 229398 150518
rect 229634 150282 229718 150518
rect 229954 150282 230038 150518
rect 230274 150282 230358 150518
rect 230594 150282 235716 150518
rect 0 150240 235716 150282
rect 0 139318 235716 139360
rect 0 139082 122 139318
rect 358 139082 442 139318
rect 678 139082 762 139318
rect 998 139082 1082 139318
rect 1318 139082 1402 139318
rect 1638 139082 1722 139318
rect 1958 139082 2042 139318
rect 2278 139082 2362 139318
rect 2598 139082 2682 139318
rect 2918 139082 3002 139318
rect 3238 139082 3322 139318
rect 3558 139082 3642 139318
rect 3878 139082 231838 139318
rect 232074 139082 232158 139318
rect 232394 139082 232478 139318
rect 232714 139082 232798 139318
rect 233034 139082 233118 139318
rect 233354 139082 233438 139318
rect 233674 139082 233758 139318
rect 233994 139082 234078 139318
rect 234314 139082 234398 139318
rect 234634 139082 234718 139318
rect 234954 139082 235038 139318
rect 235274 139082 235358 139318
rect 235594 139082 235716 139318
rect 0 139040 235716 139082
rect 0 128118 235716 128160
rect 0 127882 5122 128118
rect 5358 127882 5442 128118
rect 5678 127882 5762 128118
rect 5998 127882 6082 128118
rect 6318 127882 6402 128118
rect 6638 127882 6722 128118
rect 6958 127882 7042 128118
rect 7278 127882 7362 128118
rect 7598 127882 7682 128118
rect 7918 127882 8002 128118
rect 8238 127882 8322 128118
rect 8558 127882 8642 128118
rect 8878 127882 25549 128118
rect 25785 127882 66882 128118
rect 67118 127882 109549 128118
rect 109785 127882 150882 128118
rect 151118 127882 193549 128118
rect 193785 127882 226838 128118
rect 227074 127882 227158 128118
rect 227394 127882 227478 128118
rect 227714 127882 227798 128118
rect 228034 127882 228118 128118
rect 228354 127882 228438 128118
rect 228674 127882 228758 128118
rect 228994 127882 229078 128118
rect 229314 127882 229398 128118
rect 229634 127882 229718 128118
rect 229954 127882 230038 128118
rect 230274 127882 230358 128118
rect 230594 127882 235716 128118
rect 0 127840 235716 127882
rect 0 116918 235716 116960
rect 0 116682 122 116918
rect 358 116682 442 116918
rect 678 116682 762 116918
rect 998 116682 1082 116918
rect 1318 116682 1402 116918
rect 1638 116682 1722 116918
rect 1958 116682 2042 116918
rect 2278 116682 2362 116918
rect 2598 116682 2682 116918
rect 2918 116682 3002 116918
rect 3238 116682 3322 116918
rect 3558 116682 3642 116918
rect 3878 116682 30215 116918
rect 30451 116682 114215 116918
rect 114451 116682 198215 116918
rect 198451 116682 231838 116918
rect 232074 116682 232158 116918
rect 232394 116682 232478 116918
rect 232714 116682 232798 116918
rect 233034 116682 233118 116918
rect 233354 116682 233438 116918
rect 233674 116682 233758 116918
rect 233994 116682 234078 116918
rect 234314 116682 234398 116918
rect 234634 116682 234718 116918
rect 234954 116682 235038 116918
rect 235274 116682 235358 116918
rect 235594 116682 235716 116918
rect 0 116640 235716 116682
rect 61900 111282 134164 111324
rect 61900 111046 61942 111282
rect 62178 111046 108310 111282
rect 108546 111046 133886 111282
rect 134122 111046 134164 111282
rect 61900 111004 134164 111046
rect 0 105718 235716 105760
rect 0 105482 5122 105718
rect 5358 105482 5442 105718
rect 5678 105482 5762 105718
rect 5998 105482 6082 105718
rect 6318 105482 6402 105718
rect 6638 105482 6722 105718
rect 6958 105482 7042 105718
rect 7278 105482 7362 105718
rect 7598 105482 7682 105718
rect 7918 105482 8002 105718
rect 8238 105482 8322 105718
rect 8558 105482 8642 105718
rect 8878 105482 226838 105718
rect 227074 105482 227158 105718
rect 227394 105482 227478 105718
rect 227714 105482 227798 105718
rect 228034 105482 228118 105718
rect 228354 105482 228438 105718
rect 228674 105482 228758 105718
rect 228994 105482 229078 105718
rect 229314 105482 229398 105718
rect 229634 105482 229718 105718
rect 229954 105482 230038 105718
rect 230274 105482 230358 105718
rect 230594 105482 235716 105718
rect 0 105440 235716 105482
rect 193644 97002 209972 97044
rect 193644 96766 193686 97002
rect 193922 96766 209694 97002
rect 209930 96766 209972 97002
rect 193644 96724 209972 96766
rect 0 94518 235716 94560
rect 0 94282 122 94518
rect 358 94282 442 94518
rect 678 94282 762 94518
rect 998 94282 1082 94518
rect 1318 94282 1402 94518
rect 1638 94282 1722 94518
rect 1958 94282 2042 94518
rect 2278 94282 2362 94518
rect 2598 94282 2682 94518
rect 2918 94282 3002 94518
rect 3238 94282 3322 94518
rect 3558 94282 3642 94518
rect 3878 94282 32215 94518
rect 32451 94282 75506 94518
rect 75742 94282 116215 94518
rect 116451 94282 159506 94518
rect 159742 94282 200215 94518
rect 200451 94282 231838 94518
rect 232074 94282 232158 94518
rect 232394 94282 232478 94518
rect 232714 94282 232798 94518
rect 233034 94282 233118 94518
rect 233354 94282 233438 94518
rect 233674 94282 233758 94518
rect 233994 94282 234078 94518
rect 234314 94282 234398 94518
rect 234634 94282 234718 94518
rect 234954 94282 235038 94518
rect 235274 94282 235358 94518
rect 235594 94282 235716 94518
rect 0 94240 235716 94282
rect 0 83318 235716 83360
rect 0 83082 5122 83318
rect 5358 83082 5442 83318
rect 5678 83082 5762 83318
rect 5998 83082 6082 83318
rect 6318 83082 6402 83318
rect 6638 83082 6722 83318
rect 6958 83082 7042 83318
rect 7278 83082 7362 83318
rect 7598 83082 7682 83318
rect 7918 83082 8002 83318
rect 8238 83082 8322 83318
rect 8558 83082 8642 83318
rect 8878 83082 29549 83318
rect 29785 83082 60146 83318
rect 60382 83082 113549 83318
rect 113785 83082 144146 83318
rect 144382 83082 197549 83318
rect 197785 83082 226838 83318
rect 227074 83082 227158 83318
rect 227394 83082 227478 83318
rect 227714 83082 227798 83318
rect 228034 83082 228118 83318
rect 228354 83082 228438 83318
rect 228674 83082 228758 83318
rect 228994 83082 229078 83318
rect 229314 83082 229398 83318
rect 229634 83082 229718 83318
rect 229954 83082 230038 83318
rect 230274 83082 230358 83318
rect 230594 83082 235716 83318
rect 0 83040 235716 83082
rect 25468 76602 41980 76644
rect 25468 76366 25510 76602
rect 25746 76366 41702 76602
rect 41938 76366 41980 76602
rect 25468 76324 41980 76366
rect 0 72118 235716 72160
rect 0 71882 122 72118
rect 358 71882 442 72118
rect 678 71882 762 72118
rect 998 71882 1082 72118
rect 1318 71882 1402 72118
rect 1638 71882 1722 72118
rect 1958 71882 2042 72118
rect 2278 71882 2362 72118
rect 2598 71882 2682 72118
rect 2918 71882 3002 72118
rect 3238 71882 3322 72118
rect 3558 71882 3642 72118
rect 3878 71882 32215 72118
rect 32451 71882 75506 72118
rect 75742 71882 116215 72118
rect 116451 71882 159506 72118
rect 159742 71882 200215 72118
rect 200451 71882 231838 72118
rect 232074 71882 232158 72118
rect 232394 71882 232478 72118
rect 232714 71882 232798 72118
rect 233034 71882 233118 72118
rect 233354 71882 233438 72118
rect 233674 71882 233758 72118
rect 233994 71882 234078 72118
rect 234314 71882 234398 72118
rect 234634 71882 234718 72118
rect 234954 71882 235038 72118
rect 235274 71882 235358 72118
rect 235594 71882 235716 72118
rect 0 71840 235716 71882
rect 25652 69802 41980 69844
rect 25652 69566 25694 69802
rect 25930 69566 41702 69802
rect 41938 69566 41980 69802
rect 25652 69524 41980 69566
rect 0 60918 235716 60960
rect 0 60682 5122 60918
rect 5358 60682 5442 60918
rect 5678 60682 5762 60918
rect 5998 60682 6082 60918
rect 6318 60682 6402 60918
rect 6638 60682 6722 60918
rect 6958 60682 7042 60918
rect 7278 60682 7362 60918
rect 7598 60682 7682 60918
rect 7918 60682 8002 60918
rect 8238 60682 8322 60918
rect 8558 60682 8642 60918
rect 8878 60682 226838 60918
rect 227074 60682 227158 60918
rect 227394 60682 227478 60918
rect 227714 60682 227798 60918
rect 228034 60682 228118 60918
rect 228354 60682 228438 60918
rect 228674 60682 228758 60918
rect 228994 60682 229078 60918
rect 229314 60682 229398 60918
rect 229634 60682 229718 60918
rect 229954 60682 230038 60918
rect 230274 60682 230358 60918
rect 230594 60682 235716 60918
rect 0 60640 235716 60682
rect 0 49718 235716 49760
rect 0 49482 122 49718
rect 358 49482 442 49718
rect 678 49482 762 49718
rect 998 49482 1082 49718
rect 1318 49482 1402 49718
rect 1638 49482 1722 49718
rect 1958 49482 2042 49718
rect 2278 49482 2362 49718
rect 2598 49482 2682 49718
rect 2918 49482 3002 49718
rect 3238 49482 3322 49718
rect 3558 49482 3642 49718
rect 3878 49482 231838 49718
rect 232074 49482 232158 49718
rect 232394 49482 232478 49718
rect 232714 49482 232798 49718
rect 233034 49482 233118 49718
rect 233354 49482 233438 49718
rect 233674 49482 233758 49718
rect 233994 49482 234078 49718
rect 234314 49482 234398 49718
rect 234634 49482 234718 49718
rect 234954 49482 235038 49718
rect 235274 49482 235358 49718
rect 235594 49482 235716 49718
rect 0 49440 235716 49482
rect 211308 45322 214020 45364
rect 211308 45086 211350 45322
rect 211586 45086 213742 45322
rect 213978 45086 214020 45322
rect 211308 45044 214020 45086
rect 0 38518 235716 38560
rect 0 38282 5122 38518
rect 5358 38282 5442 38518
rect 5678 38282 5762 38518
rect 5998 38282 6082 38518
rect 6318 38282 6402 38518
rect 6638 38282 6722 38518
rect 6958 38282 7042 38518
rect 7278 38282 7362 38518
rect 7598 38282 7682 38518
rect 7918 38282 8002 38518
rect 8238 38282 8322 38518
rect 8558 38282 8642 38518
rect 8878 38282 25549 38518
rect 25785 38282 66882 38518
rect 67118 38282 109549 38518
rect 109785 38282 150882 38518
rect 151118 38282 193549 38518
rect 193785 38282 226838 38518
rect 227074 38282 227158 38518
rect 227394 38282 227478 38518
rect 227714 38282 227798 38518
rect 228034 38282 228118 38518
rect 228354 38282 228438 38518
rect 228674 38282 228758 38518
rect 228994 38282 229078 38518
rect 229314 38282 229398 38518
rect 229634 38282 229718 38518
rect 229954 38282 230038 38518
rect 230274 38282 230358 38518
rect 230594 38282 235716 38518
rect 0 38240 235716 38282
rect 212596 35122 214020 35164
rect 212596 34886 212638 35122
rect 212874 34886 213742 35122
rect 213978 34886 214020 35122
rect 212596 34844 214020 34886
rect 0 27318 235716 27360
rect 0 27082 122 27318
rect 358 27082 442 27318
rect 678 27082 762 27318
rect 998 27082 1082 27318
rect 1318 27082 1402 27318
rect 1638 27082 1722 27318
rect 1958 27082 2042 27318
rect 2278 27082 2362 27318
rect 2598 27082 2682 27318
rect 2918 27082 3002 27318
rect 3238 27082 3322 27318
rect 3558 27082 3642 27318
rect 3878 27082 30215 27318
rect 30451 27082 71882 27318
rect 72118 27082 114215 27318
rect 114451 27082 155882 27318
rect 156118 27082 198215 27318
rect 198451 27082 231838 27318
rect 232074 27082 232158 27318
rect 232394 27082 232478 27318
rect 232714 27082 232798 27318
rect 233034 27082 233118 27318
rect 233354 27082 233438 27318
rect 233674 27082 233758 27318
rect 233994 27082 234078 27318
rect 234314 27082 234398 27318
rect 234634 27082 234718 27318
rect 234954 27082 235038 27318
rect 235274 27082 235358 27318
rect 235594 27082 235716 27318
rect 0 27040 235716 27082
rect 19580 22882 54124 22924
rect 19580 22646 19622 22882
rect 19858 22646 53846 22882
rect 54082 22646 54124 22882
rect 19580 22604 54124 22646
rect 173772 22202 185316 22244
rect 173772 21966 173814 22202
rect 174050 21966 185038 22202
rect 185274 21966 185316 22202
rect 173772 21924 185316 21966
rect 88948 20842 101228 20884
rect 88948 20606 88990 20842
rect 89226 20606 100950 20842
rect 101186 20606 101228 20842
rect 88948 20564 101228 20606
rect 172852 20842 185316 20884
rect 172852 20606 172894 20842
rect 173130 20606 185038 20842
rect 185274 20606 185316 20842
rect 172852 20564 185316 20606
rect 89684 20162 101228 20204
rect 89684 19926 89726 20162
rect 89962 19926 100950 20162
rect 101186 19926 101228 20162
rect 89684 19884 101228 19926
rect 173220 20162 185684 20204
rect 173220 19926 173262 20162
rect 173498 19926 185406 20162
rect 185642 19926 185684 20162
rect 173220 19884 185684 19926
rect 0 16118 235716 16160
rect 0 15882 5122 16118
rect 5358 15882 5442 16118
rect 5678 15882 5762 16118
rect 5998 15882 6082 16118
rect 6318 15882 6402 16118
rect 6638 15882 6722 16118
rect 6958 15882 7042 16118
rect 7278 15882 7362 16118
rect 7598 15882 7682 16118
rect 7918 15882 8002 16118
rect 8238 15882 8322 16118
rect 8558 15882 8642 16118
rect 8878 15882 226838 16118
rect 227074 15882 227158 16118
rect 227394 15882 227478 16118
rect 227714 15882 227798 16118
rect 228034 15882 228118 16118
rect 228354 15882 228438 16118
rect 228674 15882 228758 16118
rect 228994 15882 229078 16118
rect 229314 15882 229398 16118
rect 229634 15882 229718 16118
rect 229954 15882 230038 16118
rect 230274 15882 230358 16118
rect 230594 15882 235716 16118
rect 0 15840 235716 15882
rect 5000 8878 230716 9000
rect 5000 8642 5122 8878
rect 5358 8642 5442 8878
rect 5678 8642 5762 8878
rect 5998 8642 6082 8878
rect 6318 8642 6402 8878
rect 6638 8642 6722 8878
rect 6958 8642 7042 8878
rect 7278 8642 7362 8878
rect 7598 8642 7682 8878
rect 7918 8642 8002 8878
rect 8238 8642 8322 8878
rect 8558 8642 8642 8878
rect 8878 8642 226838 8878
rect 227074 8642 227158 8878
rect 227394 8642 227478 8878
rect 227714 8642 227798 8878
rect 228034 8642 228118 8878
rect 228354 8642 228438 8878
rect 228674 8642 228758 8878
rect 228994 8642 229078 8878
rect 229314 8642 229398 8878
rect 229634 8642 229718 8878
rect 229954 8642 230038 8878
rect 230274 8642 230358 8878
rect 230594 8642 230716 8878
rect 5000 8558 230716 8642
rect 5000 8322 5122 8558
rect 5358 8322 5442 8558
rect 5678 8322 5762 8558
rect 5998 8322 6082 8558
rect 6318 8322 6402 8558
rect 6638 8322 6722 8558
rect 6958 8322 7042 8558
rect 7278 8322 7362 8558
rect 7598 8322 7682 8558
rect 7918 8322 8002 8558
rect 8238 8322 8322 8558
rect 8558 8322 8642 8558
rect 8878 8322 226838 8558
rect 227074 8322 227158 8558
rect 227394 8322 227478 8558
rect 227714 8322 227798 8558
rect 228034 8322 228118 8558
rect 228354 8322 228438 8558
rect 228674 8322 228758 8558
rect 228994 8322 229078 8558
rect 229314 8322 229398 8558
rect 229634 8322 229718 8558
rect 229954 8322 230038 8558
rect 230274 8322 230358 8558
rect 230594 8322 230716 8558
rect 5000 8238 230716 8322
rect 5000 8002 5122 8238
rect 5358 8002 5442 8238
rect 5678 8002 5762 8238
rect 5998 8002 6082 8238
rect 6318 8002 6402 8238
rect 6638 8002 6722 8238
rect 6958 8002 7042 8238
rect 7278 8002 7362 8238
rect 7598 8002 7682 8238
rect 7918 8002 8002 8238
rect 8238 8002 8322 8238
rect 8558 8002 8642 8238
rect 8878 8002 226838 8238
rect 227074 8002 227158 8238
rect 227394 8002 227478 8238
rect 227714 8002 227798 8238
rect 228034 8002 228118 8238
rect 228354 8002 228438 8238
rect 228674 8002 228758 8238
rect 228994 8002 229078 8238
rect 229314 8002 229398 8238
rect 229634 8002 229718 8238
rect 229954 8002 230038 8238
rect 230274 8002 230358 8238
rect 230594 8002 230716 8238
rect 5000 7918 230716 8002
rect 5000 7682 5122 7918
rect 5358 7682 5442 7918
rect 5678 7682 5762 7918
rect 5998 7682 6082 7918
rect 6318 7682 6402 7918
rect 6638 7682 6722 7918
rect 6958 7682 7042 7918
rect 7278 7682 7362 7918
rect 7598 7682 7682 7918
rect 7918 7682 8002 7918
rect 8238 7682 8322 7918
rect 8558 7682 8642 7918
rect 8878 7682 226838 7918
rect 227074 7682 227158 7918
rect 227394 7682 227478 7918
rect 227714 7682 227798 7918
rect 228034 7682 228118 7918
rect 228354 7682 228438 7918
rect 228674 7682 228758 7918
rect 228994 7682 229078 7918
rect 229314 7682 229398 7918
rect 229634 7682 229718 7918
rect 229954 7682 230038 7918
rect 230274 7682 230358 7918
rect 230594 7682 230716 7918
rect 5000 7598 230716 7682
rect 5000 7362 5122 7598
rect 5358 7362 5442 7598
rect 5678 7362 5762 7598
rect 5998 7362 6082 7598
rect 6318 7362 6402 7598
rect 6638 7362 6722 7598
rect 6958 7362 7042 7598
rect 7278 7362 7362 7598
rect 7598 7362 7682 7598
rect 7918 7362 8002 7598
rect 8238 7362 8322 7598
rect 8558 7362 8642 7598
rect 8878 7362 226838 7598
rect 227074 7362 227158 7598
rect 227394 7362 227478 7598
rect 227714 7362 227798 7598
rect 228034 7362 228118 7598
rect 228354 7362 228438 7598
rect 228674 7362 228758 7598
rect 228994 7362 229078 7598
rect 229314 7362 229398 7598
rect 229634 7362 229718 7598
rect 229954 7362 230038 7598
rect 230274 7362 230358 7598
rect 230594 7362 230716 7598
rect 5000 7278 230716 7362
rect 5000 7042 5122 7278
rect 5358 7042 5442 7278
rect 5678 7042 5762 7278
rect 5998 7042 6082 7278
rect 6318 7042 6402 7278
rect 6638 7042 6722 7278
rect 6958 7042 7042 7278
rect 7278 7042 7362 7278
rect 7598 7042 7682 7278
rect 7918 7042 8002 7278
rect 8238 7042 8322 7278
rect 8558 7042 8642 7278
rect 8878 7042 226838 7278
rect 227074 7042 227158 7278
rect 227394 7042 227478 7278
rect 227714 7042 227798 7278
rect 228034 7042 228118 7278
rect 228354 7042 228438 7278
rect 228674 7042 228758 7278
rect 228994 7042 229078 7278
rect 229314 7042 229398 7278
rect 229634 7042 229718 7278
rect 229954 7042 230038 7278
rect 230274 7042 230358 7278
rect 230594 7042 230716 7278
rect 5000 6958 230716 7042
rect 5000 6722 5122 6958
rect 5358 6722 5442 6958
rect 5678 6722 5762 6958
rect 5998 6722 6082 6958
rect 6318 6722 6402 6958
rect 6638 6722 6722 6958
rect 6958 6722 7042 6958
rect 7278 6722 7362 6958
rect 7598 6722 7682 6958
rect 7918 6722 8002 6958
rect 8238 6722 8322 6958
rect 8558 6722 8642 6958
rect 8878 6722 226838 6958
rect 227074 6722 227158 6958
rect 227394 6722 227478 6958
rect 227714 6722 227798 6958
rect 228034 6722 228118 6958
rect 228354 6722 228438 6958
rect 228674 6722 228758 6958
rect 228994 6722 229078 6958
rect 229314 6722 229398 6958
rect 229634 6722 229718 6958
rect 229954 6722 230038 6958
rect 230274 6722 230358 6958
rect 230594 6722 230716 6958
rect 5000 6638 230716 6722
rect 5000 6402 5122 6638
rect 5358 6402 5442 6638
rect 5678 6402 5762 6638
rect 5998 6402 6082 6638
rect 6318 6402 6402 6638
rect 6638 6402 6722 6638
rect 6958 6402 7042 6638
rect 7278 6402 7362 6638
rect 7598 6402 7682 6638
rect 7918 6402 8002 6638
rect 8238 6402 8322 6638
rect 8558 6402 8642 6638
rect 8878 6402 226838 6638
rect 227074 6402 227158 6638
rect 227394 6402 227478 6638
rect 227714 6402 227798 6638
rect 228034 6402 228118 6638
rect 228354 6402 228438 6638
rect 228674 6402 228758 6638
rect 228994 6402 229078 6638
rect 229314 6402 229398 6638
rect 229634 6402 229718 6638
rect 229954 6402 230038 6638
rect 230274 6402 230358 6638
rect 230594 6402 230716 6638
rect 5000 6318 230716 6402
rect 5000 6082 5122 6318
rect 5358 6082 5442 6318
rect 5678 6082 5762 6318
rect 5998 6082 6082 6318
rect 6318 6082 6402 6318
rect 6638 6082 6722 6318
rect 6958 6082 7042 6318
rect 7278 6082 7362 6318
rect 7598 6082 7682 6318
rect 7918 6082 8002 6318
rect 8238 6082 8322 6318
rect 8558 6082 8642 6318
rect 8878 6082 226838 6318
rect 227074 6082 227158 6318
rect 227394 6082 227478 6318
rect 227714 6082 227798 6318
rect 228034 6082 228118 6318
rect 228354 6082 228438 6318
rect 228674 6082 228758 6318
rect 228994 6082 229078 6318
rect 229314 6082 229398 6318
rect 229634 6082 229718 6318
rect 229954 6082 230038 6318
rect 230274 6082 230358 6318
rect 230594 6082 230716 6318
rect 5000 5998 230716 6082
rect 5000 5762 5122 5998
rect 5358 5762 5442 5998
rect 5678 5762 5762 5998
rect 5998 5762 6082 5998
rect 6318 5762 6402 5998
rect 6638 5762 6722 5998
rect 6958 5762 7042 5998
rect 7278 5762 7362 5998
rect 7598 5762 7682 5998
rect 7918 5762 8002 5998
rect 8238 5762 8322 5998
rect 8558 5762 8642 5998
rect 8878 5762 226838 5998
rect 227074 5762 227158 5998
rect 227394 5762 227478 5998
rect 227714 5762 227798 5998
rect 228034 5762 228118 5998
rect 228354 5762 228438 5998
rect 228674 5762 228758 5998
rect 228994 5762 229078 5998
rect 229314 5762 229398 5998
rect 229634 5762 229718 5998
rect 229954 5762 230038 5998
rect 230274 5762 230358 5998
rect 230594 5762 230716 5998
rect 5000 5678 230716 5762
rect 5000 5442 5122 5678
rect 5358 5442 5442 5678
rect 5678 5442 5762 5678
rect 5998 5442 6082 5678
rect 6318 5442 6402 5678
rect 6638 5442 6722 5678
rect 6958 5442 7042 5678
rect 7278 5442 7362 5678
rect 7598 5442 7682 5678
rect 7918 5442 8002 5678
rect 8238 5442 8322 5678
rect 8558 5442 8642 5678
rect 8878 5442 226838 5678
rect 227074 5442 227158 5678
rect 227394 5442 227478 5678
rect 227714 5442 227798 5678
rect 228034 5442 228118 5678
rect 228354 5442 228438 5678
rect 228674 5442 228758 5678
rect 228994 5442 229078 5678
rect 229314 5442 229398 5678
rect 229634 5442 229718 5678
rect 229954 5442 230038 5678
rect 230274 5442 230358 5678
rect 230594 5442 230716 5678
rect 5000 5358 230716 5442
rect 5000 5122 5122 5358
rect 5358 5122 5442 5358
rect 5678 5122 5762 5358
rect 5998 5122 6082 5358
rect 6318 5122 6402 5358
rect 6638 5122 6722 5358
rect 6958 5122 7042 5358
rect 7278 5122 7362 5358
rect 7598 5122 7682 5358
rect 7918 5122 8002 5358
rect 8238 5122 8322 5358
rect 8558 5122 8642 5358
rect 8878 5122 226838 5358
rect 227074 5122 227158 5358
rect 227394 5122 227478 5358
rect 227714 5122 227798 5358
rect 228034 5122 228118 5358
rect 228354 5122 228438 5358
rect 228674 5122 228758 5358
rect 228994 5122 229078 5358
rect 229314 5122 229398 5358
rect 229634 5122 229718 5358
rect 229954 5122 230038 5358
rect 230274 5122 230358 5358
rect 230594 5122 230716 5358
rect 5000 5000 230716 5122
rect 0 3878 235716 4000
rect 0 3642 122 3878
rect 358 3642 442 3878
rect 678 3642 762 3878
rect 998 3642 1082 3878
rect 1318 3642 1402 3878
rect 1638 3642 1722 3878
rect 1958 3642 2042 3878
rect 2278 3642 2362 3878
rect 2598 3642 2682 3878
rect 2918 3642 3002 3878
rect 3238 3642 3322 3878
rect 3558 3642 3642 3878
rect 3878 3642 231838 3878
rect 232074 3642 232158 3878
rect 232394 3642 232478 3878
rect 232714 3642 232798 3878
rect 233034 3642 233118 3878
rect 233354 3642 233438 3878
rect 233674 3642 233758 3878
rect 233994 3642 234078 3878
rect 234314 3642 234398 3878
rect 234634 3642 234718 3878
rect 234954 3642 235038 3878
rect 235274 3642 235358 3878
rect 235594 3642 235716 3878
rect 0 3558 235716 3642
rect 0 3322 122 3558
rect 358 3322 442 3558
rect 678 3322 762 3558
rect 998 3322 1082 3558
rect 1318 3322 1402 3558
rect 1638 3322 1722 3558
rect 1958 3322 2042 3558
rect 2278 3322 2362 3558
rect 2598 3322 2682 3558
rect 2918 3322 3002 3558
rect 3238 3322 3322 3558
rect 3558 3322 3642 3558
rect 3878 3322 231838 3558
rect 232074 3322 232158 3558
rect 232394 3322 232478 3558
rect 232714 3322 232798 3558
rect 233034 3322 233118 3558
rect 233354 3322 233438 3558
rect 233674 3322 233758 3558
rect 233994 3322 234078 3558
rect 234314 3322 234398 3558
rect 234634 3322 234718 3558
rect 234954 3322 235038 3558
rect 235274 3322 235358 3558
rect 235594 3322 235716 3558
rect 0 3238 235716 3322
rect 0 3002 122 3238
rect 358 3002 442 3238
rect 678 3002 762 3238
rect 998 3002 1082 3238
rect 1318 3002 1402 3238
rect 1638 3002 1722 3238
rect 1958 3002 2042 3238
rect 2278 3002 2362 3238
rect 2598 3002 2682 3238
rect 2918 3002 3002 3238
rect 3238 3002 3322 3238
rect 3558 3002 3642 3238
rect 3878 3002 231838 3238
rect 232074 3002 232158 3238
rect 232394 3002 232478 3238
rect 232714 3002 232798 3238
rect 233034 3002 233118 3238
rect 233354 3002 233438 3238
rect 233674 3002 233758 3238
rect 233994 3002 234078 3238
rect 234314 3002 234398 3238
rect 234634 3002 234718 3238
rect 234954 3002 235038 3238
rect 235274 3002 235358 3238
rect 235594 3002 235716 3238
rect 0 2918 235716 3002
rect 0 2682 122 2918
rect 358 2682 442 2918
rect 678 2682 762 2918
rect 998 2682 1082 2918
rect 1318 2682 1402 2918
rect 1638 2682 1722 2918
rect 1958 2682 2042 2918
rect 2278 2682 2362 2918
rect 2598 2682 2682 2918
rect 2918 2682 3002 2918
rect 3238 2682 3322 2918
rect 3558 2682 3642 2918
rect 3878 2682 231838 2918
rect 232074 2682 232158 2918
rect 232394 2682 232478 2918
rect 232714 2682 232798 2918
rect 233034 2682 233118 2918
rect 233354 2682 233438 2918
rect 233674 2682 233758 2918
rect 233994 2682 234078 2918
rect 234314 2682 234398 2918
rect 234634 2682 234718 2918
rect 234954 2682 235038 2918
rect 235274 2682 235358 2918
rect 235594 2682 235716 2918
rect 0 2598 235716 2682
rect 0 2362 122 2598
rect 358 2362 442 2598
rect 678 2362 762 2598
rect 998 2362 1082 2598
rect 1318 2362 1402 2598
rect 1638 2362 1722 2598
rect 1958 2362 2042 2598
rect 2278 2362 2362 2598
rect 2598 2362 2682 2598
rect 2918 2362 3002 2598
rect 3238 2362 3322 2598
rect 3558 2362 3642 2598
rect 3878 2362 231838 2598
rect 232074 2362 232158 2598
rect 232394 2362 232478 2598
rect 232714 2362 232798 2598
rect 233034 2362 233118 2598
rect 233354 2362 233438 2598
rect 233674 2362 233758 2598
rect 233994 2362 234078 2598
rect 234314 2362 234398 2598
rect 234634 2362 234718 2598
rect 234954 2362 235038 2598
rect 235274 2362 235358 2598
rect 235594 2362 235716 2598
rect 0 2278 235716 2362
rect 0 2042 122 2278
rect 358 2042 442 2278
rect 678 2042 762 2278
rect 998 2042 1082 2278
rect 1318 2042 1402 2278
rect 1638 2042 1722 2278
rect 1958 2042 2042 2278
rect 2278 2042 2362 2278
rect 2598 2042 2682 2278
rect 2918 2042 3002 2278
rect 3238 2042 3322 2278
rect 3558 2042 3642 2278
rect 3878 2042 231838 2278
rect 232074 2042 232158 2278
rect 232394 2042 232478 2278
rect 232714 2042 232798 2278
rect 233034 2042 233118 2278
rect 233354 2042 233438 2278
rect 233674 2042 233758 2278
rect 233994 2042 234078 2278
rect 234314 2042 234398 2278
rect 234634 2042 234718 2278
rect 234954 2042 235038 2278
rect 235274 2042 235358 2278
rect 235594 2042 235716 2278
rect 0 1958 235716 2042
rect 0 1722 122 1958
rect 358 1722 442 1958
rect 678 1722 762 1958
rect 998 1722 1082 1958
rect 1318 1722 1402 1958
rect 1638 1722 1722 1958
rect 1958 1722 2042 1958
rect 2278 1722 2362 1958
rect 2598 1722 2682 1958
rect 2918 1722 3002 1958
rect 3238 1722 3322 1958
rect 3558 1722 3642 1958
rect 3878 1722 231838 1958
rect 232074 1722 232158 1958
rect 232394 1722 232478 1958
rect 232714 1722 232798 1958
rect 233034 1722 233118 1958
rect 233354 1722 233438 1958
rect 233674 1722 233758 1958
rect 233994 1722 234078 1958
rect 234314 1722 234398 1958
rect 234634 1722 234718 1958
rect 234954 1722 235038 1958
rect 235274 1722 235358 1958
rect 235594 1722 235716 1958
rect 0 1638 235716 1722
rect 0 1402 122 1638
rect 358 1402 442 1638
rect 678 1402 762 1638
rect 998 1402 1082 1638
rect 1318 1402 1402 1638
rect 1638 1402 1722 1638
rect 1958 1402 2042 1638
rect 2278 1402 2362 1638
rect 2598 1402 2682 1638
rect 2918 1402 3002 1638
rect 3238 1402 3322 1638
rect 3558 1402 3642 1638
rect 3878 1402 231838 1638
rect 232074 1402 232158 1638
rect 232394 1402 232478 1638
rect 232714 1402 232798 1638
rect 233034 1402 233118 1638
rect 233354 1402 233438 1638
rect 233674 1402 233758 1638
rect 233994 1402 234078 1638
rect 234314 1402 234398 1638
rect 234634 1402 234718 1638
rect 234954 1402 235038 1638
rect 235274 1402 235358 1638
rect 235594 1402 235716 1638
rect 0 1318 235716 1402
rect 0 1082 122 1318
rect 358 1082 442 1318
rect 678 1082 762 1318
rect 998 1082 1082 1318
rect 1318 1082 1402 1318
rect 1638 1082 1722 1318
rect 1958 1082 2042 1318
rect 2278 1082 2362 1318
rect 2598 1082 2682 1318
rect 2918 1082 3002 1318
rect 3238 1082 3322 1318
rect 3558 1082 3642 1318
rect 3878 1082 231838 1318
rect 232074 1082 232158 1318
rect 232394 1082 232478 1318
rect 232714 1082 232798 1318
rect 233034 1082 233118 1318
rect 233354 1082 233438 1318
rect 233674 1082 233758 1318
rect 233994 1082 234078 1318
rect 234314 1082 234398 1318
rect 234634 1082 234718 1318
rect 234954 1082 235038 1318
rect 235274 1082 235358 1318
rect 235594 1082 235716 1318
rect 0 998 235716 1082
rect 0 762 122 998
rect 358 762 442 998
rect 678 762 762 998
rect 998 762 1082 998
rect 1318 762 1402 998
rect 1638 762 1722 998
rect 1958 762 2042 998
rect 2278 762 2362 998
rect 2598 762 2682 998
rect 2918 762 3002 998
rect 3238 762 3322 998
rect 3558 762 3642 998
rect 3878 762 231838 998
rect 232074 762 232158 998
rect 232394 762 232478 998
rect 232714 762 232798 998
rect 233034 762 233118 998
rect 233354 762 233438 998
rect 233674 762 233758 998
rect 233994 762 234078 998
rect 234314 762 234398 998
rect 234634 762 234718 998
rect 234954 762 235038 998
rect 235274 762 235358 998
rect 235594 762 235716 998
rect 0 678 235716 762
rect 0 442 122 678
rect 358 442 442 678
rect 678 442 762 678
rect 998 442 1082 678
rect 1318 442 1402 678
rect 1638 442 1722 678
rect 1958 442 2042 678
rect 2278 442 2362 678
rect 2598 442 2682 678
rect 2918 442 3002 678
rect 3238 442 3322 678
rect 3558 442 3642 678
rect 3878 442 231838 678
rect 232074 442 232158 678
rect 232394 442 232478 678
rect 232714 442 232798 678
rect 233034 442 233118 678
rect 233354 442 233438 678
rect 233674 442 233758 678
rect 233994 442 234078 678
rect 234314 442 234398 678
rect 234634 442 234718 678
rect 234954 442 235038 678
rect 235274 442 235358 678
rect 235594 442 235716 678
rect 0 358 235716 442
rect 0 122 122 358
rect 358 122 442 358
rect 678 122 762 358
rect 998 122 1082 358
rect 1318 122 1402 358
rect 1638 122 1722 358
rect 1958 122 2042 358
rect 2278 122 2362 358
rect 2598 122 2682 358
rect 2918 122 3002 358
rect 3238 122 3322 358
rect 3558 122 3642 358
rect 3878 122 231838 358
rect 232074 122 232158 358
rect 232394 122 232478 358
rect 232714 122 232798 358
rect 233034 122 233118 358
rect 233354 122 233438 358
rect 233674 122 233758 358
rect 233994 122 234078 358
rect 234314 122 234398 358
rect 234634 122 234718 358
rect 234954 122 235038 358
rect 235274 122 235358 358
rect 235594 122 235716 358
rect 0 0 235716 122
use grid_clb  grid_clb_1__1_
timestamp 1605016838
transform 1 0 55896 0 1 59824
box 0 0 40000 40000
use sb_0__0_  sb_0__0_
timestamp 1605016838
transform 1 0 19896 0 1 18824
box 0 0 28000 27720
use cby_0__1_  cby_0__1_
timestamp 1605016838
transform 1 0 25896 0 1 59824
box 0 0 16000 40000
use cbx_1__0_  cbx_1__0_
timestamp 1605016838
transform 1 0 60896 0 1 20824
box 0 0 30000 24000
use grid_clb  grid_clb_2__1_
timestamp 1605016838
transform 1 0 139896 0 1 59824
box 0 0 40000 40000
use sb_1__0_  sb_1__0_
timestamp 1605016838
transform 1 0 103896 0 1 18824
box 0 0 28000 28000
use cby_1__1_  cby_1__1_
timestamp 1605016838
transform 1 0 109896 0 1 59824
box 0 0 16000 40000
use cbx_1__0_  cbx_2__0_
timestamp 1605016838
transform 1 0 144896 0 1 20824
box 0 0 30000 24000
use sb_2__0_  sb_2__0_
timestamp 1605016838
transform 1 0 187896 0 1 18824
box 0 0 27679 28000
use cby_2__1_  cby_2__1_
timestamp 1605016838
transform 1 0 193896 0 1 59824
box 0 0 16000 40000
use sb_0__1_  sb_0__1_
timestamp 1605016838
transform 1 0 19896 0 1 112824
box 0 0 28000 28000
use cbx_1__1_  cbx_1__1_
timestamp 1605016838
transform 1 0 60896 0 1 114824
box 0 0 30000 24000
use sb_1__1_  sb_1__1_
timestamp 1605016838
transform 1 0 103896 0 1 112824
box 0 0 28000 28000
use cbx_1__1_  cbx_2__1_
timestamp 1605016838
transform 1 0 144896 0 1 114824
box 0 0 30000 24000
use sb_2__1_  sb_2__1_
timestamp 1605016838
transform 1 0 187896 0 1 112824
box 0 0 28000 28000
use grid_clb  grid_clb_1__2_
timestamp 1605016838
transform 1 0 55896 0 1 153824
box 0 0 40000 40000
use cby_0__1_  cby_0__2_
timestamp 1605016838
transform 1 0 25896 0 1 153824
box 0 0 16000 40000
use grid_clb  grid_clb_2__2_
timestamp 1605016838
transform 1 0 139896 0 1 153824
box 0 0 40000 40000
use cby_1__1_  cby_1__2_
timestamp 1605016838
transform 1 0 109896 0 1 153824
box 0 0 16000 40000
use cby_2__1_  cby_2__2_
timestamp 1605016838
transform 1 0 193896 0 1 153824
box 0 0 16000 40000
use sb_0__2_  sb_0__2_
timestamp 1605016838
transform 1 0 19895 0 1 206824
box 1 0 27712 28000
use cbx_1__2_  cbx_1__2_
timestamp 1605016838
transform 1 0 60896 0 1 208824
box 0 0 30000 24000
use sb_1__2_  sb_1__2_
timestamp 1605016838
transform 1 0 103896 0 1 206824
box 0 0 28000 28000
use cbx_1__2_  cbx_2__2_
timestamp 1605016838
transform 1 0 144896 0 1 208824
box 0 0 30000 24000
use sb_2__2_  sb_2__2_
timestamp 1605016838
transform 1 0 187896 0 1 206824
box 0 0 28000 27736
<< labels >>
rlabel metal3 s 9896 20528 10376 20648 6 Test_en
port 0 nsew default input
rlabel metal3 s 225416 21888 225896 22008 6 ccff_head
port 1 nsew default input
rlabel metal3 s 9896 209296 10376 209416 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 9896 44056 10376 44176 6 clk
port 3 nsew default input
rlabel metal2 s 27854 244344 27910 244824 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[0]
port 4 nsew default tristate
rlabel metal2 s 120866 8824 120922 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[10]
port 5 nsew default tristate
rlabel metal2 s 126846 8824 126902 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[11]
port 6 nsew default tristate
rlabel metal2 s 132826 8824 132882 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[12]
port 7 nsew default tristate
rlabel metal2 s 138806 8824 138862 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[13]
port 8 nsew default tristate
rlabel metal2 s 144786 8824 144842 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[14]
port 9 nsew default tristate
rlabel metal2 s 150858 8824 150914 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[15]
port 10 nsew default tristate
rlabel metal3 s 9896 67720 10376 67840 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[16]
port 11 nsew default tristate
rlabel metal3 s 9896 138440 10376 138560 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[17]
port 12 nsew default tristate
rlabel metal2 s 63826 244344 63882 244824 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[1]
port 13 nsew default tristate
rlabel metal3 s 225416 100496 225896 100616 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[2]
port 14 nsew default tristate
rlabel metal3 s 225416 126744 225896 126864 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[3]
port 15 nsew default tristate
rlabel metal2 s 12858 8824 12914 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[4]
port 16 nsew default tristate
rlabel metal2 s 18838 8824 18894 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[5]
port 17 nsew default tristate
rlabel metal2 s 24818 8824 24874 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[6]
port 18 nsew default tristate
rlabel metal2 s 30798 8824 30854 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[7]
port 19 nsew default tristate
rlabel metal2 s 36778 8824 36834 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[8]
port 20 nsew default tristate
rlabel metal2 s 42850 8824 42906 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[9]
port 21 nsew default tristate
rlabel metal2 s 99798 244344 99854 244824 6 gfpga_pad_EMBEDDED_IO_SOC_IN[0]
port 22 nsew default input
rlabel metal2 s 156838 8824 156894 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[10]
port 23 nsew default input
rlabel metal2 s 162818 8824 162874 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[11]
port 24 nsew default input
rlabel metal2 s 168798 8824 168854 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[12]
port 25 nsew default input
rlabel metal2 s 174870 8824 174926 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[13]
port 26 nsew default input
rlabel metal2 s 180850 8824 180906 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[14]
port 27 nsew default input
rlabel metal2 s 186830 8824 186886 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[15]
port 28 nsew default input
rlabel metal3 s 9896 91248 10376 91368 6 gfpga_pad_EMBEDDED_IO_SOC_IN[16]
port 29 nsew default input
rlabel metal3 s 9896 162104 10376 162224 6 gfpga_pad_EMBEDDED_IO_SOC_IN[17]
port 30 nsew default input
rlabel metal2 s 135862 244344 135918 244824 6 gfpga_pad_EMBEDDED_IO_SOC_IN[1]
port 31 nsew default input
rlabel metal3 s 225416 152856 225896 152976 6 gfpga_pad_EMBEDDED_IO_SOC_IN[2]
port 32 nsew default input
rlabel metal3 s 225416 179104 225896 179224 6 gfpga_pad_EMBEDDED_IO_SOC_IN[3]
port 33 nsew default input
rlabel metal2 s 48830 8824 48886 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[4]
port 34 nsew default input
rlabel metal2 s 54810 8824 54866 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[5]
port 35 nsew default input
rlabel metal2 s 60790 8824 60846 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[6]
port 36 nsew default input
rlabel metal2 s 66862 8824 66918 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[7]
port 37 nsew default input
rlabel metal2 s 72842 8824 72898 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[8]
port 38 nsew default input
rlabel metal2 s 78822 8824 78878 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[9]
port 39 nsew default input
rlabel metal2 s 171834 244344 171890 244824 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[0]
port 40 nsew default tristate
rlabel metal2 s 192810 8824 192866 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[10]
port 41 nsew default tristate
rlabel metal2 s 198790 8824 198846 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[11]
port 42 nsew default tristate
rlabel metal2 s 204862 8824 204918 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[12]
port 43 nsew default tristate
rlabel metal2 s 210842 8824 210898 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[13]
port 44 nsew default tristate
rlabel metal2 s 216822 8824 216878 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[14]
port 45 nsew default tristate
rlabel metal2 s 222802 8824 222858 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[15]
port 46 nsew default tristate
rlabel metal3 s 9896 114912 10376 115032 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[16]
port 47 nsew default tristate
rlabel metal3 s 9896 185632 10376 185752 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[17]
port 48 nsew default tristate
rlabel metal2 s 207806 244344 207862 244824 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[1]
port 49 nsew default tristate
rlabel metal3 s 225416 205352 225896 205472 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[2]
port 50 nsew default tristate
rlabel metal3 s 225416 231600 225896 231720 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[3]
port 51 nsew default tristate
rlabel metal2 s 84802 8824 84858 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[4]
port 52 nsew default tristate
rlabel metal2 s 90782 8824 90838 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[5]
port 53 nsew default tristate
rlabel metal2 s 96854 8824 96910 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[6]
port 54 nsew default tristate
rlabel metal2 s 102834 8824 102890 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[7]
port 55 nsew default tristate
rlabel metal2 s 108814 8824 108870 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[8]
port 56 nsew default tristate
rlabel metal2 s 114794 8824 114850 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[9]
port 57 nsew default tristate
rlabel metal3 s 225416 74248 225896 74368 6 prog_clk
port 58 nsew default input
rlabel metal3 s 225416 48000 225896 48120 6 sc_head
port 59 nsew default input
rlabel metal3 s 9896 232824 10376 232944 6 sc_tail
port 60 nsew default tristate
rlabel metal5 s 5000 5000 230716 9000 8 VPWR
port 61 nsew default input
rlabel metal5 s 0 0 235716 4000 8 VGND
port 62 nsew default input
<< properties >>
string FIXED_BBOX 0 0 235716 253200
<< end >>
