magic
tech sky130A
magscale 1 2
timestamp 1606928374
<< locali >>
rect 4445 12291 4479 12393
rect 6653 8347 6687 8585
rect 9505 7905 9597 7939
rect 9505 7735 9539 7905
<< viali >>
rect 1961 14569 1995 14603
rect 2697 14569 2731 14603
rect 1777 14433 1811 14467
rect 2513 14433 2547 14467
rect 3249 14433 3283 14467
rect 15485 14433 15519 14467
rect 3433 14229 3467 14263
rect 15669 14229 15703 14263
rect 3341 14025 3375 14059
rect 7021 14025 7055 14059
rect 1593 13957 1627 13991
rect 14657 13957 14691 13991
rect 2237 13889 2271 13923
rect 2053 13821 2087 13855
rect 3157 13821 3191 13855
rect 6009 13821 6043 13855
rect 6837 13821 6871 13855
rect 13461 13821 13495 13855
rect 14473 13821 14507 13855
rect 15577 13821 15611 13855
rect 1961 13685 1995 13719
rect 6193 13685 6227 13719
rect 13645 13685 13679 13719
rect 15761 13685 15795 13719
rect 1685 13481 1719 13515
rect 2697 13413 2731 13447
rect 1501 13345 1535 13379
rect 2605 13345 2639 13379
rect 15336 13345 15370 13379
rect 17877 13345 17911 13379
rect 2789 13277 2823 13311
rect 4077 13277 4111 13311
rect 17233 13277 17267 13311
rect 2237 13141 2271 13175
rect 15439 13141 15473 13175
rect 18061 13141 18095 13175
rect 1501 12937 1535 12971
rect 2145 12801 2179 12835
rect 4537 12801 4571 12835
rect 6101 12801 6135 12835
rect 8493 12801 8527 12835
rect 1869 12733 1903 12767
rect 2697 12733 2731 12767
rect 8033 12733 8067 12767
rect 12484 12733 12518 12767
rect 13128 12733 13162 12767
rect 15276 12733 15310 12767
rect 16221 12733 16255 12767
rect 17233 12733 17267 12767
rect 2942 12665 2976 12699
rect 1961 12597 1995 12631
rect 4077 12597 4111 12631
rect 5549 12597 5583 12631
rect 5917 12597 5951 12631
rect 6009 12597 6043 12631
rect 6837 12597 6871 12631
rect 12587 12597 12621 12631
rect 13231 12597 13265 12631
rect 15347 12597 15381 12631
rect 16405 12597 16439 12631
rect 17417 12597 17451 12631
rect 2237 12393 2271 12427
rect 4445 12393 4479 12427
rect 5917 12393 5951 12427
rect 4782 12325 4816 12359
rect 8585 12325 8619 12359
rect 1501 12257 1535 12291
rect 2605 12257 2639 12291
rect 4445 12257 4479 12291
rect 4537 12257 4571 12291
rect 6644 12257 6678 12291
rect 12300 12257 12334 12291
rect 13312 12257 13346 12291
rect 14264 12257 14298 12291
rect 15577 12257 15611 12291
rect 16405 12257 16439 12291
rect 17141 12257 17175 12291
rect 17877 12257 17911 12291
rect 2697 12189 2731 12223
rect 2789 12189 2823 12223
rect 6377 12189 6411 12223
rect 8677 12189 8711 12223
rect 8769 12189 8803 12223
rect 1685 12121 1719 12155
rect 17325 12121 17359 12155
rect 7757 12053 7791 12087
rect 8217 12053 8251 12087
rect 12403 12053 12437 12087
rect 13415 12053 13449 12087
rect 14335 12053 14369 12087
rect 15761 12053 15795 12087
rect 16589 12053 16623 12087
rect 18061 12053 18095 12087
rect 4905 11849 4939 11883
rect 8769 11849 8803 11883
rect 16681 11781 16715 11815
rect 2881 11713 2915 11747
rect 6009 11713 6043 11747
rect 6193 11713 6227 11747
rect 9321 11713 9355 11747
rect 13461 11713 13495 11747
rect 13645 11713 13679 11747
rect 15669 11713 15703 11747
rect 1593 11645 1627 11679
rect 3525 11645 3559 11679
rect 3792 11645 3826 11679
rect 6837 11645 6871 11679
rect 14381 11645 14415 11679
rect 16497 11645 16531 11679
rect 17233 11645 17267 11679
rect 2697 11577 2731 11611
rect 5917 11577 5951 11611
rect 7082 11577 7116 11611
rect 15485 11577 15519 11611
rect 1777 11509 1811 11543
rect 2329 11509 2363 11543
rect 2789 11509 2823 11543
rect 5549 11509 5583 11543
rect 8217 11509 8251 11543
rect 9137 11509 9171 11543
rect 9229 11509 9263 11543
rect 11161 11509 11195 11543
rect 13001 11509 13035 11543
rect 13369 11509 13403 11543
rect 14565 11509 14599 11543
rect 15117 11509 15151 11543
rect 15577 11509 15611 11543
rect 17417 11509 17451 11543
rect 1501 11305 1535 11339
rect 1869 11305 1903 11339
rect 2697 11305 2731 11339
rect 6009 11305 6043 11339
rect 14657 11305 14691 11339
rect 15761 11305 15795 11339
rect 16957 11305 16991 11339
rect 3157 11237 3191 11271
rect 7840 11237 7874 11271
rect 16129 11237 16163 11271
rect 3065 11169 3099 11203
rect 4721 11169 4755 11203
rect 5917 11169 5951 11203
rect 6837 11169 6871 11203
rect 7580 11169 7614 11203
rect 10032 11169 10066 11203
rect 10876 11169 10910 11203
rect 12900 11169 12934 11203
rect 14473 11169 14507 11203
rect 16221 11169 16255 11203
rect 17325 11169 17359 11203
rect 1961 11101 1995 11135
rect 2145 11101 2179 11135
rect 3341 11101 3375 11135
rect 4813 11101 4847 11135
rect 4997 11101 5031 11135
rect 6193 11101 6227 11135
rect 10609 11101 10643 11135
rect 12633 11101 12667 11135
rect 16313 11101 16347 11135
rect 17417 11101 17451 11135
rect 17509 11101 17543 11135
rect 7021 11033 7055 11067
rect 10103 11033 10137 11067
rect 4353 10965 4387 10999
rect 5549 10965 5583 10999
rect 8953 10965 8987 10999
rect 11989 10965 12023 10999
rect 14013 10965 14047 10999
rect 6837 10761 6871 10795
rect 16773 10761 16807 10795
rect 5089 10625 5123 10659
rect 5273 10625 5307 10659
rect 7389 10625 7423 10659
rect 8953 10625 8987 10659
rect 11253 10625 11287 10659
rect 11437 10625 11471 10659
rect 13093 10625 13127 10659
rect 13829 10625 13863 10659
rect 17417 10625 17451 10659
rect 1685 10557 1719 10591
rect 2421 10557 2455 10591
rect 4997 10557 5031 10591
rect 5825 10557 5859 10591
rect 7205 10557 7239 10591
rect 8033 10557 8067 10591
rect 16037 10557 16071 10591
rect 17141 10557 17175 10591
rect 17233 10557 17267 10591
rect 2688 10489 2722 10523
rect 6101 10489 6135 10523
rect 9220 10489 9254 10523
rect 12817 10489 12851 10523
rect 14096 10489 14130 10523
rect 1869 10421 1903 10455
rect 3801 10421 3835 10455
rect 4629 10421 4663 10455
rect 7297 10421 7331 10455
rect 8217 10421 8251 10455
rect 10333 10421 10367 10455
rect 10793 10421 10827 10455
rect 11161 10421 11195 10455
rect 12449 10421 12483 10455
rect 12909 10421 12943 10455
rect 15209 10421 15243 10455
rect 16221 10421 16255 10455
rect 1593 10217 1627 10251
rect 1961 10217 1995 10251
rect 2789 10217 2823 10251
rect 5365 10217 5399 10251
rect 9873 10217 9907 10251
rect 10241 10217 10275 10251
rect 11069 10217 11103 10251
rect 12633 10217 12667 10251
rect 13461 10217 13495 10251
rect 17233 10217 17267 10251
rect 17601 10217 17635 10251
rect 5733 10149 5767 10183
rect 7840 10149 7874 10183
rect 11529 10149 11563 10183
rect 13921 10149 13955 10183
rect 2053 10081 2087 10115
rect 3157 10081 3191 10115
rect 4445 10081 4479 10115
rect 6561 10081 6595 10115
rect 11437 10081 11471 10115
rect 13829 10081 13863 10115
rect 15393 10081 15427 10115
rect 15660 10081 15694 10115
rect 2237 10013 2271 10047
rect 3249 10013 3283 10047
rect 3341 10013 3375 10047
rect 4537 10013 4571 10047
rect 4721 10013 4755 10047
rect 5825 10013 5859 10047
rect 6009 10013 6043 10047
rect 6745 10013 6779 10047
rect 7573 10013 7607 10047
rect 10333 10013 10367 10047
rect 10425 10013 10459 10047
rect 11621 10013 11655 10047
rect 12725 10013 12759 10047
rect 12817 10013 12851 10047
rect 14013 10013 14047 10047
rect 17693 10013 17727 10047
rect 17785 10013 17819 10047
rect 8953 9945 8987 9979
rect 12265 9945 12299 9979
rect 4077 9877 4111 9911
rect 16773 9877 16807 9911
rect 3709 9673 3743 9707
rect 12449 9673 12483 9707
rect 3249 9605 3283 9639
rect 4997 9605 5031 9639
rect 5273 9605 5307 9639
rect 8309 9605 8343 9639
rect 10793 9605 10827 9639
rect 15577 9605 15611 9639
rect 4261 9537 4295 9571
rect 5733 9537 5767 9571
rect 5917 9537 5951 9571
rect 6929 9537 6963 9571
rect 9321 9537 9355 9571
rect 10241 9537 10275 9571
rect 10425 9537 10459 9571
rect 11437 9537 11471 9571
rect 13001 9537 13035 9571
rect 14197 9537 14231 9571
rect 17325 9537 17359 9571
rect 1869 9469 1903 9503
rect 5181 9469 5215 9503
rect 6653 9469 6687 9503
rect 7196 9469 7230 9503
rect 11161 9469 11195 9503
rect 11253 9469 11287 9503
rect 12909 9469 12943 9503
rect 16037 9469 16071 9503
rect 17141 9469 17175 9503
rect 2136 9401 2170 9435
rect 4169 9401 4203 9435
rect 5641 9401 5675 9435
rect 14464 9401 14498 9435
rect 4077 9333 4111 9367
rect 6469 9333 6503 9367
rect 8769 9333 8803 9367
rect 9137 9333 9171 9367
rect 9229 9333 9263 9367
rect 9781 9333 9815 9367
rect 10149 9333 10183 9367
rect 12817 9333 12851 9367
rect 16221 9333 16255 9367
rect 16773 9333 16807 9367
rect 17233 9333 17267 9367
rect 2973 9129 3007 9163
rect 5917 9129 5951 9163
rect 7113 9129 7147 9163
rect 7481 9129 7515 9163
rect 7573 9129 7607 9163
rect 8401 9129 8435 9163
rect 12357 9129 12391 9163
rect 13001 9129 13035 9163
rect 14197 9129 14231 9163
rect 16681 9129 16715 9163
rect 17601 9129 17635 9163
rect 1860 9061 1894 9095
rect 6285 9061 6319 9095
rect 8769 9061 8803 9095
rect 10057 9061 10091 9095
rect 13369 9061 13403 9095
rect 1593 8993 1627 9027
rect 4077 8993 4111 9027
rect 4344 8993 4378 9027
rect 6377 8993 6411 9027
rect 10517 8993 10551 9027
rect 10977 8993 11011 9027
rect 11244 8993 11278 9027
rect 14381 8993 14415 9027
rect 14473 8993 14507 9027
rect 15568 8993 15602 9027
rect 17509 8993 17543 9027
rect 6561 8925 6595 8959
rect 7665 8925 7699 8959
rect 8861 8925 8895 8959
rect 9045 8925 9079 8959
rect 10149 8925 10183 8959
rect 10333 8925 10367 8959
rect 13461 8925 13495 8959
rect 13645 8925 13679 8959
rect 15301 8925 15335 8959
rect 17693 8925 17727 8959
rect 9689 8857 9723 8891
rect 17141 8857 17175 8891
rect 5457 8789 5491 8823
rect 10701 8789 10735 8823
rect 14657 8789 14691 8823
rect 4261 8585 4295 8619
rect 6653 8585 6687 8619
rect 7389 8585 7423 8619
rect 14013 8585 14047 8619
rect 16405 8585 16439 8619
rect 1869 8517 1903 8551
rect 2513 8449 2547 8483
rect 3525 8449 3559 8483
rect 3709 8449 3743 8483
rect 4905 8449 4939 8483
rect 6009 8449 6043 8483
rect 2329 8381 2363 8415
rect 3433 8381 3467 8415
rect 7021 8517 7055 8551
rect 15945 8517 15979 8551
rect 7849 8449 7883 8483
rect 8033 8449 8067 8483
rect 10425 8449 10459 8483
rect 12909 8449 12943 8483
rect 13093 8449 13127 8483
rect 14565 8449 14599 8483
rect 16957 8449 16991 8483
rect 6837 8381 6871 8415
rect 8585 8381 8619 8415
rect 10333 8381 10367 8415
rect 13829 8381 13863 8415
rect 14832 8381 14866 8415
rect 4629 8313 4663 8347
rect 5825 8313 5859 8347
rect 5917 8313 5951 8347
rect 6653 8313 6687 8347
rect 10692 8313 10726 8347
rect 12817 8313 12851 8347
rect 13277 8313 13311 8347
rect 16865 8313 16899 8347
rect 2237 8245 2271 8279
rect 3065 8245 3099 8279
rect 4721 8245 4755 8279
rect 5457 8245 5491 8279
rect 7757 8245 7791 8279
rect 11805 8245 11839 8279
rect 12449 8245 12483 8279
rect 16773 8245 16807 8279
rect 3065 8041 3099 8075
rect 12081 8041 12115 8075
rect 15853 8041 15887 8075
rect 15945 8041 15979 8075
rect 16681 8041 16715 8075
rect 3157 7973 3191 8007
rect 12173 7973 12207 8007
rect 17141 7973 17175 8007
rect 1685 7905 1719 7939
rect 4905 7905 4939 7939
rect 6000 7905 6034 7939
rect 7941 7905 7975 7939
rect 8033 7905 8067 7939
rect 8769 7905 8803 7939
rect 9597 7905 9631 7939
rect 9945 7905 9979 7939
rect 13277 7905 13311 7939
rect 13369 7905 13403 7939
rect 14289 7905 14323 7939
rect 14473 7905 14507 7939
rect 17049 7905 17083 7939
rect 17877 7905 17911 7939
rect 3341 7837 3375 7871
rect 4997 7837 5031 7871
rect 5181 7837 5215 7871
rect 5733 7837 5767 7871
rect 8125 7837 8159 7871
rect 1869 7769 1903 7803
rect 8953 7769 8987 7803
rect 9689 7837 9723 7871
rect 12265 7837 12299 7871
rect 13461 7837 13495 7871
rect 16129 7837 16163 7871
rect 17233 7837 17267 7871
rect 2697 7701 2731 7735
rect 4537 7701 4571 7735
rect 7113 7701 7147 7735
rect 7573 7701 7607 7735
rect 9505 7701 9539 7735
rect 11069 7701 11103 7735
rect 11713 7701 11747 7735
rect 12909 7701 12943 7735
rect 14105 7701 14139 7735
rect 14657 7701 14691 7735
rect 15485 7701 15519 7735
rect 18061 7701 18095 7735
rect 2237 7497 2271 7531
rect 4261 7497 4295 7531
rect 5457 7497 5491 7531
rect 7205 7497 7239 7531
rect 15117 7497 15151 7531
rect 1685 7429 1719 7463
rect 9781 7429 9815 7463
rect 2789 7361 2823 7395
rect 4721 7361 4755 7395
rect 4905 7361 4939 7395
rect 6009 7361 6043 7395
rect 7849 7361 7883 7395
rect 13093 7361 13127 7395
rect 13737 7361 13771 7395
rect 15577 7361 15611 7395
rect 1501 7293 1535 7327
rect 2605 7293 2639 7327
rect 2697 7293 2731 7327
rect 3433 7293 3467 7327
rect 5825 7293 5859 7327
rect 7573 7293 7607 7327
rect 8401 7293 8435 7327
rect 10425 7293 10459 7327
rect 7665 7225 7699 7259
rect 8646 7225 8680 7259
rect 10670 7225 10704 7259
rect 12817 7225 12851 7259
rect 14004 7225 14038 7259
rect 15844 7225 15878 7259
rect 3617 7157 3651 7191
rect 4629 7157 4663 7191
rect 5917 7157 5951 7191
rect 11805 7157 11839 7191
rect 12449 7157 12483 7191
rect 12909 7157 12943 7191
rect 16957 7157 16991 7191
rect 1593 6953 1627 6987
rect 1961 6953 1995 6987
rect 5457 6953 5491 6987
rect 7481 6953 7515 6987
rect 8309 6953 8343 6987
rect 8677 6953 8711 6987
rect 10701 6953 10735 6987
rect 14381 6953 14415 6987
rect 15301 6953 15335 6987
rect 17049 6953 17083 6987
rect 3157 6885 3191 6919
rect 3249 6885 3283 6919
rect 9689 6885 9723 6919
rect 17141 6885 17175 6919
rect 4333 6817 4367 6851
rect 6285 6817 6319 6851
rect 10793 6817 10827 6851
rect 11796 6817 11830 6851
rect 13369 6817 13403 6851
rect 15669 6817 15703 6851
rect 17877 6817 17911 6851
rect 2053 6749 2087 6783
rect 2237 6749 2271 6783
rect 3341 6749 3375 6783
rect 4077 6749 4111 6783
rect 6377 6749 6411 6783
rect 6561 6749 6595 6783
rect 7573 6749 7607 6783
rect 7665 6749 7699 6783
rect 8769 6749 8803 6783
rect 8953 6749 8987 6783
rect 10885 6749 10919 6783
rect 11529 6749 11563 6783
rect 14473 6749 14507 6783
rect 14565 6749 14599 6783
rect 15761 6749 15795 6783
rect 15853 6749 15887 6783
rect 17233 6749 17267 6783
rect 2789 6681 2823 6715
rect 5917 6681 5951 6715
rect 7113 6681 7147 6715
rect 10333 6681 10367 6715
rect 16681 6681 16715 6715
rect 12909 6613 12943 6647
rect 14013 6613 14047 6647
rect 18061 6613 18095 6647
rect 3801 6409 3835 6443
rect 6837 6409 6871 6443
rect 8125 6409 8159 6443
rect 16037 6409 16071 6443
rect 1869 6341 1903 6375
rect 7481 6273 7515 6307
rect 8677 6273 8711 6307
rect 9321 6273 9355 6307
rect 11621 6273 11655 6307
rect 11805 6273 11839 6307
rect 12909 6273 12943 6307
rect 13001 6273 13035 6307
rect 16589 6273 16623 6307
rect 1685 6205 1719 6239
rect 2421 6205 2455 6239
rect 4445 6205 4479 6239
rect 4712 6205 4746 6239
rect 6469 6205 6503 6239
rect 7297 6205 7331 6239
rect 8493 6205 8527 6239
rect 8585 6205 8619 6239
rect 9588 6205 9622 6239
rect 12817 6205 12851 6239
rect 14197 6205 14231 6239
rect 17233 6205 17267 6239
rect 2688 6137 2722 6171
rect 7205 6137 7239 6171
rect 11529 6137 11563 6171
rect 14442 6137 14476 6171
rect 16405 6137 16439 6171
rect 5825 6069 5859 6103
rect 6285 6069 6319 6103
rect 10701 6069 10735 6103
rect 11161 6069 11195 6103
rect 12449 6069 12483 6103
rect 15577 6069 15611 6103
rect 16497 6069 16531 6103
rect 17417 6069 17451 6103
rect 3157 5865 3191 5899
rect 3249 5865 3283 5899
rect 4077 5865 4111 5899
rect 8861 5865 8895 5899
rect 17877 5865 17911 5899
rect 6552 5797 6586 5831
rect 11621 5797 11655 5831
rect 11713 5797 11747 5831
rect 12633 5797 12667 5831
rect 13360 5797 13394 5831
rect 16589 5797 16623 5831
rect 1777 5729 1811 5763
rect 4445 5729 4479 5763
rect 5549 5729 5583 5763
rect 6285 5729 6319 5763
rect 8769 5729 8803 5763
rect 9945 5729 9979 5763
rect 15485 5729 15519 5763
rect 16681 5729 16715 5763
rect 17785 5729 17819 5763
rect 1961 5661 1995 5695
rect 3433 5661 3467 5695
rect 4537 5661 4571 5695
rect 4629 5661 4663 5695
rect 8401 5661 8435 5695
rect 9689 5661 9723 5695
rect 13093 5661 13127 5695
rect 16773 5661 16807 5695
rect 17969 5661 18003 5695
rect 2789 5593 2823 5627
rect 14473 5593 14507 5627
rect 5733 5525 5767 5559
rect 7665 5525 7699 5559
rect 11069 5525 11103 5559
rect 15669 5525 15703 5559
rect 16221 5525 16255 5559
rect 17417 5525 17451 5559
rect 1869 5321 1903 5355
rect 3709 5321 3743 5355
rect 9505 5321 9539 5355
rect 15485 5321 15519 5355
rect 16681 5321 16715 5355
rect 6285 5253 6319 5287
rect 7297 5253 7331 5287
rect 11989 5253 12023 5287
rect 12633 5253 12667 5287
rect 4353 5185 4387 5219
rect 10149 5185 10183 5219
rect 13277 5185 13311 5219
rect 14289 5185 14323 5219
rect 16129 5185 16163 5219
rect 17233 5185 17267 5219
rect 1685 5117 1719 5151
rect 2615 5117 2649 5151
rect 4077 5117 4111 5151
rect 4905 5117 4939 5151
rect 6837 5117 6871 5151
rect 7205 5117 7239 5151
rect 8125 5117 8159 5151
rect 10416 5117 10450 5151
rect 12173 5117 12207 5151
rect 12449 5117 12483 5151
rect 14749 5117 14783 5151
rect 15853 5117 15887 5151
rect 17049 5117 17083 5151
rect 2881 5049 2915 5083
rect 5150 5049 5184 5083
rect 8392 5049 8426 5083
rect 13369 5049 13403 5083
rect 15945 5049 15979 5083
rect 4169 4981 4203 5015
rect 11529 4981 11563 5015
rect 14933 4981 14967 5015
rect 17141 4981 17175 5015
rect 1869 4777 1903 4811
rect 2605 4777 2639 4811
rect 5641 4777 5675 4811
rect 9045 4777 9079 4811
rect 9689 4777 9723 4811
rect 16865 4777 16899 4811
rect 17233 4777 17267 4811
rect 11805 4709 11839 4743
rect 11897 4709 11931 4743
rect 13737 4709 13771 4743
rect 13829 4709 13863 4743
rect 15485 4709 15519 4743
rect 17325 4709 17359 4743
rect 1685 4641 1719 4675
rect 2421 4641 2455 4675
rect 3157 4641 3191 4675
rect 4813 4641 4847 4675
rect 4905 4641 4939 4675
rect 6009 4641 6043 4675
rect 6101 4641 6135 4675
rect 6929 4641 6963 4675
rect 7932 4641 7966 4675
rect 10701 4641 10735 4675
rect 5089 4573 5123 4607
rect 6193 4573 6227 4607
rect 7665 4573 7699 4607
rect 10333 4573 10367 4607
rect 12817 4573 12851 4607
rect 14749 4573 14783 4607
rect 15393 4573 15427 4607
rect 15669 4573 15703 4607
rect 17509 4573 17543 4607
rect 3341 4437 3375 4471
rect 4445 4437 4479 4471
rect 7113 4437 7147 4471
rect 10793 4437 10827 4471
rect 1869 4233 1903 4267
rect 3985 4233 4019 4267
rect 9505 4233 9539 4267
rect 9045 4165 9079 4199
rect 4445 4097 4479 4131
rect 4629 4097 4663 4131
rect 5641 4097 5675 4131
rect 5825 4097 5859 4131
rect 6837 4097 6871 4131
rect 12909 4097 12943 4131
rect 13737 4097 13771 4131
rect 14933 4097 14967 4131
rect 16129 4097 16163 4131
rect 17141 4097 17175 4131
rect 1685 4029 1719 4063
rect 2421 4029 2455 4063
rect 3157 4029 3191 4063
rect 9413 4029 9447 4063
rect 10241 4029 10275 4063
rect 5549 3961 5583 3995
rect 7104 3961 7138 3995
rect 10508 3961 10542 3995
rect 13001 3961 13035 3995
rect 14473 3961 14507 3995
rect 14565 3961 14599 3995
rect 16221 3961 16255 3995
rect 2605 3893 2639 3927
rect 3341 3893 3375 3927
rect 4353 3893 4387 3927
rect 5181 3893 5215 3927
rect 8217 3893 8251 3927
rect 11621 3893 11655 3927
rect 7297 3689 7331 3723
rect 7757 3689 7791 3723
rect 8861 3689 8895 3723
rect 16865 3689 16899 3723
rect 6184 3621 6218 3655
rect 11437 3621 11471 3655
rect 13001 3621 13035 3655
rect 15485 3621 15519 3655
rect 16405 3621 16439 3655
rect 17233 3621 17267 3655
rect 1685 3553 1719 3587
rect 2697 3553 2731 3587
rect 4077 3553 4111 3587
rect 4344 3553 4378 3587
rect 8769 3553 8803 3587
rect 10425 3553 10459 3587
rect 14473 3553 14507 3587
rect 2973 3485 3007 3519
rect 5917 3485 5951 3519
rect 10793 3485 10827 3519
rect 11345 3485 11379 3519
rect 11713 3485 11747 3519
rect 12909 3485 12943 3519
rect 13461 3485 13495 3519
rect 15393 3485 15427 3519
rect 17325 3485 17359 3519
rect 17509 3485 17543 3519
rect 5457 3417 5491 3451
rect 8401 3417 8435 3451
rect 10057 3417 10091 3451
rect 1869 3349 1903 3383
rect 14657 3349 14691 3383
rect 5457 3145 5491 3179
rect 17417 3145 17451 3179
rect 6193 3077 6227 3111
rect 4445 3009 4479 3043
rect 11345 3009 11379 3043
rect 12541 3009 12575 3043
rect 14105 3009 14139 3043
rect 14933 3009 14967 3043
rect 16497 3009 16531 3043
rect 1501 2941 1535 2975
rect 2421 2941 2455 2975
rect 3341 2941 3375 2975
rect 4261 2941 4295 2975
rect 5273 2941 5307 2975
rect 6009 2941 6043 2975
rect 6837 2941 6871 2975
rect 7205 2941 7239 2975
rect 8068 2941 8102 2975
rect 17233 2941 17267 2975
rect 1777 2873 1811 2907
rect 2697 2873 2731 2907
rect 3617 2873 3651 2907
rect 8769 2873 8803 2907
rect 8861 2873 8895 2907
rect 9781 2873 9815 2907
rect 10333 2873 10367 2907
rect 10425 2873 10459 2907
rect 12633 2873 12667 2907
rect 13553 2873 13587 2907
rect 14197 2873 14231 2907
rect 15669 2873 15703 2907
rect 15761 2873 15795 2907
rect 7297 2805 7331 2839
rect 8171 2805 8205 2839
rect 2697 2601 2731 2635
rect 3433 2601 3467 2635
rect 6285 2601 6319 2635
rect 16221 2601 16255 2635
rect 16957 2601 16991 2635
rect 17693 2601 17727 2635
rect 10241 2533 10275 2567
rect 10333 2533 10367 2567
rect 11253 2533 11287 2567
rect 13921 2533 13955 2567
rect 14841 2533 14875 2567
rect 1593 2465 1627 2499
rect 2513 2465 2547 2499
rect 3249 2465 3283 2499
rect 4077 2465 4111 2499
rect 4813 2465 4847 2499
rect 6101 2465 6135 2499
rect 7297 2465 7331 2499
rect 7665 2465 7699 2499
rect 8493 2465 8527 2499
rect 11805 2465 11839 2499
rect 13001 2465 13035 2499
rect 16037 2465 16071 2499
rect 16773 2465 16807 2499
rect 17509 2465 17543 2499
rect 1777 2397 1811 2431
rect 13829 2397 13863 2431
rect 6929 2329 6963 2363
rect 8125 2329 8159 2363
rect 4261 2261 4295 2295
rect 4997 2261 5031 2295
rect 8585 2261 8619 2295
rect 11989 2261 12023 2295
rect 13185 2261 13219 2295
<< metal1 >>
rect 3602 15240 3608 15292
rect 3660 15280 3666 15292
rect 5626 15280 5632 15292
rect 3660 15252 5632 15280
rect 3660 15240 3666 15252
rect 5626 15240 5632 15252
rect 5684 15240 5690 15292
rect 12066 15172 12072 15224
rect 12124 15212 12130 15224
rect 15930 15212 15936 15224
rect 12124 15184 15936 15212
rect 12124 15172 12130 15184
rect 15930 15172 15936 15184
rect 15988 15172 15994 15224
rect 3510 14764 3516 14816
rect 3568 14804 3574 14816
rect 8754 14804 8760 14816
rect 3568 14776 8760 14804
rect 3568 14764 3574 14776
rect 8754 14764 8760 14776
rect 8812 14764 8818 14816
rect 1104 14714 18860 14736
rect 1104 14662 6912 14714
rect 6964 14662 6976 14714
rect 7028 14662 7040 14714
rect 7092 14662 7104 14714
rect 7156 14662 12843 14714
rect 12895 14662 12907 14714
rect 12959 14662 12971 14714
rect 13023 14662 13035 14714
rect 13087 14662 18860 14714
rect 1104 14640 18860 14662
rect 1578 14560 1584 14612
rect 1636 14600 1642 14612
rect 1949 14603 2007 14609
rect 1949 14600 1961 14603
rect 1636 14572 1961 14600
rect 1636 14560 1642 14572
rect 1949 14569 1961 14572
rect 1995 14569 2007 14603
rect 1949 14563 2007 14569
rect 2222 14560 2228 14612
rect 2280 14600 2286 14612
rect 2685 14603 2743 14609
rect 2685 14600 2697 14603
rect 2280 14572 2697 14600
rect 2280 14560 2286 14572
rect 2685 14569 2697 14572
rect 2731 14569 2743 14603
rect 2685 14563 2743 14569
rect 14918 14532 14924 14544
rect 2516 14504 14924 14532
rect 2516 14473 2544 14504
rect 14918 14492 14924 14504
rect 14976 14492 14982 14544
rect 17034 14532 17040 14544
rect 15028 14504 17040 14532
rect 1765 14467 1823 14473
rect 1765 14433 1777 14467
rect 1811 14433 1823 14467
rect 1765 14427 1823 14433
rect 2501 14467 2559 14473
rect 2501 14433 2513 14467
rect 2547 14433 2559 14467
rect 2501 14427 2559 14433
rect 3237 14467 3295 14473
rect 3237 14433 3249 14467
rect 3283 14464 3295 14467
rect 9582 14464 9588 14476
rect 3283 14436 9588 14464
rect 3283 14433 3295 14436
rect 3237 14427 3295 14433
rect 1780 14396 1808 14427
rect 9582 14424 9588 14436
rect 9640 14464 9646 14476
rect 15028 14464 15056 14504
rect 17034 14492 17040 14504
rect 17092 14492 17098 14544
rect 15470 14464 15476 14476
rect 9640 14436 15056 14464
rect 15431 14436 15476 14464
rect 9640 14424 9646 14436
rect 15470 14424 15476 14436
rect 15528 14464 15534 14476
rect 15746 14464 15752 14476
rect 15528 14436 15752 14464
rect 15528 14424 15534 14436
rect 15746 14424 15752 14436
rect 15804 14424 15810 14476
rect 13722 14396 13728 14408
rect 1780 14368 13728 14396
rect 13722 14356 13728 14368
rect 13780 14356 13786 14408
rect 3252 14300 3556 14328
rect 1670 14220 1676 14272
rect 1728 14260 1734 14272
rect 3252 14260 3280 14300
rect 3418 14260 3424 14272
rect 1728 14232 3280 14260
rect 3379 14232 3424 14260
rect 1728 14220 1734 14232
rect 3418 14220 3424 14232
rect 3476 14220 3482 14272
rect 3528 14260 3556 14300
rect 15562 14260 15568 14272
rect 3528 14232 15568 14260
rect 15562 14220 15568 14232
rect 15620 14220 15626 14272
rect 15654 14220 15660 14272
rect 15712 14260 15718 14272
rect 15712 14232 15757 14260
rect 15712 14220 15718 14232
rect 1104 14170 18860 14192
rect 1104 14118 3947 14170
rect 3999 14118 4011 14170
rect 4063 14118 4075 14170
rect 4127 14118 4139 14170
rect 4191 14118 9878 14170
rect 9930 14118 9942 14170
rect 9994 14118 10006 14170
rect 10058 14118 10070 14170
rect 10122 14118 15808 14170
rect 15860 14118 15872 14170
rect 15924 14118 15936 14170
rect 15988 14118 16000 14170
rect 16052 14118 18860 14170
rect 1104 14096 18860 14118
rect 2866 14016 2872 14068
rect 2924 14056 2930 14068
rect 3329 14059 3387 14065
rect 3329 14056 3341 14059
rect 2924 14028 3341 14056
rect 2924 14016 2930 14028
rect 3329 14025 3341 14028
rect 3375 14025 3387 14059
rect 3329 14019 3387 14025
rect 3510 14016 3516 14068
rect 3568 14056 3574 14068
rect 5534 14056 5540 14068
rect 3568 14028 5540 14056
rect 3568 14016 3574 14028
rect 5534 14016 5540 14028
rect 5592 14016 5598 14068
rect 6914 14016 6920 14068
rect 6972 14056 6978 14068
rect 7009 14059 7067 14065
rect 7009 14056 7021 14059
rect 6972 14028 7021 14056
rect 6972 14016 6978 14028
rect 7009 14025 7021 14028
rect 7055 14025 7067 14059
rect 7009 14019 7067 14025
rect 1581 13991 1639 13997
rect 1581 13957 1593 13991
rect 1627 13988 1639 13991
rect 2038 13988 2044 14000
rect 1627 13960 2044 13988
rect 1627 13957 1639 13960
rect 1581 13951 1639 13957
rect 2038 13948 2044 13960
rect 2096 13948 2102 14000
rect 4614 13988 4620 14000
rect 2240 13960 4620 13988
rect 2240 13929 2268 13960
rect 4614 13948 4620 13960
rect 4672 13948 4678 14000
rect 13538 13948 13544 14000
rect 13596 13988 13602 14000
rect 14645 13991 14703 13997
rect 14645 13988 14657 13991
rect 13596 13960 14657 13988
rect 13596 13948 13602 13960
rect 14645 13957 14657 13960
rect 14691 13957 14703 13991
rect 14645 13951 14703 13957
rect 2225 13923 2283 13929
rect 2225 13889 2237 13923
rect 2271 13889 2283 13923
rect 13354 13920 13360 13932
rect 2225 13883 2283 13889
rect 3160 13892 13360 13920
rect 1486 13812 1492 13864
rect 1544 13852 1550 13864
rect 3160 13861 3188 13892
rect 13354 13880 13360 13892
rect 13412 13880 13418 13932
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 1544 13824 2053 13852
rect 1544 13812 1550 13824
rect 2041 13821 2053 13824
rect 2087 13821 2099 13855
rect 2041 13815 2099 13821
rect 3145 13855 3203 13861
rect 3145 13821 3157 13855
rect 3191 13821 3203 13855
rect 3145 13815 3203 13821
rect 5997 13855 6055 13861
rect 5997 13821 6009 13855
rect 6043 13852 6055 13855
rect 6086 13852 6092 13864
rect 6043 13824 6092 13852
rect 6043 13821 6055 13824
rect 5997 13815 6055 13821
rect 6086 13812 6092 13824
rect 6144 13812 6150 13864
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6196 13824 6837 13852
rect 290 13744 296 13796
rect 348 13784 354 13796
rect 3418 13784 3424 13796
rect 348 13756 3424 13784
rect 348 13744 354 13756
rect 3418 13744 3424 13756
rect 3476 13744 3482 13796
rect 5902 13744 5908 13796
rect 5960 13784 5966 13796
rect 6196 13784 6224 13824
rect 6825 13821 6837 13824
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 13449 13855 13507 13861
rect 13449 13821 13461 13855
rect 13495 13852 13507 13855
rect 14366 13852 14372 13864
rect 13495 13824 14372 13852
rect 13495 13821 13507 13824
rect 13449 13815 13507 13821
rect 14366 13812 14372 13824
rect 14424 13812 14430 13864
rect 14461 13855 14519 13861
rect 14461 13821 14473 13855
rect 14507 13852 14519 13855
rect 15102 13852 15108 13864
rect 14507 13824 15108 13852
rect 14507 13821 14519 13824
rect 14461 13815 14519 13821
rect 15102 13812 15108 13824
rect 15160 13812 15166 13864
rect 15565 13855 15623 13861
rect 15565 13821 15577 13855
rect 15611 13852 15623 13855
rect 16390 13852 16396 13864
rect 15611 13824 16396 13852
rect 15611 13821 15623 13824
rect 15565 13815 15623 13821
rect 16390 13812 16396 13824
rect 16448 13812 16454 13864
rect 5960 13756 6224 13784
rect 5960 13744 5966 13756
rect 7374 13744 7380 13796
rect 7432 13784 7438 13796
rect 9030 13784 9036 13796
rect 7432 13756 9036 13784
rect 7432 13744 7438 13756
rect 9030 13744 9036 13756
rect 9088 13744 9094 13796
rect 9306 13744 9312 13796
rect 9364 13784 9370 13796
rect 10318 13784 10324 13796
rect 9364 13756 10324 13784
rect 9364 13744 9370 13756
rect 10318 13744 10324 13756
rect 10376 13744 10382 13796
rect 11330 13744 11336 13796
rect 11388 13784 11394 13796
rect 11882 13784 11888 13796
rect 11388 13756 11888 13784
rect 11388 13744 11394 13756
rect 11882 13744 11888 13756
rect 11940 13744 11946 13796
rect 11974 13744 11980 13796
rect 12032 13784 12038 13796
rect 15654 13784 15660 13796
rect 12032 13756 12664 13784
rect 12032 13744 12038 13756
rect 1946 13716 1952 13728
rect 1907 13688 1952 13716
rect 1946 13676 1952 13688
rect 2004 13676 2010 13728
rect 6178 13716 6184 13728
rect 6139 13688 6184 13716
rect 6178 13676 6184 13688
rect 6236 13676 6242 13728
rect 11238 13676 11244 13728
rect 11296 13716 11302 13728
rect 11790 13716 11796 13728
rect 11296 13688 11796 13716
rect 11296 13676 11302 13688
rect 11790 13676 11796 13688
rect 11848 13676 11854 13728
rect 12636 13716 12664 13756
rect 13315 13756 15660 13784
rect 13315 13716 13343 13756
rect 15654 13744 15660 13756
rect 15712 13744 15718 13796
rect 13630 13716 13636 13728
rect 12636 13688 13343 13716
rect 13591 13688 13636 13716
rect 13630 13676 13636 13688
rect 13688 13676 13694 13728
rect 15286 13676 15292 13728
rect 15344 13716 15350 13728
rect 15749 13719 15807 13725
rect 15749 13716 15761 13719
rect 15344 13688 15761 13716
rect 15344 13676 15350 13688
rect 15749 13685 15761 13688
rect 15795 13685 15807 13719
rect 15749 13679 15807 13685
rect 1104 13626 18860 13648
rect 1104 13574 6912 13626
rect 6964 13574 6976 13626
rect 7028 13574 7040 13626
rect 7092 13574 7104 13626
rect 7156 13574 12843 13626
rect 12895 13574 12907 13626
rect 12959 13574 12971 13626
rect 13023 13574 13035 13626
rect 13087 13574 18860 13626
rect 1104 13552 18860 13574
rect 934 13472 940 13524
rect 992 13512 998 13524
rect 1673 13515 1731 13521
rect 1673 13512 1685 13515
rect 992 13484 1685 13512
rect 992 13472 998 13484
rect 1673 13481 1685 13484
rect 1719 13481 1731 13515
rect 1673 13475 1731 13481
rect 4798 13472 4804 13524
rect 4856 13512 4862 13524
rect 11974 13512 11980 13524
rect 4856 13484 11980 13512
rect 4856 13472 4862 13484
rect 11974 13472 11980 13484
rect 12032 13472 12038 13524
rect 13538 13512 13544 13524
rect 12084 13484 13544 13512
rect 1578 13404 1584 13456
rect 1636 13444 1642 13456
rect 2685 13447 2743 13453
rect 2685 13444 2697 13447
rect 1636 13416 2697 13444
rect 1636 13404 1642 13416
rect 2685 13413 2697 13416
rect 2731 13444 2743 13447
rect 2731 13416 4200 13444
rect 2731 13413 2743 13416
rect 2685 13407 2743 13413
rect 1489 13379 1547 13385
rect 1489 13345 1501 13379
rect 1535 13345 1547 13379
rect 1489 13339 1547 13345
rect 2593 13379 2651 13385
rect 2593 13345 2605 13379
rect 2639 13376 2651 13379
rect 2639 13348 3188 13376
rect 2639 13345 2651 13348
rect 2593 13339 2651 13345
rect 1504 13240 1532 13339
rect 2774 13308 2780 13320
rect 2735 13280 2780 13308
rect 2774 13268 2780 13280
rect 2832 13268 2838 13320
rect 3160 13240 3188 13348
rect 3234 13268 3240 13320
rect 3292 13308 3298 13320
rect 4065 13311 4123 13317
rect 4065 13308 4077 13311
rect 3292 13280 4077 13308
rect 3292 13268 3298 13280
rect 4065 13277 4077 13280
rect 4111 13277 4123 13311
rect 4172 13308 4200 13416
rect 4246 13404 4252 13456
rect 4304 13444 4310 13456
rect 12084 13444 12112 13484
rect 13538 13472 13544 13484
rect 13596 13472 13602 13524
rect 14918 13472 14924 13524
rect 14976 13512 14982 13524
rect 18966 13512 18972 13524
rect 14976 13484 18972 13512
rect 14976 13472 14982 13484
rect 18966 13472 18972 13484
rect 19024 13472 19030 13524
rect 18322 13444 18328 13456
rect 4304 13416 12112 13444
rect 17144 13416 18328 13444
rect 4304 13404 4310 13416
rect 15102 13336 15108 13388
rect 15160 13376 15166 13388
rect 15324 13379 15382 13385
rect 15324 13376 15336 13379
rect 15160 13348 15336 13376
rect 15160 13336 15166 13348
rect 15324 13345 15336 13348
rect 15370 13345 15382 13379
rect 15324 13339 15382 13345
rect 11974 13308 11980 13320
rect 4172 13280 11980 13308
rect 4065 13271 4123 13277
rect 11974 13268 11980 13280
rect 12032 13268 12038 13320
rect 13538 13268 13544 13320
rect 13596 13308 13602 13320
rect 13722 13308 13728 13320
rect 13596 13280 13728 13308
rect 13596 13268 13602 13280
rect 13722 13268 13728 13280
rect 13780 13308 13786 13320
rect 17144 13308 17172 13416
rect 18322 13404 18328 13416
rect 18380 13404 18386 13456
rect 17770 13336 17776 13388
rect 17828 13376 17834 13388
rect 17865 13379 17923 13385
rect 17865 13376 17877 13379
rect 17828 13348 17877 13376
rect 17828 13336 17834 13348
rect 17865 13345 17877 13348
rect 17911 13345 17923 13379
rect 17865 13339 17923 13345
rect 13780 13280 17172 13308
rect 17221 13311 17279 13317
rect 13780 13268 13786 13280
rect 17221 13277 17233 13311
rect 17267 13308 17279 13311
rect 17586 13308 17592 13320
rect 17267 13280 17592 13308
rect 17267 13277 17279 13280
rect 17221 13271 17279 13277
rect 17586 13268 17592 13280
rect 17644 13268 17650 13320
rect 4522 13240 4528 13252
rect 1504 13212 2544 13240
rect 3160 13212 4528 13240
rect 1854 13132 1860 13184
rect 1912 13172 1918 13184
rect 2225 13175 2283 13181
rect 2225 13172 2237 13175
rect 1912 13144 2237 13172
rect 1912 13132 1918 13144
rect 2225 13141 2237 13144
rect 2271 13141 2283 13175
rect 2516 13172 2544 13212
rect 4522 13200 4528 13212
rect 4580 13200 4586 13252
rect 11422 13200 11428 13252
rect 11480 13240 11486 13252
rect 17678 13240 17684 13252
rect 11480 13212 17684 13240
rect 11480 13200 11486 13212
rect 17678 13200 17684 13212
rect 17736 13200 17742 13252
rect 8110 13172 8116 13184
rect 2516 13144 8116 13172
rect 2225 13135 2283 13141
rect 8110 13132 8116 13144
rect 8168 13132 8174 13184
rect 10226 13132 10232 13184
rect 10284 13172 10290 13184
rect 12618 13172 12624 13184
rect 10284 13144 12624 13172
rect 10284 13132 10290 13144
rect 12618 13132 12624 13144
rect 12676 13132 12682 13184
rect 13814 13132 13820 13184
rect 13872 13172 13878 13184
rect 14642 13172 14648 13184
rect 13872 13144 14648 13172
rect 13872 13132 13878 13144
rect 14642 13132 14648 13144
rect 14700 13132 14706 13184
rect 15194 13132 15200 13184
rect 15252 13172 15258 13184
rect 15427 13175 15485 13181
rect 15427 13172 15439 13175
rect 15252 13144 15439 13172
rect 15252 13132 15258 13144
rect 15427 13141 15439 13144
rect 15473 13141 15485 13175
rect 15427 13135 15485 13141
rect 18049 13175 18107 13181
rect 18049 13141 18061 13175
rect 18095 13172 18107 13175
rect 18598 13172 18604 13184
rect 18095 13144 18604 13172
rect 18095 13141 18107 13144
rect 18049 13135 18107 13141
rect 18598 13132 18604 13144
rect 18656 13132 18662 13184
rect 1104 13082 18860 13104
rect 1104 13030 3947 13082
rect 3999 13030 4011 13082
rect 4063 13030 4075 13082
rect 4127 13030 4139 13082
rect 4191 13030 9878 13082
rect 9930 13030 9942 13082
rect 9994 13030 10006 13082
rect 10058 13030 10070 13082
rect 10122 13030 15808 13082
rect 15860 13030 15872 13082
rect 15924 13030 15936 13082
rect 15988 13030 16000 13082
rect 16052 13030 18860 13082
rect 1104 13008 18860 13030
rect 1489 12971 1547 12977
rect 1489 12937 1501 12971
rect 1535 12968 1547 12971
rect 1946 12968 1952 12980
rect 1535 12940 1952 12968
rect 1535 12937 1547 12940
rect 1489 12931 1547 12937
rect 1946 12928 1952 12940
rect 2004 12928 2010 12980
rect 5442 12928 5448 12980
rect 5500 12968 5506 12980
rect 15286 12968 15292 12980
rect 5500 12940 12388 12968
rect 5500 12928 5506 12940
rect 12360 12900 12388 12940
rect 12912 12940 15292 12968
rect 12912 12900 12940 12940
rect 15286 12928 15292 12940
rect 15344 12928 15350 12980
rect 13630 12900 13636 12912
rect 12360 12872 12940 12900
rect 13004 12872 13636 12900
rect 2130 12832 2136 12844
rect 2043 12804 2136 12832
rect 2130 12792 2136 12804
rect 2188 12832 2194 12844
rect 4522 12832 4528 12844
rect 2188 12804 2452 12832
rect 4483 12804 4528 12832
rect 2188 12792 2194 12804
rect 1854 12764 1860 12776
rect 1815 12736 1860 12764
rect 1854 12724 1860 12736
rect 1912 12724 1918 12776
rect 1946 12588 1952 12640
rect 2004 12628 2010 12640
rect 2424 12628 2452 12804
rect 4522 12792 4528 12804
rect 4580 12792 4586 12844
rect 6086 12832 6092 12844
rect 6047 12804 6092 12832
rect 6086 12792 6092 12804
rect 6144 12792 6150 12844
rect 8478 12832 8484 12844
rect 8439 12804 8484 12832
rect 8478 12792 8484 12804
rect 8536 12792 8542 12844
rect 8754 12792 8760 12844
rect 8812 12832 8818 12844
rect 13004 12832 13032 12872
rect 13630 12860 13636 12872
rect 13688 12860 13694 12912
rect 13722 12860 13728 12912
rect 13780 12900 13786 12912
rect 19610 12900 19616 12912
rect 13780 12872 19616 12900
rect 13780 12860 13786 12872
rect 19610 12860 19616 12872
rect 19668 12860 19674 12912
rect 8812 12804 13032 12832
rect 8812 12792 8818 12804
rect 13354 12792 13360 12844
rect 13412 12832 13418 12844
rect 13740 12832 13768 12860
rect 13412 12804 13768 12832
rect 13412 12792 13418 12804
rect 2685 12767 2743 12773
rect 2685 12733 2697 12767
rect 2731 12764 2743 12767
rect 2731 12736 3096 12764
rect 2731 12733 2743 12736
rect 2685 12727 2743 12733
rect 3068 12708 3096 12736
rect 3510 12724 3516 12776
rect 3568 12764 3574 12776
rect 4706 12764 4712 12776
rect 3568 12736 4712 12764
rect 3568 12724 3574 12736
rect 4706 12724 4712 12736
rect 4764 12724 4770 12776
rect 8018 12764 8024 12776
rect 7979 12736 8024 12764
rect 8018 12724 8024 12736
rect 8076 12724 8082 12776
rect 8110 12724 8116 12776
rect 8168 12764 8174 12776
rect 8168 12736 10180 12764
rect 8168 12724 8174 12736
rect 2774 12656 2780 12708
rect 2832 12696 2838 12708
rect 2930 12699 2988 12705
rect 2930 12696 2942 12699
rect 2832 12668 2942 12696
rect 2832 12656 2838 12668
rect 2930 12665 2942 12668
rect 2976 12665 2988 12699
rect 2930 12659 2988 12665
rect 3050 12656 3056 12708
rect 3108 12656 3114 12708
rect 10152 12696 10180 12736
rect 10594 12724 10600 12776
rect 10652 12764 10658 12776
rect 12472 12767 12530 12773
rect 12472 12764 12484 12767
rect 10652 12736 12484 12764
rect 10652 12724 10658 12736
rect 12472 12733 12484 12736
rect 12518 12733 12530 12767
rect 13116 12767 13174 12773
rect 13116 12764 13128 12767
rect 12472 12727 12530 12733
rect 12728 12736 13128 12764
rect 11422 12696 11428 12708
rect 10152 12668 11428 12696
rect 11422 12656 11428 12668
rect 11480 12656 11486 12708
rect 11698 12656 11704 12708
rect 11756 12696 11762 12708
rect 12728 12696 12756 12736
rect 13116 12733 13128 12736
rect 13162 12733 13174 12767
rect 13116 12727 13174 12733
rect 13262 12724 13268 12776
rect 13320 12724 13326 12776
rect 15264 12767 15322 12773
rect 15264 12733 15276 12767
rect 15310 12764 15322 12767
rect 15470 12764 15476 12776
rect 15310 12736 15476 12764
rect 15310 12733 15322 12736
rect 15264 12727 15322 12733
rect 15470 12724 15476 12736
rect 15528 12724 15534 12776
rect 16206 12764 16212 12776
rect 16167 12736 16212 12764
rect 16206 12724 16212 12736
rect 16264 12724 16270 12776
rect 16574 12724 16580 12776
rect 16632 12764 16638 12776
rect 17221 12767 17279 12773
rect 17221 12764 17233 12767
rect 16632 12736 17233 12764
rect 16632 12724 16638 12736
rect 17221 12733 17233 12736
rect 17267 12733 17279 12767
rect 17221 12727 17279 12733
rect 13280 12696 13308 12724
rect 11756 12668 12756 12696
rect 13096 12668 13308 12696
rect 11756 12656 11762 12668
rect 4065 12631 4123 12637
rect 4065 12628 4077 12631
rect 2004 12600 2049 12628
rect 2424 12600 4077 12628
rect 2004 12588 2010 12600
rect 4065 12597 4077 12600
rect 4111 12628 4123 12631
rect 4338 12628 4344 12640
rect 4111 12600 4344 12628
rect 4111 12597 4123 12600
rect 4065 12591 4123 12597
rect 4338 12588 4344 12600
rect 4396 12588 4402 12640
rect 5537 12631 5595 12637
rect 5537 12597 5549 12631
rect 5583 12628 5595 12631
rect 5718 12628 5724 12640
rect 5583 12600 5724 12628
rect 5583 12597 5595 12600
rect 5537 12591 5595 12597
rect 5718 12588 5724 12600
rect 5776 12588 5782 12640
rect 5810 12588 5816 12640
rect 5868 12628 5874 12640
rect 5905 12631 5963 12637
rect 5905 12628 5917 12631
rect 5868 12600 5917 12628
rect 5868 12588 5874 12600
rect 5905 12597 5917 12600
rect 5951 12597 5963 12631
rect 5905 12591 5963 12597
rect 5994 12588 6000 12640
rect 6052 12628 6058 12640
rect 6825 12631 6883 12637
rect 6052 12600 6097 12628
rect 6052 12588 6058 12600
rect 6825 12597 6837 12631
rect 6871 12628 6883 12631
rect 7282 12628 7288 12640
rect 6871 12600 7288 12628
rect 6871 12597 6883 12600
rect 6825 12591 6883 12597
rect 7282 12588 7288 12600
rect 7340 12588 7346 12640
rect 12575 12631 12633 12637
rect 12575 12597 12587 12631
rect 12621 12628 12633 12631
rect 13096 12628 13124 12668
rect 12621 12600 13124 12628
rect 13219 12631 13277 12637
rect 12621 12597 12633 12600
rect 12575 12591 12633 12597
rect 13219 12597 13231 12631
rect 13265 12628 13277 12631
rect 13354 12628 13360 12640
rect 13265 12600 13360 12628
rect 13265 12597 13277 12600
rect 13219 12591 13277 12597
rect 13354 12588 13360 12600
rect 13412 12588 13418 12640
rect 15378 12637 15384 12640
rect 15335 12631 15384 12637
rect 15335 12597 15347 12631
rect 15381 12597 15384 12631
rect 15335 12591 15384 12597
rect 15378 12588 15384 12591
rect 15436 12588 15442 12640
rect 16393 12631 16451 12637
rect 16393 12597 16405 12631
rect 16439 12628 16451 12631
rect 17218 12628 17224 12640
rect 16439 12600 17224 12628
rect 16439 12597 16451 12600
rect 16393 12591 16451 12597
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 17405 12631 17463 12637
rect 17405 12597 17417 12631
rect 17451 12628 17463 12631
rect 18138 12628 18144 12640
rect 17451 12600 18144 12628
rect 17451 12597 17463 12600
rect 17405 12591 17463 12597
rect 18138 12588 18144 12600
rect 18196 12588 18202 12640
rect 1104 12538 18860 12560
rect 1104 12486 6912 12538
rect 6964 12486 6976 12538
rect 7028 12486 7040 12538
rect 7092 12486 7104 12538
rect 7156 12486 12843 12538
rect 12895 12486 12907 12538
rect 12959 12486 12971 12538
rect 13023 12486 13035 12538
rect 13087 12486 18860 12538
rect 1104 12464 18860 12486
rect 1946 12384 1952 12436
rect 2004 12424 2010 12436
rect 2225 12427 2283 12433
rect 2225 12424 2237 12427
rect 2004 12396 2237 12424
rect 2004 12384 2010 12396
rect 2225 12393 2237 12396
rect 2271 12393 2283 12427
rect 2225 12387 2283 12393
rect 2958 12384 2964 12436
rect 3016 12424 3022 12436
rect 4433 12427 4491 12433
rect 4433 12424 4445 12427
rect 3016 12396 4445 12424
rect 3016 12384 3022 12396
rect 4433 12393 4445 12396
rect 4479 12393 4491 12427
rect 5905 12427 5963 12433
rect 4433 12387 4491 12393
rect 4540 12396 5856 12424
rect 4540 12356 4568 12396
rect 1504 12328 4568 12356
rect 1504 12297 1532 12328
rect 4614 12316 4620 12368
rect 4672 12356 4678 12368
rect 4770 12359 4828 12365
rect 4770 12356 4782 12359
rect 4672 12328 4782 12356
rect 4672 12316 4678 12328
rect 4770 12325 4782 12328
rect 4816 12325 4828 12359
rect 5828 12356 5856 12396
rect 5905 12393 5917 12427
rect 5951 12424 5963 12427
rect 6086 12424 6092 12436
rect 5951 12396 6092 12424
rect 5951 12393 5963 12396
rect 5905 12387 5963 12393
rect 6086 12384 6092 12396
rect 6144 12424 6150 12436
rect 6546 12424 6552 12436
rect 6144 12396 6552 12424
rect 6144 12384 6150 12396
rect 6546 12384 6552 12396
rect 6604 12384 6610 12436
rect 11514 12384 11520 12436
rect 11572 12424 11578 12436
rect 11572 12396 15608 12424
rect 11572 12384 11578 12396
rect 6270 12356 6276 12368
rect 5828 12328 6276 12356
rect 4770 12319 4828 12325
rect 6270 12316 6276 12328
rect 6328 12316 6334 12368
rect 8573 12359 8631 12365
rect 8573 12356 8585 12359
rect 6564 12328 8585 12356
rect 1489 12291 1547 12297
rect 1489 12257 1501 12291
rect 1535 12257 1547 12291
rect 1489 12251 1547 12257
rect 2406 12248 2412 12300
rect 2464 12288 2470 12300
rect 2593 12291 2651 12297
rect 2593 12288 2605 12291
rect 2464 12260 2605 12288
rect 2464 12248 2470 12260
rect 2593 12257 2605 12260
rect 2639 12288 2651 12291
rect 4246 12288 4252 12300
rect 2639 12260 4252 12288
rect 2639 12257 2651 12260
rect 2593 12251 2651 12257
rect 4246 12248 4252 12260
rect 4304 12248 4310 12300
rect 4433 12291 4491 12297
rect 4433 12257 4445 12291
rect 4479 12288 4491 12291
rect 4522 12288 4528 12300
rect 4479 12260 4528 12288
rect 4479 12257 4491 12260
rect 4433 12251 4491 12257
rect 4522 12248 4528 12260
rect 4580 12248 4586 12300
rect 6564 12288 6592 12328
rect 8573 12325 8585 12328
rect 8619 12356 8631 12359
rect 9122 12356 9128 12368
rect 8619 12328 9128 12356
rect 8619 12325 8631 12328
rect 8573 12319 8631 12325
rect 9122 12316 9128 12328
rect 9180 12316 9186 12368
rect 6638 12297 6644 12300
rect 4632 12260 6592 12288
rect 2314 12180 2320 12232
rect 2372 12220 2378 12232
rect 2685 12223 2743 12229
rect 2685 12220 2697 12223
rect 2372 12192 2697 12220
rect 2372 12180 2378 12192
rect 2685 12189 2697 12192
rect 2731 12189 2743 12223
rect 2685 12183 2743 12189
rect 2774 12180 2780 12232
rect 2832 12220 2838 12232
rect 2832 12192 2877 12220
rect 2832 12180 2838 12192
rect 3050 12180 3056 12232
rect 3108 12220 3114 12232
rect 3418 12220 3424 12232
rect 3108 12192 3424 12220
rect 3108 12180 3114 12192
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 4062 12180 4068 12232
rect 4120 12220 4126 12232
rect 4632 12220 4660 12260
rect 6632 12251 6644 12297
rect 6696 12288 6702 12300
rect 6696 12260 6732 12288
rect 6638 12248 6644 12251
rect 6696 12248 6702 12260
rect 7650 12248 7656 12300
rect 7708 12288 7714 12300
rect 9398 12288 9404 12300
rect 7708 12260 9404 12288
rect 7708 12248 7714 12260
rect 9398 12248 9404 12260
rect 9456 12248 9462 12300
rect 11606 12248 11612 12300
rect 11664 12288 11670 12300
rect 12288 12291 12346 12297
rect 12288 12288 12300 12291
rect 11664 12260 12300 12288
rect 11664 12248 11670 12260
rect 12288 12257 12300 12260
rect 12334 12257 12346 12291
rect 12288 12251 12346 12257
rect 12526 12248 12532 12300
rect 12584 12288 12590 12300
rect 13300 12291 13358 12297
rect 13300 12288 13312 12291
rect 12584 12260 13312 12288
rect 12584 12248 12590 12260
rect 13300 12257 13312 12260
rect 13346 12257 13358 12291
rect 13300 12251 13358 12257
rect 14252 12291 14310 12297
rect 14252 12257 14264 12291
rect 14298 12288 14310 12291
rect 14734 12288 14740 12300
rect 14298 12260 14740 12288
rect 14298 12257 14310 12260
rect 14252 12251 14310 12257
rect 14734 12248 14740 12260
rect 14792 12248 14798 12300
rect 15580 12297 15608 12396
rect 15565 12291 15623 12297
rect 15565 12257 15577 12291
rect 15611 12257 15623 12291
rect 15565 12251 15623 12257
rect 16393 12291 16451 12297
rect 16393 12257 16405 12291
rect 16439 12257 16451 12291
rect 17126 12288 17132 12300
rect 17087 12260 17132 12288
rect 16393 12251 16451 12257
rect 4120 12192 4660 12220
rect 4120 12180 4126 12192
rect 6086 12180 6092 12232
rect 6144 12220 6150 12232
rect 6362 12220 6368 12232
rect 6144 12192 6368 12220
rect 6144 12180 6150 12192
rect 6362 12180 6368 12192
rect 6420 12180 6426 12232
rect 8662 12220 8668 12232
rect 8623 12192 8668 12220
rect 8662 12180 8668 12192
rect 8720 12180 8726 12232
rect 8754 12180 8760 12232
rect 8812 12220 8818 12232
rect 8812 12192 8857 12220
rect 8812 12180 8818 12192
rect 9306 12180 9312 12232
rect 9364 12220 9370 12232
rect 15286 12220 15292 12232
rect 9364 12192 15292 12220
rect 9364 12180 9370 12192
rect 15286 12180 15292 12192
rect 15344 12180 15350 12232
rect 1673 12155 1731 12161
rect 1673 12121 1685 12155
rect 1719 12152 1731 12155
rect 1719 12124 2360 12152
rect 1719 12121 1731 12124
rect 1673 12115 1731 12121
rect 2332 12084 2360 12124
rect 3602 12112 3608 12164
rect 3660 12152 3666 12164
rect 3878 12152 3884 12164
rect 3660 12124 3884 12152
rect 3660 12112 3666 12124
rect 3878 12112 3884 12124
rect 3936 12112 3942 12164
rect 9398 12112 9404 12164
rect 9456 12152 9462 12164
rect 13906 12152 13912 12164
rect 9456 12124 13912 12152
rect 9456 12112 9462 12124
rect 13906 12112 13912 12124
rect 13964 12112 13970 12164
rect 13998 12112 14004 12164
rect 14056 12152 14062 12164
rect 16408 12152 16436 12251
rect 17126 12248 17132 12260
rect 17184 12248 17190 12300
rect 17862 12288 17868 12300
rect 17823 12260 17868 12288
rect 17862 12248 17868 12260
rect 17920 12248 17926 12300
rect 14056 12124 16436 12152
rect 17313 12155 17371 12161
rect 14056 12112 14062 12124
rect 17313 12121 17325 12155
rect 17359 12152 17371 12155
rect 19150 12152 19156 12164
rect 17359 12124 19156 12152
rect 17359 12121 17371 12124
rect 17313 12115 17371 12121
rect 19150 12112 19156 12124
rect 19208 12112 19214 12164
rect 3050 12084 3056 12096
rect 2332 12056 3056 12084
rect 3050 12044 3056 12056
rect 3108 12044 3114 12096
rect 3326 12044 3332 12096
rect 3384 12084 3390 12096
rect 5994 12084 6000 12096
rect 3384 12056 6000 12084
rect 3384 12044 3390 12056
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 6730 12044 6736 12096
rect 6788 12084 6794 12096
rect 7745 12087 7803 12093
rect 7745 12084 7757 12087
rect 6788 12056 7757 12084
rect 6788 12044 6794 12056
rect 7745 12053 7757 12056
rect 7791 12053 7803 12087
rect 7745 12047 7803 12053
rect 8110 12044 8116 12096
rect 8168 12084 8174 12096
rect 8205 12087 8263 12093
rect 8205 12084 8217 12087
rect 8168 12056 8217 12084
rect 8168 12044 8174 12056
rect 8205 12053 8217 12056
rect 8251 12053 8263 12087
rect 8205 12047 8263 12053
rect 12250 12044 12256 12096
rect 12308 12084 12314 12096
rect 12391 12087 12449 12093
rect 12391 12084 12403 12087
rect 12308 12056 12403 12084
rect 12308 12044 12314 12056
rect 12391 12053 12403 12056
rect 12437 12084 12449 12087
rect 12437 12056 12493 12084
rect 12437 12053 12449 12056
rect 12391 12047 12449 12053
rect 12710 12044 12716 12096
rect 12768 12084 12774 12096
rect 13403 12087 13461 12093
rect 13403 12084 13415 12087
rect 12768 12056 13415 12084
rect 12768 12044 12774 12056
rect 13403 12053 13415 12056
rect 13449 12053 13461 12087
rect 13403 12047 13461 12053
rect 14323 12087 14381 12093
rect 14323 12053 14335 12087
rect 14369 12084 14381 12087
rect 14550 12084 14556 12096
rect 14369 12056 14556 12084
rect 14369 12053 14381 12056
rect 14323 12047 14381 12053
rect 14550 12044 14556 12056
rect 14608 12044 14614 12096
rect 15749 12087 15807 12093
rect 15749 12053 15761 12087
rect 15795 12084 15807 12087
rect 16114 12084 16120 12096
rect 15795 12056 16120 12084
rect 15795 12053 15807 12056
rect 15749 12047 15807 12053
rect 16114 12044 16120 12056
rect 16172 12044 16178 12096
rect 16577 12087 16635 12093
rect 16577 12053 16589 12087
rect 16623 12084 16635 12087
rect 17770 12084 17776 12096
rect 16623 12056 17776 12084
rect 16623 12053 16635 12056
rect 16577 12047 16635 12053
rect 17770 12044 17776 12056
rect 17828 12044 17834 12096
rect 18046 12084 18052 12096
rect 18007 12056 18052 12084
rect 18046 12044 18052 12056
rect 18104 12044 18110 12096
rect 1104 11994 18860 12016
rect 1104 11942 3947 11994
rect 3999 11942 4011 11994
rect 4063 11942 4075 11994
rect 4127 11942 4139 11994
rect 4191 11942 9878 11994
rect 9930 11942 9942 11994
rect 9994 11942 10006 11994
rect 10058 11942 10070 11994
rect 10122 11942 15808 11994
rect 15860 11942 15872 11994
rect 15924 11942 15936 11994
rect 15988 11942 16000 11994
rect 16052 11942 18860 11994
rect 1104 11920 18860 11942
rect 4614 11840 4620 11892
rect 4672 11880 4678 11892
rect 4893 11883 4951 11889
rect 4893 11880 4905 11883
rect 4672 11852 4905 11880
rect 4672 11840 4678 11852
rect 4893 11849 4905 11852
rect 4939 11849 4951 11883
rect 4893 11843 4951 11849
rect 5810 11840 5816 11892
rect 5868 11880 5874 11892
rect 5868 11852 7880 11880
rect 5868 11840 5874 11852
rect 2682 11772 2688 11824
rect 2740 11812 2746 11824
rect 3142 11812 3148 11824
rect 2740 11784 3148 11812
rect 2740 11772 2746 11784
rect 3142 11772 3148 11784
rect 3200 11772 3206 11824
rect 3510 11772 3516 11824
rect 3568 11772 3574 11824
rect 2774 11704 2780 11756
rect 2832 11744 2838 11756
rect 2869 11747 2927 11753
rect 2869 11744 2881 11747
rect 2832 11716 2881 11744
rect 2832 11704 2838 11716
rect 2869 11713 2881 11716
rect 2915 11744 2927 11747
rect 3528 11744 3556 11772
rect 2915 11716 3556 11744
rect 2915 11713 2927 11716
rect 2869 11707 2927 11713
rect 5350 11704 5356 11756
rect 5408 11744 5414 11756
rect 5810 11744 5816 11756
rect 5408 11716 5816 11744
rect 5408 11704 5414 11716
rect 5810 11704 5816 11716
rect 5868 11704 5874 11756
rect 5997 11747 6055 11753
rect 5997 11713 6009 11747
rect 6043 11744 6055 11747
rect 6086 11744 6092 11756
rect 6043 11716 6092 11744
rect 6043 11713 6055 11716
rect 5997 11707 6055 11713
rect 6086 11704 6092 11716
rect 6144 11704 6150 11756
rect 6181 11747 6239 11753
rect 6181 11713 6193 11747
rect 6227 11744 6239 11747
rect 6730 11744 6736 11756
rect 6227 11716 6736 11744
rect 6227 11713 6239 11716
rect 6181 11707 6239 11713
rect 6730 11704 6736 11716
rect 6788 11704 6794 11756
rect 1578 11676 1584 11688
rect 1539 11648 1584 11676
rect 1578 11636 1584 11648
rect 1636 11636 1642 11688
rect 2958 11636 2964 11688
rect 3016 11676 3022 11688
rect 3513 11679 3571 11685
rect 3513 11676 3525 11679
rect 3016 11648 3525 11676
rect 3016 11636 3022 11648
rect 3513 11645 3525 11648
rect 3559 11645 3571 11679
rect 3513 11639 3571 11645
rect 3780 11679 3838 11685
rect 3780 11645 3792 11679
rect 3826 11676 3838 11679
rect 4338 11676 4344 11688
rect 3826 11648 4344 11676
rect 3826 11645 3838 11648
rect 3780 11639 3838 11645
rect 4338 11636 4344 11648
rect 4396 11636 4402 11688
rect 6362 11636 6368 11688
rect 6420 11676 6426 11688
rect 6825 11679 6883 11685
rect 6825 11676 6837 11679
rect 6420 11648 6837 11676
rect 6420 11636 6426 11648
rect 6825 11645 6837 11648
rect 6871 11645 6883 11679
rect 7852 11676 7880 11852
rect 8662 11840 8668 11892
rect 8720 11880 8726 11892
rect 8757 11883 8815 11889
rect 8757 11880 8769 11883
rect 8720 11852 8769 11880
rect 8720 11840 8726 11852
rect 8757 11849 8769 11852
rect 8803 11849 8815 11883
rect 8757 11843 8815 11849
rect 8846 11840 8852 11892
rect 8904 11880 8910 11892
rect 8904 11852 13216 11880
rect 8904 11840 8910 11852
rect 13188 11812 13216 11852
rect 13262 11840 13268 11892
rect 13320 11880 13326 11892
rect 13538 11880 13544 11892
rect 13320 11852 13544 11880
rect 13320 11840 13326 11852
rect 13538 11840 13544 11852
rect 13596 11840 13602 11892
rect 13906 11840 13912 11892
rect 13964 11880 13970 11892
rect 16758 11880 16764 11892
rect 13964 11852 16764 11880
rect 13964 11840 13970 11852
rect 16758 11840 16764 11852
rect 16816 11840 16822 11892
rect 16298 11812 16304 11824
rect 13188 11784 16304 11812
rect 16298 11772 16304 11784
rect 16356 11772 16362 11824
rect 16669 11815 16727 11821
rect 16669 11781 16681 11815
rect 16715 11812 16727 11815
rect 19610 11812 19616 11824
rect 16715 11784 19616 11812
rect 16715 11781 16727 11784
rect 16669 11775 16727 11781
rect 19610 11772 19616 11784
rect 19668 11772 19674 11824
rect 9306 11744 9312 11756
rect 9267 11716 9312 11744
rect 9306 11704 9312 11716
rect 9364 11704 9370 11756
rect 12342 11704 12348 11756
rect 12400 11744 12406 11756
rect 13449 11747 13507 11753
rect 13449 11744 13461 11747
rect 12400 11716 13461 11744
rect 12400 11704 12406 11716
rect 13449 11713 13461 11716
rect 13495 11713 13507 11747
rect 13630 11744 13636 11756
rect 13591 11716 13636 11744
rect 13449 11707 13507 11713
rect 13630 11704 13636 11716
rect 13688 11704 13694 11756
rect 15654 11744 15660 11756
rect 14292 11716 15516 11744
rect 15615 11716 15660 11744
rect 14292 11676 14320 11716
rect 7852 11648 14320 11676
rect 14369 11679 14427 11685
rect 6825 11639 6883 11645
rect 14369 11645 14381 11679
rect 14415 11645 14427 11679
rect 15488 11676 15516 11716
rect 15654 11704 15660 11716
rect 15712 11704 15718 11756
rect 16850 11744 16856 11756
rect 16316 11716 16856 11744
rect 16316 11676 16344 11716
rect 16850 11704 16856 11716
rect 16908 11704 16914 11756
rect 16482 11676 16488 11688
rect 15488 11648 16344 11676
rect 16443 11648 16488 11676
rect 14369 11639 14427 11645
rect 2222 11568 2228 11620
rect 2280 11608 2286 11620
rect 2685 11611 2743 11617
rect 2685 11608 2697 11611
rect 2280 11580 2697 11608
rect 2280 11568 2286 11580
rect 2685 11577 2697 11580
rect 2731 11608 2743 11611
rect 2731 11580 3464 11608
rect 2731 11577 2743 11580
rect 2685 11571 2743 11577
rect 1762 11540 1768 11552
rect 1723 11512 1768 11540
rect 1762 11500 1768 11512
rect 1820 11500 1826 11552
rect 1854 11500 1860 11552
rect 1912 11540 1918 11552
rect 2317 11543 2375 11549
rect 2317 11540 2329 11543
rect 1912 11512 2329 11540
rect 1912 11500 1918 11512
rect 2317 11509 2329 11512
rect 2363 11509 2375 11543
rect 2317 11503 2375 11509
rect 2774 11500 2780 11552
rect 2832 11540 2838 11552
rect 3436 11540 3464 11580
rect 5626 11568 5632 11620
rect 5684 11608 5690 11620
rect 5905 11611 5963 11617
rect 5905 11608 5917 11611
rect 5684 11580 5917 11608
rect 5684 11568 5690 11580
rect 5905 11577 5917 11580
rect 5951 11608 5963 11611
rect 5951 11580 6684 11608
rect 5951 11577 5963 11580
rect 5905 11571 5963 11577
rect 4430 11540 4436 11552
rect 2832 11512 2877 11540
rect 3436 11512 4436 11540
rect 2832 11500 2838 11512
rect 4430 11500 4436 11512
rect 4488 11500 4494 11552
rect 5534 11540 5540 11552
rect 5495 11512 5540 11540
rect 5534 11500 5540 11512
rect 5592 11500 5598 11552
rect 6656 11540 6684 11580
rect 6730 11568 6736 11620
rect 6788 11608 6794 11620
rect 7070 11611 7128 11617
rect 7070 11608 7082 11611
rect 6788 11580 7082 11608
rect 6788 11568 6794 11580
rect 7070 11577 7082 11580
rect 7116 11577 7128 11611
rect 13906 11608 13912 11620
rect 7070 11571 7128 11577
rect 7944 11580 13912 11608
rect 7944 11540 7972 11580
rect 13906 11568 13912 11580
rect 13964 11568 13970 11620
rect 14090 11568 14096 11620
rect 14148 11608 14154 11620
rect 14384 11608 14412 11639
rect 16482 11636 16488 11648
rect 16540 11636 16546 11688
rect 16758 11636 16764 11688
rect 16816 11676 16822 11688
rect 17221 11679 17279 11685
rect 17221 11676 17233 11679
rect 16816 11648 17233 11676
rect 16816 11636 16822 11648
rect 17221 11645 17233 11648
rect 17267 11676 17279 11679
rect 17954 11676 17960 11688
rect 17267 11648 17960 11676
rect 17267 11645 17279 11648
rect 17221 11639 17279 11645
rect 17954 11636 17960 11648
rect 18012 11636 18018 11688
rect 14148 11580 14412 11608
rect 15473 11611 15531 11617
rect 14148 11568 14154 11580
rect 15473 11577 15485 11611
rect 15519 11608 15531 11611
rect 16942 11608 16948 11620
rect 15519 11580 16948 11608
rect 15519 11577 15531 11580
rect 15473 11571 15531 11577
rect 16942 11568 16948 11580
rect 17000 11568 17006 11620
rect 8202 11540 8208 11552
rect 6656 11512 7972 11540
rect 8163 11512 8208 11540
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 8846 11500 8852 11552
rect 8904 11540 8910 11552
rect 9125 11543 9183 11549
rect 9125 11540 9137 11543
rect 8904 11512 9137 11540
rect 8904 11500 8910 11512
rect 9125 11509 9137 11512
rect 9171 11509 9183 11543
rect 9125 11503 9183 11509
rect 9214 11500 9220 11552
rect 9272 11540 9278 11552
rect 11146 11540 11152 11552
rect 9272 11512 9317 11540
rect 11107 11512 11152 11540
rect 9272 11500 9278 11512
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 12158 11500 12164 11552
rect 12216 11540 12222 11552
rect 12526 11540 12532 11552
rect 12216 11512 12532 11540
rect 12216 11500 12222 11512
rect 12526 11500 12532 11512
rect 12584 11500 12590 11552
rect 12989 11543 13047 11549
rect 12989 11509 13001 11543
rect 13035 11540 13047 11543
rect 13170 11540 13176 11552
rect 13035 11512 13176 11540
rect 13035 11509 13047 11512
rect 12989 11503 13047 11509
rect 13170 11500 13176 11512
rect 13228 11500 13234 11552
rect 13354 11540 13360 11552
rect 13315 11512 13360 11540
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 14274 11500 14280 11552
rect 14332 11540 14338 11552
rect 14553 11543 14611 11549
rect 14553 11540 14565 11543
rect 14332 11512 14565 11540
rect 14332 11500 14338 11512
rect 14553 11509 14565 11512
rect 14599 11509 14611 11543
rect 15102 11540 15108 11552
rect 15063 11512 15108 11540
rect 14553 11503 14611 11509
rect 15102 11500 15108 11512
rect 15160 11500 15166 11552
rect 15565 11543 15623 11549
rect 15565 11509 15577 11543
rect 15611 11540 15623 11543
rect 15746 11540 15752 11552
rect 15611 11512 15752 11540
rect 15611 11509 15623 11512
rect 15565 11503 15623 11509
rect 15746 11500 15752 11512
rect 15804 11500 15810 11552
rect 17405 11543 17463 11549
rect 17405 11509 17417 11543
rect 17451 11540 17463 11543
rect 17494 11540 17500 11552
rect 17451 11512 17500 11540
rect 17451 11509 17463 11512
rect 17405 11503 17463 11509
rect 17494 11500 17500 11512
rect 17552 11500 17558 11552
rect 1104 11450 18860 11472
rect 1104 11398 6912 11450
rect 6964 11398 6976 11450
rect 7028 11398 7040 11450
rect 7092 11398 7104 11450
rect 7156 11398 12843 11450
rect 12895 11398 12907 11450
rect 12959 11398 12971 11450
rect 13023 11398 13035 11450
rect 13087 11398 18860 11450
rect 1104 11376 18860 11398
rect 1486 11336 1492 11348
rect 1447 11308 1492 11336
rect 1486 11296 1492 11308
rect 1544 11296 1550 11348
rect 1854 11336 1860 11348
rect 1815 11308 1860 11336
rect 1854 11296 1860 11308
rect 1912 11296 1918 11348
rect 2685 11339 2743 11345
rect 2685 11305 2697 11339
rect 2731 11336 2743 11339
rect 2774 11336 2780 11348
rect 2731 11308 2780 11336
rect 2731 11305 2743 11308
rect 2685 11299 2743 11305
rect 2774 11296 2780 11308
rect 2832 11296 2838 11348
rect 5534 11296 5540 11348
rect 5592 11336 5598 11348
rect 5997 11339 6055 11345
rect 5997 11336 6009 11339
rect 5592 11308 6009 11336
rect 5592 11296 5598 11308
rect 5997 11305 6009 11308
rect 6043 11305 6055 11339
rect 14366 11336 14372 11348
rect 5997 11299 6055 11305
rect 6104 11308 14372 11336
rect 3142 11268 3148 11280
rect 3055 11240 3148 11268
rect 3142 11228 3148 11240
rect 3200 11268 3206 11280
rect 6104 11268 6132 11308
rect 14366 11296 14372 11308
rect 14424 11296 14430 11348
rect 14645 11339 14703 11345
rect 14645 11305 14657 11339
rect 14691 11305 14703 11339
rect 15746 11336 15752 11348
rect 15707 11308 15752 11336
rect 14645 11299 14703 11305
rect 7828 11271 7886 11277
rect 7828 11268 7840 11271
rect 3200 11240 6132 11268
rect 6196 11240 7840 11268
rect 3200 11228 3206 11240
rect 3053 11203 3111 11209
rect 3053 11169 3065 11203
rect 3099 11169 3111 11203
rect 3053 11163 3111 11169
rect 4709 11203 4767 11209
rect 4709 11169 4721 11203
rect 4755 11200 4767 11203
rect 5258 11200 5264 11212
rect 4755 11172 5264 11200
rect 4755 11169 4767 11172
rect 4709 11163 4767 11169
rect 1578 11092 1584 11144
rect 1636 11132 1642 11144
rect 1949 11135 2007 11141
rect 1949 11132 1961 11135
rect 1636 11104 1961 11132
rect 1636 11092 1642 11104
rect 1949 11101 1961 11104
rect 1995 11101 2007 11135
rect 2130 11132 2136 11144
rect 2091 11104 2136 11132
rect 1949 11095 2007 11101
rect 2130 11092 2136 11104
rect 2188 11092 2194 11144
rect 3068 11132 3096 11163
rect 5258 11160 5264 11172
rect 5316 11160 5322 11212
rect 5902 11200 5908 11212
rect 5863 11172 5908 11200
rect 5902 11160 5908 11172
rect 5960 11160 5966 11212
rect 3142 11132 3148 11144
rect 3068 11104 3148 11132
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 3326 11132 3332 11144
rect 3287 11104 3332 11132
rect 3326 11092 3332 11104
rect 3384 11092 3390 11144
rect 4798 11132 4804 11144
rect 4759 11104 4804 11132
rect 4798 11092 4804 11104
rect 4856 11092 4862 11144
rect 6196 11141 6224 11240
rect 7828 11237 7840 11240
rect 7874 11268 7886 11271
rect 8202 11268 8208 11280
rect 7874 11240 8208 11268
rect 7874 11237 7886 11240
rect 7828 11231 7886 11237
rect 8202 11228 8208 11240
rect 8260 11228 8266 11280
rect 8294 11228 8300 11280
rect 8352 11268 8358 11280
rect 9214 11268 9220 11280
rect 8352 11240 9220 11268
rect 8352 11228 8358 11240
rect 9214 11228 9220 11240
rect 9272 11228 9278 11280
rect 12066 11228 12072 11280
rect 12124 11268 12130 11280
rect 13354 11268 13360 11280
rect 12124 11240 13360 11268
rect 12124 11228 12130 11240
rect 13354 11228 13360 11240
rect 13412 11228 13418 11280
rect 14660 11268 14688 11299
rect 15746 11296 15752 11308
rect 15804 11296 15810 11348
rect 16758 11336 16764 11348
rect 16040 11308 16764 11336
rect 16040 11268 16068 11308
rect 16758 11296 16764 11308
rect 16816 11296 16822 11348
rect 16942 11336 16948 11348
rect 16903 11308 16948 11336
rect 16942 11296 16948 11308
rect 17000 11296 17006 11348
rect 14660 11240 16068 11268
rect 16117 11271 16175 11277
rect 16117 11237 16129 11271
rect 16163 11268 16175 11271
rect 17034 11268 17040 11280
rect 16163 11240 17040 11268
rect 16163 11237 16175 11240
rect 16117 11231 16175 11237
rect 17034 11228 17040 11240
rect 17092 11228 17098 11280
rect 6825 11203 6883 11209
rect 6825 11169 6837 11203
rect 6871 11200 6883 11203
rect 7190 11200 7196 11212
rect 6871 11172 7196 11200
rect 6871 11169 6883 11172
rect 6825 11163 6883 11169
rect 7190 11160 7196 11172
rect 7248 11160 7254 11212
rect 7565 11200 7571 11212
rect 7526 11172 7571 11200
rect 7565 11160 7571 11172
rect 7623 11160 7629 11212
rect 10020 11203 10078 11209
rect 10020 11169 10032 11203
rect 10066 11200 10078 11203
rect 10686 11200 10692 11212
rect 10066 11172 10692 11200
rect 10066 11169 10078 11172
rect 10020 11163 10078 11169
rect 10686 11160 10692 11172
rect 10744 11160 10750 11212
rect 10870 11209 10876 11212
rect 10864 11200 10876 11209
rect 10831 11172 10876 11200
rect 10864 11163 10876 11172
rect 10870 11160 10876 11163
rect 10928 11160 10934 11212
rect 12888 11203 12946 11209
rect 12888 11169 12900 11203
rect 12934 11200 12946 11203
rect 13630 11200 13636 11212
rect 12934 11172 13636 11200
rect 12934 11169 12946 11172
rect 12888 11163 12946 11169
rect 13630 11160 13636 11172
rect 13688 11160 13694 11212
rect 14461 11203 14519 11209
rect 14461 11169 14473 11203
rect 14507 11200 14519 11203
rect 14826 11200 14832 11212
rect 14507 11172 14832 11200
rect 14507 11169 14519 11172
rect 14461 11163 14519 11169
rect 14826 11160 14832 11172
rect 14884 11160 14890 11212
rect 16209 11203 16267 11209
rect 16209 11169 16221 11203
rect 16255 11200 16267 11203
rect 16390 11200 16396 11212
rect 16255 11172 16396 11200
rect 16255 11169 16267 11172
rect 16209 11163 16267 11169
rect 16390 11160 16396 11172
rect 16448 11160 16454 11212
rect 17310 11200 17316 11212
rect 17271 11172 17316 11200
rect 17310 11160 17316 11172
rect 17368 11160 17374 11212
rect 4985 11135 5043 11141
rect 4985 11101 4997 11135
rect 5031 11132 5043 11135
rect 6181 11135 6239 11141
rect 6181 11132 6193 11135
rect 5031 11104 6193 11132
rect 5031 11101 5043 11104
rect 4985 11095 5043 11101
rect 6181 11101 6193 11104
rect 6227 11101 6239 11135
rect 6181 11095 6239 11101
rect 10226 11092 10232 11144
rect 10284 11132 10290 11144
rect 10597 11135 10655 11141
rect 10597 11132 10609 11135
rect 10284 11104 10609 11132
rect 10284 11092 10290 11104
rect 10597 11101 10609 11104
rect 10643 11101 10655 11135
rect 10597 11095 10655 11101
rect 11698 11092 11704 11144
rect 11756 11132 11762 11144
rect 11882 11132 11888 11144
rect 11756 11104 11888 11132
rect 11756 11092 11762 11104
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 12621 11135 12679 11141
rect 12621 11101 12633 11135
rect 12667 11101 12679 11135
rect 12621 11095 12679 11101
rect 16301 11135 16359 11141
rect 16301 11101 16313 11135
rect 16347 11132 16359 11135
rect 16666 11132 16672 11144
rect 16347 11104 16672 11132
rect 16347 11101 16359 11104
rect 16301 11095 16359 11101
rect 4172 11036 4476 11064
rect 2314 10956 2320 11008
rect 2372 10996 2378 11008
rect 4172 10996 4200 11036
rect 4338 10996 4344 11008
rect 2372 10968 4200 10996
rect 4299 10968 4344 10996
rect 2372 10956 2378 10968
rect 4338 10956 4344 10968
rect 4396 10956 4402 11008
rect 4448 10996 4476 11036
rect 5368 11036 5672 11064
rect 5368 10996 5396 11036
rect 5534 10996 5540 11008
rect 4448 10968 5396 10996
rect 5495 10968 5540 10996
rect 5534 10956 5540 10968
rect 5592 10956 5598 11008
rect 5644 10996 5672 11036
rect 5994 11024 6000 11076
rect 6052 11064 6058 11076
rect 6362 11064 6368 11076
rect 6052 11036 6368 11064
rect 6052 11024 6058 11036
rect 6362 11024 6368 11036
rect 6420 11024 6426 11076
rect 6638 11024 6644 11076
rect 6696 11064 6702 11076
rect 7009 11067 7067 11073
rect 7009 11064 7021 11067
rect 6696 11036 7021 11064
rect 6696 11024 6702 11036
rect 7009 11033 7021 11036
rect 7055 11033 7067 11067
rect 10091 11067 10149 11073
rect 7009 11027 7067 11033
rect 8772 11036 9076 11064
rect 8772 10996 8800 11036
rect 8938 10996 8944 11008
rect 5644 10968 8800 10996
rect 8899 10968 8944 10996
rect 8938 10956 8944 10968
rect 8996 10956 9002 11008
rect 9048 10996 9076 11036
rect 10091 11033 10103 11067
rect 10137 11064 10149 11067
rect 10502 11064 10508 11076
rect 10137 11036 10508 11064
rect 10137 11033 10149 11036
rect 10091 11027 10149 11033
rect 10502 11024 10508 11036
rect 10560 11024 10566 11076
rect 12636 11064 12664 11095
rect 16666 11092 16672 11104
rect 16724 11092 16730 11144
rect 17402 11132 17408 11144
rect 17363 11104 17408 11132
rect 17402 11092 17408 11104
rect 17460 11092 17466 11144
rect 17497 11135 17555 11141
rect 17497 11101 17509 11135
rect 17543 11101 17555 11135
rect 17497 11095 17555 11101
rect 16684 11064 16712 11092
rect 17512 11064 17540 11095
rect 11532 11036 12664 11064
rect 13648 11036 14136 11064
rect 16684 11036 17540 11064
rect 10410 10996 10416 11008
rect 9048 10968 10416 10996
rect 10410 10956 10416 10968
rect 10468 10956 10474 11008
rect 10778 10956 10784 11008
rect 10836 10996 10842 11008
rect 11532 10996 11560 11036
rect 10836 10968 11560 10996
rect 10836 10956 10842 10968
rect 11606 10956 11612 11008
rect 11664 10996 11670 11008
rect 11977 10999 12035 11005
rect 11977 10996 11989 10999
rect 11664 10968 11989 10996
rect 11664 10956 11670 10968
rect 11977 10965 11989 10968
rect 12023 10965 12035 10999
rect 11977 10959 12035 10965
rect 12618 10956 12624 11008
rect 12676 10996 12682 11008
rect 13648 10996 13676 11036
rect 12676 10968 13676 10996
rect 12676 10956 12682 10968
rect 13814 10956 13820 11008
rect 13872 10996 13878 11008
rect 14001 10999 14059 11005
rect 14001 10996 14013 10999
rect 13872 10968 14013 10996
rect 13872 10956 13878 10968
rect 14001 10965 14013 10968
rect 14047 10965 14059 10999
rect 14108 10996 14136 11036
rect 16942 10996 16948 11008
rect 14108 10968 16948 10996
rect 14001 10959 14059 10965
rect 16942 10956 16948 10968
rect 17000 10996 17006 11008
rect 17862 10996 17868 11008
rect 17000 10968 17868 10996
rect 17000 10956 17006 10968
rect 17862 10956 17868 10968
rect 17920 10956 17926 11008
rect 1104 10906 18860 10928
rect 1104 10854 3947 10906
rect 3999 10854 4011 10906
rect 4063 10854 4075 10906
rect 4127 10854 4139 10906
rect 4191 10854 9878 10906
rect 9930 10854 9942 10906
rect 9994 10854 10006 10906
rect 10058 10854 10070 10906
rect 10122 10854 15808 10906
rect 15860 10854 15872 10906
rect 15924 10854 15936 10906
rect 15988 10854 16000 10906
rect 16052 10854 18860 10906
rect 1104 10832 18860 10854
rect 1688 10764 4292 10792
rect 1688 10597 1716 10764
rect 1673 10591 1731 10597
rect 1673 10557 1685 10591
rect 1719 10557 1731 10591
rect 2406 10588 2412 10600
rect 2367 10560 2412 10588
rect 1673 10551 1731 10557
rect 2406 10548 2412 10560
rect 2464 10548 2470 10600
rect 2516 10560 2820 10588
rect 2516 10520 2544 10560
rect 2792 10532 2820 10560
rect 3142 10548 3148 10600
rect 3200 10588 3206 10600
rect 3878 10588 3884 10600
rect 3200 10560 3884 10588
rect 3200 10548 3206 10560
rect 3878 10548 3884 10560
rect 3936 10548 3942 10600
rect 4264 10588 4292 10764
rect 4430 10752 4436 10804
rect 4488 10792 4494 10804
rect 5442 10792 5448 10804
rect 4488 10764 5448 10792
rect 4488 10752 4494 10764
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 5902 10752 5908 10804
rect 5960 10792 5966 10804
rect 6825 10795 6883 10801
rect 6825 10792 6837 10795
rect 5960 10764 6837 10792
rect 5960 10752 5966 10764
rect 6825 10761 6837 10764
rect 6871 10761 6883 10795
rect 6825 10755 6883 10761
rect 7098 10752 7104 10804
rect 7156 10792 7162 10804
rect 7742 10792 7748 10804
rect 7156 10764 7748 10792
rect 7156 10752 7162 10764
rect 7742 10752 7748 10764
rect 7800 10752 7806 10804
rect 10226 10792 10232 10804
rect 8956 10764 10232 10792
rect 8386 10724 8392 10736
rect 5276 10696 8392 10724
rect 4338 10616 4344 10668
rect 4396 10656 4402 10668
rect 5276 10665 5304 10696
rect 8386 10684 8392 10696
rect 8444 10684 8450 10736
rect 5077 10659 5135 10665
rect 5077 10656 5089 10659
rect 4396 10628 5089 10656
rect 4396 10616 4402 10628
rect 5077 10625 5089 10628
rect 5123 10625 5135 10659
rect 5077 10619 5135 10625
rect 5261 10659 5319 10665
rect 5261 10625 5273 10659
rect 5307 10625 5319 10659
rect 5261 10619 5319 10625
rect 5994 10616 6000 10668
rect 6052 10656 6058 10668
rect 6730 10656 6736 10668
rect 6052 10628 6736 10656
rect 6052 10616 6058 10628
rect 6730 10616 6736 10628
rect 6788 10656 6794 10668
rect 8956 10665 8984 10764
rect 10226 10752 10232 10764
rect 10284 10792 10290 10804
rect 10778 10792 10784 10804
rect 10284 10764 10784 10792
rect 10284 10752 10290 10764
rect 10778 10752 10784 10764
rect 10836 10792 10842 10804
rect 14182 10792 14188 10804
rect 10836 10764 14188 10792
rect 10836 10752 10842 10764
rect 10870 10684 10876 10736
rect 10928 10724 10934 10736
rect 10928 10696 11468 10724
rect 10928 10684 10934 10696
rect 7377 10659 7435 10665
rect 7377 10656 7389 10659
rect 6788 10628 7389 10656
rect 6788 10616 6794 10628
rect 7377 10625 7389 10628
rect 7423 10625 7435 10659
rect 8941 10659 8999 10665
rect 7377 10619 7435 10625
rect 7484 10628 8892 10656
rect 4985 10591 5043 10597
rect 4264 10560 4936 10588
rect 1872 10492 2544 10520
rect 2676 10523 2734 10529
rect 1872 10461 1900 10492
rect 2676 10489 2688 10523
rect 2722 10489 2734 10523
rect 2676 10483 2734 10489
rect 1857 10455 1915 10461
rect 1857 10421 1869 10455
rect 1903 10421 1915 10455
rect 2700 10452 2728 10483
rect 2774 10480 2780 10532
rect 2832 10480 2838 10532
rect 2866 10480 2872 10532
rect 2924 10520 2930 10532
rect 4908 10520 4936 10560
rect 4985 10557 4997 10591
rect 5031 10588 5043 10591
rect 5534 10588 5540 10600
rect 5031 10560 5540 10588
rect 5031 10557 5043 10560
rect 4985 10551 5043 10557
rect 5534 10548 5540 10560
rect 5592 10548 5598 10600
rect 5810 10588 5816 10600
rect 5771 10560 5816 10588
rect 5810 10548 5816 10560
rect 5868 10548 5874 10600
rect 7098 10588 7104 10600
rect 5920 10560 7104 10588
rect 5920 10520 5948 10560
rect 7098 10548 7104 10560
rect 7156 10548 7162 10600
rect 7193 10591 7251 10597
rect 7193 10557 7205 10591
rect 7239 10588 7251 10591
rect 7282 10588 7288 10600
rect 7239 10560 7288 10588
rect 7239 10557 7251 10560
rect 7193 10551 7251 10557
rect 7282 10548 7288 10560
rect 7340 10548 7346 10600
rect 6086 10520 6092 10532
rect 2924 10492 4752 10520
rect 4908 10492 5948 10520
rect 6047 10492 6092 10520
rect 2924 10480 2930 10492
rect 3326 10452 3332 10464
rect 2700 10424 3332 10452
rect 1857 10415 1915 10421
rect 3326 10412 3332 10424
rect 3384 10412 3390 10464
rect 3510 10412 3516 10464
rect 3568 10452 3574 10464
rect 3789 10455 3847 10461
rect 3789 10452 3801 10455
rect 3568 10424 3801 10452
rect 3568 10412 3574 10424
rect 3789 10421 3801 10424
rect 3835 10421 3847 10455
rect 3789 10415 3847 10421
rect 4246 10412 4252 10464
rect 4304 10452 4310 10464
rect 4617 10455 4675 10461
rect 4617 10452 4629 10455
rect 4304 10424 4629 10452
rect 4304 10412 4310 10424
rect 4617 10421 4629 10424
rect 4663 10421 4675 10455
rect 4724 10452 4752 10492
rect 6086 10480 6092 10492
rect 6144 10480 6150 10532
rect 7484 10520 7512 10628
rect 8021 10591 8079 10597
rect 8021 10557 8033 10591
rect 8067 10588 8079 10591
rect 8662 10588 8668 10600
rect 8067 10560 8668 10588
rect 8067 10557 8079 10560
rect 8021 10551 8079 10557
rect 8662 10548 8668 10560
rect 8720 10548 8726 10600
rect 8864 10588 8892 10628
rect 8941 10625 8953 10659
rect 8987 10625 8999 10659
rect 8941 10619 8999 10625
rect 10410 10616 10416 10668
rect 10468 10656 10474 10668
rect 11238 10656 11244 10668
rect 10468 10628 11244 10656
rect 10468 10616 10474 10628
rect 11238 10616 11244 10628
rect 11296 10616 11302 10668
rect 11440 10665 11468 10696
rect 12066 10684 12072 10736
rect 12124 10724 12130 10736
rect 12342 10724 12348 10736
rect 12124 10696 12348 10724
rect 12124 10684 12130 10696
rect 12342 10684 12348 10696
rect 12400 10684 12406 10736
rect 12636 10696 12848 10724
rect 11425 10659 11483 10665
rect 11425 10625 11437 10659
rect 11471 10656 11483 10659
rect 12636 10656 12664 10696
rect 11471 10628 12664 10656
rect 12820 10656 12848 10696
rect 13081 10659 13139 10665
rect 13081 10656 13093 10659
rect 12820 10628 13093 10656
rect 11471 10625 11483 10628
rect 11425 10619 11483 10625
rect 13081 10625 13093 10628
rect 13127 10656 13139 10659
rect 13446 10656 13452 10668
rect 13127 10628 13452 10656
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 13446 10616 13452 10628
rect 13504 10616 13510 10668
rect 13556 10656 13584 10764
rect 14182 10752 14188 10764
rect 14240 10752 14246 10804
rect 16761 10795 16819 10801
rect 16761 10761 16773 10795
rect 16807 10792 16819 10795
rect 17402 10792 17408 10804
rect 16807 10764 17408 10792
rect 16807 10761 16819 10764
rect 16761 10755 16819 10761
rect 17402 10752 17408 10764
rect 17460 10752 17466 10804
rect 13817 10659 13875 10665
rect 13817 10656 13829 10659
rect 13556 10628 13829 10656
rect 13817 10625 13829 10628
rect 13863 10625 13875 10659
rect 17402 10656 17408 10668
rect 17363 10628 17408 10656
rect 13817 10619 13875 10625
rect 17402 10616 17408 10628
rect 17460 10616 17466 10668
rect 12618 10588 12624 10600
rect 8864 10560 12624 10588
rect 12618 10548 12624 10560
rect 12676 10548 12682 10600
rect 16025 10591 16083 10597
rect 16025 10588 16037 10591
rect 13924 10560 16037 10588
rect 6196 10492 7512 10520
rect 9208 10523 9266 10529
rect 6196 10452 6224 10492
rect 9208 10489 9220 10523
rect 9254 10520 9266 10523
rect 11606 10520 11612 10532
rect 9254 10492 11612 10520
rect 9254 10489 9266 10492
rect 9208 10483 9266 10489
rect 11606 10480 11612 10492
rect 11664 10480 11670 10532
rect 11698 10480 11704 10532
rect 11756 10520 11762 10532
rect 12805 10523 12863 10529
rect 12805 10520 12817 10523
rect 11756 10492 12817 10520
rect 11756 10480 11762 10492
rect 12805 10489 12817 10492
rect 12851 10520 12863 10523
rect 13924 10520 13952 10560
rect 16025 10557 16037 10560
rect 16071 10557 16083 10591
rect 16025 10551 16083 10557
rect 16942 10548 16948 10600
rect 17000 10588 17006 10600
rect 17129 10591 17187 10597
rect 17129 10588 17141 10591
rect 17000 10560 17141 10588
rect 17000 10548 17006 10560
rect 17129 10557 17141 10560
rect 17175 10557 17187 10591
rect 17129 10551 17187 10557
rect 17221 10591 17279 10597
rect 17221 10557 17233 10591
rect 17267 10588 17279 10591
rect 18322 10588 18328 10600
rect 17267 10560 18328 10588
rect 17267 10557 17279 10560
rect 17221 10551 17279 10557
rect 12851 10492 13952 10520
rect 14084 10523 14142 10529
rect 12851 10489 12863 10492
rect 12805 10483 12863 10489
rect 14084 10489 14096 10523
rect 14130 10520 14142 10523
rect 15654 10520 15660 10532
rect 14130 10492 15660 10520
rect 14130 10489 14142 10492
rect 14084 10483 14142 10489
rect 15654 10480 15660 10492
rect 15712 10480 15718 10532
rect 15838 10480 15844 10532
rect 15896 10520 15902 10532
rect 17236 10520 17264 10551
rect 18322 10548 18328 10560
rect 18380 10548 18386 10600
rect 15896 10492 17264 10520
rect 15896 10480 15902 10492
rect 4724 10424 6224 10452
rect 4617 10415 4675 10421
rect 6270 10412 6276 10464
rect 6328 10452 6334 10464
rect 7285 10455 7343 10461
rect 7285 10452 7297 10455
rect 6328 10424 7297 10452
rect 6328 10412 6334 10424
rect 7285 10421 7297 10424
rect 7331 10421 7343 10455
rect 7285 10415 7343 10421
rect 7834 10412 7840 10464
rect 7892 10452 7898 10464
rect 8205 10455 8263 10461
rect 8205 10452 8217 10455
rect 7892 10424 8217 10452
rect 7892 10412 7898 10424
rect 8205 10421 8217 10424
rect 8251 10421 8263 10455
rect 8205 10415 8263 10421
rect 10321 10455 10379 10461
rect 10321 10421 10333 10455
rect 10367 10452 10379 10455
rect 10410 10452 10416 10464
rect 10367 10424 10416 10452
rect 10367 10421 10379 10424
rect 10321 10415 10379 10421
rect 10410 10412 10416 10424
rect 10468 10412 10474 10464
rect 10778 10452 10784 10464
rect 10739 10424 10784 10452
rect 10778 10412 10784 10424
rect 10836 10412 10842 10464
rect 11054 10412 11060 10464
rect 11112 10452 11118 10464
rect 11149 10455 11207 10461
rect 11149 10452 11161 10455
rect 11112 10424 11161 10452
rect 11112 10412 11118 10424
rect 11149 10421 11161 10424
rect 11195 10452 11207 10455
rect 12066 10452 12072 10464
rect 11195 10424 12072 10452
rect 11195 10421 11207 10424
rect 11149 10415 11207 10421
rect 12066 10412 12072 10424
rect 12124 10412 12130 10464
rect 12437 10455 12495 10461
rect 12437 10421 12449 10455
rect 12483 10452 12495 10455
rect 12618 10452 12624 10464
rect 12483 10424 12624 10452
rect 12483 10421 12495 10424
rect 12437 10415 12495 10421
rect 12618 10412 12624 10424
rect 12676 10412 12682 10464
rect 12897 10455 12955 10461
rect 12897 10421 12909 10455
rect 12943 10452 12955 10455
rect 13446 10452 13452 10464
rect 12943 10424 13452 10452
rect 12943 10421 12955 10424
rect 12897 10415 12955 10421
rect 13446 10412 13452 10424
rect 13504 10412 13510 10464
rect 13630 10412 13636 10464
rect 13688 10452 13694 10464
rect 15197 10455 15255 10461
rect 15197 10452 15209 10455
rect 13688 10424 15209 10452
rect 13688 10412 13694 10424
rect 15197 10421 15209 10424
rect 15243 10421 15255 10455
rect 15197 10415 15255 10421
rect 15470 10412 15476 10464
rect 15528 10452 15534 10464
rect 16209 10455 16267 10461
rect 16209 10452 16221 10455
rect 15528 10424 16221 10452
rect 15528 10412 15534 10424
rect 16209 10421 16221 10424
rect 16255 10421 16267 10455
rect 16209 10415 16267 10421
rect 1104 10362 18860 10384
rect 1104 10310 6912 10362
rect 6964 10310 6976 10362
rect 7028 10310 7040 10362
rect 7092 10310 7104 10362
rect 7156 10310 12843 10362
rect 12895 10310 12907 10362
rect 12959 10310 12971 10362
rect 13023 10310 13035 10362
rect 13087 10310 18860 10362
rect 1104 10288 18860 10310
rect 1578 10248 1584 10260
rect 1539 10220 1584 10248
rect 1578 10208 1584 10220
rect 1636 10208 1642 10260
rect 1949 10251 2007 10257
rect 1949 10217 1961 10251
rect 1995 10248 2007 10251
rect 2777 10251 2835 10257
rect 2777 10248 2789 10251
rect 1995 10220 2789 10248
rect 1995 10217 2007 10220
rect 1949 10211 2007 10217
rect 2777 10217 2789 10220
rect 2823 10217 2835 10251
rect 2777 10211 2835 10217
rect 4798 10208 4804 10260
rect 4856 10248 4862 10260
rect 5353 10251 5411 10257
rect 5353 10248 5365 10251
rect 4856 10220 5365 10248
rect 4856 10208 4862 10220
rect 5353 10217 5365 10220
rect 5399 10217 5411 10251
rect 5353 10211 5411 10217
rect 5810 10208 5816 10260
rect 5868 10248 5874 10260
rect 9861 10251 9919 10257
rect 9861 10248 9873 10251
rect 5868 10220 9873 10248
rect 5868 10208 5874 10220
rect 9861 10217 9873 10220
rect 9907 10217 9919 10251
rect 9861 10211 9919 10217
rect 10229 10251 10287 10257
rect 10229 10217 10241 10251
rect 10275 10248 10287 10251
rect 11057 10251 11115 10257
rect 11057 10248 11069 10251
rect 10275 10220 11069 10248
rect 10275 10217 10287 10220
rect 10229 10211 10287 10217
rect 11057 10217 11069 10220
rect 11103 10217 11115 10251
rect 12618 10248 12624 10260
rect 12579 10220 12624 10248
rect 11057 10211 11115 10217
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 13446 10248 13452 10260
rect 13407 10220 13452 10248
rect 13446 10208 13452 10220
rect 13504 10208 13510 10260
rect 14182 10208 14188 10260
rect 14240 10248 14246 10260
rect 17221 10251 17279 10257
rect 14240 10220 15424 10248
rect 14240 10208 14246 10220
rect 2406 10140 2412 10192
rect 2464 10180 2470 10192
rect 2958 10180 2964 10192
rect 2464 10152 2964 10180
rect 2464 10140 2470 10152
rect 2958 10140 2964 10152
rect 3016 10140 3022 10192
rect 5721 10183 5779 10189
rect 5721 10149 5733 10183
rect 5767 10180 5779 10183
rect 7282 10180 7288 10192
rect 5767 10152 7288 10180
rect 5767 10149 5779 10152
rect 5721 10143 5779 10149
rect 7282 10140 7288 10152
rect 7340 10140 7346 10192
rect 7828 10183 7886 10189
rect 7828 10149 7840 10183
rect 7874 10180 7886 10183
rect 8386 10180 8392 10192
rect 7874 10152 8392 10180
rect 7874 10149 7886 10152
rect 7828 10143 7886 10149
rect 8386 10140 8392 10152
rect 8444 10180 8450 10192
rect 8938 10180 8944 10192
rect 8444 10152 8944 10180
rect 8444 10140 8450 10152
rect 8938 10140 8944 10152
rect 8996 10140 9002 10192
rect 10778 10140 10784 10192
rect 10836 10180 10842 10192
rect 11517 10183 11575 10189
rect 11517 10180 11529 10183
rect 10836 10152 11529 10180
rect 10836 10140 10842 10152
rect 11517 10149 11529 10152
rect 11563 10149 11575 10183
rect 11517 10143 11575 10149
rect 12802 10140 12808 10192
rect 12860 10180 12866 10192
rect 13909 10183 13967 10189
rect 13909 10180 13921 10183
rect 12860 10152 13921 10180
rect 12860 10140 12866 10152
rect 13909 10149 13921 10152
rect 13955 10180 13967 10183
rect 15286 10180 15292 10192
rect 13955 10152 15292 10180
rect 13955 10149 13967 10152
rect 13909 10143 13967 10149
rect 15286 10140 15292 10152
rect 15344 10140 15350 10192
rect 2041 10115 2099 10121
rect 2041 10081 2053 10115
rect 2087 10112 2099 10115
rect 3050 10112 3056 10124
rect 2087 10084 3056 10112
rect 2087 10081 2099 10084
rect 2041 10075 2099 10081
rect 3050 10072 3056 10084
rect 3108 10072 3114 10124
rect 3145 10115 3203 10121
rect 3145 10081 3157 10115
rect 3191 10112 3203 10115
rect 4430 10112 4436 10124
rect 3191 10084 4200 10112
rect 4391 10084 4436 10112
rect 3191 10081 3203 10084
rect 3145 10075 3203 10081
rect 2225 10047 2283 10053
rect 2225 10013 2237 10047
rect 2271 10013 2283 10047
rect 2225 10007 2283 10013
rect 2240 9976 2268 10007
rect 2590 10004 2596 10056
rect 2648 10044 2654 10056
rect 3237 10047 3295 10053
rect 3237 10044 3249 10047
rect 2648 10016 3249 10044
rect 2648 10004 2654 10016
rect 3237 10013 3249 10016
rect 3283 10013 3295 10047
rect 3237 10007 3295 10013
rect 3326 10004 3332 10056
rect 3384 10044 3390 10056
rect 3384 10016 3429 10044
rect 3384 10004 3390 10016
rect 3510 9976 3516 9988
rect 2240 9948 3516 9976
rect 3510 9936 3516 9948
rect 3568 9936 3574 9988
rect 2866 9868 2872 9920
rect 2924 9908 2930 9920
rect 4065 9911 4123 9917
rect 4065 9908 4077 9911
rect 2924 9880 4077 9908
rect 2924 9868 2930 9880
rect 4065 9877 4077 9880
rect 4111 9877 4123 9911
rect 4172 9908 4200 10084
rect 4430 10072 4436 10084
rect 4488 10072 4494 10124
rect 6270 10072 6276 10124
rect 6328 10112 6334 10124
rect 6549 10115 6607 10121
rect 6549 10112 6561 10115
rect 6328 10084 6561 10112
rect 6328 10072 6334 10084
rect 6549 10081 6561 10084
rect 6595 10081 6607 10115
rect 6549 10075 6607 10081
rect 7466 10072 7472 10124
rect 7524 10112 7530 10124
rect 10134 10112 10140 10124
rect 7524 10084 10140 10112
rect 7524 10072 7530 10084
rect 10134 10072 10140 10084
rect 10192 10072 10198 10124
rect 10226 10072 10232 10124
rect 10284 10112 10290 10124
rect 10594 10112 10600 10124
rect 10284 10084 10600 10112
rect 10284 10072 10290 10084
rect 10594 10072 10600 10084
rect 10652 10072 10658 10124
rect 11054 10072 11060 10124
rect 11112 10112 11118 10124
rect 11425 10115 11483 10121
rect 11425 10112 11437 10115
rect 11112 10084 11437 10112
rect 11112 10072 11118 10084
rect 11425 10081 11437 10084
rect 11471 10081 11483 10115
rect 11425 10075 11483 10081
rect 13817 10115 13875 10121
rect 13817 10081 13829 10115
rect 13863 10112 13875 10115
rect 15010 10112 15016 10124
rect 13863 10084 15016 10112
rect 13863 10081 13875 10084
rect 13817 10075 13875 10081
rect 15010 10072 15016 10084
rect 15068 10072 15074 10124
rect 15396 10121 15424 10220
rect 17221 10217 17233 10251
rect 17267 10248 17279 10251
rect 17310 10248 17316 10260
rect 17267 10220 17316 10248
rect 17267 10217 17279 10220
rect 17221 10211 17279 10217
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 17586 10248 17592 10260
rect 17547 10220 17592 10248
rect 17586 10208 17592 10220
rect 17644 10208 17650 10260
rect 18414 10248 18420 10260
rect 17696 10220 18420 10248
rect 15838 10180 15844 10192
rect 15488 10152 15844 10180
rect 15381 10115 15439 10121
rect 15381 10081 15393 10115
rect 15427 10081 15439 10115
rect 15381 10075 15439 10081
rect 4522 10044 4528 10056
rect 4483 10016 4528 10044
rect 4522 10004 4528 10016
rect 4580 10004 4586 10056
rect 4706 10044 4712 10056
rect 4667 10016 4712 10044
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 5810 10044 5816 10056
rect 5771 10016 5816 10044
rect 5810 10004 5816 10016
rect 5868 10004 5874 10056
rect 5994 10044 6000 10056
rect 5955 10016 6000 10044
rect 5994 10004 6000 10016
rect 6052 10004 6058 10056
rect 6730 10044 6736 10056
rect 6691 10016 6736 10044
rect 6730 10004 6736 10016
rect 6788 10004 6794 10056
rect 7558 10044 7564 10056
rect 7471 10016 7564 10044
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 10321 10047 10379 10053
rect 10321 10013 10333 10047
rect 10367 10013 10379 10047
rect 10321 10007 10379 10013
rect 6914 9936 6920 9988
rect 6972 9976 6978 9988
rect 7576 9976 7604 10004
rect 6972 9948 7604 9976
rect 8941 9979 8999 9985
rect 6972 9936 6978 9948
rect 8941 9945 8953 9979
rect 8987 9976 8999 9979
rect 9306 9976 9312 9988
rect 8987 9948 9312 9976
rect 8987 9945 8999 9948
rect 8941 9939 8999 9945
rect 9306 9936 9312 9948
rect 9364 9936 9370 9988
rect 9398 9936 9404 9988
rect 9456 9976 9462 9988
rect 9766 9976 9772 9988
rect 9456 9948 9772 9976
rect 9456 9936 9462 9948
rect 9766 9936 9772 9948
rect 9824 9936 9830 9988
rect 10336 9976 10364 10007
rect 10410 10004 10416 10056
rect 10468 10044 10474 10056
rect 11606 10044 11612 10056
rect 10468 10016 10513 10044
rect 11567 10016 11612 10044
rect 10468 10004 10474 10016
rect 11606 10004 11612 10016
rect 11664 10004 11670 10056
rect 12710 10044 12716 10056
rect 12671 10016 12716 10044
rect 12710 10004 12716 10016
rect 12768 10004 12774 10056
rect 12802 10004 12808 10056
rect 12860 10044 12866 10056
rect 14001 10047 14059 10053
rect 12860 10016 12905 10044
rect 12860 10004 12866 10016
rect 14001 10013 14013 10047
rect 14047 10013 14059 10047
rect 15488 10044 15516 10152
rect 15838 10140 15844 10152
rect 15896 10140 15902 10192
rect 15648 10115 15706 10121
rect 15648 10081 15660 10115
rect 15694 10112 15706 10115
rect 16574 10112 16580 10124
rect 15694 10084 16580 10112
rect 15694 10081 15706 10084
rect 15648 10075 15706 10081
rect 16574 10072 16580 10084
rect 16632 10112 16638 10124
rect 17402 10112 17408 10124
rect 16632 10084 17408 10112
rect 16632 10072 16638 10084
rect 14001 10007 14059 10013
rect 15304 10016 15516 10044
rect 12253 9979 12311 9985
rect 12253 9976 12265 9979
rect 10336 9948 12265 9976
rect 12253 9945 12265 9948
rect 12299 9945 12311 9979
rect 12253 9939 12311 9945
rect 13630 9936 13636 9988
rect 13688 9976 13694 9988
rect 14016 9976 14044 10007
rect 15304 9988 15332 10016
rect 13688 9948 14044 9976
rect 13688 9936 13694 9948
rect 15286 9936 15292 9988
rect 15344 9936 15350 9988
rect 6730 9908 6736 9920
rect 4172 9880 6736 9908
rect 4065 9871 4123 9877
rect 6730 9868 6736 9880
rect 6788 9868 6794 9920
rect 9490 9868 9496 9920
rect 9548 9908 9554 9920
rect 15102 9908 15108 9920
rect 9548 9880 15108 9908
rect 9548 9868 9554 9880
rect 15102 9868 15108 9880
rect 15160 9868 15166 9920
rect 16666 9868 16672 9920
rect 16724 9908 16730 9920
rect 16761 9911 16819 9917
rect 16761 9908 16773 9911
rect 16724 9880 16773 9908
rect 16724 9868 16730 9880
rect 16761 9877 16773 9880
rect 16807 9877 16819 9911
rect 16868 9908 16896 10084
rect 17402 10072 17408 10084
rect 17460 10072 17466 10124
rect 17586 10004 17592 10056
rect 17644 10044 17650 10056
rect 17696 10053 17724 10220
rect 18414 10208 18420 10220
rect 18472 10208 18478 10260
rect 17681 10047 17739 10053
rect 17681 10044 17693 10047
rect 17644 10016 17693 10044
rect 17644 10004 17650 10016
rect 17681 10013 17693 10016
rect 17727 10013 17739 10047
rect 17681 10007 17739 10013
rect 17773 10047 17831 10053
rect 17773 10013 17785 10047
rect 17819 10013 17831 10047
rect 17773 10007 17831 10013
rect 17788 9908 17816 10007
rect 16868 9880 17816 9908
rect 16761 9871 16819 9877
rect 1104 9818 18860 9840
rect 1104 9766 3947 9818
rect 3999 9766 4011 9818
rect 4063 9766 4075 9818
rect 4127 9766 4139 9818
rect 4191 9766 9878 9818
rect 9930 9766 9942 9818
rect 9994 9766 10006 9818
rect 10058 9766 10070 9818
rect 10122 9766 15808 9818
rect 15860 9766 15872 9818
rect 15924 9766 15936 9818
rect 15988 9766 16000 9818
rect 16052 9766 18860 9818
rect 1104 9744 18860 9766
rect 3050 9664 3056 9716
rect 3108 9704 3114 9716
rect 3697 9707 3755 9713
rect 3697 9704 3709 9707
rect 3108 9676 3709 9704
rect 3108 9664 3114 9676
rect 3697 9673 3709 9676
rect 3743 9673 3755 9707
rect 3697 9667 3755 9673
rect 3804 9676 4292 9704
rect 3237 9639 3295 9645
rect 3237 9605 3249 9639
rect 3283 9636 3295 9639
rect 3326 9636 3332 9648
rect 3283 9608 3332 9636
rect 3283 9605 3295 9608
rect 3237 9599 3295 9605
rect 3326 9596 3332 9608
rect 3384 9636 3390 9648
rect 3804 9636 3832 9676
rect 3384 9608 3832 9636
rect 3384 9596 3390 9608
rect 2958 9528 2964 9580
rect 3016 9528 3022 9580
rect 4264 9577 4292 9676
rect 5442 9664 5448 9716
rect 5500 9704 5506 9716
rect 11698 9704 11704 9716
rect 5500 9676 11704 9704
rect 5500 9664 5506 9676
rect 11698 9664 11704 9676
rect 11756 9664 11762 9716
rect 12437 9707 12495 9713
rect 12437 9673 12449 9707
rect 12483 9704 12495 9707
rect 12710 9704 12716 9716
rect 12483 9676 12716 9704
rect 12483 9673 12495 9676
rect 12437 9667 12495 9673
rect 12710 9664 12716 9676
rect 12768 9664 12774 9716
rect 15286 9704 15292 9716
rect 14200 9676 15292 9704
rect 4985 9639 5043 9645
rect 4985 9605 4997 9639
rect 5031 9605 5043 9639
rect 5258 9636 5264 9648
rect 5219 9608 5264 9636
rect 4985 9599 5043 9605
rect 4249 9571 4307 9577
rect 4249 9537 4261 9571
rect 4295 9537 4307 9571
rect 4249 9531 4307 9537
rect 5000 9568 5028 9599
rect 5258 9596 5264 9608
rect 5316 9596 5322 9648
rect 8297 9639 8355 9645
rect 5368 9608 6960 9636
rect 5368 9568 5396 9608
rect 6932 9580 6960 9608
rect 8297 9605 8309 9639
rect 8343 9636 8355 9639
rect 8754 9636 8760 9648
rect 8343 9608 8760 9636
rect 8343 9605 8355 9608
rect 8297 9599 8355 9605
rect 8754 9596 8760 9608
rect 8812 9596 8818 9648
rect 9122 9596 9128 9648
rect 9180 9636 9186 9648
rect 10781 9639 10839 9645
rect 9180 9608 10732 9636
rect 9180 9596 9186 9608
rect 5718 9568 5724 9580
rect 5000 9540 5396 9568
rect 5679 9540 5724 9568
rect 1578 9460 1584 9512
rect 1636 9500 1642 9512
rect 1857 9503 1915 9509
rect 1857 9500 1869 9503
rect 1636 9472 1869 9500
rect 1636 9460 1642 9472
rect 1857 9469 1869 9472
rect 1903 9500 1915 9503
rect 2976 9500 3004 9528
rect 4062 9500 4068 9512
rect 1903 9472 4068 9500
rect 1903 9469 1915 9472
rect 1857 9463 1915 9469
rect 4062 9460 4068 9472
rect 4120 9500 4126 9512
rect 5000 9500 5028 9540
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 5905 9571 5963 9577
rect 5905 9537 5917 9571
rect 5951 9568 5963 9571
rect 5994 9568 6000 9580
rect 5951 9540 6000 9568
rect 5951 9537 5963 9540
rect 5905 9531 5963 9537
rect 5994 9528 6000 9540
rect 6052 9528 6058 9580
rect 6914 9568 6920 9580
rect 6875 9540 6920 9568
rect 6914 9528 6920 9540
rect 6972 9528 6978 9580
rect 9306 9568 9312 9580
rect 9267 9540 9312 9568
rect 9306 9528 9312 9540
rect 9364 9528 9370 9580
rect 9490 9528 9496 9580
rect 9548 9568 9554 9580
rect 10229 9571 10287 9577
rect 10229 9568 10241 9571
rect 9548 9540 10241 9568
rect 9548 9528 9554 9540
rect 10229 9537 10241 9540
rect 10275 9537 10287 9571
rect 10229 9531 10287 9537
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9568 10471 9571
rect 10594 9568 10600 9580
rect 10459 9540 10600 9568
rect 10459 9537 10471 9540
rect 10413 9531 10471 9537
rect 10594 9528 10600 9540
rect 10652 9528 10658 9580
rect 10704 9568 10732 9608
rect 10781 9605 10793 9639
rect 10827 9636 10839 9639
rect 11054 9636 11060 9648
rect 10827 9608 11060 9636
rect 10827 9605 10839 9608
rect 10781 9599 10839 9605
rect 11054 9596 11060 9608
rect 11112 9596 11118 9648
rect 14200 9636 14228 9676
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 11225 9608 14228 9636
rect 15565 9639 15623 9645
rect 11225 9568 11253 9608
rect 15565 9605 15577 9639
rect 15611 9636 15623 9639
rect 15654 9636 15660 9648
rect 15611 9608 15660 9636
rect 15611 9605 15623 9608
rect 15565 9599 15623 9605
rect 15654 9596 15660 9608
rect 15712 9596 15718 9648
rect 10704 9540 11253 9568
rect 11425 9571 11483 9577
rect 11425 9537 11437 9571
rect 11471 9568 11483 9571
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 11471 9540 13001 9568
rect 11471 9537 11483 9540
rect 11425 9531 11483 9537
rect 12989 9537 13001 9540
rect 13035 9568 13047 9571
rect 13814 9568 13820 9580
rect 13035 9540 13820 9568
rect 13035 9537 13047 9540
rect 12989 9531 13047 9537
rect 13814 9528 13820 9540
rect 13872 9528 13878 9580
rect 14182 9568 14188 9580
rect 14143 9540 14188 9568
rect 14182 9528 14188 9540
rect 14240 9528 14246 9580
rect 16850 9528 16856 9580
rect 16908 9568 16914 9580
rect 16908 9540 17172 9568
rect 16908 9528 16914 9540
rect 4120 9472 5028 9500
rect 5169 9503 5227 9509
rect 4120 9460 4126 9472
rect 5169 9469 5181 9503
rect 5215 9500 5227 9503
rect 6270 9500 6276 9512
rect 5215 9472 6276 9500
rect 5215 9469 5227 9472
rect 5169 9463 5227 9469
rect 6270 9460 6276 9472
rect 6328 9460 6334 9512
rect 6641 9503 6699 9509
rect 6641 9469 6653 9503
rect 6687 9469 6699 9503
rect 6641 9463 6699 9469
rect 7184 9503 7242 9509
rect 7184 9469 7196 9503
rect 7230 9500 7242 9503
rect 8202 9500 8208 9512
rect 7230 9472 8208 9500
rect 7230 9469 7242 9472
rect 7184 9463 7242 9469
rect 2124 9435 2182 9441
rect 2124 9401 2136 9435
rect 2170 9432 2182 9435
rect 2958 9432 2964 9444
rect 2170 9404 2964 9432
rect 2170 9401 2182 9404
rect 2124 9395 2182 9401
rect 2958 9392 2964 9404
rect 3016 9392 3022 9444
rect 4154 9432 4160 9444
rect 4115 9404 4160 9432
rect 4154 9392 4160 9404
rect 4212 9392 4218 9444
rect 5626 9432 5632 9444
rect 5539 9404 5632 9432
rect 5626 9392 5632 9404
rect 5684 9432 5690 9444
rect 6656 9432 6684 9463
rect 8202 9460 8208 9472
rect 8260 9500 8266 9512
rect 9324 9500 9352 9528
rect 8260 9472 9352 9500
rect 9508 9472 9812 9500
rect 8260 9460 8266 9472
rect 9508 9432 9536 9472
rect 9784 9432 9812 9472
rect 10042 9460 10048 9512
rect 10100 9500 10106 9512
rect 11146 9500 11152 9512
rect 10100 9472 11015 9500
rect 11107 9472 11152 9500
rect 10100 9460 10106 9472
rect 10987 9432 11015 9472
rect 11146 9460 11152 9472
rect 11204 9460 11210 9512
rect 11241 9503 11299 9509
rect 11241 9469 11253 9503
rect 11287 9500 11299 9503
rect 11974 9500 11980 9512
rect 11287 9472 11980 9500
rect 11287 9469 11299 9472
rect 11241 9463 11299 9469
rect 11974 9460 11980 9472
rect 12032 9460 12038 9512
rect 12897 9503 12955 9509
rect 12897 9469 12909 9503
rect 12943 9500 12955 9503
rect 13170 9500 13176 9512
rect 12943 9472 13176 9500
rect 12943 9469 12955 9472
rect 12897 9463 12955 9469
rect 13170 9460 13176 9472
rect 13228 9460 13234 9512
rect 13354 9460 13360 9512
rect 13412 9500 13418 9512
rect 17144 9509 17172 9540
rect 17218 9528 17224 9580
rect 17276 9568 17282 9580
rect 17313 9571 17371 9577
rect 17313 9568 17325 9571
rect 17276 9540 17325 9568
rect 17276 9528 17282 9540
rect 17313 9537 17325 9540
rect 17359 9537 17371 9571
rect 17313 9531 17371 9537
rect 16025 9503 16083 9509
rect 16025 9500 16037 9503
rect 13412 9472 16037 9500
rect 13412 9460 13418 9472
rect 16025 9469 16037 9472
rect 16071 9469 16083 9503
rect 16025 9463 16083 9469
rect 17129 9503 17187 9509
rect 17129 9469 17141 9503
rect 17175 9469 17187 9503
rect 17129 9463 17187 9469
rect 12158 9432 12164 9444
rect 5684 9404 6592 9432
rect 6656 9404 9536 9432
rect 9591 9404 9720 9432
rect 9784 9404 10907 9432
rect 10987 9404 12164 9432
rect 5684 9392 5690 9404
rect 2682 9324 2688 9376
rect 2740 9364 2746 9376
rect 3050 9364 3056 9376
rect 2740 9336 3056 9364
rect 2740 9324 2746 9336
rect 3050 9324 3056 9336
rect 3108 9324 3114 9376
rect 4065 9367 4123 9373
rect 4065 9333 4077 9367
rect 4111 9364 4123 9367
rect 4798 9364 4804 9376
rect 4111 9336 4804 9364
rect 4111 9333 4123 9336
rect 4065 9327 4123 9333
rect 4798 9324 4804 9336
rect 4856 9364 4862 9376
rect 5442 9364 5448 9376
rect 4856 9336 5448 9364
rect 4856 9324 4862 9336
rect 5442 9324 5448 9336
rect 5500 9324 5506 9376
rect 6270 9324 6276 9376
rect 6328 9364 6334 9376
rect 6454 9364 6460 9376
rect 6328 9336 6460 9364
rect 6328 9324 6334 9336
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 6564 9364 6592 9404
rect 7926 9364 7932 9376
rect 6564 9336 7932 9364
rect 7926 9324 7932 9336
rect 7984 9324 7990 9376
rect 8754 9364 8760 9376
rect 8715 9336 8760 9364
rect 8754 9324 8760 9336
rect 8812 9324 8818 9376
rect 8846 9324 8852 9376
rect 8904 9364 8910 9376
rect 9125 9367 9183 9373
rect 9125 9364 9137 9367
rect 8904 9336 9137 9364
rect 8904 9324 8910 9336
rect 9125 9333 9137 9336
rect 9171 9333 9183 9367
rect 9125 9327 9183 9333
rect 9217 9367 9275 9373
rect 9217 9333 9229 9367
rect 9263 9364 9275 9367
rect 9591 9364 9619 9404
rect 9692 9376 9720 9404
rect 9263 9336 9619 9364
rect 9263 9333 9275 9336
rect 9217 9327 9275 9333
rect 9674 9324 9680 9376
rect 9732 9324 9738 9376
rect 9769 9367 9827 9373
rect 9769 9333 9781 9367
rect 9815 9364 9827 9367
rect 10042 9364 10048 9376
rect 9815 9336 10048 9364
rect 9815 9333 9827 9336
rect 9769 9327 9827 9333
rect 10042 9324 10048 9336
rect 10100 9324 10106 9376
rect 10137 9367 10195 9373
rect 10137 9333 10149 9367
rect 10183 9364 10195 9367
rect 10318 9364 10324 9376
rect 10183 9336 10324 9364
rect 10183 9333 10195 9336
rect 10137 9327 10195 9333
rect 10318 9324 10324 9336
rect 10376 9324 10382 9376
rect 10879 9364 10907 9404
rect 12158 9392 12164 9404
rect 12216 9392 12222 9444
rect 14452 9435 14510 9441
rect 14452 9401 14464 9435
rect 14498 9432 14510 9435
rect 16666 9432 16672 9444
rect 14498 9404 16672 9432
rect 14498 9401 14510 9404
rect 14452 9395 14510 9401
rect 16666 9392 16672 9404
rect 16724 9392 16730 9444
rect 11238 9364 11244 9376
rect 10879 9336 11244 9364
rect 11238 9324 11244 9336
rect 11296 9324 11302 9376
rect 12805 9367 12863 9373
rect 12805 9333 12817 9367
rect 12851 9364 12863 9367
rect 13170 9364 13176 9376
rect 12851 9336 13176 9364
rect 12851 9333 12863 9336
rect 12805 9327 12863 9333
rect 13170 9324 13176 9336
rect 13228 9324 13234 9376
rect 13814 9324 13820 9376
rect 13872 9364 13878 9376
rect 14366 9364 14372 9376
rect 13872 9336 14372 9364
rect 13872 9324 13878 9336
rect 14366 9324 14372 9336
rect 14424 9364 14430 9376
rect 15286 9364 15292 9376
rect 14424 9336 15292 9364
rect 14424 9324 14430 9336
rect 15286 9324 15292 9336
rect 15344 9324 15350 9376
rect 16206 9364 16212 9376
rect 16167 9336 16212 9364
rect 16206 9324 16212 9336
rect 16264 9324 16270 9376
rect 16758 9364 16764 9376
rect 16719 9336 16764 9364
rect 16758 9324 16764 9336
rect 16816 9324 16822 9376
rect 16850 9324 16856 9376
rect 16908 9364 16914 9376
rect 17221 9367 17279 9373
rect 17221 9364 17233 9367
rect 16908 9336 17233 9364
rect 16908 9324 16914 9336
rect 17221 9333 17233 9336
rect 17267 9333 17279 9367
rect 17221 9327 17279 9333
rect 1104 9274 18860 9296
rect 1104 9222 6912 9274
rect 6964 9222 6976 9274
rect 7028 9222 7040 9274
rect 7092 9222 7104 9274
rect 7156 9222 12843 9274
rect 12895 9222 12907 9274
rect 12959 9222 12971 9274
rect 13023 9222 13035 9274
rect 13087 9222 18860 9274
rect 1104 9200 18860 9222
rect 2958 9160 2964 9172
rect 2919 9132 2964 9160
rect 2958 9120 2964 9132
rect 3016 9120 3022 9172
rect 5810 9120 5816 9172
rect 5868 9160 5874 9172
rect 5905 9163 5963 9169
rect 5905 9160 5917 9163
rect 5868 9132 5917 9160
rect 5868 9120 5874 9132
rect 5905 9129 5917 9132
rect 5951 9129 5963 9163
rect 5905 9123 5963 9129
rect 7101 9163 7159 9169
rect 7101 9129 7113 9163
rect 7147 9160 7159 9163
rect 7282 9160 7288 9172
rect 7147 9132 7288 9160
rect 7147 9129 7159 9132
rect 7101 9123 7159 9129
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 7466 9160 7472 9172
rect 7427 9132 7472 9160
rect 7466 9120 7472 9132
rect 7524 9120 7530 9172
rect 7561 9163 7619 9169
rect 7561 9129 7573 9163
rect 7607 9160 7619 9163
rect 7926 9160 7932 9172
rect 7607 9132 7932 9160
rect 7607 9129 7619 9132
rect 7561 9123 7619 9129
rect 7926 9120 7932 9132
rect 7984 9120 7990 9172
rect 8389 9163 8447 9169
rect 8389 9129 8401 9163
rect 8435 9160 8447 9163
rect 8846 9160 8852 9172
rect 8435 9132 8852 9160
rect 8435 9129 8447 9132
rect 8389 9123 8447 9129
rect 8846 9120 8852 9132
rect 8904 9120 8910 9172
rect 10594 9120 10600 9172
rect 10652 9160 10658 9172
rect 12345 9163 12403 9169
rect 12345 9160 12357 9163
rect 10652 9132 12357 9160
rect 10652 9120 10658 9132
rect 12345 9129 12357 9132
rect 12391 9129 12403 9163
rect 12345 9123 12403 9129
rect 12989 9163 13047 9169
rect 12989 9129 13001 9163
rect 13035 9160 13047 9163
rect 13170 9160 13176 9172
rect 13035 9132 13176 9160
rect 13035 9129 13047 9132
rect 12989 9123 13047 9129
rect 1848 9095 1906 9101
rect 1848 9061 1860 9095
rect 1894 9092 1906 9095
rect 2682 9092 2688 9104
rect 1894 9064 2688 9092
rect 1894 9061 1906 9064
rect 1848 9055 1906 9061
rect 2682 9052 2688 9064
rect 2740 9052 2746 9104
rect 3970 9052 3976 9104
rect 4028 9092 4034 9104
rect 5718 9092 5724 9104
rect 4028 9064 5724 9092
rect 4028 9052 4034 9064
rect 5718 9052 5724 9064
rect 5776 9092 5782 9104
rect 6270 9092 6276 9104
rect 5776 9064 6132 9092
rect 6231 9064 6276 9092
rect 5776 9052 5782 9064
rect 1578 9024 1584 9036
rect 1539 8996 1584 9024
rect 1578 8984 1584 8996
rect 1636 8984 1642 9036
rect 4062 9024 4068 9036
rect 4023 8996 4068 9024
rect 4062 8984 4068 8996
rect 4120 8984 4126 9036
rect 4332 9027 4390 9033
rect 4332 8993 4344 9027
rect 4378 9024 4390 9027
rect 4890 9024 4896 9036
rect 4378 8996 4896 9024
rect 4378 8993 4390 8996
rect 4332 8987 4390 8993
rect 4890 8984 4896 8996
rect 4948 8984 4954 9036
rect 6104 9024 6132 9064
rect 6270 9052 6276 9064
rect 6328 9092 6334 9104
rect 8757 9095 8815 9101
rect 8757 9092 8769 9095
rect 6328 9064 8769 9092
rect 6328 9052 6334 9064
rect 8757 9061 8769 9064
rect 8803 9092 8815 9095
rect 9674 9092 9680 9104
rect 8803 9064 9680 9092
rect 8803 9061 8815 9064
rect 8757 9055 8815 9061
rect 9674 9052 9680 9064
rect 9732 9052 9738 9104
rect 9766 9052 9772 9104
rect 9824 9092 9830 9104
rect 10045 9095 10103 9101
rect 10045 9092 10057 9095
rect 9824 9064 10057 9092
rect 9824 9052 9830 9064
rect 10045 9061 10057 9064
rect 10091 9061 10103 9095
rect 12360 9092 12388 9123
rect 13170 9120 13176 9132
rect 13228 9120 13234 9172
rect 14182 9160 14188 9172
rect 14143 9132 14188 9160
rect 14182 9120 14188 9132
rect 14240 9120 14246 9172
rect 16574 9120 16580 9172
rect 16632 9160 16638 9172
rect 16669 9163 16727 9169
rect 16669 9160 16681 9163
rect 16632 9132 16681 9160
rect 16632 9120 16638 9132
rect 16669 9129 16681 9132
rect 16715 9129 16727 9163
rect 16669 9123 16727 9129
rect 16758 9120 16764 9172
rect 16816 9160 16822 9172
rect 17589 9163 17647 9169
rect 17589 9160 17601 9163
rect 16816 9132 17601 9160
rect 16816 9120 16822 9132
rect 17589 9129 17601 9132
rect 17635 9129 17647 9163
rect 17589 9123 17647 9129
rect 13078 9092 13084 9104
rect 12360 9064 13084 9092
rect 10045 9055 10103 9061
rect 13078 9052 13084 9064
rect 13136 9052 13142 9104
rect 13357 9095 13415 9101
rect 13357 9061 13369 9095
rect 13403 9092 13415 9095
rect 13403 9064 13768 9092
rect 13403 9061 13415 9064
rect 13357 9055 13415 9061
rect 6365 9027 6423 9033
rect 6365 9024 6377 9027
rect 6104 8996 6377 9024
rect 6365 8993 6377 8996
rect 6411 9024 6423 9027
rect 10505 9027 10563 9033
rect 6411 8996 8524 9024
rect 6411 8993 6423 8996
rect 6365 8987 6423 8993
rect 6546 8956 6552 8968
rect 6459 8928 6552 8956
rect 6546 8916 6552 8928
rect 6604 8916 6610 8968
rect 7653 8959 7711 8965
rect 7653 8925 7665 8959
rect 7699 8925 7711 8959
rect 8496 8956 8524 8996
rect 9048 8996 10364 9024
rect 9048 8965 9076 8996
rect 8849 8959 8907 8965
rect 8849 8956 8861 8959
rect 8496 8928 8861 8956
rect 7653 8919 7711 8925
rect 8849 8925 8861 8928
rect 8895 8925 8907 8959
rect 8849 8919 8907 8925
rect 9033 8959 9091 8965
rect 9033 8925 9045 8959
rect 9079 8925 9091 8959
rect 9033 8919 9091 8925
rect 6564 8888 6592 8916
rect 7668 8888 7696 8919
rect 6564 8860 7696 8888
rect 8864 8832 8892 8919
rect 9398 8916 9404 8968
rect 9456 8956 9462 8968
rect 10336 8965 10364 8996
rect 10505 8993 10517 9027
rect 10551 9024 10563 9027
rect 10686 9024 10692 9036
rect 10551 8996 10692 9024
rect 10551 8993 10563 8996
rect 10505 8987 10563 8993
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 10870 8984 10876 9036
rect 10928 9024 10934 9036
rect 10965 9027 11023 9033
rect 10965 9024 10977 9027
rect 10928 8996 10977 9024
rect 10928 8984 10934 8996
rect 10965 8993 10977 8996
rect 11011 8993 11023 9027
rect 11232 9027 11290 9033
rect 11232 9024 11244 9027
rect 10965 8987 11023 8993
rect 11072 8996 11244 9024
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 9456 8928 10149 8956
rect 9456 8916 9462 8928
rect 10137 8925 10149 8928
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 10321 8959 10379 8965
rect 10321 8925 10333 8959
rect 10367 8956 10379 8959
rect 11072 8956 11100 8996
rect 11232 8993 11244 8996
rect 11278 9024 11290 9027
rect 11698 9024 11704 9036
rect 11278 8996 11704 9024
rect 11278 8993 11290 8996
rect 11232 8987 11290 8993
rect 11698 8984 11704 8996
rect 11756 8984 11762 9036
rect 12342 8984 12348 9036
rect 12400 9024 12406 9036
rect 13372 9024 13400 9055
rect 12400 8996 13400 9024
rect 12400 8984 12406 8996
rect 10367 8928 11100 8956
rect 10367 8925 10379 8928
rect 10321 8919 10379 8925
rect 13354 8916 13360 8968
rect 13412 8956 13418 8968
rect 13449 8959 13507 8965
rect 13449 8956 13461 8959
rect 13412 8928 13461 8956
rect 13412 8916 13418 8928
rect 13449 8925 13461 8928
rect 13495 8925 13507 8959
rect 13630 8956 13636 8968
rect 13591 8928 13636 8956
rect 13449 8919 13507 8925
rect 13630 8916 13636 8928
rect 13688 8916 13694 8968
rect 9677 8891 9735 8897
rect 9677 8857 9689 8891
rect 9723 8888 9735 8891
rect 13740 8888 13768 9064
rect 13906 9052 13912 9104
rect 13964 9092 13970 9104
rect 13964 9064 14504 9092
rect 13964 9052 13970 9064
rect 14476 9033 14504 9064
rect 16206 9052 16212 9104
rect 16264 9092 16270 9104
rect 18506 9092 18512 9104
rect 16264 9064 18512 9092
rect 16264 9052 16270 9064
rect 18506 9052 18512 9064
rect 18564 9052 18570 9104
rect 14369 9027 14427 9033
rect 14369 9024 14381 9027
rect 13924 8996 14381 9024
rect 13924 8968 13952 8996
rect 14369 8993 14381 8996
rect 14415 8993 14427 9027
rect 14369 8987 14427 8993
rect 14461 9027 14519 9033
rect 14461 8993 14473 9027
rect 14507 8993 14519 9027
rect 14461 8987 14519 8993
rect 15556 9027 15614 9033
rect 15556 8993 15568 9027
rect 15602 9024 15614 9027
rect 16666 9024 16672 9036
rect 15602 8996 16672 9024
rect 15602 8993 15614 8996
rect 15556 8987 15614 8993
rect 16666 8984 16672 8996
rect 16724 8984 16730 9036
rect 17497 9027 17555 9033
rect 17497 8993 17509 9027
rect 17543 9024 17555 9027
rect 18322 9024 18328 9036
rect 17543 8996 18328 9024
rect 17543 8993 17555 8996
rect 17497 8987 17555 8993
rect 18322 8984 18328 8996
rect 18380 8984 18386 9036
rect 13906 8916 13912 8968
rect 13964 8916 13970 8968
rect 14182 8916 14188 8968
rect 14240 8956 14246 8968
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 14240 8928 15301 8956
rect 14240 8916 14246 8928
rect 15289 8925 15301 8928
rect 15335 8925 15347 8959
rect 15289 8919 15347 8925
rect 16574 8916 16580 8968
rect 16632 8956 16638 8968
rect 17681 8959 17739 8965
rect 17681 8956 17693 8959
rect 16632 8928 17693 8956
rect 16632 8916 16638 8928
rect 17681 8925 17693 8928
rect 17727 8925 17739 8959
rect 17681 8919 17739 8925
rect 9723 8860 11015 8888
rect 13740 8860 15332 8888
rect 9723 8857 9735 8860
rect 9677 8851 9735 8857
rect 2682 8780 2688 8832
rect 2740 8820 2746 8832
rect 4706 8820 4712 8832
rect 2740 8792 4712 8820
rect 2740 8780 2746 8792
rect 4706 8780 4712 8792
rect 4764 8820 4770 8832
rect 5445 8823 5503 8829
rect 5445 8820 5457 8823
rect 4764 8792 5457 8820
rect 4764 8780 4770 8792
rect 5445 8789 5457 8792
rect 5491 8789 5503 8823
rect 5445 8783 5503 8789
rect 7926 8780 7932 8832
rect 7984 8820 7990 8832
rect 8478 8820 8484 8832
rect 7984 8792 8484 8820
rect 7984 8780 7990 8792
rect 8478 8780 8484 8792
rect 8536 8780 8542 8832
rect 8846 8780 8852 8832
rect 8904 8780 8910 8832
rect 9490 8780 9496 8832
rect 9548 8820 9554 8832
rect 10689 8823 10747 8829
rect 10689 8820 10701 8823
rect 9548 8792 10701 8820
rect 9548 8780 9554 8792
rect 10689 8789 10701 8792
rect 10735 8789 10747 8823
rect 10987 8820 11015 8860
rect 12894 8820 12900 8832
rect 10987 8792 12900 8820
rect 10689 8783 10747 8789
rect 12894 8780 12900 8792
rect 12952 8780 12958 8832
rect 14645 8823 14703 8829
rect 14645 8789 14657 8823
rect 14691 8820 14703 8823
rect 15194 8820 15200 8832
rect 14691 8792 15200 8820
rect 14691 8789 14703 8792
rect 14645 8783 14703 8789
rect 15194 8780 15200 8792
rect 15252 8780 15258 8832
rect 15304 8820 15332 8860
rect 17034 8848 17040 8900
rect 17092 8888 17098 8900
rect 17129 8891 17187 8897
rect 17129 8888 17141 8891
rect 17092 8860 17141 8888
rect 17092 8848 17098 8860
rect 17129 8857 17141 8860
rect 17175 8857 17187 8891
rect 17129 8851 17187 8857
rect 17862 8820 17868 8832
rect 15304 8792 17868 8820
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 1104 8730 18860 8752
rect 1104 8678 3947 8730
rect 3999 8678 4011 8730
rect 4063 8678 4075 8730
rect 4127 8678 4139 8730
rect 4191 8678 9878 8730
rect 9930 8678 9942 8730
rect 9994 8678 10006 8730
rect 10058 8678 10070 8730
rect 10122 8678 15808 8730
rect 15860 8678 15872 8730
rect 15924 8678 15936 8730
rect 15988 8678 16000 8730
rect 16052 8678 18860 8730
rect 1104 8656 18860 8678
rect 4249 8619 4307 8625
rect 4249 8585 4261 8619
rect 4295 8616 4307 8619
rect 4522 8616 4528 8628
rect 4295 8588 4528 8616
rect 4295 8585 4307 8588
rect 4249 8579 4307 8585
rect 4522 8576 4528 8588
rect 4580 8576 4586 8628
rect 5534 8576 5540 8628
rect 5592 8616 5598 8628
rect 6641 8619 6699 8625
rect 6641 8616 6653 8619
rect 5592 8588 6653 8616
rect 5592 8576 5598 8588
rect 6641 8585 6653 8588
rect 6687 8616 6699 8619
rect 7190 8616 7196 8628
rect 6687 8588 7196 8616
rect 6687 8585 6699 8588
rect 6641 8579 6699 8585
rect 7190 8576 7196 8588
rect 7248 8576 7254 8628
rect 7377 8619 7435 8625
rect 7377 8585 7389 8619
rect 7423 8616 7435 8619
rect 8294 8616 8300 8628
rect 7423 8588 8300 8616
rect 7423 8585 7435 8588
rect 7377 8579 7435 8585
rect 8294 8576 8300 8588
rect 8352 8576 8358 8628
rect 12342 8616 12348 8628
rect 9876 8588 12348 8616
rect 1578 8508 1584 8560
rect 1636 8548 1642 8560
rect 1857 8551 1915 8557
rect 1857 8548 1869 8551
rect 1636 8520 1869 8548
rect 1636 8508 1642 8520
rect 1857 8517 1869 8520
rect 1903 8517 1915 8551
rect 1857 8511 1915 8517
rect 2130 8508 2136 8560
rect 2188 8548 2194 8560
rect 7009 8551 7067 8557
rect 7009 8548 7021 8551
rect 2188 8520 7021 8548
rect 2188 8508 2194 8520
rect 7009 8517 7021 8520
rect 7055 8517 7067 8551
rect 7009 8511 7067 8517
rect 2501 8483 2559 8489
rect 2501 8449 2513 8483
rect 2547 8480 2559 8483
rect 2958 8480 2964 8492
rect 2547 8452 2964 8480
rect 2547 8449 2559 8452
rect 2501 8443 2559 8449
rect 2958 8440 2964 8452
rect 3016 8440 3022 8492
rect 3513 8483 3571 8489
rect 3513 8449 3525 8483
rect 3559 8480 3571 8483
rect 3602 8480 3608 8492
rect 3559 8452 3608 8480
rect 3559 8449 3571 8452
rect 3513 8443 3571 8449
rect 2317 8415 2375 8421
rect 2317 8381 2329 8415
rect 2363 8412 2375 8415
rect 2866 8412 2872 8424
rect 2363 8384 2872 8412
rect 2363 8381 2375 8384
rect 2317 8375 2375 8381
rect 2866 8372 2872 8384
rect 2924 8372 2930 8424
rect 3050 8372 3056 8424
rect 3108 8412 3114 8424
rect 3421 8415 3479 8421
rect 3421 8412 3433 8415
rect 3108 8384 3433 8412
rect 3108 8372 3114 8384
rect 3421 8381 3433 8384
rect 3467 8381 3479 8415
rect 3421 8375 3479 8381
rect 2406 8304 2412 8356
rect 2464 8344 2470 8356
rect 3528 8344 3556 8443
rect 3602 8440 3608 8452
rect 3660 8440 3666 8492
rect 3697 8483 3755 8489
rect 3697 8449 3709 8483
rect 3743 8480 3755 8483
rect 4522 8480 4528 8492
rect 3743 8452 4528 8480
rect 3743 8449 3755 8452
rect 3697 8443 3755 8449
rect 4522 8440 4528 8452
rect 4580 8480 4586 8492
rect 4890 8480 4896 8492
rect 4580 8452 4896 8480
rect 4580 8440 4586 8452
rect 4890 8440 4896 8452
rect 4948 8440 4954 8492
rect 5994 8440 6000 8492
rect 6052 8480 6058 8492
rect 6052 8452 6097 8480
rect 6052 8440 6058 8452
rect 6730 8440 6736 8492
rect 6788 8480 6794 8492
rect 6788 8452 7236 8480
rect 6788 8440 6794 8452
rect 4338 8372 4344 8424
rect 4396 8412 4402 8424
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 4396 8384 6837 8412
rect 4396 8372 4402 8384
rect 6825 8381 6837 8384
rect 6871 8381 6883 8415
rect 7208 8412 7236 8452
rect 7282 8440 7288 8492
rect 7340 8480 7346 8492
rect 7558 8480 7564 8492
rect 7340 8452 7564 8480
rect 7340 8440 7346 8452
rect 7558 8440 7564 8452
rect 7616 8480 7622 8492
rect 7837 8483 7895 8489
rect 7837 8480 7849 8483
rect 7616 8452 7849 8480
rect 7616 8440 7622 8452
rect 7837 8449 7849 8452
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 8021 8483 8079 8489
rect 8021 8449 8033 8483
rect 8067 8480 8079 8483
rect 8202 8480 8208 8492
rect 8067 8452 8208 8480
rect 8067 8449 8079 8452
rect 8021 8443 8079 8449
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 8573 8415 8631 8421
rect 8573 8412 8585 8415
rect 7208 8384 7788 8412
rect 6825 8375 6883 8381
rect 2464 8316 3556 8344
rect 4617 8347 4675 8353
rect 2464 8304 2470 8316
rect 4617 8313 4629 8347
rect 4663 8344 4675 8347
rect 4663 8316 5488 8344
rect 4663 8313 4675 8316
rect 4617 8307 4675 8313
rect 2222 8276 2228 8288
rect 2183 8248 2228 8276
rect 2222 8236 2228 8248
rect 2280 8236 2286 8288
rect 3050 8276 3056 8288
rect 3011 8248 3056 8276
rect 3050 8236 3056 8248
rect 3108 8236 3114 8288
rect 4709 8279 4767 8285
rect 4709 8245 4721 8279
rect 4755 8276 4767 8279
rect 5074 8276 5080 8288
rect 4755 8248 5080 8276
rect 4755 8245 4767 8248
rect 4709 8239 4767 8245
rect 5074 8236 5080 8248
rect 5132 8236 5138 8288
rect 5460 8285 5488 8316
rect 5626 8304 5632 8356
rect 5684 8344 5690 8356
rect 5813 8347 5871 8353
rect 5813 8344 5825 8347
rect 5684 8316 5825 8344
rect 5684 8304 5690 8316
rect 5813 8313 5825 8316
rect 5859 8313 5871 8347
rect 5813 8307 5871 8313
rect 5905 8347 5963 8353
rect 5905 8313 5917 8347
rect 5951 8344 5963 8347
rect 6641 8347 6699 8353
rect 6641 8344 6653 8347
rect 5951 8316 6653 8344
rect 5951 8313 5963 8316
rect 5905 8307 5963 8313
rect 6641 8313 6653 8316
rect 6687 8313 6699 8347
rect 6840 8344 6868 8375
rect 7558 8344 7564 8356
rect 6840 8316 7564 8344
rect 6641 8307 6699 8313
rect 5445 8279 5503 8285
rect 5445 8245 5457 8279
rect 5491 8245 5503 8279
rect 5828 8276 5856 8307
rect 7558 8304 7564 8316
rect 7616 8304 7622 8356
rect 7466 8276 7472 8288
rect 5828 8248 7472 8276
rect 5445 8239 5503 8245
rect 7466 8236 7472 8248
rect 7524 8236 7530 8288
rect 7760 8285 7788 8384
rect 8496 8384 8585 8412
rect 7926 8304 7932 8356
rect 7984 8344 7990 8356
rect 8496 8344 8524 8384
rect 8573 8381 8585 8384
rect 8619 8381 8631 8415
rect 9876 8412 9904 8588
rect 12342 8576 12348 8588
rect 12400 8576 12406 8628
rect 13354 8576 13360 8628
rect 13412 8616 13418 8628
rect 14001 8619 14059 8625
rect 13412 8588 13952 8616
rect 13412 8576 13418 8588
rect 10244 8520 10456 8548
rect 10244 8480 10272 8520
rect 10428 8489 10456 8520
rect 12066 8508 12072 8560
rect 12124 8548 12130 8560
rect 13924 8548 13952 8588
rect 14001 8585 14013 8619
rect 14047 8616 14059 8619
rect 15286 8616 15292 8628
rect 14047 8588 15292 8616
rect 14047 8585 14059 8588
rect 14001 8579 14059 8585
rect 15286 8576 15292 8588
rect 15344 8576 15350 8628
rect 16390 8616 16396 8628
rect 16351 8588 16396 8616
rect 16390 8576 16396 8588
rect 16448 8576 16454 8628
rect 17034 8576 17040 8628
rect 17092 8616 17098 8628
rect 17954 8616 17960 8628
rect 17092 8588 17960 8616
rect 17092 8576 17098 8588
rect 17954 8576 17960 8588
rect 18012 8576 18018 8628
rect 14090 8548 14096 8560
rect 12124 8520 13860 8548
rect 13924 8520 14096 8548
rect 12124 8508 12130 8520
rect 9968 8452 10272 8480
rect 10413 8483 10471 8489
rect 9968 8424 9996 8452
rect 10413 8449 10425 8483
rect 10459 8449 10471 8483
rect 12894 8480 12900 8492
rect 12855 8452 12900 8480
rect 10413 8443 10471 8449
rect 12894 8440 12900 8452
rect 12952 8440 12958 8492
rect 13078 8480 13084 8492
rect 13039 8452 13084 8480
rect 13078 8440 13084 8452
rect 13136 8440 13142 8492
rect 8573 8375 8631 8381
rect 8772 8384 9904 8412
rect 8772 8344 8800 8384
rect 9950 8372 9956 8424
rect 10008 8372 10014 8424
rect 10321 8415 10379 8421
rect 10321 8381 10333 8415
rect 10367 8412 10379 8415
rect 11238 8412 11244 8424
rect 10367 8384 11244 8412
rect 10367 8381 10379 8384
rect 10321 8375 10379 8381
rect 11238 8372 11244 8384
rect 11296 8412 11302 8424
rect 13832 8421 13860 8520
rect 14090 8508 14096 8520
rect 14148 8508 14154 8560
rect 15933 8551 15991 8557
rect 15933 8517 15945 8551
rect 15979 8548 15991 8551
rect 16666 8548 16672 8560
rect 15979 8520 16672 8548
rect 15979 8517 15991 8520
rect 15933 8511 15991 8517
rect 16666 8508 16672 8520
rect 16724 8548 16730 8560
rect 17218 8548 17224 8560
rect 16724 8520 17224 8548
rect 16724 8508 16730 8520
rect 17218 8508 17224 8520
rect 17276 8508 17282 8560
rect 14182 8440 14188 8492
rect 14240 8480 14246 8492
rect 14553 8483 14611 8489
rect 14553 8480 14565 8483
rect 14240 8452 14565 8480
rect 14240 8440 14246 8452
rect 14553 8449 14565 8452
rect 14599 8449 14611 8483
rect 14553 8443 14611 8449
rect 16574 8440 16580 8492
rect 16632 8480 16638 8492
rect 16945 8483 17003 8489
rect 16945 8480 16957 8483
rect 16632 8452 16957 8480
rect 16632 8440 16638 8452
rect 16945 8449 16957 8452
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 13817 8415 13875 8421
rect 11296 8384 13391 8412
rect 11296 8372 11302 8384
rect 10686 8353 10692 8356
rect 7984 8316 8524 8344
rect 8680 8316 8800 8344
rect 7984 8304 7990 8316
rect 7745 8279 7803 8285
rect 7745 8245 7757 8279
rect 7791 8276 7803 8279
rect 8680 8276 8708 8316
rect 10680 8307 10692 8353
rect 10744 8344 10750 8356
rect 12802 8344 12808 8356
rect 10744 8316 10780 8344
rect 12763 8316 12808 8344
rect 10686 8304 10692 8307
rect 10744 8304 10750 8316
rect 12802 8304 12808 8316
rect 12860 8344 12866 8356
rect 13265 8347 13323 8353
rect 13265 8344 13277 8347
rect 12860 8316 13277 8344
rect 12860 8304 12866 8316
rect 13265 8313 13277 8316
rect 13311 8313 13323 8347
rect 13363 8344 13391 8384
rect 13817 8381 13829 8415
rect 13863 8381 13875 8415
rect 13817 8375 13875 8381
rect 14820 8415 14878 8421
rect 14820 8381 14832 8415
rect 14866 8412 14878 8415
rect 15838 8412 15844 8424
rect 14866 8384 15844 8412
rect 14866 8381 14878 8384
rect 14820 8375 14878 8381
rect 15838 8372 15844 8384
rect 15896 8372 15902 8424
rect 14090 8344 14096 8356
rect 13363 8316 14096 8344
rect 13265 8307 13323 8313
rect 14090 8304 14096 8316
rect 14148 8304 14154 8356
rect 15194 8304 15200 8356
rect 15252 8344 15258 8356
rect 15746 8344 15752 8356
rect 15252 8316 15752 8344
rect 15252 8304 15258 8316
rect 15746 8304 15752 8316
rect 15804 8304 15810 8356
rect 16666 8304 16672 8356
rect 16724 8344 16730 8356
rect 16853 8347 16911 8353
rect 16853 8344 16865 8347
rect 16724 8316 16865 8344
rect 16724 8304 16730 8316
rect 16853 8313 16865 8316
rect 16899 8313 16911 8347
rect 16853 8307 16911 8313
rect 7791 8248 8708 8276
rect 7791 8245 7803 8248
rect 7745 8239 7803 8245
rect 8846 8236 8852 8288
rect 8904 8276 8910 8288
rect 11238 8276 11244 8288
rect 8904 8248 11244 8276
rect 8904 8236 8910 8248
rect 11238 8236 11244 8248
rect 11296 8236 11302 8288
rect 11698 8236 11704 8288
rect 11756 8276 11762 8288
rect 11793 8279 11851 8285
rect 11793 8276 11805 8279
rect 11756 8248 11805 8276
rect 11756 8236 11762 8248
rect 11793 8245 11805 8248
rect 11839 8245 11851 8279
rect 11793 8239 11851 8245
rect 12434 8236 12440 8288
rect 12492 8276 12498 8288
rect 16758 8276 16764 8288
rect 12492 8248 12537 8276
rect 16719 8248 16764 8276
rect 12492 8236 12498 8248
rect 16758 8236 16764 8248
rect 16816 8236 16822 8288
rect 1104 8186 18860 8208
rect 1104 8134 6912 8186
rect 6964 8134 6976 8186
rect 7028 8134 7040 8186
rect 7092 8134 7104 8186
rect 7156 8134 12843 8186
rect 12895 8134 12907 8186
rect 12959 8134 12971 8186
rect 13023 8134 13035 8186
rect 13087 8134 18860 8186
rect 1104 8112 18860 8134
rect 3053 8075 3111 8081
rect 3053 8041 3065 8075
rect 3099 8072 3111 8075
rect 3234 8072 3240 8084
rect 3099 8044 3240 8072
rect 3099 8041 3111 8044
rect 3053 8035 3111 8041
rect 3234 8032 3240 8044
rect 3292 8032 3298 8084
rect 4614 8032 4620 8084
rect 4672 8072 4678 8084
rect 4672 8044 6408 8072
rect 4672 8032 4678 8044
rect 3145 8007 3203 8013
rect 3145 7973 3157 8007
rect 3191 8004 3203 8007
rect 4338 8004 4344 8016
rect 3191 7976 4344 8004
rect 3191 7973 3203 7976
rect 3145 7967 3203 7973
rect 4338 7964 4344 7976
rect 4396 7964 4402 8016
rect 6270 8004 6276 8016
rect 4816 7976 6276 8004
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 4816 7936 4844 7976
rect 6270 7964 6276 7976
rect 6328 7964 6334 8016
rect 6380 8004 6408 8044
rect 7466 8032 7472 8084
rect 7524 8072 7530 8084
rect 9398 8072 9404 8084
rect 7524 8044 9404 8072
rect 7524 8032 7530 8044
rect 9398 8032 9404 8044
rect 9456 8032 9462 8084
rect 12069 8075 12127 8081
rect 12069 8041 12081 8075
rect 12115 8072 12127 8075
rect 12434 8072 12440 8084
rect 12115 8044 12440 8072
rect 12115 8041 12127 8044
rect 12069 8035 12127 8041
rect 12434 8032 12440 8044
rect 12492 8032 12498 8084
rect 13814 8032 13820 8084
rect 13872 8072 13878 8084
rect 15841 8075 15899 8081
rect 15841 8072 15853 8075
rect 13872 8044 15853 8072
rect 13872 8032 13878 8044
rect 15841 8041 15853 8044
rect 15887 8041 15899 8075
rect 15841 8035 15899 8041
rect 15933 8075 15991 8081
rect 15933 8041 15945 8075
rect 15979 8072 15991 8075
rect 16022 8072 16028 8084
rect 15979 8044 16028 8072
rect 15979 8041 15991 8044
rect 15933 8035 15991 8041
rect 16022 8032 16028 8044
rect 16080 8032 16086 8084
rect 16669 8075 16727 8081
rect 16669 8041 16681 8075
rect 16715 8072 16727 8075
rect 16758 8072 16764 8084
rect 16715 8044 16764 8072
rect 16715 8041 16727 8044
rect 16669 8035 16727 8041
rect 16758 8032 16764 8044
rect 16816 8032 16822 8084
rect 10042 8004 10048 8016
rect 6380 7976 8708 8004
rect 5994 7945 6000 7948
rect 1719 7908 4844 7936
rect 4893 7939 4951 7945
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 4893 7905 4905 7939
rect 4939 7936 4951 7939
rect 5988 7936 6000 7945
rect 4939 7908 5120 7936
rect 4939 7905 4951 7908
rect 4893 7899 4951 7905
rect 3329 7871 3387 7877
rect 3329 7837 3341 7871
rect 3375 7868 3387 7871
rect 4522 7868 4528 7880
rect 3375 7840 4528 7868
rect 3375 7837 3387 7840
rect 3329 7831 3387 7837
rect 4522 7828 4528 7840
rect 4580 7828 4586 7880
rect 4706 7828 4712 7880
rect 4764 7868 4770 7880
rect 4985 7871 5043 7877
rect 4985 7868 4997 7871
rect 4764 7840 4997 7868
rect 4764 7828 4770 7840
rect 4985 7837 4997 7840
rect 5031 7837 5043 7871
rect 4985 7831 5043 7837
rect 1857 7803 1915 7809
rect 1857 7769 1869 7803
rect 1903 7800 1915 7803
rect 3694 7800 3700 7812
rect 1903 7772 3700 7800
rect 1903 7769 1915 7772
rect 1857 7763 1915 7769
rect 3694 7760 3700 7772
rect 3752 7760 3758 7812
rect 5092 7800 5120 7908
rect 5184 7908 6000 7936
rect 5184 7877 5212 7908
rect 5988 7899 6000 7908
rect 5994 7896 6000 7899
rect 6052 7896 6058 7948
rect 7190 7896 7196 7948
rect 7248 7936 7254 7948
rect 7929 7939 7987 7945
rect 7929 7936 7941 7939
rect 7248 7908 7941 7936
rect 7248 7896 7254 7908
rect 7929 7905 7941 7908
rect 7975 7905 7987 7939
rect 7929 7899 7987 7905
rect 8021 7939 8079 7945
rect 8021 7905 8033 7939
rect 8067 7936 8079 7939
rect 8294 7936 8300 7948
rect 8067 7908 8300 7936
rect 8067 7905 8079 7908
rect 8021 7899 8079 7905
rect 8294 7896 8300 7908
rect 8352 7896 8358 7948
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 5350 7828 5356 7880
rect 5408 7868 5414 7880
rect 5721 7871 5779 7877
rect 5721 7868 5733 7871
rect 5408 7840 5733 7868
rect 5408 7828 5414 7840
rect 5721 7837 5733 7840
rect 5767 7837 5779 7871
rect 5721 7831 5779 7837
rect 8113 7871 8171 7877
rect 8113 7837 8125 7871
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 5442 7800 5448 7812
rect 4448 7772 5448 7800
rect 2590 7692 2596 7744
rect 2648 7732 2654 7744
rect 2685 7735 2743 7741
rect 2685 7732 2697 7735
rect 2648 7704 2697 7732
rect 2648 7692 2654 7704
rect 2685 7701 2697 7704
rect 2731 7701 2743 7735
rect 2685 7695 2743 7701
rect 3142 7692 3148 7744
rect 3200 7732 3206 7744
rect 4448 7732 4476 7772
rect 5442 7760 5448 7772
rect 5500 7760 5506 7812
rect 3200 7704 4476 7732
rect 4525 7735 4583 7741
rect 3200 7692 3206 7704
rect 4525 7701 4537 7735
rect 4571 7732 4583 7735
rect 4706 7732 4712 7744
rect 4571 7704 4712 7732
rect 4571 7701 4583 7704
rect 4525 7695 4583 7701
rect 4706 7692 4712 7704
rect 4764 7692 4770 7744
rect 4890 7692 4896 7744
rect 4948 7732 4954 7744
rect 7101 7735 7159 7741
rect 7101 7732 7113 7735
rect 4948 7704 7113 7732
rect 4948 7692 4954 7704
rect 7101 7701 7113 7704
rect 7147 7701 7159 7735
rect 7558 7732 7564 7744
rect 7519 7704 7564 7732
rect 7101 7695 7159 7701
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 8128 7732 8156 7831
rect 8202 7828 8208 7880
rect 8260 7868 8266 7880
rect 8478 7868 8484 7880
rect 8260 7840 8484 7868
rect 8260 7828 8266 7840
rect 8478 7828 8484 7840
rect 8536 7828 8542 7880
rect 8680 7868 8708 7976
rect 8864 7976 10048 8004
rect 8864 7948 8892 7976
rect 10042 7964 10048 7976
rect 10100 7964 10106 8016
rect 10870 7964 10876 8016
rect 10928 8004 10934 8016
rect 11698 8004 11704 8016
rect 10928 7976 11704 8004
rect 10928 7964 10934 7976
rect 11698 7964 11704 7976
rect 11756 7964 11762 8016
rect 12158 8004 12164 8016
rect 12119 7976 12164 8004
rect 12158 7964 12164 7976
rect 12216 7964 12222 8016
rect 17129 8007 17187 8013
rect 17129 8004 17141 8007
rect 12360 7976 17141 8004
rect 8757 7939 8815 7945
rect 8757 7905 8769 7939
rect 8803 7936 8815 7939
rect 8846 7936 8852 7948
rect 8803 7908 8852 7936
rect 8803 7905 8815 7908
rect 8757 7899 8815 7905
rect 8846 7896 8852 7908
rect 8904 7896 8910 7948
rect 9585 7939 9643 7945
rect 9585 7905 9597 7939
rect 9631 7936 9643 7939
rect 9933 7939 9991 7945
rect 9933 7936 9945 7939
rect 9631 7908 9945 7936
rect 9631 7905 9643 7908
rect 9585 7899 9643 7905
rect 9933 7905 9945 7908
rect 9979 7905 9991 7939
rect 9933 7899 9991 7905
rect 12360 7880 12388 7976
rect 17129 7973 17141 7976
rect 17175 7973 17187 8007
rect 17129 7967 17187 7973
rect 13265 7939 13323 7945
rect 13265 7905 13277 7939
rect 13311 7905 13323 7939
rect 13265 7899 13323 7905
rect 13357 7939 13415 7945
rect 13357 7905 13369 7939
rect 13403 7936 13415 7939
rect 13630 7936 13636 7948
rect 13403 7908 13636 7936
rect 13403 7905 13415 7908
rect 13357 7899 13415 7905
rect 9122 7868 9128 7880
rect 8680 7840 9128 7868
rect 9122 7828 9128 7840
rect 9180 7828 9186 7880
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7837 9735 7871
rect 9677 7831 9735 7837
rect 12253 7871 12311 7877
rect 12253 7837 12265 7871
rect 12299 7837 12311 7871
rect 12253 7831 12311 7837
rect 8941 7803 8999 7809
rect 8220 7772 8677 7800
rect 8220 7732 8248 7772
rect 8128 7704 8248 7732
rect 8649 7744 8677 7772
rect 8941 7769 8953 7803
rect 8987 7800 8999 7803
rect 9306 7800 9312 7812
rect 8987 7772 9312 7800
rect 8987 7769 8999 7772
rect 8941 7763 8999 7769
rect 9306 7760 9312 7772
rect 9364 7760 9370 7812
rect 9692 7744 9720 7831
rect 11238 7760 11244 7812
rect 11296 7800 11302 7812
rect 11296 7772 11827 7800
rect 11296 7760 11302 7772
rect 8649 7704 8668 7744
rect 8662 7692 8668 7704
rect 8720 7692 8726 7744
rect 9490 7732 9496 7744
rect 9451 7704 9496 7732
rect 9490 7692 9496 7704
rect 9548 7692 9554 7744
rect 9674 7692 9680 7744
rect 9732 7692 9738 7744
rect 10686 7692 10692 7744
rect 10744 7732 10750 7744
rect 11057 7735 11115 7741
rect 11057 7732 11069 7735
rect 10744 7704 11069 7732
rect 10744 7692 10750 7704
rect 11057 7701 11069 7704
rect 11103 7701 11115 7735
rect 11698 7732 11704 7744
rect 11659 7704 11704 7732
rect 11057 7695 11115 7701
rect 11698 7692 11704 7704
rect 11756 7692 11762 7744
rect 11799 7732 11827 7772
rect 12066 7760 12072 7812
rect 12124 7800 12130 7812
rect 12268 7800 12296 7831
rect 12342 7828 12348 7880
rect 12400 7828 12406 7880
rect 12434 7828 12440 7880
rect 12492 7868 12498 7880
rect 13280 7868 13308 7899
rect 13630 7896 13636 7908
rect 13688 7896 13694 7948
rect 14090 7896 14096 7948
rect 14148 7936 14154 7948
rect 14277 7939 14335 7945
rect 14277 7936 14289 7939
rect 14148 7908 14289 7936
rect 14148 7896 14154 7908
rect 14277 7905 14289 7908
rect 14323 7905 14335 7939
rect 14277 7899 14335 7905
rect 14461 7939 14519 7945
rect 14461 7905 14473 7939
rect 14507 7905 14519 7939
rect 14461 7899 14519 7905
rect 12492 7840 13308 7868
rect 13449 7871 13507 7877
rect 12492 7828 12498 7840
rect 13449 7837 13461 7871
rect 13495 7837 13507 7871
rect 13449 7831 13507 7837
rect 12124 7772 12296 7800
rect 12360 7772 13032 7800
rect 12124 7760 12130 7772
rect 12360 7732 12388 7772
rect 11799 7704 12388 7732
rect 12710 7692 12716 7744
rect 12768 7732 12774 7744
rect 12897 7735 12955 7741
rect 12897 7732 12909 7735
rect 12768 7704 12909 7732
rect 12768 7692 12774 7704
rect 12897 7701 12909 7704
rect 12943 7701 12955 7735
rect 13004 7732 13032 7772
rect 13170 7760 13176 7812
rect 13228 7800 13234 7812
rect 13464 7800 13492 7831
rect 14476 7800 14504 7899
rect 16206 7896 16212 7948
rect 16264 7936 16270 7948
rect 17037 7939 17095 7945
rect 17037 7936 17049 7939
rect 16264 7908 17049 7936
rect 16264 7896 16270 7908
rect 17037 7905 17049 7908
rect 17083 7905 17095 7939
rect 17144 7936 17172 7967
rect 17865 7939 17923 7945
rect 17865 7936 17877 7939
rect 17144 7908 17877 7936
rect 17037 7899 17095 7905
rect 17865 7905 17877 7908
rect 17911 7905 17923 7939
rect 17865 7899 17923 7905
rect 15102 7828 15108 7880
rect 15160 7868 15166 7880
rect 15838 7868 15844 7880
rect 15160 7840 15844 7868
rect 15160 7828 15166 7840
rect 15838 7828 15844 7840
rect 15896 7828 15902 7880
rect 16117 7871 16175 7877
rect 16117 7837 16129 7871
rect 16163 7868 16175 7871
rect 16574 7868 16580 7880
rect 16163 7840 16580 7868
rect 16163 7837 16175 7840
rect 16117 7831 16175 7837
rect 16574 7828 16580 7840
rect 16632 7828 16638 7880
rect 16850 7800 16856 7812
rect 13228 7772 13492 7800
rect 13556 7772 16856 7800
rect 13228 7760 13234 7772
rect 13556 7732 13584 7772
rect 16850 7760 16856 7772
rect 16908 7760 16914 7812
rect 17052 7800 17080 7899
rect 17218 7828 17224 7880
rect 17276 7868 17282 7880
rect 17276 7840 17321 7868
rect 17276 7828 17282 7840
rect 17402 7800 17408 7812
rect 17052 7772 17408 7800
rect 17402 7760 17408 7772
rect 17460 7760 17466 7812
rect 13004 7704 13584 7732
rect 12897 7695 12955 7701
rect 13906 7692 13912 7744
rect 13964 7732 13970 7744
rect 14093 7735 14151 7741
rect 14093 7732 14105 7735
rect 13964 7704 14105 7732
rect 13964 7692 13970 7704
rect 14093 7701 14105 7704
rect 14139 7701 14151 7735
rect 14093 7695 14151 7701
rect 14645 7735 14703 7741
rect 14645 7701 14657 7735
rect 14691 7732 14703 7735
rect 15286 7732 15292 7744
rect 14691 7704 15292 7732
rect 14691 7701 14703 7704
rect 14645 7695 14703 7701
rect 15286 7692 15292 7704
rect 15344 7692 15350 7744
rect 15473 7735 15531 7741
rect 15473 7701 15485 7735
rect 15519 7732 15531 7735
rect 16390 7732 16396 7744
rect 15519 7704 16396 7732
rect 15519 7701 15531 7704
rect 15473 7695 15531 7701
rect 16390 7692 16396 7704
rect 16448 7692 16454 7744
rect 18049 7735 18107 7741
rect 18049 7701 18061 7735
rect 18095 7732 18107 7735
rect 18874 7732 18880 7744
rect 18095 7704 18880 7732
rect 18095 7701 18107 7704
rect 18049 7695 18107 7701
rect 18874 7692 18880 7704
rect 18932 7692 18938 7744
rect 1104 7642 18860 7664
rect 1104 7590 3947 7642
rect 3999 7590 4011 7642
rect 4063 7590 4075 7642
rect 4127 7590 4139 7642
rect 4191 7590 9878 7642
rect 9930 7590 9942 7642
rect 9994 7590 10006 7642
rect 10058 7590 10070 7642
rect 10122 7590 15808 7642
rect 15860 7590 15872 7642
rect 15924 7590 15936 7642
rect 15988 7590 16000 7642
rect 16052 7590 18860 7642
rect 1104 7568 18860 7590
rect 2222 7528 2228 7540
rect 2183 7500 2228 7528
rect 2222 7488 2228 7500
rect 2280 7488 2286 7540
rect 2958 7488 2964 7540
rect 3016 7528 3022 7540
rect 3602 7528 3608 7540
rect 3016 7500 3608 7528
rect 3016 7488 3022 7500
rect 3602 7488 3608 7500
rect 3660 7488 3666 7540
rect 4249 7531 4307 7537
rect 4249 7497 4261 7531
rect 4295 7528 4307 7531
rect 4430 7528 4436 7540
rect 4295 7500 4436 7528
rect 4295 7497 4307 7500
rect 4249 7491 4307 7497
rect 4430 7488 4436 7500
rect 4488 7488 4494 7540
rect 5074 7488 5080 7540
rect 5132 7528 5138 7540
rect 5445 7531 5503 7537
rect 5445 7528 5457 7531
rect 5132 7500 5457 7528
rect 5132 7488 5138 7500
rect 5445 7497 5457 7500
rect 5491 7497 5503 7531
rect 5445 7491 5503 7497
rect 5810 7488 5816 7540
rect 5868 7528 5874 7540
rect 6730 7528 6736 7540
rect 5868 7500 6736 7528
rect 5868 7488 5874 7500
rect 6730 7488 6736 7500
rect 6788 7488 6794 7540
rect 7190 7528 7196 7540
rect 7151 7500 7196 7528
rect 7190 7488 7196 7500
rect 7248 7488 7254 7540
rect 14090 7528 14096 7540
rect 8404 7500 11468 7528
rect 1673 7463 1731 7469
rect 1673 7429 1685 7463
rect 1719 7460 1731 7463
rect 3234 7460 3240 7472
rect 1719 7432 3240 7460
rect 1719 7429 1731 7432
rect 1673 7423 1731 7429
rect 3234 7420 3240 7432
rect 3292 7420 3298 7472
rect 8404 7460 8432 7500
rect 3436 7432 8432 7460
rect 2498 7352 2504 7404
rect 2556 7392 2562 7404
rect 2777 7395 2835 7401
rect 2777 7392 2789 7395
rect 2556 7364 2789 7392
rect 2556 7352 2562 7364
rect 2777 7361 2789 7364
rect 2823 7361 2835 7395
rect 2777 7355 2835 7361
rect 1489 7327 1547 7333
rect 1489 7293 1501 7327
rect 1535 7293 1547 7327
rect 2590 7324 2596 7336
rect 2551 7296 2596 7324
rect 1489 7287 1547 7293
rect 1504 7256 1532 7287
rect 2590 7284 2596 7296
rect 2648 7284 2654 7336
rect 2685 7327 2743 7333
rect 2685 7293 2697 7327
rect 2731 7324 2743 7327
rect 3050 7324 3056 7336
rect 2731 7296 3056 7324
rect 2731 7293 2743 7296
rect 2685 7287 2743 7293
rect 3050 7284 3056 7296
rect 3108 7284 3114 7336
rect 3436 7333 3464 7432
rect 9490 7420 9496 7472
rect 9548 7460 9554 7472
rect 9769 7463 9827 7469
rect 9769 7460 9781 7463
rect 9548 7432 9781 7460
rect 9548 7420 9554 7432
rect 9769 7429 9781 7432
rect 9815 7429 9827 7463
rect 9769 7423 9827 7429
rect 4706 7392 4712 7404
rect 4667 7364 4712 7392
rect 4706 7352 4712 7364
rect 4764 7352 4770 7404
rect 4890 7392 4896 7404
rect 4851 7364 4896 7392
rect 4890 7352 4896 7364
rect 4948 7352 4954 7404
rect 5442 7352 5448 7404
rect 5500 7392 5506 7404
rect 5994 7392 6000 7404
rect 5500 7364 6000 7392
rect 5500 7352 5506 7364
rect 5994 7352 6000 7364
rect 6052 7352 6058 7404
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7392 7895 7395
rect 7883 7364 8524 7392
rect 7883 7361 7895 7364
rect 7837 7355 7895 7361
rect 3421 7327 3479 7333
rect 3421 7293 3433 7327
rect 3467 7293 3479 7327
rect 5626 7324 5632 7336
rect 3421 7287 3479 7293
rect 4080 7296 5632 7324
rect 4080 7256 4108 7296
rect 5626 7284 5632 7296
rect 5684 7284 5690 7336
rect 5813 7327 5871 7333
rect 5813 7293 5825 7327
rect 5859 7324 5871 7327
rect 6270 7324 6276 7336
rect 5859 7296 6276 7324
rect 5859 7293 5871 7296
rect 5813 7287 5871 7293
rect 6270 7284 6276 7296
rect 6328 7284 6334 7336
rect 6362 7284 6368 7336
rect 6420 7324 6426 7336
rect 7561 7327 7619 7333
rect 7561 7324 7573 7327
rect 6420 7296 7573 7324
rect 6420 7284 6426 7296
rect 7561 7293 7573 7296
rect 7607 7293 7619 7327
rect 7561 7287 7619 7293
rect 8389 7327 8447 7333
rect 8389 7293 8401 7327
rect 8435 7293 8447 7327
rect 8496 7324 8524 7364
rect 9398 7352 9404 7404
rect 9456 7392 9462 7404
rect 11440 7392 11468 7500
rect 13740 7500 14096 7528
rect 12158 7420 12164 7472
rect 12216 7460 12222 7472
rect 12216 7432 13676 7460
rect 12216 7420 12222 7432
rect 13081 7395 13139 7401
rect 9456 7364 10548 7392
rect 11440 7364 12940 7392
rect 9456 7352 9462 7364
rect 9490 7324 9496 7336
rect 8496 7296 9496 7324
rect 8389 7287 8447 7293
rect 1504 7228 4108 7256
rect 4154 7216 4160 7268
rect 4212 7256 4218 7268
rect 7653 7259 7711 7265
rect 7653 7256 7665 7259
rect 4212 7228 7665 7256
rect 4212 7216 4218 7228
rect 7653 7225 7665 7228
rect 7699 7225 7711 7259
rect 7653 7219 7711 7225
rect 3602 7188 3608 7200
rect 3563 7160 3608 7188
rect 3602 7148 3608 7160
rect 3660 7148 3666 7200
rect 4614 7188 4620 7200
rect 4575 7160 4620 7188
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 5718 7148 5724 7200
rect 5776 7188 5782 7200
rect 5905 7191 5963 7197
rect 5905 7188 5917 7191
rect 5776 7160 5917 7188
rect 5776 7148 5782 7160
rect 5905 7157 5917 7160
rect 5951 7157 5963 7191
rect 5905 7151 5963 7157
rect 6362 7148 6368 7200
rect 6420 7188 6426 7200
rect 7282 7188 7288 7200
rect 6420 7160 7288 7188
rect 6420 7148 6426 7160
rect 7282 7148 7288 7160
rect 7340 7148 7346 7200
rect 8404 7188 8432 7287
rect 9490 7284 9496 7296
rect 9548 7284 9554 7336
rect 9674 7284 9680 7336
rect 9732 7324 9738 7336
rect 10042 7324 10048 7336
rect 9732 7296 10048 7324
rect 9732 7284 9738 7296
rect 10042 7284 10048 7296
rect 10100 7324 10106 7336
rect 10413 7327 10471 7333
rect 10413 7324 10425 7327
rect 10100 7296 10425 7324
rect 10100 7284 10106 7296
rect 10413 7293 10425 7296
rect 10459 7293 10471 7327
rect 10520 7324 10548 7364
rect 12158 7324 12164 7336
rect 10520 7296 12164 7324
rect 10413 7287 10471 7293
rect 12158 7284 12164 7296
rect 12216 7284 12222 7336
rect 8570 7216 8576 7268
rect 8628 7265 8634 7268
rect 8628 7259 8692 7265
rect 8628 7225 8646 7259
rect 8680 7225 8692 7259
rect 8628 7219 8692 7225
rect 8628 7216 8634 7219
rect 10594 7216 10600 7268
rect 10652 7265 10658 7268
rect 10652 7259 10716 7265
rect 10652 7225 10670 7259
rect 10704 7225 10716 7259
rect 12805 7259 12863 7265
rect 12805 7256 12817 7259
rect 10652 7219 10716 7225
rect 10796 7228 12817 7256
rect 10652 7216 10658 7219
rect 9674 7188 9680 7200
rect 8404 7160 9680 7188
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 9858 7148 9864 7200
rect 9916 7188 9922 7200
rect 10796 7188 10824 7228
rect 12805 7225 12817 7228
rect 12851 7225 12863 7259
rect 12805 7219 12863 7225
rect 9916 7160 10824 7188
rect 11793 7191 11851 7197
rect 9916 7148 9922 7160
rect 11793 7157 11805 7191
rect 11839 7188 11851 7191
rect 12066 7188 12072 7200
rect 11839 7160 12072 7188
rect 11839 7157 11851 7160
rect 11793 7151 11851 7157
rect 12066 7148 12072 7160
rect 12124 7148 12130 7200
rect 12434 7148 12440 7200
rect 12492 7188 12498 7200
rect 12912 7197 12940 7364
rect 13081 7361 13093 7395
rect 13127 7392 13139 7395
rect 13170 7392 13176 7404
rect 13127 7364 13176 7392
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 13170 7352 13176 7364
rect 13228 7352 13234 7404
rect 13648 7324 13676 7432
rect 13740 7401 13768 7500
rect 14090 7488 14096 7500
rect 14148 7528 14154 7540
rect 15102 7528 15108 7540
rect 14148 7500 14688 7528
rect 15063 7500 15108 7528
rect 14148 7488 14154 7500
rect 14660 7460 14688 7500
rect 15102 7488 15108 7500
rect 15160 7488 15166 7540
rect 15286 7488 15292 7540
rect 15344 7528 15350 7540
rect 18414 7528 18420 7540
rect 15344 7500 18420 7528
rect 15344 7488 15350 7500
rect 18414 7488 18420 7500
rect 18472 7488 18478 7540
rect 14660 7432 15608 7460
rect 15580 7401 15608 7432
rect 13725 7395 13783 7401
rect 13725 7361 13737 7395
rect 13771 7361 13783 7395
rect 13725 7355 13783 7361
rect 15565 7395 15623 7401
rect 15565 7361 15577 7395
rect 15611 7361 15623 7395
rect 15565 7355 15623 7361
rect 16206 7324 16212 7336
rect 13648 7296 16212 7324
rect 16206 7284 16212 7296
rect 16264 7284 16270 7336
rect 13992 7259 14050 7265
rect 13992 7225 14004 7259
rect 14038 7256 14050 7259
rect 15832 7259 15890 7265
rect 14038 7228 15700 7256
rect 14038 7225 14050 7228
rect 13992 7219 14050 7225
rect 12897 7191 12955 7197
rect 12492 7160 12537 7188
rect 12492 7148 12498 7160
rect 12897 7157 12909 7191
rect 12943 7188 12955 7191
rect 13630 7188 13636 7200
rect 12943 7160 13636 7188
rect 12943 7157 12955 7160
rect 12897 7151 12955 7157
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 15672 7188 15700 7228
rect 15832 7225 15844 7259
rect 15878 7256 15890 7259
rect 16574 7256 16580 7268
rect 15878 7228 16580 7256
rect 15878 7225 15890 7228
rect 15832 7219 15890 7225
rect 16574 7216 16580 7228
rect 16632 7216 16638 7268
rect 16206 7188 16212 7200
rect 15672 7160 16212 7188
rect 16206 7148 16212 7160
rect 16264 7188 16270 7200
rect 16945 7191 17003 7197
rect 16945 7188 16957 7191
rect 16264 7160 16957 7188
rect 16264 7148 16270 7160
rect 16945 7157 16957 7160
rect 16991 7157 17003 7191
rect 16945 7151 17003 7157
rect 1104 7098 18860 7120
rect 1104 7046 6912 7098
rect 6964 7046 6976 7098
rect 7028 7046 7040 7098
rect 7092 7046 7104 7098
rect 7156 7046 12843 7098
rect 12895 7046 12907 7098
rect 12959 7046 12971 7098
rect 13023 7046 13035 7098
rect 13087 7046 18860 7098
rect 1104 7024 18860 7046
rect 1581 6987 1639 6993
rect 1581 6953 1593 6987
rect 1627 6984 1639 6987
rect 1762 6984 1768 6996
rect 1627 6956 1768 6984
rect 1627 6953 1639 6956
rect 1581 6947 1639 6953
rect 1762 6944 1768 6956
rect 1820 6944 1826 6996
rect 1949 6987 2007 6993
rect 1949 6953 1961 6987
rect 1995 6984 2007 6987
rect 5442 6984 5448 6996
rect 1995 6956 5304 6984
rect 5403 6956 5448 6984
rect 1995 6953 2007 6956
rect 1949 6947 2007 6953
rect 3050 6876 3056 6928
rect 3108 6916 3114 6928
rect 3145 6919 3203 6925
rect 3145 6916 3157 6919
rect 3108 6888 3157 6916
rect 3108 6876 3114 6888
rect 3145 6885 3157 6888
rect 3191 6885 3203 6919
rect 3145 6879 3203 6885
rect 3237 6919 3295 6925
rect 3237 6885 3249 6919
rect 3283 6916 3295 6919
rect 5276 6916 5304 6956
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 7469 6987 7527 6993
rect 5552 6956 6500 6984
rect 5552 6916 5580 6956
rect 3283 6888 5212 6916
rect 5276 6888 5580 6916
rect 6472 6916 6500 6956
rect 7469 6953 7481 6987
rect 7515 6984 7527 6987
rect 7650 6984 7656 6996
rect 7515 6956 7656 6984
rect 7515 6953 7527 6956
rect 7469 6947 7527 6953
rect 7650 6944 7656 6956
rect 7708 6944 7714 6996
rect 8294 6984 8300 6996
rect 8255 6956 8300 6984
rect 8294 6944 8300 6956
rect 8352 6944 8358 6996
rect 8478 6944 8484 6996
rect 8536 6984 8542 6996
rect 8665 6987 8723 6993
rect 8665 6984 8677 6987
rect 8536 6956 8677 6984
rect 8536 6944 8542 6956
rect 8665 6953 8677 6956
rect 8711 6953 8723 6987
rect 8665 6947 8723 6953
rect 9398 6944 9404 6996
rect 9456 6984 9462 6996
rect 10689 6987 10747 6993
rect 10689 6984 10701 6987
rect 9456 6956 10701 6984
rect 9456 6944 9462 6956
rect 10689 6953 10701 6956
rect 10735 6953 10747 6987
rect 11054 6984 11060 6996
rect 10689 6947 10747 6953
rect 10796 6956 11060 6984
rect 9122 6916 9128 6928
rect 6472 6888 9128 6916
rect 3283 6885 3295 6888
rect 3237 6879 3295 6885
rect 2958 6808 2964 6860
rect 3016 6848 3022 6860
rect 3252 6848 3280 6879
rect 3016 6820 3280 6848
rect 3016 6808 3022 6820
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 3476 6820 3740 6848
rect 3476 6808 3482 6820
rect 1670 6740 1676 6792
rect 1728 6780 1734 6792
rect 2041 6783 2099 6789
rect 2041 6780 2053 6783
rect 1728 6752 2053 6780
rect 1728 6740 1734 6752
rect 2041 6749 2053 6752
rect 2087 6749 2099 6783
rect 2222 6780 2228 6792
rect 2183 6752 2228 6780
rect 2041 6743 2099 6749
rect 2222 6740 2228 6752
rect 2280 6740 2286 6792
rect 3326 6740 3332 6792
rect 3384 6780 3390 6792
rect 3712 6780 3740 6820
rect 3786 6808 3792 6860
rect 3844 6848 3850 6860
rect 4321 6851 4379 6857
rect 4321 6848 4333 6851
rect 3844 6820 4333 6848
rect 3844 6808 3850 6820
rect 4321 6817 4333 6820
rect 4367 6817 4379 6851
rect 5184 6848 5212 6888
rect 9122 6876 9128 6888
rect 9180 6876 9186 6928
rect 9677 6919 9735 6925
rect 9677 6885 9689 6919
rect 9723 6916 9735 6919
rect 9858 6916 9864 6928
rect 9723 6888 9864 6916
rect 9723 6885 9735 6888
rect 9677 6879 9735 6885
rect 9858 6876 9864 6888
rect 9916 6876 9922 6928
rect 9950 6876 9956 6928
rect 10008 6916 10014 6928
rect 10796 6916 10824 6956
rect 11054 6944 11060 6956
rect 11112 6944 11118 6996
rect 12342 6944 12348 6996
rect 12400 6984 12406 6996
rect 13354 6984 13360 6996
rect 12400 6956 13360 6984
rect 12400 6944 12406 6956
rect 13354 6944 13360 6956
rect 13412 6944 13418 6996
rect 14366 6984 14372 6996
rect 14327 6956 14372 6984
rect 14366 6944 14372 6956
rect 14424 6944 14430 6996
rect 15289 6987 15347 6993
rect 15289 6953 15301 6987
rect 15335 6953 15347 6987
rect 15289 6947 15347 6953
rect 15304 6916 15332 6947
rect 15654 6944 15660 6996
rect 15712 6984 15718 6996
rect 17037 6987 17095 6993
rect 17037 6984 17049 6987
rect 15712 6956 17049 6984
rect 15712 6944 15718 6956
rect 17037 6953 17049 6956
rect 17083 6953 17095 6987
rect 17037 6947 17095 6953
rect 10008 6888 10824 6916
rect 10980 6888 15332 6916
rect 15396 6888 15792 6916
rect 10008 6876 10014 6888
rect 6270 6848 6276 6860
rect 5184 6820 6031 6848
rect 6231 6820 6276 6848
rect 4321 6811 4379 6817
rect 4065 6783 4123 6789
rect 4065 6780 4077 6783
rect 3384 6752 3429 6780
rect 3712 6752 4077 6780
rect 3384 6740 3390 6752
rect 4065 6749 4077 6752
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 2777 6715 2835 6721
rect 2777 6681 2789 6715
rect 2823 6712 2835 6715
rect 3970 6712 3976 6724
rect 2823 6684 3976 6712
rect 2823 6681 2835 6684
rect 2777 6675 2835 6681
rect 3970 6672 3976 6684
rect 4028 6672 4034 6724
rect 5905 6715 5963 6721
rect 5905 6712 5917 6715
rect 5000 6684 5917 6712
rect 2682 6604 2688 6656
rect 2740 6644 2746 6656
rect 5000 6644 5028 6684
rect 5905 6681 5917 6684
rect 5951 6681 5963 6715
rect 5905 6675 5963 6681
rect 2740 6616 5028 6644
rect 6003 6644 6031 6820
rect 6270 6808 6276 6820
rect 6328 6808 6334 6860
rect 10134 6808 10140 6860
rect 10192 6848 10198 6860
rect 10781 6851 10839 6857
rect 10781 6848 10793 6851
rect 10192 6820 10793 6848
rect 10192 6808 10198 6820
rect 10781 6817 10793 6820
rect 10827 6817 10839 6851
rect 10781 6811 10839 6817
rect 6365 6783 6423 6789
rect 6365 6749 6377 6783
rect 6411 6749 6423 6783
rect 6546 6780 6552 6792
rect 6507 6752 6552 6780
rect 6365 6743 6423 6749
rect 6380 6712 6408 6743
rect 6546 6740 6552 6752
rect 6604 6740 6610 6792
rect 7561 6783 7619 6789
rect 7561 6749 7573 6783
rect 7607 6749 7619 6783
rect 7561 6743 7619 6749
rect 7101 6715 7159 6721
rect 7101 6712 7113 6715
rect 6380 6684 7113 6712
rect 7101 6681 7113 6684
rect 7147 6681 7159 6715
rect 7101 6675 7159 6681
rect 7466 6672 7472 6724
rect 7524 6712 7530 6724
rect 7576 6712 7604 6743
rect 7650 6740 7656 6792
rect 7708 6780 7714 6792
rect 7708 6752 7753 6780
rect 7708 6740 7714 6752
rect 8110 6740 8116 6792
rect 8168 6780 8174 6792
rect 8757 6783 8815 6789
rect 8757 6780 8769 6783
rect 8168 6752 8769 6780
rect 8168 6740 8174 6752
rect 8757 6749 8769 6752
rect 8803 6749 8815 6783
rect 8757 6743 8815 6749
rect 8941 6783 8999 6789
rect 8941 6749 8953 6783
rect 8987 6780 8999 6783
rect 9490 6780 9496 6792
rect 8987 6752 9496 6780
rect 8987 6749 8999 6752
rect 8941 6743 8999 6749
rect 9490 6740 9496 6752
rect 9548 6740 9554 6792
rect 10594 6780 10600 6792
rect 9876 6752 10600 6780
rect 7524 6684 7604 6712
rect 7524 6672 7530 6684
rect 8202 6672 8208 6724
rect 8260 6712 8266 6724
rect 9876 6712 9904 6752
rect 10594 6740 10600 6752
rect 10652 6740 10658 6792
rect 10870 6780 10876 6792
rect 10831 6752 10876 6780
rect 10870 6740 10876 6752
rect 10928 6740 10934 6792
rect 8260 6684 9904 6712
rect 8260 6672 8266 6684
rect 9950 6672 9956 6724
rect 10008 6672 10014 6724
rect 10042 6672 10048 6724
rect 10100 6672 10106 6724
rect 10318 6712 10324 6724
rect 10279 6684 10324 6712
rect 10318 6672 10324 6684
rect 10376 6672 10382 6724
rect 10686 6672 10692 6724
rect 10744 6712 10750 6724
rect 10980 6712 11008 6888
rect 11784 6851 11842 6857
rect 11784 6817 11796 6851
rect 11830 6848 11842 6851
rect 12066 6848 12072 6860
rect 11830 6820 12072 6848
rect 11830 6817 11842 6820
rect 11784 6811 11842 6817
rect 12066 6808 12072 6820
rect 12124 6808 12130 6860
rect 13357 6851 13415 6857
rect 13357 6817 13369 6851
rect 13403 6848 13415 6851
rect 13814 6848 13820 6860
rect 13403 6820 13820 6848
rect 13403 6817 13415 6820
rect 13357 6811 13415 6817
rect 13814 6808 13820 6820
rect 13872 6808 13878 6860
rect 15396 6848 15424 6888
rect 15654 6848 15660 6860
rect 13924 6820 15424 6848
rect 15615 6820 15660 6848
rect 11517 6783 11575 6789
rect 11517 6780 11529 6783
rect 10744 6684 11008 6712
rect 11072 6752 11529 6780
rect 10744 6672 10750 6684
rect 9968 6644 9996 6672
rect 6003 6616 9996 6644
rect 10060 6644 10088 6672
rect 11072 6644 11100 6752
rect 11517 6749 11529 6752
rect 11563 6749 11575 6783
rect 11517 6743 11575 6749
rect 13170 6740 13176 6792
rect 13228 6780 13234 6792
rect 13924 6780 13952 6820
rect 15654 6808 15660 6820
rect 15712 6808 15718 6860
rect 15764 6848 15792 6888
rect 16850 6876 16856 6928
rect 16908 6916 16914 6928
rect 17129 6919 17187 6925
rect 17129 6916 17141 6919
rect 16908 6888 17141 6916
rect 16908 6876 16914 6888
rect 17129 6885 17141 6888
rect 17175 6885 17187 6919
rect 17129 6879 17187 6885
rect 17865 6851 17923 6857
rect 17865 6848 17877 6851
rect 15764 6820 17877 6848
rect 17865 6817 17877 6820
rect 17911 6817 17923 6851
rect 17865 6811 17923 6817
rect 13228 6752 13952 6780
rect 13228 6740 13234 6752
rect 14090 6740 14096 6792
rect 14148 6780 14154 6792
rect 14461 6783 14519 6789
rect 14461 6780 14473 6783
rect 14148 6752 14473 6780
rect 14148 6740 14154 6752
rect 14461 6749 14473 6752
rect 14507 6749 14519 6783
rect 14461 6743 14519 6749
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6749 14611 6783
rect 14553 6743 14611 6749
rect 10060 6616 11100 6644
rect 2740 6604 2746 6616
rect 12158 6604 12164 6656
rect 12216 6644 12222 6656
rect 12897 6647 12955 6653
rect 12897 6644 12909 6647
rect 12216 6616 12909 6644
rect 12216 6604 12222 6616
rect 12897 6613 12909 6616
rect 12943 6644 12955 6647
rect 13354 6644 13360 6656
rect 12943 6616 13360 6644
rect 12943 6613 12955 6616
rect 12897 6607 12955 6613
rect 13354 6604 13360 6616
rect 13412 6604 13418 6656
rect 13998 6644 14004 6656
rect 13959 6616 14004 6644
rect 13998 6604 14004 6616
rect 14056 6604 14062 6656
rect 14366 6604 14372 6656
rect 14424 6644 14430 6656
rect 14568 6644 14596 6743
rect 15470 6740 15476 6792
rect 15528 6780 15534 6792
rect 15749 6783 15807 6789
rect 15749 6780 15761 6783
rect 15528 6752 15761 6780
rect 15528 6740 15534 6752
rect 15749 6749 15761 6752
rect 15795 6749 15807 6783
rect 15749 6743 15807 6749
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 15102 6672 15108 6724
rect 15160 6712 15166 6724
rect 15856 6712 15884 6743
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 17276 6752 17321 6780
rect 17276 6740 17282 6752
rect 16666 6712 16672 6724
rect 15160 6684 15884 6712
rect 16627 6684 16672 6712
rect 15160 6672 15166 6684
rect 16666 6672 16672 6684
rect 16724 6672 16730 6724
rect 18046 6644 18052 6656
rect 14424 6616 14596 6644
rect 18007 6616 18052 6644
rect 14424 6604 14430 6616
rect 18046 6604 18052 6616
rect 18104 6604 18110 6656
rect 1104 6554 18860 6576
rect 1104 6502 3947 6554
rect 3999 6502 4011 6554
rect 4063 6502 4075 6554
rect 4127 6502 4139 6554
rect 4191 6502 9878 6554
rect 9930 6502 9942 6554
rect 9994 6502 10006 6554
rect 10058 6502 10070 6554
rect 10122 6502 15808 6554
rect 15860 6502 15872 6554
rect 15924 6502 15936 6554
rect 15988 6502 16000 6554
rect 16052 6502 18860 6554
rect 1104 6480 18860 6502
rect 2222 6400 2228 6452
rect 2280 6440 2286 6452
rect 2774 6440 2780 6452
rect 2280 6412 2780 6440
rect 2280 6400 2286 6412
rect 2774 6400 2780 6412
rect 2832 6400 2838 6452
rect 3786 6440 3792 6452
rect 3747 6412 3792 6440
rect 3786 6400 3792 6412
rect 3844 6400 3850 6452
rect 6270 6400 6276 6452
rect 6328 6440 6334 6452
rect 6825 6443 6883 6449
rect 6825 6440 6837 6443
rect 6328 6412 6837 6440
rect 6328 6400 6334 6412
rect 6825 6409 6837 6412
rect 6871 6409 6883 6443
rect 8110 6440 8116 6452
rect 8071 6412 8116 6440
rect 6825 6403 6883 6409
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 9674 6440 9680 6452
rect 9324 6412 9680 6440
rect 1854 6372 1860 6384
rect 1815 6344 1860 6372
rect 1854 6332 1860 6344
rect 1912 6332 1918 6384
rect 5534 6332 5540 6384
rect 5592 6372 5598 6384
rect 8478 6372 8484 6384
rect 5592 6344 8484 6372
rect 5592 6332 5598 6344
rect 8478 6332 8484 6344
rect 8536 6332 8542 6384
rect 8570 6332 8576 6384
rect 8628 6372 8634 6384
rect 8628 6344 8708 6372
rect 8628 6332 8634 6344
rect 6270 6264 6276 6316
rect 6328 6304 6334 6316
rect 7469 6307 7527 6313
rect 7469 6304 7481 6307
rect 6328 6276 7481 6304
rect 6328 6264 6334 6276
rect 7469 6273 7481 6276
rect 7515 6304 7527 6307
rect 7650 6304 7656 6316
rect 7515 6276 7656 6304
rect 7515 6273 7527 6276
rect 7469 6267 7527 6273
rect 7650 6264 7656 6276
rect 7708 6264 7714 6316
rect 7742 6264 7748 6316
rect 7800 6264 7806 6316
rect 8680 6313 8708 6344
rect 9324 6313 9352 6412
rect 9674 6400 9680 6412
rect 9732 6400 9738 6452
rect 10318 6400 10324 6452
rect 10376 6440 10382 6452
rect 11606 6440 11612 6452
rect 10376 6412 11612 6440
rect 10376 6400 10382 6412
rect 11606 6400 11612 6412
rect 11664 6400 11670 6452
rect 11716 6412 15240 6440
rect 10594 6332 10600 6384
rect 10652 6372 10658 6384
rect 11716 6372 11744 6412
rect 12158 6372 12164 6384
rect 10652 6344 11744 6372
rect 11808 6344 12164 6372
rect 10652 6332 10658 6344
rect 8665 6307 8723 6313
rect 8665 6273 8677 6307
rect 8711 6273 8723 6307
rect 8665 6267 8723 6273
rect 9309 6307 9367 6313
rect 9309 6273 9321 6307
rect 9355 6273 9367 6307
rect 9309 6267 9367 6273
rect 11609 6307 11667 6313
rect 11609 6273 11621 6307
rect 11655 6304 11667 6307
rect 11698 6304 11704 6316
rect 11655 6276 11704 6304
rect 11655 6273 11667 6276
rect 11609 6267 11667 6273
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 11808 6313 11836 6344
rect 12158 6332 12164 6344
rect 12216 6332 12222 6384
rect 11793 6307 11851 6313
rect 11793 6273 11805 6307
rect 11839 6273 11851 6307
rect 11793 6267 11851 6273
rect 12710 6264 12716 6316
rect 12768 6304 12774 6316
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 12768 6276 12909 6304
rect 12768 6264 12774 6276
rect 12897 6273 12909 6276
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 12989 6307 13047 6313
rect 12989 6273 13001 6307
rect 13035 6273 13047 6307
rect 12989 6267 13047 6273
rect 1670 6236 1676 6248
rect 1631 6208 1676 6236
rect 1670 6196 1676 6208
rect 1728 6196 1734 6248
rect 2409 6239 2467 6245
rect 2409 6205 2421 6239
rect 2455 6205 2467 6239
rect 4430 6236 4436 6248
rect 4391 6208 4436 6236
rect 2409 6199 2467 6205
rect 2424 6100 2452 6199
rect 4430 6196 4436 6208
rect 4488 6196 4494 6248
rect 4706 6245 4712 6248
rect 4700 6236 4712 6245
rect 4619 6208 4712 6236
rect 4700 6199 4712 6208
rect 4764 6236 4770 6248
rect 6288 6236 6316 6264
rect 6454 6236 6460 6248
rect 4764 6208 6316 6236
rect 6415 6208 6460 6236
rect 4706 6196 4712 6199
rect 4764 6196 4770 6208
rect 6454 6196 6460 6208
rect 6512 6196 6518 6248
rect 7285 6239 7343 6245
rect 7285 6205 7297 6239
rect 7331 6236 7343 6239
rect 7760 6236 7788 6264
rect 7331 6208 7788 6236
rect 7331 6205 7343 6208
rect 7285 6199 7343 6205
rect 8386 6196 8392 6248
rect 8444 6236 8450 6248
rect 8481 6239 8539 6245
rect 8481 6236 8493 6239
rect 8444 6208 8493 6236
rect 8444 6196 8450 6208
rect 8481 6205 8493 6208
rect 8527 6205 8539 6239
rect 8481 6199 8539 6205
rect 8573 6239 8631 6245
rect 8573 6205 8585 6239
rect 8619 6236 8631 6239
rect 8754 6236 8760 6248
rect 8619 6208 8760 6236
rect 8619 6205 8631 6208
rect 8573 6199 8631 6205
rect 8754 6196 8760 6208
rect 8812 6196 8818 6248
rect 9576 6239 9634 6245
rect 9576 6205 9588 6239
rect 9622 6236 9634 6239
rect 10410 6236 10416 6248
rect 9622 6208 10416 6236
rect 9622 6205 9634 6208
rect 9576 6199 9634 6205
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 10594 6196 10600 6248
rect 10652 6236 10658 6248
rect 10778 6236 10784 6248
rect 10652 6208 10784 6236
rect 10652 6196 10658 6208
rect 10778 6196 10784 6208
rect 10836 6196 10842 6248
rect 12434 6196 12440 6248
rect 12492 6236 12498 6248
rect 12805 6239 12863 6245
rect 12805 6236 12817 6239
rect 12492 6208 12817 6236
rect 12492 6196 12498 6208
rect 12805 6205 12817 6208
rect 12851 6205 12863 6239
rect 12805 6199 12863 6205
rect 2676 6171 2734 6177
rect 2676 6137 2688 6171
rect 2722 6168 2734 6171
rect 4614 6168 4620 6180
rect 2722 6140 4620 6168
rect 2722 6137 2734 6140
rect 2676 6131 2734 6137
rect 4614 6128 4620 6140
rect 4672 6168 4678 6180
rect 6546 6168 6552 6180
rect 4672 6140 6552 6168
rect 4672 6128 4678 6140
rect 3418 6100 3424 6112
rect 2424 6072 3424 6100
rect 3418 6060 3424 6072
rect 3476 6100 3482 6112
rect 4430 6100 4436 6112
rect 3476 6072 4436 6100
rect 3476 6060 3482 6072
rect 4430 6060 4436 6072
rect 4488 6060 4494 6112
rect 5828 6109 5856 6140
rect 6546 6128 6552 6140
rect 6604 6128 6610 6180
rect 7193 6171 7251 6177
rect 7193 6137 7205 6171
rect 7239 6168 7251 6171
rect 7742 6168 7748 6180
rect 7239 6140 7748 6168
rect 7239 6137 7251 6140
rect 7193 6131 7251 6137
rect 7742 6128 7748 6140
rect 7800 6128 7806 6180
rect 8294 6128 8300 6180
rect 8352 6168 8358 6180
rect 11517 6171 11575 6177
rect 8352 6140 11192 6168
rect 8352 6128 8358 6140
rect 5813 6103 5871 6109
rect 5813 6069 5825 6103
rect 5859 6069 5871 6103
rect 5813 6063 5871 6069
rect 5994 6060 6000 6112
rect 6052 6100 6058 6112
rect 6273 6103 6331 6109
rect 6273 6100 6285 6103
rect 6052 6072 6285 6100
rect 6052 6060 6058 6072
rect 6273 6069 6285 6072
rect 6319 6069 6331 6103
rect 6273 6063 6331 6069
rect 7374 6060 7380 6112
rect 7432 6100 7438 6112
rect 11164 6109 11192 6140
rect 11517 6137 11529 6171
rect 11563 6168 11575 6171
rect 11563 6140 12020 6168
rect 11563 6137 11575 6140
rect 11517 6131 11575 6137
rect 10689 6103 10747 6109
rect 10689 6100 10701 6103
rect 7432 6072 10701 6100
rect 7432 6060 7438 6072
rect 10689 6069 10701 6072
rect 10735 6069 10747 6103
rect 10689 6063 10747 6069
rect 11149 6103 11207 6109
rect 11149 6069 11161 6103
rect 11195 6069 11207 6103
rect 11992 6100 12020 6140
rect 12066 6128 12072 6180
rect 12124 6168 12130 6180
rect 13004 6168 13032 6267
rect 14182 6236 14188 6248
rect 14143 6208 14188 6236
rect 14182 6196 14188 6208
rect 14240 6196 14246 6248
rect 15212 6236 15240 6412
rect 15654 6400 15660 6452
rect 15712 6440 15718 6452
rect 16025 6443 16083 6449
rect 16025 6440 16037 6443
rect 15712 6412 16037 6440
rect 15712 6400 15718 6412
rect 16025 6409 16037 6412
rect 16071 6409 16083 6443
rect 16025 6403 16083 6409
rect 16574 6400 16580 6452
rect 16632 6440 16638 6452
rect 17218 6440 17224 6452
rect 16632 6412 17224 6440
rect 16632 6400 16638 6412
rect 17218 6400 17224 6412
rect 17276 6400 17282 6452
rect 15746 6332 15752 6384
rect 15804 6372 15810 6384
rect 18322 6372 18328 6384
rect 15804 6344 18328 6372
rect 15804 6332 15810 6344
rect 18322 6332 18328 6344
rect 18380 6332 18386 6384
rect 16206 6264 16212 6316
rect 16264 6304 16270 6316
rect 16577 6307 16635 6313
rect 16577 6304 16589 6307
rect 16264 6276 16589 6304
rect 16264 6264 16270 6276
rect 16577 6273 16589 6276
rect 16623 6273 16635 6307
rect 16577 6267 16635 6273
rect 17221 6239 17279 6245
rect 17221 6236 17233 6239
rect 15212 6208 17233 6236
rect 17221 6205 17233 6208
rect 17267 6205 17279 6239
rect 17221 6199 17279 6205
rect 12124 6140 13032 6168
rect 12124 6128 12130 6140
rect 14366 6128 14372 6180
rect 14424 6177 14430 6180
rect 14424 6171 14488 6177
rect 14424 6137 14442 6171
rect 14476 6137 14488 6171
rect 16390 6168 16396 6180
rect 16351 6140 16396 6168
rect 14424 6131 14488 6137
rect 14424 6128 14430 6131
rect 16390 6128 16396 6140
rect 16448 6128 16454 6180
rect 12437 6103 12495 6109
rect 12437 6100 12449 6103
rect 11992 6072 12449 6100
rect 11149 6063 11207 6069
rect 12437 6069 12449 6072
rect 12483 6069 12495 6103
rect 12437 6063 12495 6069
rect 15565 6103 15623 6109
rect 15565 6069 15577 6103
rect 15611 6100 15623 6103
rect 15654 6100 15660 6112
rect 15611 6072 15660 6100
rect 15611 6069 15623 6072
rect 15565 6063 15623 6069
rect 15654 6060 15660 6072
rect 15712 6060 15718 6112
rect 16485 6103 16543 6109
rect 16485 6069 16497 6103
rect 16531 6100 16543 6103
rect 16666 6100 16672 6112
rect 16531 6072 16672 6100
rect 16531 6069 16543 6072
rect 16485 6063 16543 6069
rect 16666 6060 16672 6072
rect 16724 6060 16730 6112
rect 17402 6100 17408 6112
rect 17363 6072 17408 6100
rect 17402 6060 17408 6072
rect 17460 6060 17466 6112
rect 17586 6060 17592 6112
rect 17644 6100 17650 6112
rect 17770 6100 17776 6112
rect 17644 6072 17776 6100
rect 17644 6060 17650 6072
rect 17770 6060 17776 6072
rect 17828 6060 17834 6112
rect 1104 6010 18860 6032
rect 1104 5958 6912 6010
rect 6964 5958 6976 6010
rect 7028 5958 7040 6010
rect 7092 5958 7104 6010
rect 7156 5958 12843 6010
rect 12895 5958 12907 6010
rect 12959 5958 12971 6010
rect 13023 5958 13035 6010
rect 13087 5958 18860 6010
rect 1104 5936 18860 5958
rect 2682 5856 2688 5908
rect 2740 5896 2746 5908
rect 3145 5899 3203 5905
rect 3145 5896 3157 5899
rect 2740 5868 3157 5896
rect 2740 5856 2746 5868
rect 3145 5865 3157 5868
rect 3191 5865 3203 5899
rect 3145 5859 3203 5865
rect 3237 5899 3295 5905
rect 3237 5865 3249 5899
rect 3283 5896 3295 5899
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 3283 5868 4077 5896
rect 3283 5865 3295 5868
rect 3237 5859 3295 5865
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 8570 5896 8576 5908
rect 4065 5859 4123 5865
rect 6472 5868 8576 5896
rect 2774 5788 2780 5840
rect 2832 5828 2838 5840
rect 3326 5828 3332 5840
rect 2832 5800 3332 5828
rect 2832 5788 2838 5800
rect 3326 5788 3332 5800
rect 3384 5828 3390 5840
rect 6472 5828 6500 5868
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 8846 5896 8852 5908
rect 8759 5868 8852 5896
rect 8846 5856 8852 5868
rect 8904 5896 8910 5908
rect 8904 5868 11744 5896
rect 8904 5856 8910 5868
rect 3384 5800 6500 5828
rect 6540 5831 6598 5837
rect 3384 5788 3390 5800
rect 6540 5797 6552 5831
rect 6586 5828 6598 5831
rect 7374 5828 7380 5840
rect 6586 5800 7380 5828
rect 6586 5797 6598 5800
rect 6540 5791 6598 5797
rect 7374 5788 7380 5800
rect 7432 5788 7438 5840
rect 10686 5828 10692 5840
rect 7484 5800 10692 5828
rect 1765 5763 1823 5769
rect 1765 5729 1777 5763
rect 1811 5760 1823 5763
rect 4430 5760 4436 5772
rect 1811 5732 2820 5760
rect 4391 5732 4436 5760
rect 1811 5729 1823 5732
rect 1765 5723 1823 5729
rect 1946 5692 1952 5704
rect 1907 5664 1952 5692
rect 1946 5652 1952 5664
rect 2004 5652 2010 5704
rect 2792 5633 2820 5732
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 5534 5760 5540 5772
rect 5495 5732 5540 5760
rect 5534 5720 5540 5732
rect 5592 5720 5598 5772
rect 5994 5760 6000 5772
rect 5828 5732 6000 5760
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5692 3479 5695
rect 3786 5692 3792 5704
rect 3467 5664 3792 5692
rect 3467 5661 3479 5664
rect 3421 5655 3479 5661
rect 3786 5652 3792 5664
rect 3844 5652 3850 5704
rect 4338 5652 4344 5704
rect 4396 5692 4402 5704
rect 4525 5695 4583 5701
rect 4525 5692 4537 5695
rect 4396 5664 4537 5692
rect 4396 5652 4402 5664
rect 4525 5661 4537 5664
rect 4571 5661 4583 5695
rect 4525 5655 4583 5661
rect 4614 5652 4620 5704
rect 4672 5692 4678 5704
rect 4672 5664 4717 5692
rect 4672 5652 4678 5664
rect 4890 5652 4896 5704
rect 4948 5692 4954 5704
rect 5350 5692 5356 5704
rect 4948 5664 5356 5692
rect 4948 5652 4954 5664
rect 5350 5652 5356 5664
rect 5408 5692 5414 5704
rect 5828 5692 5856 5732
rect 5994 5720 6000 5732
rect 6052 5760 6058 5772
rect 6273 5763 6331 5769
rect 6273 5760 6285 5763
rect 6052 5732 6285 5760
rect 6052 5720 6058 5732
rect 6273 5729 6285 5732
rect 6319 5729 6331 5763
rect 7484 5760 7512 5800
rect 10686 5788 10692 5800
rect 10744 5788 10750 5840
rect 11330 5788 11336 5840
rect 11388 5828 11394 5840
rect 11716 5837 11744 5868
rect 12066 5856 12072 5908
rect 12124 5896 12130 5908
rect 12124 5868 13952 5896
rect 12124 5856 12130 5868
rect 11609 5831 11667 5837
rect 11609 5828 11621 5831
rect 11388 5800 11621 5828
rect 11388 5788 11394 5800
rect 11609 5797 11621 5800
rect 11655 5797 11667 5831
rect 11609 5791 11667 5797
rect 11701 5831 11759 5837
rect 11701 5797 11713 5831
rect 11747 5828 11759 5831
rect 11974 5828 11980 5840
rect 11747 5800 11980 5828
rect 11747 5797 11759 5800
rect 11701 5791 11759 5797
rect 11974 5788 11980 5800
rect 12032 5788 12038 5840
rect 12621 5831 12679 5837
rect 12621 5797 12633 5831
rect 12667 5828 12679 5831
rect 13170 5828 13176 5840
rect 12667 5800 13176 5828
rect 12667 5797 12679 5800
rect 12621 5791 12679 5797
rect 13170 5788 13176 5800
rect 13228 5788 13234 5840
rect 13354 5837 13360 5840
rect 13348 5791 13360 5837
rect 13412 5828 13418 5840
rect 13924 5828 13952 5868
rect 13998 5856 14004 5908
rect 14056 5896 14062 5908
rect 17865 5899 17923 5905
rect 17865 5896 17877 5899
rect 14056 5868 17877 5896
rect 14056 5856 14062 5868
rect 17865 5865 17877 5868
rect 17911 5865 17923 5899
rect 17865 5859 17923 5865
rect 16574 5828 16580 5840
rect 13412 5800 13448 5828
rect 13924 5800 16580 5828
rect 13354 5788 13360 5791
rect 13412 5788 13418 5800
rect 16574 5788 16580 5800
rect 16632 5788 16638 5840
rect 6273 5723 6331 5729
rect 6380 5732 7512 5760
rect 8757 5763 8815 5769
rect 6380 5692 6408 5732
rect 8757 5729 8769 5763
rect 8803 5760 8815 5763
rect 9490 5760 9496 5772
rect 8803 5732 9496 5760
rect 8803 5729 8815 5732
rect 8757 5723 8815 5729
rect 9490 5720 9496 5732
rect 9548 5760 9554 5772
rect 9933 5763 9991 5769
rect 9933 5760 9945 5763
rect 9548 5732 9945 5760
rect 9548 5720 9554 5732
rect 9933 5729 9945 5732
rect 9979 5729 9991 5763
rect 9933 5723 9991 5729
rect 10318 5720 10324 5772
rect 10376 5760 10382 5772
rect 14182 5760 14188 5772
rect 10376 5732 10732 5760
rect 10376 5720 10382 5732
rect 10704 5704 10732 5732
rect 13096 5732 14188 5760
rect 5408 5664 5856 5692
rect 6288 5664 6408 5692
rect 8389 5695 8447 5701
rect 5408 5652 5414 5664
rect 2777 5627 2835 5633
rect 2777 5593 2789 5627
rect 2823 5593 2835 5627
rect 6288 5624 6316 5664
rect 8389 5661 8401 5695
rect 8435 5692 8447 5695
rect 9030 5692 9036 5704
rect 8435 5664 9036 5692
rect 8435 5661 8447 5664
rect 8389 5655 8447 5661
rect 9030 5652 9036 5664
rect 9088 5652 9094 5704
rect 9674 5692 9680 5704
rect 9635 5664 9680 5692
rect 9674 5652 9680 5664
rect 9732 5652 9738 5704
rect 10686 5652 10692 5704
rect 10744 5652 10750 5704
rect 11974 5652 11980 5704
rect 12032 5692 12038 5704
rect 13096 5701 13124 5732
rect 14182 5720 14188 5732
rect 14240 5720 14246 5772
rect 14734 5720 14740 5772
rect 14792 5760 14798 5772
rect 15473 5763 15531 5769
rect 15473 5760 15485 5763
rect 14792 5732 15485 5760
rect 14792 5720 14798 5732
rect 15473 5729 15485 5732
rect 15519 5729 15531 5763
rect 15473 5723 15531 5729
rect 13081 5695 13139 5701
rect 13081 5692 13093 5695
rect 12032 5664 13093 5692
rect 12032 5652 12038 5664
rect 13081 5661 13093 5664
rect 13127 5661 13139 5695
rect 15488 5692 15516 5723
rect 15654 5720 15660 5772
rect 15712 5760 15718 5772
rect 16669 5763 16727 5769
rect 15712 5732 16528 5760
rect 15712 5720 15718 5732
rect 15746 5692 15752 5704
rect 15488 5664 15752 5692
rect 13081 5655 13139 5661
rect 15746 5652 15752 5664
rect 15804 5652 15810 5704
rect 16206 5652 16212 5704
rect 16264 5692 16270 5704
rect 16390 5692 16396 5704
rect 16264 5664 16396 5692
rect 16264 5652 16270 5664
rect 16390 5652 16396 5664
rect 16448 5652 16454 5704
rect 16500 5692 16528 5732
rect 16669 5729 16681 5763
rect 16715 5760 16727 5763
rect 16850 5760 16856 5772
rect 16715 5732 16856 5760
rect 16715 5729 16727 5732
rect 16669 5723 16727 5729
rect 16850 5720 16856 5732
rect 16908 5720 16914 5772
rect 17770 5760 17776 5772
rect 17731 5732 17776 5760
rect 17770 5720 17776 5732
rect 17828 5720 17834 5772
rect 16761 5695 16819 5701
rect 16761 5692 16773 5695
rect 16500 5664 16773 5692
rect 16761 5661 16773 5664
rect 16807 5692 16819 5695
rect 17218 5692 17224 5704
rect 16807 5664 17224 5692
rect 16807 5661 16819 5664
rect 16761 5655 16819 5661
rect 17218 5652 17224 5664
rect 17276 5692 17282 5704
rect 17957 5695 18015 5701
rect 17957 5692 17969 5695
rect 17276 5664 17969 5692
rect 17276 5652 17282 5664
rect 17957 5661 17969 5664
rect 18003 5661 18015 5695
rect 17957 5655 18015 5661
rect 8110 5624 8116 5636
rect 2777 5587 2835 5593
rect 5644 5596 6316 5624
rect 7484 5596 8116 5624
rect 3418 5516 3424 5568
rect 3476 5556 3482 5568
rect 5644 5556 5672 5596
rect 3476 5528 5672 5556
rect 5721 5559 5779 5565
rect 3476 5516 3482 5528
rect 5721 5525 5733 5559
rect 5767 5556 5779 5559
rect 7484 5556 7512 5596
rect 8110 5584 8116 5596
rect 8168 5584 8174 5636
rect 8938 5624 8944 5636
rect 8404 5596 8944 5624
rect 7650 5556 7656 5568
rect 5767 5528 7512 5556
rect 7611 5528 7656 5556
rect 5767 5525 5779 5528
rect 5721 5519 5779 5525
rect 7650 5516 7656 5528
rect 7708 5516 7714 5568
rect 8018 5516 8024 5568
rect 8076 5556 8082 5568
rect 8404 5556 8432 5596
rect 8938 5584 8944 5596
rect 8996 5584 9002 5636
rect 10778 5584 10784 5636
rect 10836 5624 10842 5636
rect 12066 5624 12072 5636
rect 10836 5596 12072 5624
rect 10836 5584 10842 5596
rect 12066 5584 12072 5596
rect 12124 5584 12130 5636
rect 14366 5584 14372 5636
rect 14424 5624 14430 5636
rect 14461 5627 14519 5633
rect 14461 5624 14473 5627
rect 14424 5596 14473 5624
rect 14424 5584 14430 5596
rect 14461 5593 14473 5596
rect 14507 5624 14519 5627
rect 17494 5624 17500 5636
rect 14507 5596 17500 5624
rect 14507 5593 14519 5596
rect 14461 5587 14519 5593
rect 17494 5584 17500 5596
rect 17552 5584 17558 5636
rect 8076 5528 8432 5556
rect 8076 5516 8082 5528
rect 8478 5516 8484 5568
rect 8536 5556 8542 5568
rect 10318 5556 10324 5568
rect 8536 5528 10324 5556
rect 8536 5516 8542 5528
rect 10318 5516 10324 5528
rect 10376 5516 10382 5568
rect 10410 5516 10416 5568
rect 10468 5556 10474 5568
rect 11057 5559 11115 5565
rect 11057 5556 11069 5559
rect 10468 5528 11069 5556
rect 10468 5516 10474 5528
rect 11057 5525 11069 5528
rect 11103 5525 11115 5559
rect 11057 5519 11115 5525
rect 12710 5516 12716 5568
rect 12768 5556 12774 5568
rect 14090 5556 14096 5568
rect 12768 5528 14096 5556
rect 12768 5516 12774 5528
rect 14090 5516 14096 5528
rect 14148 5516 14154 5568
rect 15654 5556 15660 5568
rect 15615 5528 15660 5556
rect 15654 5516 15660 5528
rect 15712 5516 15718 5568
rect 16206 5556 16212 5568
rect 16167 5528 16212 5556
rect 16206 5516 16212 5528
rect 16264 5516 16270 5568
rect 17402 5556 17408 5568
rect 17363 5528 17408 5556
rect 17402 5516 17408 5528
rect 17460 5516 17466 5568
rect 1104 5466 18860 5488
rect 1104 5414 3947 5466
rect 3999 5414 4011 5466
rect 4063 5414 4075 5466
rect 4127 5414 4139 5466
rect 4191 5414 9878 5466
rect 9930 5414 9942 5466
rect 9994 5414 10006 5466
rect 10058 5414 10070 5466
rect 10122 5414 15808 5466
rect 15860 5414 15872 5466
rect 15924 5414 15936 5466
rect 15988 5414 16000 5466
rect 16052 5414 18860 5466
rect 1104 5392 18860 5414
rect 1854 5352 1860 5364
rect 1815 5324 1860 5352
rect 1854 5312 1860 5324
rect 1912 5312 1918 5364
rect 3697 5355 3755 5361
rect 3697 5321 3709 5355
rect 3743 5352 3755 5355
rect 4430 5352 4436 5364
rect 3743 5324 4436 5352
rect 3743 5321 3755 5324
rect 3697 5315 3755 5321
rect 4430 5312 4436 5324
rect 4488 5312 4494 5364
rect 8294 5352 8300 5364
rect 4908 5324 8300 5352
rect 4908 5284 4936 5324
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 9490 5352 9496 5364
rect 9451 5324 9496 5352
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 10778 5352 10784 5364
rect 9600 5324 10784 5352
rect 6270 5284 6276 5296
rect 2608 5256 4936 5284
rect 6231 5256 6276 5284
rect 2608 5157 2636 5256
rect 6270 5244 6276 5256
rect 6328 5244 6334 5296
rect 7282 5284 7288 5296
rect 7243 5256 7288 5284
rect 7282 5244 7288 5256
rect 7340 5244 7346 5296
rect 8018 5244 8024 5296
rect 8076 5244 8082 5296
rect 2866 5176 2872 5228
rect 2924 5216 2930 5228
rect 4341 5219 4399 5225
rect 2924 5188 4108 5216
rect 2924 5176 2930 5188
rect 4080 5157 4108 5188
rect 4341 5185 4353 5219
rect 4387 5216 4399 5219
rect 4706 5216 4712 5228
rect 4387 5188 4712 5216
rect 4387 5185 4399 5188
rect 4341 5179 4399 5185
rect 4706 5176 4712 5188
rect 4764 5176 4770 5228
rect 5994 5176 6000 5228
rect 6052 5216 6058 5228
rect 8036 5216 8064 5244
rect 6052 5188 8064 5216
rect 6052 5176 6058 5188
rect 1673 5151 1731 5157
rect 1673 5117 1685 5151
rect 1719 5117 1731 5151
rect 1673 5111 1731 5117
rect 2603 5151 2661 5157
rect 2603 5117 2615 5151
rect 2649 5117 2661 5151
rect 2603 5111 2661 5117
rect 4065 5151 4123 5157
rect 4065 5117 4077 5151
rect 4111 5117 4123 5151
rect 4065 5111 4123 5117
rect 1688 5012 1716 5111
rect 2866 5080 2872 5092
rect 2827 5052 2872 5080
rect 2866 5040 2872 5052
rect 2924 5040 2930 5092
rect 4080 5080 4108 5111
rect 4522 5108 4528 5160
rect 4580 5148 4586 5160
rect 4890 5148 4896 5160
rect 4580 5120 4896 5148
rect 4580 5108 4586 5120
rect 4890 5108 4896 5120
rect 4948 5108 4954 5160
rect 5000 5120 6684 5148
rect 5000 5080 5028 5120
rect 4080 5052 5028 5080
rect 5074 5040 5080 5092
rect 5132 5089 5138 5092
rect 5132 5083 5196 5089
rect 5132 5049 5150 5083
rect 5184 5049 5196 5083
rect 6656 5080 6684 5120
rect 6730 5108 6736 5160
rect 6788 5148 6794 5160
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6788 5120 6837 5148
rect 6788 5108 6794 5120
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 7193 5151 7251 5157
rect 7193 5117 7205 5151
rect 7239 5148 7251 5151
rect 7374 5148 7380 5160
rect 7239 5120 7380 5148
rect 7239 5117 7251 5120
rect 7193 5111 7251 5117
rect 7374 5108 7380 5120
rect 7432 5108 7438 5160
rect 8018 5108 8024 5160
rect 8076 5148 8082 5160
rect 8113 5151 8171 5157
rect 8113 5148 8125 5151
rect 8076 5120 8125 5148
rect 8076 5108 8082 5120
rect 8113 5117 8125 5120
rect 8159 5117 8171 5151
rect 9600 5148 9628 5324
rect 10778 5312 10784 5324
rect 10836 5312 10842 5364
rect 15470 5352 15476 5364
rect 15431 5324 15476 5352
rect 15470 5312 15476 5324
rect 15528 5312 15534 5364
rect 16666 5352 16672 5364
rect 16627 5324 16672 5352
rect 16666 5312 16672 5324
rect 16724 5312 16730 5364
rect 11974 5284 11980 5296
rect 11164 5256 11980 5284
rect 9674 5176 9680 5228
rect 9732 5216 9738 5228
rect 10137 5219 10195 5225
rect 10137 5216 10149 5219
rect 9732 5188 10149 5216
rect 9732 5176 9738 5188
rect 10137 5185 10149 5188
rect 10183 5185 10195 5219
rect 10137 5179 10195 5185
rect 8113 5111 8171 5117
rect 8312 5120 9628 5148
rect 8312 5080 8340 5120
rect 6656 5052 8340 5080
rect 8380 5083 8438 5089
rect 5132 5043 5196 5049
rect 8380 5049 8392 5083
rect 8426 5080 8438 5083
rect 9030 5080 9036 5092
rect 8426 5052 9036 5080
rect 8426 5049 8438 5052
rect 8380 5043 8438 5049
rect 5132 5040 5138 5043
rect 9030 5040 9036 5052
rect 9088 5040 9094 5092
rect 10152 5080 10180 5179
rect 10410 5157 10416 5160
rect 10404 5148 10416 5157
rect 10371 5120 10416 5148
rect 10404 5111 10416 5120
rect 10410 5108 10416 5111
rect 10468 5108 10474 5160
rect 11164 5148 11192 5256
rect 11974 5244 11980 5256
rect 12032 5244 12038 5296
rect 12434 5284 12440 5296
rect 12176 5256 12440 5284
rect 12176 5157 12204 5256
rect 12434 5244 12440 5256
rect 12492 5244 12498 5296
rect 12621 5287 12679 5293
rect 12621 5253 12633 5287
rect 12667 5284 12679 5287
rect 13998 5284 14004 5296
rect 12667 5256 14004 5284
rect 12667 5253 12679 5256
rect 12621 5247 12679 5253
rect 13998 5244 14004 5256
rect 14056 5244 14062 5296
rect 13265 5219 13323 5225
rect 13265 5185 13277 5219
rect 13311 5216 13323 5219
rect 13630 5216 13636 5228
rect 13311 5188 13636 5216
rect 13311 5185 13323 5188
rect 13265 5179 13323 5185
rect 13630 5176 13636 5188
rect 13688 5176 13694 5228
rect 14277 5219 14335 5225
rect 14277 5185 14289 5219
rect 14323 5216 14335 5219
rect 14458 5216 14464 5228
rect 14323 5188 14464 5216
rect 14323 5185 14335 5188
rect 14277 5179 14335 5185
rect 14458 5176 14464 5188
rect 14516 5176 14522 5228
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5216 16175 5219
rect 16390 5216 16396 5228
rect 16163 5188 16396 5216
rect 16163 5185 16175 5188
rect 16117 5179 16175 5185
rect 16390 5176 16396 5188
rect 16448 5176 16454 5228
rect 17218 5216 17224 5228
rect 17179 5188 17224 5216
rect 17218 5176 17224 5188
rect 17276 5176 17282 5228
rect 10796 5120 11192 5148
rect 12161 5151 12219 5157
rect 10318 5080 10324 5092
rect 10152 5052 10324 5080
rect 10318 5040 10324 5052
rect 10376 5080 10382 5092
rect 10796 5080 10824 5120
rect 12161 5117 12173 5151
rect 12207 5117 12219 5151
rect 12161 5111 12219 5117
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5148 12495 5151
rect 12710 5148 12716 5160
rect 12483 5120 12716 5148
rect 12483 5117 12495 5120
rect 12437 5111 12495 5117
rect 12710 5108 12716 5120
rect 12768 5108 12774 5160
rect 14737 5151 14795 5157
rect 14737 5117 14749 5151
rect 14783 5117 14795 5151
rect 14737 5111 14795 5117
rect 15841 5151 15899 5157
rect 15841 5117 15853 5151
rect 15887 5148 15899 5151
rect 16206 5148 16212 5160
rect 15887 5120 16212 5148
rect 15887 5117 15899 5120
rect 15841 5111 15899 5117
rect 10376 5052 10824 5080
rect 10376 5040 10382 5052
rect 13262 5040 13268 5092
rect 13320 5080 13326 5092
rect 13357 5083 13415 5089
rect 13357 5080 13369 5083
rect 13320 5052 13369 5080
rect 13320 5040 13326 5052
rect 13357 5049 13369 5052
rect 13403 5049 13415 5083
rect 14752 5080 14780 5111
rect 16206 5108 16212 5120
rect 16264 5108 16270 5160
rect 17034 5148 17040 5160
rect 16995 5120 17040 5148
rect 17034 5108 17040 5120
rect 17092 5108 17098 5160
rect 13357 5043 13415 5049
rect 13464 5052 14780 5080
rect 15933 5083 15991 5089
rect 4062 5012 4068 5024
rect 1688 4984 4068 5012
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 4157 5015 4215 5021
rect 4157 4981 4169 5015
rect 4203 5012 4215 5015
rect 5626 5012 5632 5024
rect 4203 4984 5632 5012
rect 4203 4981 4215 4984
rect 4157 4975 4215 4981
rect 5626 4972 5632 4984
rect 5684 4972 5690 5024
rect 8202 4972 8208 5024
rect 8260 5012 8266 5024
rect 9214 5012 9220 5024
rect 8260 4984 9220 5012
rect 8260 4972 8266 4984
rect 9214 4972 9220 4984
rect 9272 5012 9278 5024
rect 9490 5012 9496 5024
rect 9272 4984 9496 5012
rect 9272 4972 9278 4984
rect 9490 4972 9496 4984
rect 9548 4972 9554 5024
rect 10686 4972 10692 5024
rect 10744 5012 10750 5024
rect 11517 5015 11575 5021
rect 11517 5012 11529 5015
rect 10744 4984 11529 5012
rect 10744 4972 10750 4984
rect 11517 4981 11529 4984
rect 11563 4981 11575 5015
rect 11517 4975 11575 4981
rect 11698 4972 11704 5024
rect 11756 5012 11762 5024
rect 13464 5012 13492 5052
rect 15933 5049 15945 5083
rect 15979 5080 15991 5083
rect 17402 5080 17408 5092
rect 15979 5052 17408 5080
rect 15979 5049 15991 5052
rect 15933 5043 15991 5049
rect 17402 5040 17408 5052
rect 17460 5040 17466 5092
rect 11756 4984 13492 5012
rect 11756 4972 11762 4984
rect 14734 4972 14740 5024
rect 14792 5012 14798 5024
rect 14921 5015 14979 5021
rect 14921 5012 14933 5015
rect 14792 4984 14933 5012
rect 14792 4972 14798 4984
rect 14921 4981 14933 4984
rect 14967 4981 14979 5015
rect 14921 4975 14979 4981
rect 16022 4972 16028 5024
rect 16080 5012 16086 5024
rect 17129 5015 17187 5021
rect 17129 5012 17141 5015
rect 16080 4984 17141 5012
rect 16080 4972 16086 4984
rect 17129 4981 17141 4984
rect 17175 4981 17187 5015
rect 17129 4975 17187 4981
rect 1104 4922 18860 4944
rect 1104 4870 6912 4922
rect 6964 4870 6976 4922
rect 7028 4870 7040 4922
rect 7092 4870 7104 4922
rect 7156 4870 12843 4922
rect 12895 4870 12907 4922
rect 12959 4870 12971 4922
rect 13023 4870 13035 4922
rect 13087 4870 18860 4922
rect 1104 4848 18860 4870
rect 1762 4768 1768 4820
rect 1820 4808 1826 4820
rect 1857 4811 1915 4817
rect 1857 4808 1869 4811
rect 1820 4780 1869 4808
rect 1820 4768 1826 4780
rect 1857 4777 1869 4780
rect 1903 4777 1915 4811
rect 1857 4771 1915 4777
rect 2593 4811 2651 4817
rect 2593 4777 2605 4811
rect 2639 4808 2651 4811
rect 2774 4808 2780 4820
rect 2639 4780 2780 4808
rect 2639 4777 2651 4780
rect 2593 4771 2651 4777
rect 2774 4768 2780 4780
rect 2832 4768 2838 4820
rect 2958 4768 2964 4820
rect 3016 4808 3022 4820
rect 3142 4808 3148 4820
rect 3016 4780 3148 4808
rect 3016 4768 3022 4780
rect 3142 4768 3148 4780
rect 3200 4768 3206 4820
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 5258 4808 5264 4820
rect 4120 4780 5264 4808
rect 4120 4768 4126 4780
rect 5258 4768 5264 4780
rect 5316 4768 5322 4820
rect 5626 4808 5632 4820
rect 5587 4780 5632 4808
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 8846 4808 8852 4820
rect 6932 4780 8852 4808
rect 2314 4740 2320 4752
rect 1688 4712 2320 4740
rect 1688 4681 1716 4712
rect 2314 4700 2320 4712
rect 2372 4700 2378 4752
rect 3160 4712 5304 4740
rect 1673 4675 1731 4681
rect 1673 4641 1685 4675
rect 1719 4641 1731 4675
rect 2406 4672 2412 4684
rect 2367 4644 2412 4672
rect 1673 4635 1731 4641
rect 2406 4632 2412 4644
rect 2464 4632 2470 4684
rect 3160 4681 3188 4712
rect 3145 4675 3203 4681
rect 3145 4641 3157 4675
rect 3191 4641 3203 4675
rect 4798 4672 4804 4684
rect 4759 4644 4804 4672
rect 3145 4635 3203 4641
rect 4798 4632 4804 4644
rect 4856 4632 4862 4684
rect 4893 4675 4951 4681
rect 4893 4641 4905 4675
rect 4939 4672 4951 4675
rect 4982 4672 4988 4684
rect 4939 4644 4988 4672
rect 4939 4641 4951 4644
rect 4893 4635 4951 4641
rect 4982 4632 4988 4644
rect 5040 4632 5046 4684
rect 5276 4672 5304 4712
rect 5534 4672 5540 4684
rect 5276 4644 5540 4672
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 5994 4672 6000 4684
rect 5955 4644 6000 4672
rect 5994 4632 6000 4644
rect 6052 4632 6058 4684
rect 6089 4675 6147 4681
rect 6089 4641 6101 4675
rect 6135 4672 6147 4675
rect 6454 4672 6460 4684
rect 6135 4644 6460 4672
rect 6135 4641 6147 4644
rect 6089 4635 6147 4641
rect 6454 4632 6460 4644
rect 6512 4632 6518 4684
rect 6932 4681 6960 4780
rect 8846 4768 8852 4780
rect 8904 4768 8910 4820
rect 9030 4808 9036 4820
rect 8991 4780 9036 4808
rect 9030 4768 9036 4780
rect 9088 4768 9094 4820
rect 9122 4768 9128 4820
rect 9180 4808 9186 4820
rect 9677 4811 9735 4817
rect 9677 4808 9689 4811
rect 9180 4780 9689 4808
rect 9180 4768 9186 4780
rect 9677 4777 9689 4780
rect 9723 4777 9735 4811
rect 9677 4771 9735 4777
rect 12434 4768 12440 4820
rect 12492 4808 12498 4820
rect 13906 4808 13912 4820
rect 12492 4780 13912 4808
rect 12492 4768 12498 4780
rect 13906 4768 13912 4780
rect 13964 4768 13970 4820
rect 14458 4768 14464 4820
rect 14516 4808 14522 4820
rect 16850 4808 16856 4820
rect 14516 4780 15599 4808
rect 16811 4780 16856 4808
rect 14516 4768 14522 4780
rect 8018 4740 8024 4752
rect 7668 4712 8024 4740
rect 6917 4675 6975 4681
rect 6917 4641 6929 4675
rect 6963 4641 6975 4675
rect 6917 4635 6975 4641
rect 5074 4604 5080 4616
rect 5035 4576 5080 4604
rect 5074 4564 5080 4576
rect 5132 4604 5138 4616
rect 5442 4604 5448 4616
rect 5132 4576 5448 4604
rect 5132 4564 5138 4576
rect 5442 4564 5448 4576
rect 5500 4604 5506 4616
rect 6181 4607 6239 4613
rect 6181 4604 6193 4607
rect 5500 4576 6193 4604
rect 5500 4564 5506 4576
rect 6181 4573 6193 4576
rect 6227 4604 6239 4607
rect 6362 4604 6368 4616
rect 6227 4576 6368 4604
rect 6227 4573 6239 4576
rect 6181 4567 6239 4573
rect 6362 4564 6368 4576
rect 6420 4564 6426 4616
rect 6822 4564 6828 4616
rect 6880 4604 6886 4616
rect 7668 4613 7696 4712
rect 8018 4700 8024 4712
rect 8076 4700 8082 4752
rect 11790 4740 11796 4752
rect 11751 4712 11796 4740
rect 11790 4700 11796 4712
rect 11848 4700 11854 4752
rect 11885 4743 11943 4749
rect 11885 4709 11897 4743
rect 11931 4740 11943 4743
rect 11974 4740 11980 4752
rect 11931 4712 11980 4740
rect 11931 4709 11943 4712
rect 11885 4703 11943 4709
rect 11974 4700 11980 4712
rect 12032 4700 12038 4752
rect 13354 4700 13360 4752
rect 13412 4740 13418 4752
rect 13725 4743 13783 4749
rect 13725 4740 13737 4743
rect 13412 4712 13737 4740
rect 13412 4700 13418 4712
rect 13725 4709 13737 4712
rect 13771 4709 13783 4743
rect 13725 4703 13783 4709
rect 13817 4743 13875 4749
rect 13817 4709 13829 4743
rect 13863 4740 13875 4743
rect 14090 4740 14096 4752
rect 13863 4712 14096 4740
rect 13863 4709 13875 4712
rect 13817 4703 13875 4709
rect 14090 4700 14096 4712
rect 14148 4740 14154 4752
rect 15010 4740 15016 4752
rect 14148 4712 15016 4740
rect 14148 4700 14154 4712
rect 15010 4700 15016 4712
rect 15068 4700 15074 4752
rect 15378 4700 15384 4752
rect 15436 4740 15442 4752
rect 15473 4743 15531 4749
rect 15473 4740 15485 4743
rect 15436 4712 15485 4740
rect 15436 4700 15442 4712
rect 15473 4709 15485 4712
rect 15519 4709 15531 4743
rect 15571 4740 15599 4780
rect 16850 4768 16856 4780
rect 16908 4768 16914 4820
rect 17221 4811 17279 4817
rect 17221 4777 17233 4811
rect 17267 4808 17279 4811
rect 18230 4808 18236 4820
rect 17267 4780 18236 4808
rect 17267 4777 17279 4780
rect 17221 4771 17279 4777
rect 17313 4743 17371 4749
rect 17313 4740 17325 4743
rect 15571 4712 17325 4740
rect 15473 4703 15531 4709
rect 17313 4709 17325 4712
rect 17359 4709 17371 4743
rect 17313 4703 17371 4709
rect 7920 4675 7978 4681
rect 7920 4641 7932 4675
rect 7966 4672 7978 4675
rect 8478 4672 8484 4684
rect 7966 4644 8484 4672
rect 7966 4641 7978 4644
rect 7920 4635 7978 4641
rect 8478 4632 8484 4644
rect 8536 4632 8542 4684
rect 10686 4672 10692 4684
rect 10647 4644 10692 4672
rect 10686 4632 10692 4644
rect 10744 4632 10750 4684
rect 16390 4632 16396 4684
rect 16448 4672 16454 4684
rect 17420 4672 17448 4780
rect 18230 4768 18236 4780
rect 18288 4768 18294 4820
rect 16448 4644 17448 4672
rect 16448 4632 16454 4644
rect 7653 4607 7711 4613
rect 7653 4604 7665 4607
rect 6880 4576 7665 4604
rect 6880 4564 6886 4576
rect 7653 4573 7665 4576
rect 7699 4573 7711 4607
rect 7653 4567 7711 4573
rect 8938 4564 8944 4616
rect 8996 4604 9002 4616
rect 10321 4607 10379 4613
rect 10321 4604 10333 4607
rect 8996 4576 10333 4604
rect 8996 4564 9002 4576
rect 10321 4573 10333 4576
rect 10367 4573 10379 4607
rect 10321 4567 10379 4573
rect 12805 4607 12863 4613
rect 12805 4573 12817 4607
rect 12851 4604 12863 4607
rect 13814 4604 13820 4616
rect 12851 4576 13820 4604
rect 12851 4573 12863 4576
rect 12805 4567 12863 4573
rect 13814 4564 13820 4576
rect 13872 4564 13878 4616
rect 14737 4607 14795 4613
rect 14737 4573 14749 4607
rect 14783 4573 14795 4607
rect 15378 4604 15384 4616
rect 15339 4576 15384 4604
rect 14737 4567 14795 4573
rect 9490 4496 9496 4548
rect 9548 4536 9554 4548
rect 14090 4536 14096 4548
rect 9548 4508 14096 4536
rect 9548 4496 9554 4508
rect 14090 4496 14096 4508
rect 14148 4496 14154 4548
rect 14752 4536 14780 4567
rect 15378 4564 15384 4576
rect 15436 4564 15442 4616
rect 15562 4564 15568 4616
rect 15620 4604 15626 4616
rect 15657 4607 15715 4613
rect 15657 4604 15669 4607
rect 15620 4576 15669 4604
rect 15620 4564 15626 4576
rect 15657 4573 15669 4576
rect 15703 4573 15715 4607
rect 15657 4567 15715 4573
rect 16666 4564 16672 4616
rect 16724 4604 16730 4616
rect 17310 4604 17316 4616
rect 16724 4576 17316 4604
rect 16724 4564 16730 4576
rect 17310 4564 17316 4576
rect 17368 4564 17374 4616
rect 17494 4604 17500 4616
rect 17455 4576 17500 4604
rect 17494 4564 17500 4576
rect 17552 4564 17558 4616
rect 17678 4536 17684 4548
rect 14752 4508 17684 4536
rect 17678 4496 17684 4508
rect 17736 4496 17742 4548
rect 3050 4428 3056 4480
rect 3108 4468 3114 4480
rect 3329 4471 3387 4477
rect 3329 4468 3341 4471
rect 3108 4440 3341 4468
rect 3108 4428 3114 4440
rect 3329 4437 3341 4440
rect 3375 4437 3387 4471
rect 4430 4468 4436 4480
rect 4391 4440 4436 4468
rect 3329 4431 3387 4437
rect 4430 4428 4436 4440
rect 4488 4428 4494 4480
rect 7101 4471 7159 4477
rect 7101 4437 7113 4471
rect 7147 4468 7159 4471
rect 9122 4468 9128 4480
rect 7147 4440 9128 4468
rect 7147 4437 7159 4440
rect 7101 4431 7159 4437
rect 9122 4428 9128 4440
rect 9180 4428 9186 4480
rect 9766 4428 9772 4480
rect 9824 4468 9830 4480
rect 10781 4471 10839 4477
rect 10781 4468 10793 4471
rect 9824 4440 10793 4468
rect 9824 4428 9830 4440
rect 10781 4437 10793 4440
rect 10827 4468 10839 4471
rect 16206 4468 16212 4480
rect 10827 4440 16212 4468
rect 10827 4437 10839 4440
rect 10781 4431 10839 4437
rect 16206 4428 16212 4440
rect 16264 4428 16270 4480
rect 1104 4378 18860 4400
rect 1104 4326 3947 4378
rect 3999 4326 4011 4378
rect 4063 4326 4075 4378
rect 4127 4326 4139 4378
rect 4191 4326 9878 4378
rect 9930 4326 9942 4378
rect 9994 4326 10006 4378
rect 10058 4326 10070 4378
rect 10122 4326 15808 4378
rect 15860 4326 15872 4378
rect 15924 4326 15936 4378
rect 15988 4326 16000 4378
rect 16052 4326 18860 4378
rect 1104 4304 18860 4326
rect 1854 4264 1860 4276
rect 1815 4236 1860 4264
rect 1854 4224 1860 4236
rect 1912 4224 1918 4276
rect 3973 4267 4031 4273
rect 3973 4233 3985 4267
rect 4019 4264 4031 4267
rect 4338 4264 4344 4276
rect 4019 4236 4344 4264
rect 4019 4233 4031 4236
rect 3973 4227 4031 4233
rect 4338 4224 4344 4236
rect 4396 4224 4402 4276
rect 4522 4224 4528 4276
rect 4580 4264 4586 4276
rect 4580 4236 6500 4264
rect 4580 4224 4586 4236
rect 4706 4196 4712 4208
rect 4632 4168 4712 4196
rect 198 4088 204 4140
rect 256 4128 262 4140
rect 1946 4128 1952 4140
rect 256 4100 1952 4128
rect 256 4088 262 4100
rect 1946 4088 1952 4100
rect 2004 4088 2010 4140
rect 4430 4128 4436 4140
rect 4391 4100 4436 4128
rect 4430 4088 4436 4100
rect 4488 4088 4494 4140
rect 4632 4137 4660 4168
rect 4706 4156 4712 4168
rect 4764 4156 4770 4208
rect 6270 4196 6276 4208
rect 5644 4168 6276 4196
rect 5644 4137 5672 4168
rect 6270 4156 6276 4168
rect 6328 4156 6334 4208
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4097 4675 4131
rect 4617 4091 4675 4097
rect 5629 4131 5687 4137
rect 5629 4097 5641 4131
rect 5675 4097 5687 4131
rect 5629 4091 5687 4097
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 6362 4128 6368 4140
rect 5859 4100 6368 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 6362 4088 6368 4100
rect 6420 4088 6426 4140
rect 6472 4128 6500 4236
rect 6546 4224 6552 4276
rect 6604 4264 6610 4276
rect 9490 4264 9496 4276
rect 6604 4236 9496 4264
rect 6604 4224 6610 4236
rect 9490 4224 9496 4236
rect 9548 4224 9554 4276
rect 10410 4264 10416 4276
rect 10152 4236 10416 4264
rect 8386 4156 8392 4208
rect 8444 4196 8450 4208
rect 8938 4196 8944 4208
rect 8444 4168 8944 4196
rect 8444 4156 8450 4168
rect 8938 4156 8944 4168
rect 8996 4196 9002 4208
rect 9033 4199 9091 4205
rect 9033 4196 9045 4199
rect 8996 4168 9045 4196
rect 8996 4156 9002 4168
rect 9033 4165 9045 4168
rect 9079 4165 9091 4199
rect 9033 4159 9091 4165
rect 6822 4128 6828 4140
rect 6472 4100 6828 4128
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 9048 4128 9076 4159
rect 10042 4128 10048 4140
rect 9048 4100 10048 4128
rect 10042 4088 10048 4100
rect 10100 4088 10106 4140
rect 1673 4063 1731 4069
rect 1673 4029 1685 4063
rect 1719 4029 1731 4063
rect 1673 4023 1731 4029
rect 2409 4063 2467 4069
rect 2409 4029 2421 4063
rect 2455 4060 2467 4063
rect 2682 4060 2688 4072
rect 2455 4032 2688 4060
rect 2455 4029 2467 4032
rect 2409 4023 2467 4029
rect 1688 3992 1716 4023
rect 2682 4020 2688 4032
rect 2740 4020 2746 4072
rect 3142 4060 3148 4072
rect 3103 4032 3148 4060
rect 3142 4020 3148 4032
rect 3200 4020 3206 4072
rect 3878 4020 3884 4072
rect 3936 4060 3942 4072
rect 5994 4060 6000 4072
rect 3936 4032 6000 4060
rect 3936 4020 3942 4032
rect 5994 4020 6000 4032
rect 6052 4020 6058 4072
rect 6270 4020 6276 4072
rect 6328 4060 6334 4072
rect 9401 4063 9459 4069
rect 6328 4032 7052 4060
rect 6328 4020 6334 4032
rect 5534 3992 5540 4004
rect 1688 3964 5304 3992
rect 5495 3964 5540 3992
rect 2593 3927 2651 3933
rect 2593 3893 2605 3927
rect 2639 3924 2651 3927
rect 2774 3924 2780 3936
rect 2639 3896 2780 3924
rect 2639 3893 2651 3896
rect 2593 3887 2651 3893
rect 2774 3884 2780 3896
rect 2832 3884 2838 3936
rect 3326 3924 3332 3936
rect 3287 3896 3332 3924
rect 3326 3884 3332 3896
rect 3384 3884 3390 3936
rect 4341 3927 4399 3933
rect 4341 3893 4353 3927
rect 4387 3924 4399 3927
rect 5169 3927 5227 3933
rect 5169 3924 5181 3927
rect 4387 3896 5181 3924
rect 4387 3893 4399 3896
rect 4341 3887 4399 3893
rect 5169 3893 5181 3896
rect 5215 3893 5227 3927
rect 5276 3924 5304 3964
rect 5534 3952 5540 3964
rect 5592 3952 5598 4004
rect 5810 3952 5816 4004
rect 5868 3992 5874 4004
rect 6546 3992 6552 4004
rect 5868 3964 6552 3992
rect 5868 3952 5874 3964
rect 6546 3952 6552 3964
rect 6604 3952 6610 4004
rect 6914 3952 6920 4004
rect 6972 3952 6978 4004
rect 6932 3924 6960 3952
rect 5276 3896 6960 3924
rect 7024 3924 7052 4032
rect 9401 4029 9413 4063
rect 9447 4060 9459 4063
rect 10152 4060 10180 4236
rect 10410 4224 10416 4236
rect 10468 4224 10474 4276
rect 13556 4168 13860 4196
rect 12897 4131 12955 4137
rect 12897 4097 12909 4131
rect 12943 4128 12955 4131
rect 13170 4128 13176 4140
rect 12943 4100 13176 4128
rect 12943 4097 12955 4100
rect 12897 4091 12955 4097
rect 13170 4088 13176 4100
rect 13228 4088 13234 4140
rect 13262 4088 13268 4140
rect 13320 4128 13326 4140
rect 13556 4128 13584 4168
rect 13722 4128 13728 4140
rect 13320 4100 13584 4128
rect 13683 4100 13728 4128
rect 13320 4088 13326 4100
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 13832 4128 13860 4168
rect 14752 4168 15056 4196
rect 14752 4128 14780 4168
rect 14918 4128 14924 4140
rect 13832 4100 14780 4128
rect 14879 4100 14924 4128
rect 14918 4088 14924 4100
rect 14976 4088 14982 4140
rect 15028 4128 15056 4168
rect 16117 4131 16175 4137
rect 16117 4128 16129 4131
rect 15028 4100 16129 4128
rect 16117 4097 16129 4100
rect 16163 4097 16175 4131
rect 17126 4128 17132 4140
rect 17087 4100 17132 4128
rect 16117 4091 16175 4097
rect 17126 4088 17132 4100
rect 17184 4088 17190 4140
rect 9447 4032 10180 4060
rect 10229 4063 10287 4069
rect 9447 4029 9459 4032
rect 9401 4023 9459 4029
rect 10229 4029 10241 4063
rect 10275 4060 10287 4063
rect 10318 4060 10324 4072
rect 10275 4032 10324 4060
rect 10275 4029 10287 4032
rect 10229 4023 10287 4029
rect 10318 4020 10324 4032
rect 10376 4020 10382 4072
rect 11882 4060 11888 4072
rect 10428 4032 11888 4060
rect 7092 3995 7150 4001
rect 7092 3961 7104 3995
rect 7138 3992 7150 3995
rect 7282 3992 7288 4004
rect 7138 3964 7288 3992
rect 7138 3961 7150 3964
rect 7092 3955 7150 3961
rect 7282 3952 7288 3964
rect 7340 3952 7346 4004
rect 10428 3992 10456 4032
rect 11882 4020 11888 4032
rect 11940 4020 11946 4072
rect 7392 3964 10456 3992
rect 10496 3995 10554 4001
rect 7392 3924 7420 3964
rect 10496 3961 10508 3995
rect 10542 3992 10554 3995
rect 10686 3992 10692 4004
rect 10542 3964 10692 3992
rect 10542 3961 10554 3964
rect 10496 3955 10554 3961
rect 10686 3952 10692 3964
rect 10744 3952 10750 4004
rect 12989 3995 13047 4001
rect 12989 3961 13001 3995
rect 13035 3992 13047 3995
rect 13538 3992 13544 4004
rect 13035 3964 13544 3992
rect 13035 3961 13047 3964
rect 12989 3955 13047 3961
rect 13538 3952 13544 3964
rect 13596 3952 13602 4004
rect 14090 3952 14096 4004
rect 14148 3992 14154 4004
rect 14461 3995 14519 4001
rect 14461 3992 14473 3995
rect 14148 3964 14473 3992
rect 14148 3952 14154 3964
rect 14461 3961 14473 3964
rect 14507 3961 14519 3995
rect 14461 3955 14519 3961
rect 14550 3952 14556 4004
rect 14608 3992 14614 4004
rect 16206 3992 16212 4004
rect 14608 3964 14653 3992
rect 16167 3964 16212 3992
rect 14608 3952 14614 3964
rect 16206 3952 16212 3964
rect 16264 3952 16270 4004
rect 7024 3896 7420 3924
rect 8205 3927 8263 3933
rect 5169 3887 5227 3893
rect 8205 3893 8217 3927
rect 8251 3924 8263 3927
rect 8478 3924 8484 3936
rect 8251 3896 8484 3924
rect 8251 3893 8263 3896
rect 8205 3887 8263 3893
rect 8478 3884 8484 3896
rect 8536 3884 8542 3936
rect 8662 3884 8668 3936
rect 8720 3924 8726 3936
rect 9306 3924 9312 3936
rect 8720 3896 9312 3924
rect 8720 3884 8726 3896
rect 9306 3884 9312 3896
rect 9364 3884 9370 3936
rect 9858 3884 9864 3936
rect 9916 3924 9922 3936
rect 11609 3927 11667 3933
rect 11609 3924 11621 3927
rect 9916 3896 11621 3924
rect 9916 3884 9922 3896
rect 11609 3893 11621 3896
rect 11655 3893 11667 3927
rect 11609 3887 11667 3893
rect 14274 3884 14280 3936
rect 14332 3924 14338 3936
rect 15654 3924 15660 3936
rect 14332 3896 15660 3924
rect 14332 3884 14338 3896
rect 15654 3884 15660 3896
rect 15712 3884 15718 3936
rect 1104 3834 18860 3856
rect 1104 3782 6912 3834
rect 6964 3782 6976 3834
rect 7028 3782 7040 3834
rect 7092 3782 7104 3834
rect 7156 3782 12843 3834
rect 12895 3782 12907 3834
rect 12959 3782 12971 3834
rect 13023 3782 13035 3834
rect 13087 3782 18860 3834
rect 1104 3760 18860 3782
rect 3878 3720 3884 3732
rect 1688 3692 3884 3720
rect 1688 3593 1716 3692
rect 3878 3680 3884 3692
rect 3936 3680 3942 3732
rect 7282 3720 7288 3732
rect 7243 3692 7288 3720
rect 7282 3680 7288 3692
rect 7340 3680 7346 3732
rect 7742 3720 7748 3732
rect 7703 3692 7748 3720
rect 7742 3680 7748 3692
rect 7800 3680 7806 3732
rect 8754 3680 8760 3732
rect 8812 3720 8818 3732
rect 8849 3723 8907 3729
rect 8849 3720 8861 3723
rect 8812 3692 8861 3720
rect 8812 3680 8818 3692
rect 8849 3689 8861 3692
rect 8895 3720 8907 3723
rect 11974 3720 11980 3732
rect 8895 3692 11980 3720
rect 8895 3689 8907 3692
rect 8849 3683 8907 3689
rect 11974 3680 11980 3692
rect 12032 3680 12038 3732
rect 12250 3680 12256 3732
rect 12308 3720 12314 3732
rect 12308 3692 13032 3720
rect 12308 3680 12314 3692
rect 4522 3652 4528 3664
rect 4080 3624 4528 3652
rect 1673 3587 1731 3593
rect 1673 3553 1685 3587
rect 1719 3553 1731 3587
rect 1673 3547 1731 3553
rect 2685 3587 2743 3593
rect 2685 3553 2697 3587
rect 2731 3584 2743 3587
rect 3602 3584 3608 3596
rect 2731 3556 3608 3584
rect 2731 3553 2743 3556
rect 2685 3547 2743 3553
rect 3602 3544 3608 3556
rect 3660 3544 3666 3596
rect 4080 3593 4108 3624
rect 4522 3612 4528 3624
rect 4580 3652 4586 3664
rect 6172 3655 6230 3661
rect 4580 3624 5120 3652
rect 4580 3612 4586 3624
rect 4065 3587 4123 3593
rect 4065 3553 4077 3587
rect 4111 3553 4123 3587
rect 4065 3547 4123 3553
rect 4332 3587 4390 3593
rect 4332 3553 4344 3587
rect 4378 3584 4390 3587
rect 4614 3584 4620 3596
rect 4378 3556 4620 3584
rect 4378 3553 4390 3556
rect 4332 3547 4390 3553
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 2961 3519 3019 3525
rect 2961 3485 2973 3519
rect 3007 3516 3019 3519
rect 3234 3516 3240 3528
rect 3007 3488 3240 3516
rect 3007 3485 3019 3488
rect 2961 3479 3019 3485
rect 3234 3476 3240 3488
rect 3292 3476 3298 3528
rect 5092 3516 5120 3624
rect 6172 3621 6184 3655
rect 6218 3652 6230 3655
rect 7374 3652 7380 3664
rect 6218 3624 7380 3652
rect 6218 3621 6230 3624
rect 6172 3615 6230 3621
rect 7374 3612 7380 3624
rect 7432 3652 7438 3664
rect 7650 3652 7656 3664
rect 7432 3624 7656 3652
rect 7432 3612 7438 3624
rect 7650 3612 7656 3624
rect 7708 3612 7714 3664
rect 8018 3612 8024 3664
rect 8076 3652 8082 3664
rect 9858 3652 9864 3664
rect 8076 3624 9864 3652
rect 8076 3612 8082 3624
rect 9858 3612 9864 3624
rect 9916 3652 9922 3664
rect 9916 3624 10456 3652
rect 9916 3612 9922 3624
rect 8757 3587 8815 3593
rect 8757 3553 8769 3587
rect 8803 3584 8815 3587
rect 9030 3584 9036 3596
rect 8803 3556 9036 3584
rect 8803 3553 8815 3556
rect 8757 3547 8815 3553
rect 9030 3544 9036 3556
rect 9088 3544 9094 3596
rect 10428 3593 10456 3624
rect 10502 3612 10508 3664
rect 10560 3652 10566 3664
rect 13004 3661 13032 3692
rect 14642 3680 14648 3732
rect 14700 3720 14706 3732
rect 15378 3720 15384 3732
rect 14700 3692 15384 3720
rect 14700 3680 14706 3692
rect 15378 3680 15384 3692
rect 15436 3680 15442 3732
rect 16853 3723 16911 3729
rect 16853 3689 16865 3723
rect 16899 3720 16911 3723
rect 17770 3720 17776 3732
rect 16899 3692 17776 3720
rect 16899 3689 16911 3692
rect 16853 3683 16911 3689
rect 17770 3680 17776 3692
rect 17828 3680 17834 3732
rect 11425 3655 11483 3661
rect 11425 3652 11437 3655
rect 10560 3624 11437 3652
rect 10560 3612 10566 3624
rect 11425 3621 11437 3624
rect 11471 3621 11483 3655
rect 11425 3615 11483 3621
rect 12989 3655 13047 3661
rect 12989 3621 13001 3655
rect 13035 3621 13047 3655
rect 12989 3615 13047 3621
rect 15194 3612 15200 3664
rect 15252 3652 15258 3664
rect 15473 3655 15531 3661
rect 15473 3652 15485 3655
rect 15252 3624 15485 3652
rect 15252 3612 15258 3624
rect 15473 3621 15485 3624
rect 15519 3621 15531 3655
rect 15473 3615 15531 3621
rect 16298 3612 16304 3664
rect 16356 3652 16362 3664
rect 16393 3655 16451 3661
rect 16393 3652 16405 3655
rect 16356 3624 16405 3652
rect 16356 3612 16362 3624
rect 16393 3621 16405 3624
rect 16439 3621 16451 3655
rect 16393 3615 16451 3621
rect 17221 3655 17279 3661
rect 17221 3621 17233 3655
rect 17267 3652 17279 3655
rect 17862 3652 17868 3664
rect 17267 3624 17868 3652
rect 17267 3621 17279 3624
rect 17221 3615 17279 3621
rect 17862 3612 17868 3624
rect 17920 3612 17926 3664
rect 10413 3587 10471 3593
rect 10413 3553 10425 3587
rect 10459 3553 10471 3587
rect 14458 3584 14464 3596
rect 14419 3556 14464 3584
rect 10413 3547 10471 3553
rect 14458 3544 14464 3556
rect 14516 3544 14522 3596
rect 5905 3519 5963 3525
rect 5905 3516 5917 3519
rect 5092 3488 5917 3516
rect 5905 3485 5917 3488
rect 5951 3485 5963 3519
rect 5905 3479 5963 3485
rect 7466 3476 7472 3528
rect 7524 3516 7530 3528
rect 10778 3516 10784 3528
rect 7524 3488 10456 3516
rect 10739 3488 10784 3516
rect 7524 3476 7530 3488
rect 10428 3460 10456 3488
rect 10778 3476 10784 3488
rect 10836 3476 10842 3528
rect 11333 3519 11391 3525
rect 11333 3485 11345 3519
rect 11379 3516 11391 3519
rect 11606 3516 11612 3528
rect 11379 3488 11612 3516
rect 11379 3485 11391 3488
rect 11333 3479 11391 3485
rect 11606 3476 11612 3488
rect 11664 3476 11670 3528
rect 11701 3519 11759 3525
rect 11701 3485 11713 3519
rect 11747 3485 11759 3519
rect 11701 3479 11759 3485
rect 5442 3448 5448 3460
rect 5403 3420 5448 3448
rect 5442 3408 5448 3420
rect 5500 3408 5506 3460
rect 8386 3448 8392 3460
rect 8347 3420 8392 3448
rect 8386 3408 8392 3420
rect 8444 3408 8450 3460
rect 9766 3448 9772 3460
rect 8772 3420 9772 3448
rect 1854 3380 1860 3392
rect 1815 3352 1860 3380
rect 1854 3340 1860 3352
rect 1912 3340 1918 3392
rect 2682 3340 2688 3392
rect 2740 3380 2746 3392
rect 6270 3380 6276 3392
rect 2740 3352 6276 3380
rect 2740 3340 2746 3352
rect 6270 3340 6276 3352
rect 6328 3340 6334 3392
rect 6546 3340 6552 3392
rect 6604 3380 6610 3392
rect 8772 3380 8800 3420
rect 9766 3408 9772 3420
rect 9824 3408 9830 3460
rect 10042 3448 10048 3460
rect 10003 3420 10048 3448
rect 10042 3408 10048 3420
rect 10100 3408 10106 3460
rect 10410 3408 10416 3460
rect 10468 3408 10474 3460
rect 11422 3408 11428 3460
rect 11480 3448 11486 3460
rect 11716 3448 11744 3479
rect 12158 3476 12164 3528
rect 12216 3516 12222 3528
rect 12897 3519 12955 3525
rect 12897 3516 12909 3519
rect 12216 3488 12909 3516
rect 12216 3476 12222 3488
rect 12897 3485 12909 3488
rect 12943 3485 12955 3519
rect 13446 3516 13452 3528
rect 13407 3488 13452 3516
rect 12897 3479 12955 3485
rect 13446 3476 13452 3488
rect 13504 3476 13510 3528
rect 15102 3476 15108 3528
rect 15160 3516 15166 3528
rect 15381 3519 15439 3525
rect 15381 3516 15393 3519
rect 15160 3488 15393 3516
rect 15160 3476 15166 3488
rect 15381 3485 15393 3488
rect 15427 3485 15439 3519
rect 15381 3479 15439 3485
rect 17313 3519 17371 3525
rect 17313 3485 17325 3519
rect 17359 3485 17371 3519
rect 17494 3516 17500 3528
rect 17455 3488 17500 3516
rect 17313 3479 17371 3485
rect 11480 3420 11744 3448
rect 11480 3408 11486 3420
rect 11790 3408 11796 3460
rect 11848 3448 11854 3460
rect 17328 3448 17356 3479
rect 17494 3476 17500 3488
rect 17552 3476 17558 3528
rect 11848 3420 17356 3448
rect 11848 3408 11854 3420
rect 6604 3352 8800 3380
rect 6604 3340 6610 3352
rect 8938 3340 8944 3392
rect 8996 3380 9002 3392
rect 10778 3380 10784 3392
rect 8996 3352 10784 3380
rect 8996 3340 9002 3352
rect 10778 3340 10784 3352
rect 10836 3340 10842 3392
rect 14645 3383 14703 3389
rect 14645 3349 14657 3383
rect 14691 3380 14703 3383
rect 15562 3380 15568 3392
rect 14691 3352 15568 3380
rect 14691 3349 14703 3352
rect 14645 3343 14703 3349
rect 15562 3340 15568 3352
rect 15620 3340 15626 3392
rect 1104 3290 18860 3312
rect 1104 3238 3947 3290
rect 3999 3238 4011 3290
rect 4063 3238 4075 3290
rect 4127 3238 4139 3290
rect 4191 3238 9878 3290
rect 9930 3238 9942 3290
rect 9994 3238 10006 3290
rect 10058 3238 10070 3290
rect 10122 3238 15808 3290
rect 15860 3238 15872 3290
rect 15924 3238 15936 3290
rect 15988 3238 16000 3290
rect 16052 3238 18860 3290
rect 1104 3216 18860 3238
rect 5445 3179 5503 3185
rect 5445 3145 5457 3179
rect 5491 3176 5503 3179
rect 9674 3176 9680 3188
rect 5491 3148 9680 3176
rect 5491 3145 5503 3148
rect 5445 3139 5503 3145
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 17402 3176 17408 3188
rect 17363 3148 17408 3176
rect 17402 3136 17408 3148
rect 17460 3136 17466 3188
rect 6181 3111 6239 3117
rect 6181 3077 6193 3111
rect 6227 3108 6239 3111
rect 9766 3108 9772 3120
rect 6227 3080 9772 3108
rect 6227 3077 6239 3080
rect 6181 3071 6239 3077
rect 9766 3068 9772 3080
rect 9824 3068 9830 3120
rect 1670 3000 1676 3052
rect 1728 3040 1734 3052
rect 4433 3043 4491 3049
rect 4433 3040 4445 3043
rect 1728 3012 4445 3040
rect 1728 3000 1734 3012
rect 4433 3009 4445 3012
rect 4479 3009 4491 3043
rect 4433 3003 4491 3009
rect 4522 3000 4528 3052
rect 4580 3040 4586 3052
rect 6086 3040 6092 3052
rect 4580 3012 6092 3040
rect 4580 3000 4586 3012
rect 6086 3000 6092 3012
rect 6144 3000 6150 3052
rect 8202 3000 8208 3052
rect 8260 3040 8266 3052
rect 10594 3040 10600 3052
rect 8260 3012 10600 3040
rect 8260 3000 8266 3012
rect 10594 3000 10600 3012
rect 10652 3000 10658 3052
rect 11146 3000 11152 3052
rect 11204 3000 11210 3052
rect 11333 3043 11391 3049
rect 11333 3009 11345 3043
rect 11379 3040 11391 3043
rect 12342 3040 12348 3052
rect 11379 3012 12348 3040
rect 11379 3009 11391 3012
rect 11333 3003 11391 3009
rect 12342 3000 12348 3012
rect 12400 3000 12406 3052
rect 12526 3040 12532 3052
rect 12487 3012 12532 3040
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 12618 3000 12624 3052
rect 12676 3040 12682 3052
rect 14093 3043 14151 3049
rect 14093 3040 14105 3043
rect 12676 3012 14105 3040
rect 12676 3000 12682 3012
rect 14093 3009 14105 3012
rect 14139 3009 14151 3043
rect 14918 3040 14924 3052
rect 14879 3012 14924 3040
rect 14093 3003 14151 3009
rect 14918 3000 14924 3012
rect 14976 3000 14982 3052
rect 16482 3040 16488 3052
rect 16443 3012 16488 3040
rect 16482 3000 16488 3012
rect 16540 3000 16546 3052
rect 1489 2975 1547 2981
rect 1489 2941 1501 2975
rect 1535 2972 1547 2975
rect 2038 2972 2044 2984
rect 1535 2944 2044 2972
rect 1535 2941 1547 2944
rect 1489 2935 1547 2941
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 2409 2975 2467 2981
rect 2409 2941 2421 2975
rect 2455 2972 2467 2975
rect 3329 2975 3387 2981
rect 2455 2944 3096 2972
rect 2455 2941 2467 2944
rect 2409 2935 2467 2941
rect 1118 2864 1124 2916
rect 1176 2904 1182 2916
rect 1765 2907 1823 2913
rect 1765 2904 1777 2907
rect 1176 2876 1777 2904
rect 1176 2864 1182 2876
rect 1765 2873 1777 2876
rect 1811 2873 1823 2907
rect 1765 2867 1823 2873
rect 2130 2864 2136 2916
rect 2188 2904 2194 2916
rect 2685 2907 2743 2913
rect 2685 2904 2697 2907
rect 2188 2876 2697 2904
rect 2188 2864 2194 2876
rect 2685 2873 2697 2876
rect 2731 2873 2743 2907
rect 2685 2867 2743 2873
rect 3068 2836 3096 2944
rect 3329 2941 3341 2975
rect 3375 2972 3387 2975
rect 3418 2972 3424 2984
rect 3375 2944 3424 2972
rect 3375 2941 3387 2944
rect 3329 2935 3387 2941
rect 3418 2932 3424 2944
rect 3476 2932 3482 2984
rect 4246 2972 4252 2984
rect 4207 2944 4252 2972
rect 4246 2932 4252 2944
rect 4304 2932 4310 2984
rect 5261 2975 5319 2981
rect 5261 2941 5273 2975
rect 5307 2972 5319 2975
rect 5810 2972 5816 2984
rect 5307 2944 5816 2972
rect 5307 2941 5319 2944
rect 5261 2935 5319 2941
rect 5810 2932 5816 2944
rect 5868 2932 5874 2984
rect 5997 2975 6055 2981
rect 5997 2941 6009 2975
rect 6043 2972 6055 2975
rect 6546 2972 6552 2984
rect 6043 2944 6552 2972
rect 6043 2941 6055 2944
rect 5997 2935 6055 2941
rect 6546 2932 6552 2944
rect 6604 2932 6610 2984
rect 6730 2932 6736 2984
rect 6788 2972 6794 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6788 2944 6837 2972
rect 6788 2932 6794 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 7193 2975 7251 2981
rect 7193 2941 7205 2975
rect 7239 2972 7251 2975
rect 7282 2972 7288 2984
rect 7239 2944 7288 2972
rect 7239 2941 7251 2944
rect 7193 2935 7251 2941
rect 7282 2932 7288 2944
rect 7340 2932 7346 2984
rect 7466 2932 7472 2984
rect 7524 2972 7530 2984
rect 8056 2975 8114 2981
rect 8056 2972 8068 2975
rect 7524 2944 8068 2972
rect 7524 2932 7530 2944
rect 8056 2941 8068 2944
rect 8102 2941 8114 2975
rect 8056 2935 8114 2941
rect 3142 2864 3148 2916
rect 3200 2904 3206 2916
rect 3605 2907 3663 2913
rect 3605 2904 3617 2907
rect 3200 2876 3617 2904
rect 3200 2864 3206 2876
rect 3605 2873 3617 2876
rect 3651 2873 3663 2907
rect 7558 2904 7564 2916
rect 3605 2867 3663 2873
rect 3712 2876 7564 2904
rect 3712 2836 3740 2876
rect 7558 2864 7564 2876
rect 7616 2864 7622 2916
rect 8570 2904 8576 2916
rect 8036 2876 8576 2904
rect 3068 2808 3740 2836
rect 7285 2839 7343 2845
rect 7285 2805 7297 2839
rect 7331 2836 7343 2839
rect 8036 2836 8064 2876
rect 8570 2864 8576 2876
rect 8628 2864 8634 2916
rect 8754 2904 8760 2916
rect 8715 2876 8760 2904
rect 8754 2864 8760 2876
rect 8812 2864 8818 2916
rect 8849 2907 8907 2913
rect 8849 2873 8861 2907
rect 8895 2873 8907 2907
rect 8849 2867 8907 2873
rect 7331 2808 8064 2836
rect 8159 2839 8217 2845
rect 7331 2805 7343 2808
rect 7285 2799 7343 2805
rect 8159 2805 8171 2839
rect 8205 2836 8217 2839
rect 8864 2836 8892 2867
rect 9582 2864 9588 2916
rect 9640 2904 9646 2916
rect 9769 2907 9827 2913
rect 9769 2904 9781 2907
rect 9640 2876 9781 2904
rect 9640 2864 9646 2876
rect 9769 2873 9781 2876
rect 9815 2873 9827 2907
rect 10318 2904 10324 2916
rect 10279 2876 10324 2904
rect 9769 2867 9827 2873
rect 10318 2864 10324 2876
rect 10376 2864 10382 2916
rect 10410 2864 10416 2916
rect 10468 2904 10474 2916
rect 11164 2904 11192 3000
rect 16574 2932 16580 2984
rect 16632 2972 16638 2984
rect 17221 2975 17279 2981
rect 17221 2972 17233 2975
rect 16632 2944 17233 2972
rect 16632 2932 16638 2944
rect 17221 2941 17233 2944
rect 17267 2941 17279 2975
rect 17221 2935 17279 2941
rect 12621 2907 12679 2913
rect 12621 2904 12633 2907
rect 10468 2876 10513 2904
rect 11164 2876 12633 2904
rect 10468 2864 10474 2876
rect 12621 2873 12633 2876
rect 12667 2873 12679 2907
rect 13538 2904 13544 2916
rect 13499 2876 13544 2904
rect 12621 2867 12679 2873
rect 13538 2864 13544 2876
rect 13596 2864 13602 2916
rect 14185 2907 14243 2913
rect 14185 2873 14197 2907
rect 14231 2873 14243 2907
rect 14185 2867 14243 2873
rect 8205 2808 8892 2836
rect 8205 2805 8217 2808
rect 8159 2799 8217 2805
rect 9214 2796 9220 2848
rect 9272 2836 9278 2848
rect 11146 2836 11152 2848
rect 9272 2808 11152 2836
rect 9272 2796 9278 2808
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 12710 2796 12716 2848
rect 12768 2836 12774 2848
rect 14200 2836 14228 2867
rect 14550 2864 14556 2916
rect 14608 2904 14614 2916
rect 15657 2907 15715 2913
rect 15657 2904 15669 2907
rect 14608 2876 15669 2904
rect 14608 2864 14614 2876
rect 15657 2873 15669 2876
rect 15703 2873 15715 2907
rect 15657 2867 15715 2873
rect 15746 2864 15752 2916
rect 15804 2904 15810 2916
rect 15804 2876 15849 2904
rect 15804 2864 15810 2876
rect 12768 2808 14228 2836
rect 12768 2796 12774 2808
rect 1104 2746 18860 2768
rect 1104 2694 6912 2746
rect 6964 2694 6976 2746
rect 7028 2694 7040 2746
rect 7092 2694 7104 2746
rect 7156 2694 12843 2746
rect 12895 2694 12907 2746
rect 12959 2694 12971 2746
rect 13023 2694 13035 2746
rect 13087 2694 18860 2746
rect 1104 2672 18860 2694
rect 2685 2635 2743 2641
rect 2685 2601 2697 2635
rect 2731 2632 2743 2635
rect 2958 2632 2964 2644
rect 2731 2604 2964 2632
rect 2731 2601 2743 2604
rect 2685 2595 2743 2601
rect 2958 2592 2964 2604
rect 3016 2592 3022 2644
rect 3418 2632 3424 2644
rect 3379 2604 3424 2632
rect 3418 2592 3424 2604
rect 3476 2592 3482 2644
rect 6273 2635 6331 2641
rect 6273 2601 6285 2635
rect 6319 2632 6331 2635
rect 8202 2632 8208 2644
rect 6319 2604 8208 2632
rect 6319 2601 6331 2604
rect 6273 2595 6331 2601
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 8754 2592 8760 2644
rect 8812 2632 8818 2644
rect 9214 2632 9220 2644
rect 8812 2604 9220 2632
rect 8812 2592 8818 2604
rect 9214 2592 9220 2604
rect 9272 2592 9278 2644
rect 16206 2632 16212 2644
rect 11164 2604 13952 2632
rect 16167 2604 16212 2632
rect 5534 2564 5540 2576
rect 4080 2536 5540 2564
rect 1578 2496 1584 2508
rect 1539 2468 1584 2496
rect 1578 2456 1584 2468
rect 1636 2456 1642 2508
rect 2498 2496 2504 2508
rect 2459 2468 2504 2496
rect 2498 2456 2504 2468
rect 2556 2456 2562 2508
rect 3050 2456 3056 2508
rect 3108 2496 3114 2508
rect 4080 2505 4108 2536
rect 5534 2524 5540 2536
rect 5592 2524 5598 2576
rect 8938 2564 8944 2576
rect 6104 2536 8944 2564
rect 3237 2499 3295 2505
rect 3237 2496 3249 2499
rect 3108 2468 3249 2496
rect 3108 2456 3114 2468
rect 3237 2465 3249 2468
rect 3283 2465 3295 2499
rect 3237 2459 3295 2465
rect 4065 2499 4123 2505
rect 4065 2465 4077 2499
rect 4111 2465 4123 2499
rect 4798 2496 4804 2508
rect 4759 2468 4804 2496
rect 4065 2459 4123 2465
rect 4798 2456 4804 2468
rect 4856 2456 4862 2508
rect 6104 2505 6132 2536
rect 8938 2524 8944 2536
rect 8996 2524 9002 2576
rect 10226 2564 10232 2576
rect 10187 2536 10232 2564
rect 10226 2524 10232 2536
rect 10284 2524 10290 2576
rect 10321 2567 10379 2573
rect 10321 2533 10333 2567
rect 10367 2564 10379 2567
rect 10502 2564 10508 2576
rect 10367 2536 10508 2564
rect 10367 2533 10379 2536
rect 10321 2527 10379 2533
rect 10502 2524 10508 2536
rect 10560 2524 10566 2576
rect 10686 2524 10692 2576
rect 10744 2564 10750 2576
rect 11164 2564 11192 2604
rect 10744 2536 11192 2564
rect 11241 2567 11299 2573
rect 10744 2524 10750 2536
rect 11241 2533 11253 2567
rect 11287 2564 11299 2567
rect 11514 2564 11520 2576
rect 11287 2536 11520 2564
rect 11287 2533 11299 2536
rect 11241 2527 11299 2533
rect 11514 2524 11520 2536
rect 11572 2524 11578 2576
rect 13924 2573 13952 2604
rect 16206 2592 16212 2604
rect 16264 2592 16270 2644
rect 16942 2632 16948 2644
rect 16903 2604 16948 2632
rect 16942 2592 16948 2604
rect 17000 2592 17006 2644
rect 17678 2632 17684 2644
rect 17639 2604 17684 2632
rect 17678 2592 17684 2604
rect 17736 2592 17742 2644
rect 13909 2567 13967 2573
rect 11624 2536 13032 2564
rect 6089 2499 6147 2505
rect 6089 2465 6101 2499
rect 6135 2465 6147 2499
rect 6089 2459 6147 2465
rect 7285 2499 7343 2505
rect 7285 2465 7297 2499
rect 7331 2496 7343 2499
rect 7374 2496 7380 2508
rect 7331 2468 7380 2496
rect 7331 2465 7343 2468
rect 7285 2459 7343 2465
rect 7374 2456 7380 2468
rect 7432 2456 7438 2508
rect 7653 2499 7711 2505
rect 7653 2465 7665 2499
rect 7699 2496 7711 2499
rect 8294 2496 8300 2508
rect 7699 2468 8300 2496
rect 7699 2465 7711 2468
rect 7653 2459 7711 2465
rect 8294 2456 8300 2468
rect 8352 2456 8358 2508
rect 8478 2496 8484 2508
rect 8439 2468 8484 2496
rect 8478 2456 8484 2468
rect 8536 2456 8542 2508
rect 11330 2456 11336 2508
rect 11388 2496 11394 2508
rect 11624 2496 11652 2536
rect 11790 2496 11796 2508
rect 11388 2468 11652 2496
rect 11751 2468 11796 2496
rect 11388 2456 11394 2468
rect 11790 2456 11796 2468
rect 11848 2456 11854 2508
rect 13004 2505 13032 2536
rect 13909 2533 13921 2567
rect 13955 2533 13967 2567
rect 14826 2564 14832 2576
rect 14787 2536 14832 2564
rect 13909 2527 13967 2533
rect 14826 2524 14832 2536
rect 14884 2524 14890 2576
rect 12989 2499 13047 2505
rect 12989 2465 13001 2499
rect 13035 2465 13047 2499
rect 16022 2496 16028 2508
rect 15983 2468 16028 2496
rect 12989 2459 13047 2465
rect 16022 2456 16028 2468
rect 16080 2456 16086 2508
rect 16758 2496 16764 2508
rect 16719 2468 16764 2496
rect 16758 2456 16764 2468
rect 16816 2456 16822 2508
rect 17494 2496 17500 2508
rect 17455 2468 17500 2496
rect 17494 2456 17500 2468
rect 17552 2456 17558 2508
rect 658 2388 664 2440
rect 716 2428 722 2440
rect 1765 2431 1823 2437
rect 1765 2428 1777 2431
rect 716 2400 1777 2428
rect 716 2388 722 2400
rect 1765 2397 1777 2400
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 11054 2388 11060 2440
rect 11112 2428 11118 2440
rect 13817 2431 13875 2437
rect 13817 2428 13829 2431
rect 11112 2400 13829 2428
rect 11112 2388 11118 2400
rect 13817 2397 13829 2400
rect 13863 2397 13875 2431
rect 13817 2391 13875 2397
rect 6730 2320 6736 2372
rect 6788 2360 6794 2372
rect 6917 2363 6975 2369
rect 6917 2360 6929 2363
rect 6788 2332 6929 2360
rect 6788 2320 6794 2332
rect 6917 2329 6929 2332
rect 6963 2360 6975 2363
rect 8113 2363 8171 2369
rect 8113 2360 8125 2363
rect 6963 2332 8125 2360
rect 6963 2329 6975 2332
rect 6917 2323 6975 2329
rect 8113 2329 8125 2332
rect 8159 2360 8171 2363
rect 8386 2360 8392 2372
rect 8159 2332 8392 2360
rect 8159 2329 8171 2332
rect 8113 2323 8171 2329
rect 8386 2320 8392 2332
rect 8444 2320 8450 2372
rect 3510 2252 3516 2304
rect 3568 2292 3574 2304
rect 4249 2295 4307 2301
rect 4249 2292 4261 2295
rect 3568 2264 4261 2292
rect 3568 2252 3574 2264
rect 4249 2261 4261 2264
rect 4295 2261 4307 2295
rect 4982 2292 4988 2304
rect 4943 2264 4988 2292
rect 4249 2255 4307 2261
rect 4982 2252 4988 2264
rect 5040 2252 5046 2304
rect 8573 2295 8631 2301
rect 8573 2261 8585 2295
rect 8619 2292 8631 2295
rect 10686 2292 10692 2304
rect 8619 2264 10692 2292
rect 8619 2261 8631 2264
rect 8573 2255 8631 2261
rect 10686 2252 10692 2264
rect 10744 2252 10750 2304
rect 11977 2295 12035 2301
rect 11977 2261 11989 2295
rect 12023 2292 12035 2295
rect 13078 2292 13084 2304
rect 12023 2264 13084 2292
rect 12023 2261 12035 2264
rect 11977 2255 12035 2261
rect 13078 2252 13084 2264
rect 13136 2252 13142 2304
rect 13173 2295 13231 2301
rect 13173 2261 13185 2295
rect 13219 2292 13231 2295
rect 16206 2292 16212 2304
rect 13219 2264 16212 2292
rect 13219 2261 13231 2264
rect 13173 2255 13231 2261
rect 16206 2252 16212 2264
rect 16264 2252 16270 2304
rect 1104 2202 18860 2224
rect 1104 2150 3947 2202
rect 3999 2150 4011 2202
rect 4063 2150 4075 2202
rect 4127 2150 4139 2202
rect 4191 2150 9878 2202
rect 9930 2150 9942 2202
rect 9994 2150 10006 2202
rect 10058 2150 10070 2202
rect 10122 2150 15808 2202
rect 15860 2150 15872 2202
rect 15924 2150 15936 2202
rect 15988 2150 16000 2202
rect 16052 2150 18860 2202
rect 1104 2128 18860 2150
rect 13078 2048 13084 2100
rect 13136 2088 13142 2100
rect 15010 2088 15016 2100
rect 13136 2060 15016 2088
rect 13136 2048 13142 2060
rect 15010 2048 15016 2060
rect 15068 2048 15074 2100
rect 5166 1300 5172 1352
rect 5224 1340 5230 1352
rect 8018 1340 8024 1352
rect 5224 1312 8024 1340
rect 5224 1300 5230 1312
rect 8018 1300 8024 1312
rect 8076 1300 8082 1352
rect 7098 1096 7104 1148
rect 7156 1136 7162 1148
rect 7926 1136 7932 1148
rect 7156 1108 7932 1136
rect 7156 1096 7162 1108
rect 7926 1096 7932 1108
rect 7984 1096 7990 1148
rect 3694 688 3700 740
rect 3752 728 3758 740
rect 4982 728 4988 740
rect 3752 700 4988 728
rect 3752 688 3758 700
rect 4982 688 4988 700
rect 5040 688 5046 740
<< via1 >>
rect 3608 15240 3660 15292
rect 5632 15240 5684 15292
rect 12072 15172 12124 15224
rect 15936 15172 15988 15224
rect 3516 14764 3568 14816
rect 8760 14764 8812 14816
rect 6912 14662 6964 14714
rect 6976 14662 7028 14714
rect 7040 14662 7092 14714
rect 7104 14662 7156 14714
rect 12843 14662 12895 14714
rect 12907 14662 12959 14714
rect 12971 14662 13023 14714
rect 13035 14662 13087 14714
rect 1584 14560 1636 14612
rect 2228 14560 2280 14612
rect 14924 14492 14976 14544
rect 9588 14424 9640 14476
rect 17040 14492 17092 14544
rect 15476 14467 15528 14476
rect 15476 14433 15485 14467
rect 15485 14433 15519 14467
rect 15519 14433 15528 14467
rect 15476 14424 15528 14433
rect 15752 14424 15804 14476
rect 13728 14356 13780 14408
rect 1676 14220 1728 14272
rect 3424 14263 3476 14272
rect 3424 14229 3433 14263
rect 3433 14229 3467 14263
rect 3467 14229 3476 14263
rect 3424 14220 3476 14229
rect 15568 14220 15620 14272
rect 15660 14263 15712 14272
rect 15660 14229 15669 14263
rect 15669 14229 15703 14263
rect 15703 14229 15712 14263
rect 15660 14220 15712 14229
rect 3947 14118 3999 14170
rect 4011 14118 4063 14170
rect 4075 14118 4127 14170
rect 4139 14118 4191 14170
rect 9878 14118 9930 14170
rect 9942 14118 9994 14170
rect 10006 14118 10058 14170
rect 10070 14118 10122 14170
rect 15808 14118 15860 14170
rect 15872 14118 15924 14170
rect 15936 14118 15988 14170
rect 16000 14118 16052 14170
rect 2872 14016 2924 14068
rect 3516 14016 3568 14068
rect 5540 14016 5592 14068
rect 6920 14016 6972 14068
rect 2044 13948 2096 14000
rect 4620 13948 4672 14000
rect 13544 13948 13596 14000
rect 1492 13812 1544 13864
rect 13360 13880 13412 13932
rect 6092 13812 6144 13864
rect 296 13744 348 13796
rect 3424 13744 3476 13796
rect 5908 13744 5960 13796
rect 14372 13812 14424 13864
rect 15108 13812 15160 13864
rect 16396 13812 16448 13864
rect 7380 13744 7432 13796
rect 9036 13744 9088 13796
rect 9312 13744 9364 13796
rect 10324 13744 10376 13796
rect 11336 13744 11388 13796
rect 11888 13744 11940 13796
rect 11980 13744 12032 13796
rect 1952 13719 2004 13728
rect 1952 13685 1961 13719
rect 1961 13685 1995 13719
rect 1995 13685 2004 13719
rect 1952 13676 2004 13685
rect 6184 13719 6236 13728
rect 6184 13685 6193 13719
rect 6193 13685 6227 13719
rect 6227 13685 6236 13719
rect 6184 13676 6236 13685
rect 11244 13676 11296 13728
rect 11796 13676 11848 13728
rect 15660 13744 15712 13796
rect 13636 13719 13688 13728
rect 13636 13685 13645 13719
rect 13645 13685 13679 13719
rect 13679 13685 13688 13719
rect 13636 13676 13688 13685
rect 15292 13676 15344 13728
rect 6912 13574 6964 13626
rect 6976 13574 7028 13626
rect 7040 13574 7092 13626
rect 7104 13574 7156 13626
rect 12843 13574 12895 13626
rect 12907 13574 12959 13626
rect 12971 13574 13023 13626
rect 13035 13574 13087 13626
rect 940 13472 992 13524
rect 4804 13472 4856 13524
rect 11980 13472 12032 13524
rect 1584 13404 1636 13456
rect 2780 13311 2832 13320
rect 2780 13277 2789 13311
rect 2789 13277 2823 13311
rect 2823 13277 2832 13311
rect 2780 13268 2832 13277
rect 3240 13268 3292 13320
rect 4252 13404 4304 13456
rect 13544 13472 13596 13524
rect 14924 13472 14976 13524
rect 18972 13472 19024 13524
rect 15108 13336 15160 13388
rect 11980 13268 12032 13320
rect 13544 13268 13596 13320
rect 13728 13268 13780 13320
rect 18328 13404 18380 13456
rect 17776 13336 17828 13388
rect 17592 13268 17644 13320
rect 1860 13132 1912 13184
rect 4528 13200 4580 13252
rect 11428 13200 11480 13252
rect 17684 13200 17736 13252
rect 8116 13132 8168 13184
rect 10232 13132 10284 13184
rect 12624 13132 12676 13184
rect 13820 13132 13872 13184
rect 14648 13132 14700 13184
rect 15200 13132 15252 13184
rect 18604 13132 18656 13184
rect 3947 13030 3999 13082
rect 4011 13030 4063 13082
rect 4075 13030 4127 13082
rect 4139 13030 4191 13082
rect 9878 13030 9930 13082
rect 9942 13030 9994 13082
rect 10006 13030 10058 13082
rect 10070 13030 10122 13082
rect 15808 13030 15860 13082
rect 15872 13030 15924 13082
rect 15936 13030 15988 13082
rect 16000 13030 16052 13082
rect 1952 12928 2004 12980
rect 5448 12928 5500 12980
rect 15292 12928 15344 12980
rect 2136 12835 2188 12844
rect 2136 12801 2145 12835
rect 2145 12801 2179 12835
rect 2179 12801 2188 12835
rect 4528 12835 4580 12844
rect 2136 12792 2188 12801
rect 1860 12767 1912 12776
rect 1860 12733 1869 12767
rect 1869 12733 1903 12767
rect 1903 12733 1912 12767
rect 1860 12724 1912 12733
rect 1952 12631 2004 12640
rect 1952 12597 1961 12631
rect 1961 12597 1995 12631
rect 1995 12597 2004 12631
rect 4528 12801 4537 12835
rect 4537 12801 4571 12835
rect 4571 12801 4580 12835
rect 4528 12792 4580 12801
rect 6092 12835 6144 12844
rect 6092 12801 6101 12835
rect 6101 12801 6135 12835
rect 6135 12801 6144 12835
rect 6092 12792 6144 12801
rect 8484 12835 8536 12844
rect 8484 12801 8493 12835
rect 8493 12801 8527 12835
rect 8527 12801 8536 12835
rect 8484 12792 8536 12801
rect 8760 12792 8812 12844
rect 13636 12860 13688 12912
rect 13728 12860 13780 12912
rect 19616 12860 19668 12912
rect 13360 12792 13412 12844
rect 3516 12724 3568 12776
rect 4712 12724 4764 12776
rect 8024 12767 8076 12776
rect 8024 12733 8033 12767
rect 8033 12733 8067 12767
rect 8067 12733 8076 12767
rect 8024 12724 8076 12733
rect 8116 12724 8168 12776
rect 2780 12656 2832 12708
rect 3056 12656 3108 12708
rect 10600 12724 10652 12776
rect 11428 12656 11480 12708
rect 11704 12656 11756 12708
rect 13268 12724 13320 12776
rect 15476 12724 15528 12776
rect 16212 12767 16264 12776
rect 16212 12733 16221 12767
rect 16221 12733 16255 12767
rect 16255 12733 16264 12767
rect 16212 12724 16264 12733
rect 16580 12724 16632 12776
rect 1952 12588 2004 12597
rect 4344 12588 4396 12640
rect 5724 12588 5776 12640
rect 5816 12588 5868 12640
rect 6000 12631 6052 12640
rect 6000 12597 6009 12631
rect 6009 12597 6043 12631
rect 6043 12597 6052 12631
rect 6000 12588 6052 12597
rect 7288 12588 7340 12640
rect 13360 12588 13412 12640
rect 15384 12588 15436 12640
rect 17224 12588 17276 12640
rect 18144 12588 18196 12640
rect 6912 12486 6964 12538
rect 6976 12486 7028 12538
rect 7040 12486 7092 12538
rect 7104 12486 7156 12538
rect 12843 12486 12895 12538
rect 12907 12486 12959 12538
rect 12971 12486 13023 12538
rect 13035 12486 13087 12538
rect 1952 12384 2004 12436
rect 2964 12384 3016 12436
rect 4620 12316 4672 12368
rect 6092 12384 6144 12436
rect 6552 12384 6604 12436
rect 11520 12384 11572 12436
rect 6276 12316 6328 12368
rect 2412 12248 2464 12300
rect 4252 12248 4304 12300
rect 4528 12291 4580 12300
rect 4528 12257 4537 12291
rect 4537 12257 4571 12291
rect 4571 12257 4580 12291
rect 4528 12248 4580 12257
rect 9128 12316 9180 12368
rect 2320 12180 2372 12232
rect 2780 12223 2832 12232
rect 2780 12189 2789 12223
rect 2789 12189 2823 12223
rect 2823 12189 2832 12223
rect 2780 12180 2832 12189
rect 3056 12180 3108 12232
rect 3424 12180 3476 12232
rect 4068 12180 4120 12232
rect 6644 12291 6696 12300
rect 6644 12257 6678 12291
rect 6678 12257 6696 12291
rect 6644 12248 6696 12257
rect 7656 12248 7708 12300
rect 9404 12248 9456 12300
rect 11612 12248 11664 12300
rect 12532 12248 12584 12300
rect 14740 12248 14792 12300
rect 17132 12291 17184 12300
rect 6092 12180 6144 12232
rect 6368 12223 6420 12232
rect 6368 12189 6377 12223
rect 6377 12189 6411 12223
rect 6411 12189 6420 12223
rect 6368 12180 6420 12189
rect 8668 12223 8720 12232
rect 8668 12189 8677 12223
rect 8677 12189 8711 12223
rect 8711 12189 8720 12223
rect 8668 12180 8720 12189
rect 8760 12223 8812 12232
rect 8760 12189 8769 12223
rect 8769 12189 8803 12223
rect 8803 12189 8812 12223
rect 8760 12180 8812 12189
rect 9312 12180 9364 12232
rect 15292 12180 15344 12232
rect 3608 12112 3660 12164
rect 3884 12112 3936 12164
rect 9404 12112 9456 12164
rect 13912 12112 13964 12164
rect 14004 12112 14056 12164
rect 17132 12257 17141 12291
rect 17141 12257 17175 12291
rect 17175 12257 17184 12291
rect 17132 12248 17184 12257
rect 17868 12291 17920 12300
rect 17868 12257 17877 12291
rect 17877 12257 17911 12291
rect 17911 12257 17920 12291
rect 17868 12248 17920 12257
rect 19156 12112 19208 12164
rect 3056 12044 3108 12096
rect 3332 12044 3384 12096
rect 6000 12044 6052 12096
rect 6736 12044 6788 12096
rect 8116 12044 8168 12096
rect 12256 12044 12308 12096
rect 12716 12044 12768 12096
rect 14556 12044 14608 12096
rect 16120 12044 16172 12096
rect 17776 12044 17828 12096
rect 18052 12087 18104 12096
rect 18052 12053 18061 12087
rect 18061 12053 18095 12087
rect 18095 12053 18104 12087
rect 18052 12044 18104 12053
rect 3947 11942 3999 11994
rect 4011 11942 4063 11994
rect 4075 11942 4127 11994
rect 4139 11942 4191 11994
rect 9878 11942 9930 11994
rect 9942 11942 9994 11994
rect 10006 11942 10058 11994
rect 10070 11942 10122 11994
rect 15808 11942 15860 11994
rect 15872 11942 15924 11994
rect 15936 11942 15988 11994
rect 16000 11942 16052 11994
rect 4620 11840 4672 11892
rect 5816 11840 5868 11892
rect 2688 11772 2740 11824
rect 3148 11772 3200 11824
rect 3516 11772 3568 11824
rect 2780 11704 2832 11756
rect 5356 11704 5408 11756
rect 5816 11704 5868 11756
rect 6092 11704 6144 11756
rect 6736 11704 6788 11756
rect 1584 11679 1636 11688
rect 1584 11645 1593 11679
rect 1593 11645 1627 11679
rect 1627 11645 1636 11679
rect 1584 11636 1636 11645
rect 2964 11636 3016 11688
rect 4344 11636 4396 11688
rect 6368 11636 6420 11688
rect 8668 11840 8720 11892
rect 8852 11840 8904 11892
rect 13268 11840 13320 11892
rect 13544 11840 13596 11892
rect 13912 11840 13964 11892
rect 16764 11840 16816 11892
rect 16304 11772 16356 11824
rect 19616 11772 19668 11824
rect 9312 11747 9364 11756
rect 9312 11713 9321 11747
rect 9321 11713 9355 11747
rect 9355 11713 9364 11747
rect 9312 11704 9364 11713
rect 12348 11704 12400 11756
rect 13636 11747 13688 11756
rect 13636 11713 13645 11747
rect 13645 11713 13679 11747
rect 13679 11713 13688 11747
rect 13636 11704 13688 11713
rect 15660 11747 15712 11756
rect 15660 11713 15669 11747
rect 15669 11713 15703 11747
rect 15703 11713 15712 11747
rect 15660 11704 15712 11713
rect 16856 11704 16908 11756
rect 16488 11679 16540 11688
rect 2228 11568 2280 11620
rect 1768 11543 1820 11552
rect 1768 11509 1777 11543
rect 1777 11509 1811 11543
rect 1811 11509 1820 11543
rect 1768 11500 1820 11509
rect 1860 11500 1912 11552
rect 2780 11543 2832 11552
rect 2780 11509 2789 11543
rect 2789 11509 2823 11543
rect 2823 11509 2832 11543
rect 5632 11568 5684 11620
rect 2780 11500 2832 11509
rect 4436 11500 4488 11552
rect 5540 11543 5592 11552
rect 5540 11509 5549 11543
rect 5549 11509 5583 11543
rect 5583 11509 5592 11543
rect 5540 11500 5592 11509
rect 6736 11568 6788 11620
rect 13912 11568 13964 11620
rect 14096 11568 14148 11620
rect 16488 11645 16497 11679
rect 16497 11645 16531 11679
rect 16531 11645 16540 11679
rect 16488 11636 16540 11645
rect 16764 11636 16816 11688
rect 17960 11636 18012 11688
rect 16948 11568 17000 11620
rect 8208 11543 8260 11552
rect 8208 11509 8217 11543
rect 8217 11509 8251 11543
rect 8251 11509 8260 11543
rect 8208 11500 8260 11509
rect 8852 11500 8904 11552
rect 9220 11543 9272 11552
rect 9220 11509 9229 11543
rect 9229 11509 9263 11543
rect 9263 11509 9272 11543
rect 11152 11543 11204 11552
rect 9220 11500 9272 11509
rect 11152 11509 11161 11543
rect 11161 11509 11195 11543
rect 11195 11509 11204 11543
rect 11152 11500 11204 11509
rect 12164 11500 12216 11552
rect 12532 11500 12584 11552
rect 13176 11500 13228 11552
rect 13360 11543 13412 11552
rect 13360 11509 13369 11543
rect 13369 11509 13403 11543
rect 13403 11509 13412 11543
rect 13360 11500 13412 11509
rect 14280 11500 14332 11552
rect 15108 11543 15160 11552
rect 15108 11509 15117 11543
rect 15117 11509 15151 11543
rect 15151 11509 15160 11543
rect 15108 11500 15160 11509
rect 15752 11500 15804 11552
rect 17500 11500 17552 11552
rect 6912 11398 6964 11450
rect 6976 11398 7028 11450
rect 7040 11398 7092 11450
rect 7104 11398 7156 11450
rect 12843 11398 12895 11450
rect 12907 11398 12959 11450
rect 12971 11398 13023 11450
rect 13035 11398 13087 11450
rect 1492 11339 1544 11348
rect 1492 11305 1501 11339
rect 1501 11305 1535 11339
rect 1535 11305 1544 11339
rect 1492 11296 1544 11305
rect 1860 11339 1912 11348
rect 1860 11305 1869 11339
rect 1869 11305 1903 11339
rect 1903 11305 1912 11339
rect 1860 11296 1912 11305
rect 2780 11296 2832 11348
rect 5540 11296 5592 11348
rect 3148 11271 3200 11280
rect 3148 11237 3157 11271
rect 3157 11237 3191 11271
rect 3191 11237 3200 11271
rect 14372 11296 14424 11348
rect 15752 11339 15804 11348
rect 3148 11228 3200 11237
rect 1584 11092 1636 11144
rect 2136 11135 2188 11144
rect 2136 11101 2145 11135
rect 2145 11101 2179 11135
rect 2179 11101 2188 11135
rect 2136 11092 2188 11101
rect 5264 11160 5316 11212
rect 5908 11203 5960 11212
rect 5908 11169 5917 11203
rect 5917 11169 5951 11203
rect 5951 11169 5960 11203
rect 5908 11160 5960 11169
rect 3148 11092 3200 11144
rect 3332 11135 3384 11144
rect 3332 11101 3341 11135
rect 3341 11101 3375 11135
rect 3375 11101 3384 11135
rect 3332 11092 3384 11101
rect 4804 11135 4856 11144
rect 4804 11101 4813 11135
rect 4813 11101 4847 11135
rect 4847 11101 4856 11135
rect 4804 11092 4856 11101
rect 8208 11228 8260 11280
rect 8300 11228 8352 11280
rect 9220 11228 9272 11280
rect 12072 11228 12124 11280
rect 13360 11228 13412 11280
rect 15752 11305 15761 11339
rect 15761 11305 15795 11339
rect 15795 11305 15804 11339
rect 15752 11296 15804 11305
rect 16764 11296 16816 11348
rect 16948 11339 17000 11348
rect 16948 11305 16957 11339
rect 16957 11305 16991 11339
rect 16991 11305 17000 11339
rect 16948 11296 17000 11305
rect 17040 11228 17092 11280
rect 7196 11160 7248 11212
rect 7571 11203 7623 11212
rect 7571 11169 7580 11203
rect 7580 11169 7614 11203
rect 7614 11169 7623 11203
rect 7571 11160 7623 11169
rect 10692 11160 10744 11212
rect 10876 11203 10928 11212
rect 10876 11169 10910 11203
rect 10910 11169 10928 11203
rect 10876 11160 10928 11169
rect 13636 11160 13688 11212
rect 14832 11160 14884 11212
rect 16396 11160 16448 11212
rect 17316 11203 17368 11212
rect 17316 11169 17325 11203
rect 17325 11169 17359 11203
rect 17359 11169 17368 11203
rect 17316 11160 17368 11169
rect 10232 11092 10284 11144
rect 11704 11092 11756 11144
rect 11888 11092 11940 11144
rect 2320 10956 2372 11008
rect 4344 10999 4396 11008
rect 4344 10965 4353 10999
rect 4353 10965 4387 10999
rect 4387 10965 4396 10999
rect 4344 10956 4396 10965
rect 5540 10999 5592 11008
rect 5540 10965 5549 10999
rect 5549 10965 5583 10999
rect 5583 10965 5592 10999
rect 5540 10956 5592 10965
rect 6000 11024 6052 11076
rect 6368 11024 6420 11076
rect 6644 11024 6696 11076
rect 8944 10999 8996 11008
rect 8944 10965 8953 10999
rect 8953 10965 8987 10999
rect 8987 10965 8996 10999
rect 8944 10956 8996 10965
rect 10508 11024 10560 11076
rect 16672 11092 16724 11144
rect 17408 11135 17460 11144
rect 17408 11101 17417 11135
rect 17417 11101 17451 11135
rect 17451 11101 17460 11135
rect 17408 11092 17460 11101
rect 10416 10956 10468 11008
rect 10784 10956 10836 11008
rect 11612 10956 11664 11008
rect 12624 10956 12676 11008
rect 13820 10956 13872 11008
rect 16948 10956 17000 11008
rect 17868 10956 17920 11008
rect 3947 10854 3999 10906
rect 4011 10854 4063 10906
rect 4075 10854 4127 10906
rect 4139 10854 4191 10906
rect 9878 10854 9930 10906
rect 9942 10854 9994 10906
rect 10006 10854 10058 10906
rect 10070 10854 10122 10906
rect 15808 10854 15860 10906
rect 15872 10854 15924 10906
rect 15936 10854 15988 10906
rect 16000 10854 16052 10906
rect 2412 10591 2464 10600
rect 2412 10557 2421 10591
rect 2421 10557 2455 10591
rect 2455 10557 2464 10591
rect 2412 10548 2464 10557
rect 3148 10548 3200 10600
rect 3884 10548 3936 10600
rect 4436 10752 4488 10804
rect 5448 10752 5500 10804
rect 5908 10752 5960 10804
rect 7104 10752 7156 10804
rect 7748 10752 7800 10804
rect 4344 10616 4396 10668
rect 8392 10684 8444 10736
rect 6000 10616 6052 10668
rect 6736 10616 6788 10668
rect 10232 10752 10284 10804
rect 10784 10752 10836 10804
rect 10876 10684 10928 10736
rect 2780 10480 2832 10532
rect 2872 10480 2924 10532
rect 5540 10548 5592 10600
rect 5816 10591 5868 10600
rect 5816 10557 5825 10591
rect 5825 10557 5859 10591
rect 5859 10557 5868 10591
rect 5816 10548 5868 10557
rect 7104 10548 7156 10600
rect 7288 10548 7340 10600
rect 6092 10523 6144 10532
rect 3332 10412 3384 10464
rect 3516 10412 3568 10464
rect 4252 10412 4304 10464
rect 6092 10489 6101 10523
rect 6101 10489 6135 10523
rect 6135 10489 6144 10523
rect 6092 10480 6144 10489
rect 8668 10548 8720 10600
rect 10416 10616 10468 10668
rect 11244 10659 11296 10668
rect 11244 10625 11253 10659
rect 11253 10625 11287 10659
rect 11287 10625 11296 10659
rect 11244 10616 11296 10625
rect 12072 10684 12124 10736
rect 12348 10684 12400 10736
rect 13452 10616 13504 10668
rect 14188 10752 14240 10804
rect 17408 10752 17460 10804
rect 17408 10659 17460 10668
rect 17408 10625 17417 10659
rect 17417 10625 17451 10659
rect 17451 10625 17460 10659
rect 17408 10616 17460 10625
rect 12624 10548 12676 10600
rect 11612 10480 11664 10532
rect 11704 10480 11756 10532
rect 16948 10548 17000 10600
rect 15660 10480 15712 10532
rect 15844 10480 15896 10532
rect 18328 10548 18380 10600
rect 6276 10412 6328 10464
rect 7840 10412 7892 10464
rect 10416 10412 10468 10464
rect 10784 10455 10836 10464
rect 10784 10421 10793 10455
rect 10793 10421 10827 10455
rect 10827 10421 10836 10455
rect 10784 10412 10836 10421
rect 11060 10412 11112 10464
rect 12072 10412 12124 10464
rect 12624 10412 12676 10464
rect 13452 10412 13504 10464
rect 13636 10412 13688 10464
rect 15476 10412 15528 10464
rect 6912 10310 6964 10362
rect 6976 10310 7028 10362
rect 7040 10310 7092 10362
rect 7104 10310 7156 10362
rect 12843 10310 12895 10362
rect 12907 10310 12959 10362
rect 12971 10310 13023 10362
rect 13035 10310 13087 10362
rect 1584 10251 1636 10260
rect 1584 10217 1593 10251
rect 1593 10217 1627 10251
rect 1627 10217 1636 10251
rect 1584 10208 1636 10217
rect 4804 10208 4856 10260
rect 5816 10208 5868 10260
rect 12624 10251 12676 10260
rect 12624 10217 12633 10251
rect 12633 10217 12667 10251
rect 12667 10217 12676 10251
rect 12624 10208 12676 10217
rect 13452 10251 13504 10260
rect 13452 10217 13461 10251
rect 13461 10217 13495 10251
rect 13495 10217 13504 10251
rect 13452 10208 13504 10217
rect 14188 10208 14240 10260
rect 2412 10140 2464 10192
rect 2964 10140 3016 10192
rect 7288 10140 7340 10192
rect 8392 10140 8444 10192
rect 8944 10140 8996 10192
rect 10784 10140 10836 10192
rect 12808 10140 12860 10192
rect 15292 10140 15344 10192
rect 3056 10072 3108 10124
rect 4436 10115 4488 10124
rect 2596 10004 2648 10056
rect 3332 10047 3384 10056
rect 3332 10013 3341 10047
rect 3341 10013 3375 10047
rect 3375 10013 3384 10047
rect 3332 10004 3384 10013
rect 3516 9936 3568 9988
rect 2872 9868 2924 9920
rect 4436 10081 4445 10115
rect 4445 10081 4479 10115
rect 4479 10081 4488 10115
rect 4436 10072 4488 10081
rect 6276 10072 6328 10124
rect 7472 10072 7524 10124
rect 10140 10072 10192 10124
rect 10232 10072 10284 10124
rect 10600 10072 10652 10124
rect 11060 10072 11112 10124
rect 15016 10072 15068 10124
rect 17316 10208 17368 10260
rect 17592 10251 17644 10260
rect 17592 10217 17601 10251
rect 17601 10217 17635 10251
rect 17635 10217 17644 10251
rect 17592 10208 17644 10217
rect 4528 10047 4580 10056
rect 4528 10013 4537 10047
rect 4537 10013 4571 10047
rect 4571 10013 4580 10047
rect 4528 10004 4580 10013
rect 4712 10047 4764 10056
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 4712 10004 4764 10013
rect 5816 10047 5868 10056
rect 5816 10013 5825 10047
rect 5825 10013 5859 10047
rect 5859 10013 5868 10047
rect 5816 10004 5868 10013
rect 6000 10047 6052 10056
rect 6000 10013 6009 10047
rect 6009 10013 6043 10047
rect 6043 10013 6052 10047
rect 6000 10004 6052 10013
rect 6736 10047 6788 10056
rect 6736 10013 6745 10047
rect 6745 10013 6779 10047
rect 6779 10013 6788 10047
rect 6736 10004 6788 10013
rect 7564 10047 7616 10056
rect 7564 10013 7573 10047
rect 7573 10013 7607 10047
rect 7607 10013 7616 10047
rect 7564 10004 7616 10013
rect 6920 9936 6972 9988
rect 9312 9936 9364 9988
rect 9404 9936 9456 9988
rect 9772 9936 9824 9988
rect 10416 10047 10468 10056
rect 10416 10013 10425 10047
rect 10425 10013 10459 10047
rect 10459 10013 10468 10047
rect 11612 10047 11664 10056
rect 10416 10004 10468 10013
rect 11612 10013 11621 10047
rect 11621 10013 11655 10047
rect 11655 10013 11664 10047
rect 11612 10004 11664 10013
rect 12716 10047 12768 10056
rect 12716 10013 12725 10047
rect 12725 10013 12759 10047
rect 12759 10013 12768 10047
rect 12716 10004 12768 10013
rect 12808 10047 12860 10056
rect 12808 10013 12817 10047
rect 12817 10013 12851 10047
rect 12851 10013 12860 10047
rect 12808 10004 12860 10013
rect 15844 10140 15896 10192
rect 16580 10072 16632 10124
rect 13636 9936 13688 9988
rect 15292 9936 15344 9988
rect 6736 9868 6788 9920
rect 9496 9868 9548 9920
rect 15108 9868 15160 9920
rect 16672 9868 16724 9920
rect 17408 10072 17460 10124
rect 17592 10004 17644 10056
rect 18420 10208 18472 10260
rect 3947 9766 3999 9818
rect 4011 9766 4063 9818
rect 4075 9766 4127 9818
rect 4139 9766 4191 9818
rect 9878 9766 9930 9818
rect 9942 9766 9994 9818
rect 10006 9766 10058 9818
rect 10070 9766 10122 9818
rect 15808 9766 15860 9818
rect 15872 9766 15924 9818
rect 15936 9766 15988 9818
rect 16000 9766 16052 9818
rect 3056 9664 3108 9716
rect 3332 9596 3384 9648
rect 2964 9528 3016 9580
rect 5448 9664 5500 9716
rect 11704 9664 11756 9716
rect 12716 9664 12768 9716
rect 5264 9639 5316 9648
rect 5264 9605 5273 9639
rect 5273 9605 5307 9639
rect 5307 9605 5316 9639
rect 5264 9596 5316 9605
rect 8760 9596 8812 9648
rect 9128 9596 9180 9648
rect 5724 9571 5776 9580
rect 1584 9460 1636 9512
rect 4068 9460 4120 9512
rect 5724 9537 5733 9571
rect 5733 9537 5767 9571
rect 5767 9537 5776 9571
rect 5724 9528 5776 9537
rect 6000 9528 6052 9580
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 9312 9571 9364 9580
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 9496 9528 9548 9580
rect 10600 9528 10652 9580
rect 11060 9596 11112 9648
rect 15292 9664 15344 9716
rect 15660 9596 15712 9648
rect 13820 9528 13872 9580
rect 14188 9571 14240 9580
rect 14188 9537 14197 9571
rect 14197 9537 14231 9571
rect 14231 9537 14240 9571
rect 14188 9528 14240 9537
rect 16856 9528 16908 9580
rect 6276 9460 6328 9512
rect 2964 9392 3016 9444
rect 4160 9435 4212 9444
rect 4160 9401 4169 9435
rect 4169 9401 4203 9435
rect 4203 9401 4212 9435
rect 4160 9392 4212 9401
rect 5632 9435 5684 9444
rect 5632 9401 5641 9435
rect 5641 9401 5675 9435
rect 5675 9401 5684 9435
rect 8208 9460 8260 9512
rect 10048 9460 10100 9512
rect 11152 9503 11204 9512
rect 11152 9469 11161 9503
rect 11161 9469 11195 9503
rect 11195 9469 11204 9503
rect 11152 9460 11204 9469
rect 11980 9460 12032 9512
rect 13176 9460 13228 9512
rect 13360 9460 13412 9512
rect 17224 9528 17276 9580
rect 5632 9392 5684 9401
rect 2688 9324 2740 9376
rect 3056 9324 3108 9376
rect 4804 9324 4856 9376
rect 5448 9324 5500 9376
rect 6276 9324 6328 9376
rect 6460 9367 6512 9376
rect 6460 9333 6469 9367
rect 6469 9333 6503 9367
rect 6503 9333 6512 9367
rect 6460 9324 6512 9333
rect 7932 9324 7984 9376
rect 8760 9367 8812 9376
rect 8760 9333 8769 9367
rect 8769 9333 8803 9367
rect 8803 9333 8812 9367
rect 8760 9324 8812 9333
rect 8852 9324 8904 9376
rect 9680 9324 9732 9376
rect 10048 9324 10100 9376
rect 10324 9324 10376 9376
rect 12164 9392 12216 9444
rect 16672 9392 16724 9444
rect 11244 9324 11296 9376
rect 13176 9324 13228 9376
rect 13820 9324 13872 9376
rect 14372 9324 14424 9376
rect 15292 9324 15344 9376
rect 16212 9367 16264 9376
rect 16212 9333 16221 9367
rect 16221 9333 16255 9367
rect 16255 9333 16264 9367
rect 16212 9324 16264 9333
rect 16764 9367 16816 9376
rect 16764 9333 16773 9367
rect 16773 9333 16807 9367
rect 16807 9333 16816 9367
rect 16764 9324 16816 9333
rect 16856 9324 16908 9376
rect 6912 9222 6964 9274
rect 6976 9222 7028 9274
rect 7040 9222 7092 9274
rect 7104 9222 7156 9274
rect 12843 9222 12895 9274
rect 12907 9222 12959 9274
rect 12971 9222 13023 9274
rect 13035 9222 13087 9274
rect 2964 9163 3016 9172
rect 2964 9129 2973 9163
rect 2973 9129 3007 9163
rect 3007 9129 3016 9163
rect 2964 9120 3016 9129
rect 5816 9120 5868 9172
rect 7288 9120 7340 9172
rect 7472 9163 7524 9172
rect 7472 9129 7481 9163
rect 7481 9129 7515 9163
rect 7515 9129 7524 9163
rect 7472 9120 7524 9129
rect 7932 9120 7984 9172
rect 8852 9120 8904 9172
rect 10600 9120 10652 9172
rect 2688 9052 2740 9104
rect 3976 9052 4028 9104
rect 5724 9052 5776 9104
rect 6276 9095 6328 9104
rect 1584 9027 1636 9036
rect 1584 8993 1593 9027
rect 1593 8993 1627 9027
rect 1627 8993 1636 9027
rect 1584 8984 1636 8993
rect 4068 9027 4120 9036
rect 4068 8993 4077 9027
rect 4077 8993 4111 9027
rect 4111 8993 4120 9027
rect 4068 8984 4120 8993
rect 4896 8984 4948 9036
rect 6276 9061 6285 9095
rect 6285 9061 6319 9095
rect 6319 9061 6328 9095
rect 6276 9052 6328 9061
rect 9680 9052 9732 9104
rect 9772 9052 9824 9104
rect 13176 9120 13228 9172
rect 14188 9163 14240 9172
rect 14188 9129 14197 9163
rect 14197 9129 14231 9163
rect 14231 9129 14240 9163
rect 14188 9120 14240 9129
rect 16580 9120 16632 9172
rect 16764 9120 16816 9172
rect 13084 9052 13136 9104
rect 6552 8959 6604 8968
rect 6552 8925 6561 8959
rect 6561 8925 6595 8959
rect 6595 8925 6604 8959
rect 6552 8916 6604 8925
rect 9404 8916 9456 8968
rect 10692 8984 10744 9036
rect 10876 8984 10928 9036
rect 11704 8984 11756 9036
rect 12348 8984 12400 9036
rect 13360 8916 13412 8968
rect 13636 8959 13688 8968
rect 13636 8925 13645 8959
rect 13645 8925 13679 8959
rect 13679 8925 13688 8959
rect 13636 8916 13688 8925
rect 13912 9052 13964 9104
rect 16212 9052 16264 9104
rect 18512 9052 18564 9104
rect 16672 8984 16724 9036
rect 18328 8984 18380 9036
rect 13912 8916 13964 8968
rect 14188 8916 14240 8968
rect 16580 8916 16632 8968
rect 2688 8780 2740 8832
rect 4712 8780 4764 8832
rect 7932 8780 7984 8832
rect 8484 8780 8536 8832
rect 8852 8780 8904 8832
rect 9496 8780 9548 8832
rect 12900 8780 12952 8832
rect 15200 8780 15252 8832
rect 17040 8848 17092 8900
rect 17868 8780 17920 8832
rect 3947 8678 3999 8730
rect 4011 8678 4063 8730
rect 4075 8678 4127 8730
rect 4139 8678 4191 8730
rect 9878 8678 9930 8730
rect 9942 8678 9994 8730
rect 10006 8678 10058 8730
rect 10070 8678 10122 8730
rect 15808 8678 15860 8730
rect 15872 8678 15924 8730
rect 15936 8678 15988 8730
rect 16000 8678 16052 8730
rect 4528 8576 4580 8628
rect 5540 8576 5592 8628
rect 7196 8576 7248 8628
rect 8300 8576 8352 8628
rect 1584 8508 1636 8560
rect 2136 8508 2188 8560
rect 2964 8440 3016 8492
rect 2872 8372 2924 8424
rect 3056 8372 3108 8424
rect 2412 8304 2464 8356
rect 3608 8440 3660 8492
rect 4528 8440 4580 8492
rect 4896 8483 4948 8492
rect 4896 8449 4905 8483
rect 4905 8449 4939 8483
rect 4939 8449 4948 8483
rect 4896 8440 4948 8449
rect 6000 8483 6052 8492
rect 6000 8449 6009 8483
rect 6009 8449 6043 8483
rect 6043 8449 6052 8483
rect 6000 8440 6052 8449
rect 6736 8440 6788 8492
rect 4344 8372 4396 8424
rect 7288 8440 7340 8492
rect 7564 8440 7616 8492
rect 8208 8440 8260 8492
rect 2228 8279 2280 8288
rect 2228 8245 2237 8279
rect 2237 8245 2271 8279
rect 2271 8245 2280 8279
rect 2228 8236 2280 8245
rect 3056 8279 3108 8288
rect 3056 8245 3065 8279
rect 3065 8245 3099 8279
rect 3099 8245 3108 8279
rect 3056 8236 3108 8245
rect 5080 8236 5132 8288
rect 5632 8304 5684 8356
rect 7564 8304 7616 8356
rect 7472 8236 7524 8288
rect 7932 8304 7984 8356
rect 12348 8576 12400 8628
rect 13360 8576 13412 8628
rect 12072 8508 12124 8560
rect 15292 8576 15344 8628
rect 16396 8619 16448 8628
rect 16396 8585 16405 8619
rect 16405 8585 16439 8619
rect 16439 8585 16448 8619
rect 16396 8576 16448 8585
rect 17040 8576 17092 8628
rect 17960 8576 18012 8628
rect 12900 8483 12952 8492
rect 12900 8449 12909 8483
rect 12909 8449 12943 8483
rect 12943 8449 12952 8483
rect 12900 8440 12952 8449
rect 13084 8483 13136 8492
rect 13084 8449 13093 8483
rect 13093 8449 13127 8483
rect 13127 8449 13136 8483
rect 13084 8440 13136 8449
rect 9956 8372 10008 8424
rect 11244 8372 11296 8424
rect 14096 8508 14148 8560
rect 16672 8508 16724 8560
rect 17224 8508 17276 8560
rect 14188 8440 14240 8492
rect 16580 8440 16632 8492
rect 10692 8347 10744 8356
rect 10692 8313 10726 8347
rect 10726 8313 10744 8347
rect 12808 8347 12860 8356
rect 10692 8304 10744 8313
rect 12808 8313 12817 8347
rect 12817 8313 12851 8347
rect 12851 8313 12860 8347
rect 12808 8304 12860 8313
rect 15844 8372 15896 8424
rect 14096 8304 14148 8356
rect 15200 8304 15252 8356
rect 15752 8304 15804 8356
rect 16672 8304 16724 8356
rect 8852 8236 8904 8288
rect 11244 8236 11296 8288
rect 11704 8236 11756 8288
rect 12440 8279 12492 8288
rect 12440 8245 12449 8279
rect 12449 8245 12483 8279
rect 12483 8245 12492 8279
rect 16764 8279 16816 8288
rect 12440 8236 12492 8245
rect 16764 8245 16773 8279
rect 16773 8245 16807 8279
rect 16807 8245 16816 8279
rect 16764 8236 16816 8245
rect 6912 8134 6964 8186
rect 6976 8134 7028 8186
rect 7040 8134 7092 8186
rect 7104 8134 7156 8186
rect 12843 8134 12895 8186
rect 12907 8134 12959 8186
rect 12971 8134 13023 8186
rect 13035 8134 13087 8186
rect 3240 8032 3292 8084
rect 4620 8032 4672 8084
rect 4344 7964 4396 8016
rect 6276 7964 6328 8016
rect 7472 8032 7524 8084
rect 9404 8032 9456 8084
rect 12440 8032 12492 8084
rect 13820 8032 13872 8084
rect 16028 8032 16080 8084
rect 16764 8032 16816 8084
rect 6000 7939 6052 7948
rect 4528 7828 4580 7880
rect 4712 7828 4764 7880
rect 3700 7760 3752 7812
rect 6000 7905 6034 7939
rect 6034 7905 6052 7939
rect 6000 7896 6052 7905
rect 7196 7896 7248 7948
rect 8300 7896 8352 7948
rect 5356 7828 5408 7880
rect 2596 7692 2648 7744
rect 3148 7692 3200 7744
rect 5448 7760 5500 7812
rect 4712 7692 4764 7744
rect 4896 7692 4948 7744
rect 7564 7735 7616 7744
rect 7564 7701 7573 7735
rect 7573 7701 7607 7735
rect 7607 7701 7616 7735
rect 7564 7692 7616 7701
rect 8208 7828 8260 7880
rect 8484 7828 8536 7880
rect 10048 7964 10100 8016
rect 10876 7964 10928 8016
rect 11704 7964 11756 8016
rect 12164 8007 12216 8016
rect 12164 7973 12173 8007
rect 12173 7973 12207 8007
rect 12207 7973 12216 8007
rect 12164 7964 12216 7973
rect 8852 7896 8904 7948
rect 9128 7828 9180 7880
rect 9312 7760 9364 7812
rect 11244 7760 11296 7812
rect 8668 7692 8720 7744
rect 9496 7735 9548 7744
rect 9496 7701 9505 7735
rect 9505 7701 9539 7735
rect 9539 7701 9548 7735
rect 9496 7692 9548 7701
rect 9680 7692 9732 7744
rect 10692 7692 10744 7744
rect 11704 7735 11756 7744
rect 11704 7701 11713 7735
rect 11713 7701 11747 7735
rect 11747 7701 11756 7735
rect 11704 7692 11756 7701
rect 12072 7760 12124 7812
rect 12348 7828 12400 7880
rect 12440 7828 12492 7880
rect 13636 7896 13688 7948
rect 14096 7896 14148 7948
rect 12716 7692 12768 7744
rect 13176 7760 13228 7812
rect 16212 7896 16264 7948
rect 15108 7828 15160 7880
rect 15844 7828 15896 7880
rect 16580 7828 16632 7880
rect 16856 7760 16908 7812
rect 17224 7871 17276 7880
rect 17224 7837 17233 7871
rect 17233 7837 17267 7871
rect 17267 7837 17276 7871
rect 17224 7828 17276 7837
rect 17408 7760 17460 7812
rect 13912 7692 13964 7744
rect 15292 7692 15344 7744
rect 16396 7692 16448 7744
rect 18880 7692 18932 7744
rect 3947 7590 3999 7642
rect 4011 7590 4063 7642
rect 4075 7590 4127 7642
rect 4139 7590 4191 7642
rect 9878 7590 9930 7642
rect 9942 7590 9994 7642
rect 10006 7590 10058 7642
rect 10070 7590 10122 7642
rect 15808 7590 15860 7642
rect 15872 7590 15924 7642
rect 15936 7590 15988 7642
rect 16000 7590 16052 7642
rect 2228 7531 2280 7540
rect 2228 7497 2237 7531
rect 2237 7497 2271 7531
rect 2271 7497 2280 7531
rect 2228 7488 2280 7497
rect 2964 7488 3016 7540
rect 3608 7488 3660 7540
rect 4436 7488 4488 7540
rect 5080 7488 5132 7540
rect 5816 7488 5868 7540
rect 6736 7488 6788 7540
rect 7196 7531 7248 7540
rect 7196 7497 7205 7531
rect 7205 7497 7239 7531
rect 7239 7497 7248 7531
rect 7196 7488 7248 7497
rect 3240 7420 3292 7472
rect 2504 7352 2556 7404
rect 2596 7327 2648 7336
rect 2596 7293 2605 7327
rect 2605 7293 2639 7327
rect 2639 7293 2648 7327
rect 2596 7284 2648 7293
rect 3056 7284 3108 7336
rect 9496 7420 9548 7472
rect 4712 7395 4764 7404
rect 4712 7361 4721 7395
rect 4721 7361 4755 7395
rect 4755 7361 4764 7395
rect 4712 7352 4764 7361
rect 4896 7395 4948 7404
rect 4896 7361 4905 7395
rect 4905 7361 4939 7395
rect 4939 7361 4948 7395
rect 4896 7352 4948 7361
rect 5448 7352 5500 7404
rect 6000 7395 6052 7404
rect 6000 7361 6009 7395
rect 6009 7361 6043 7395
rect 6043 7361 6052 7395
rect 6000 7352 6052 7361
rect 5632 7284 5684 7336
rect 6276 7284 6328 7336
rect 6368 7284 6420 7336
rect 9404 7352 9456 7404
rect 12164 7420 12216 7472
rect 4160 7216 4212 7268
rect 3608 7191 3660 7200
rect 3608 7157 3617 7191
rect 3617 7157 3651 7191
rect 3651 7157 3660 7191
rect 3608 7148 3660 7157
rect 4620 7191 4672 7200
rect 4620 7157 4629 7191
rect 4629 7157 4663 7191
rect 4663 7157 4672 7191
rect 4620 7148 4672 7157
rect 5724 7148 5776 7200
rect 6368 7148 6420 7200
rect 7288 7148 7340 7200
rect 9496 7284 9548 7336
rect 9680 7284 9732 7336
rect 10048 7284 10100 7336
rect 12164 7284 12216 7336
rect 8576 7216 8628 7268
rect 10600 7216 10652 7268
rect 9680 7148 9732 7200
rect 9864 7148 9916 7200
rect 12072 7148 12124 7200
rect 12440 7191 12492 7200
rect 12440 7157 12449 7191
rect 12449 7157 12483 7191
rect 12483 7157 12492 7191
rect 13176 7352 13228 7404
rect 14096 7488 14148 7540
rect 15108 7531 15160 7540
rect 15108 7497 15117 7531
rect 15117 7497 15151 7531
rect 15151 7497 15160 7531
rect 15108 7488 15160 7497
rect 15292 7488 15344 7540
rect 18420 7488 18472 7540
rect 16212 7284 16264 7336
rect 12440 7148 12492 7157
rect 13636 7148 13688 7200
rect 16580 7216 16632 7268
rect 16212 7148 16264 7200
rect 6912 7046 6964 7098
rect 6976 7046 7028 7098
rect 7040 7046 7092 7098
rect 7104 7046 7156 7098
rect 12843 7046 12895 7098
rect 12907 7046 12959 7098
rect 12971 7046 13023 7098
rect 13035 7046 13087 7098
rect 1768 6944 1820 6996
rect 5448 6987 5500 6996
rect 3056 6876 3108 6928
rect 5448 6953 5457 6987
rect 5457 6953 5491 6987
rect 5491 6953 5500 6987
rect 5448 6944 5500 6953
rect 7656 6944 7708 6996
rect 8300 6987 8352 6996
rect 8300 6953 8309 6987
rect 8309 6953 8343 6987
rect 8343 6953 8352 6987
rect 8300 6944 8352 6953
rect 8484 6944 8536 6996
rect 9404 6944 9456 6996
rect 2964 6808 3016 6860
rect 3424 6808 3476 6860
rect 1676 6740 1728 6792
rect 2228 6783 2280 6792
rect 2228 6749 2237 6783
rect 2237 6749 2271 6783
rect 2271 6749 2280 6783
rect 2228 6740 2280 6749
rect 3332 6783 3384 6792
rect 3332 6749 3341 6783
rect 3341 6749 3375 6783
rect 3375 6749 3384 6783
rect 3792 6808 3844 6860
rect 9128 6876 9180 6928
rect 9864 6876 9916 6928
rect 9956 6876 10008 6928
rect 11060 6944 11112 6996
rect 12348 6944 12400 6996
rect 13360 6944 13412 6996
rect 14372 6987 14424 6996
rect 14372 6953 14381 6987
rect 14381 6953 14415 6987
rect 14415 6953 14424 6987
rect 14372 6944 14424 6953
rect 15660 6944 15712 6996
rect 6276 6851 6328 6860
rect 3332 6740 3384 6749
rect 3976 6672 4028 6724
rect 2688 6604 2740 6656
rect 6276 6817 6285 6851
rect 6285 6817 6319 6851
rect 6319 6817 6328 6851
rect 6276 6808 6328 6817
rect 10140 6808 10192 6860
rect 6552 6783 6604 6792
rect 6552 6749 6561 6783
rect 6561 6749 6595 6783
rect 6595 6749 6604 6783
rect 6552 6740 6604 6749
rect 7472 6672 7524 6724
rect 7656 6783 7708 6792
rect 7656 6749 7665 6783
rect 7665 6749 7699 6783
rect 7699 6749 7708 6783
rect 7656 6740 7708 6749
rect 8116 6740 8168 6792
rect 9496 6740 9548 6792
rect 8208 6672 8260 6724
rect 10600 6740 10652 6792
rect 10876 6783 10928 6792
rect 10876 6749 10885 6783
rect 10885 6749 10919 6783
rect 10919 6749 10928 6783
rect 10876 6740 10928 6749
rect 9956 6672 10008 6724
rect 10048 6672 10100 6724
rect 10324 6715 10376 6724
rect 10324 6681 10333 6715
rect 10333 6681 10367 6715
rect 10367 6681 10376 6715
rect 10324 6672 10376 6681
rect 10692 6672 10744 6724
rect 12072 6808 12124 6860
rect 13820 6808 13872 6860
rect 15660 6851 15712 6860
rect 13176 6740 13228 6792
rect 15660 6817 15669 6851
rect 15669 6817 15703 6851
rect 15703 6817 15712 6851
rect 15660 6808 15712 6817
rect 16856 6876 16908 6928
rect 14096 6740 14148 6792
rect 12164 6604 12216 6656
rect 13360 6604 13412 6656
rect 14004 6647 14056 6656
rect 14004 6613 14013 6647
rect 14013 6613 14047 6647
rect 14047 6613 14056 6647
rect 14004 6604 14056 6613
rect 14372 6604 14424 6656
rect 15476 6740 15528 6792
rect 15108 6672 15160 6724
rect 17224 6783 17276 6792
rect 17224 6749 17233 6783
rect 17233 6749 17267 6783
rect 17267 6749 17276 6783
rect 17224 6740 17276 6749
rect 16672 6715 16724 6724
rect 16672 6681 16681 6715
rect 16681 6681 16715 6715
rect 16715 6681 16724 6715
rect 16672 6672 16724 6681
rect 18052 6647 18104 6656
rect 18052 6613 18061 6647
rect 18061 6613 18095 6647
rect 18095 6613 18104 6647
rect 18052 6604 18104 6613
rect 3947 6502 3999 6554
rect 4011 6502 4063 6554
rect 4075 6502 4127 6554
rect 4139 6502 4191 6554
rect 9878 6502 9930 6554
rect 9942 6502 9994 6554
rect 10006 6502 10058 6554
rect 10070 6502 10122 6554
rect 15808 6502 15860 6554
rect 15872 6502 15924 6554
rect 15936 6502 15988 6554
rect 16000 6502 16052 6554
rect 2228 6400 2280 6452
rect 2780 6400 2832 6452
rect 3792 6443 3844 6452
rect 3792 6409 3801 6443
rect 3801 6409 3835 6443
rect 3835 6409 3844 6443
rect 3792 6400 3844 6409
rect 6276 6400 6328 6452
rect 8116 6443 8168 6452
rect 8116 6409 8125 6443
rect 8125 6409 8159 6443
rect 8159 6409 8168 6443
rect 8116 6400 8168 6409
rect 1860 6375 1912 6384
rect 1860 6341 1869 6375
rect 1869 6341 1903 6375
rect 1903 6341 1912 6375
rect 1860 6332 1912 6341
rect 5540 6332 5592 6384
rect 8484 6332 8536 6384
rect 8576 6332 8628 6384
rect 6276 6264 6328 6316
rect 7656 6264 7708 6316
rect 7748 6264 7800 6316
rect 9680 6400 9732 6452
rect 10324 6400 10376 6452
rect 11612 6400 11664 6452
rect 10600 6332 10652 6384
rect 11704 6264 11756 6316
rect 12164 6332 12216 6384
rect 12716 6264 12768 6316
rect 1676 6239 1728 6248
rect 1676 6205 1685 6239
rect 1685 6205 1719 6239
rect 1719 6205 1728 6239
rect 1676 6196 1728 6205
rect 4436 6239 4488 6248
rect 4436 6205 4445 6239
rect 4445 6205 4479 6239
rect 4479 6205 4488 6239
rect 4436 6196 4488 6205
rect 4712 6239 4764 6248
rect 4712 6205 4746 6239
rect 4746 6205 4764 6239
rect 6460 6239 6512 6248
rect 4712 6196 4764 6205
rect 6460 6205 6469 6239
rect 6469 6205 6503 6239
rect 6503 6205 6512 6239
rect 6460 6196 6512 6205
rect 8392 6196 8444 6248
rect 8760 6196 8812 6248
rect 10416 6196 10468 6248
rect 10600 6196 10652 6248
rect 10784 6196 10836 6248
rect 12440 6196 12492 6248
rect 4620 6128 4672 6180
rect 3424 6060 3476 6112
rect 4436 6060 4488 6112
rect 6552 6128 6604 6180
rect 7748 6128 7800 6180
rect 8300 6128 8352 6180
rect 6000 6060 6052 6112
rect 7380 6060 7432 6112
rect 12072 6128 12124 6180
rect 14188 6239 14240 6248
rect 14188 6205 14197 6239
rect 14197 6205 14231 6239
rect 14231 6205 14240 6239
rect 14188 6196 14240 6205
rect 15660 6400 15712 6452
rect 16580 6400 16632 6452
rect 17224 6400 17276 6452
rect 15752 6332 15804 6384
rect 18328 6332 18380 6384
rect 16212 6264 16264 6316
rect 14372 6128 14424 6180
rect 16396 6171 16448 6180
rect 16396 6137 16405 6171
rect 16405 6137 16439 6171
rect 16439 6137 16448 6171
rect 16396 6128 16448 6137
rect 15660 6060 15712 6112
rect 16672 6060 16724 6112
rect 17408 6103 17460 6112
rect 17408 6069 17417 6103
rect 17417 6069 17451 6103
rect 17451 6069 17460 6103
rect 17408 6060 17460 6069
rect 17592 6060 17644 6112
rect 17776 6060 17828 6112
rect 6912 5958 6964 6010
rect 6976 5958 7028 6010
rect 7040 5958 7092 6010
rect 7104 5958 7156 6010
rect 12843 5958 12895 6010
rect 12907 5958 12959 6010
rect 12971 5958 13023 6010
rect 13035 5958 13087 6010
rect 2688 5856 2740 5908
rect 2780 5788 2832 5840
rect 3332 5788 3384 5840
rect 8576 5856 8628 5908
rect 8852 5899 8904 5908
rect 8852 5865 8861 5899
rect 8861 5865 8895 5899
rect 8895 5865 8904 5899
rect 8852 5856 8904 5865
rect 7380 5788 7432 5840
rect 4436 5763 4488 5772
rect 1952 5695 2004 5704
rect 1952 5661 1961 5695
rect 1961 5661 1995 5695
rect 1995 5661 2004 5695
rect 1952 5652 2004 5661
rect 4436 5729 4445 5763
rect 4445 5729 4479 5763
rect 4479 5729 4488 5763
rect 4436 5720 4488 5729
rect 5540 5763 5592 5772
rect 5540 5729 5549 5763
rect 5549 5729 5583 5763
rect 5583 5729 5592 5763
rect 5540 5720 5592 5729
rect 3792 5652 3844 5704
rect 4344 5652 4396 5704
rect 4620 5695 4672 5704
rect 4620 5661 4629 5695
rect 4629 5661 4663 5695
rect 4663 5661 4672 5695
rect 4620 5652 4672 5661
rect 4896 5652 4948 5704
rect 5356 5652 5408 5704
rect 6000 5720 6052 5772
rect 10692 5788 10744 5840
rect 11336 5788 11388 5840
rect 12072 5856 12124 5908
rect 11980 5788 12032 5840
rect 13176 5788 13228 5840
rect 13360 5831 13412 5840
rect 13360 5797 13394 5831
rect 13394 5797 13412 5831
rect 14004 5856 14056 5908
rect 16580 5831 16632 5840
rect 13360 5788 13412 5797
rect 16580 5797 16589 5831
rect 16589 5797 16623 5831
rect 16623 5797 16632 5831
rect 16580 5788 16632 5797
rect 9496 5720 9548 5772
rect 10324 5720 10376 5772
rect 9036 5652 9088 5704
rect 9680 5695 9732 5704
rect 9680 5661 9689 5695
rect 9689 5661 9723 5695
rect 9723 5661 9732 5695
rect 9680 5652 9732 5661
rect 10692 5652 10744 5704
rect 11980 5652 12032 5704
rect 14188 5720 14240 5772
rect 14740 5720 14792 5772
rect 15660 5720 15712 5772
rect 15752 5652 15804 5704
rect 16212 5652 16264 5704
rect 16396 5652 16448 5704
rect 16856 5720 16908 5772
rect 17776 5763 17828 5772
rect 17776 5729 17785 5763
rect 17785 5729 17819 5763
rect 17819 5729 17828 5763
rect 17776 5720 17828 5729
rect 17224 5652 17276 5704
rect 3424 5516 3476 5568
rect 8116 5584 8168 5636
rect 7656 5559 7708 5568
rect 7656 5525 7665 5559
rect 7665 5525 7699 5559
rect 7699 5525 7708 5559
rect 7656 5516 7708 5525
rect 8024 5516 8076 5568
rect 8944 5584 8996 5636
rect 10784 5584 10836 5636
rect 12072 5584 12124 5636
rect 14372 5584 14424 5636
rect 17500 5584 17552 5636
rect 8484 5516 8536 5568
rect 10324 5516 10376 5568
rect 10416 5516 10468 5568
rect 12716 5516 12768 5568
rect 14096 5516 14148 5568
rect 15660 5559 15712 5568
rect 15660 5525 15669 5559
rect 15669 5525 15703 5559
rect 15703 5525 15712 5559
rect 15660 5516 15712 5525
rect 16212 5559 16264 5568
rect 16212 5525 16221 5559
rect 16221 5525 16255 5559
rect 16255 5525 16264 5559
rect 16212 5516 16264 5525
rect 17408 5559 17460 5568
rect 17408 5525 17417 5559
rect 17417 5525 17451 5559
rect 17451 5525 17460 5559
rect 17408 5516 17460 5525
rect 3947 5414 3999 5466
rect 4011 5414 4063 5466
rect 4075 5414 4127 5466
rect 4139 5414 4191 5466
rect 9878 5414 9930 5466
rect 9942 5414 9994 5466
rect 10006 5414 10058 5466
rect 10070 5414 10122 5466
rect 15808 5414 15860 5466
rect 15872 5414 15924 5466
rect 15936 5414 15988 5466
rect 16000 5414 16052 5466
rect 1860 5355 1912 5364
rect 1860 5321 1869 5355
rect 1869 5321 1903 5355
rect 1903 5321 1912 5355
rect 1860 5312 1912 5321
rect 4436 5312 4488 5364
rect 8300 5312 8352 5364
rect 9496 5355 9548 5364
rect 9496 5321 9505 5355
rect 9505 5321 9539 5355
rect 9539 5321 9548 5355
rect 9496 5312 9548 5321
rect 6276 5287 6328 5296
rect 6276 5253 6285 5287
rect 6285 5253 6319 5287
rect 6319 5253 6328 5287
rect 6276 5244 6328 5253
rect 7288 5287 7340 5296
rect 7288 5253 7297 5287
rect 7297 5253 7331 5287
rect 7331 5253 7340 5287
rect 7288 5244 7340 5253
rect 8024 5244 8076 5296
rect 2872 5176 2924 5228
rect 4712 5176 4764 5228
rect 6000 5176 6052 5228
rect 2872 5083 2924 5092
rect 2872 5049 2881 5083
rect 2881 5049 2915 5083
rect 2915 5049 2924 5083
rect 2872 5040 2924 5049
rect 4528 5108 4580 5160
rect 4896 5151 4948 5160
rect 4896 5117 4905 5151
rect 4905 5117 4939 5151
rect 4939 5117 4948 5151
rect 4896 5108 4948 5117
rect 5080 5040 5132 5092
rect 6736 5108 6788 5160
rect 7380 5108 7432 5160
rect 8024 5108 8076 5160
rect 10784 5312 10836 5364
rect 15476 5355 15528 5364
rect 15476 5321 15485 5355
rect 15485 5321 15519 5355
rect 15519 5321 15528 5355
rect 15476 5312 15528 5321
rect 16672 5355 16724 5364
rect 16672 5321 16681 5355
rect 16681 5321 16715 5355
rect 16715 5321 16724 5355
rect 16672 5312 16724 5321
rect 11980 5287 12032 5296
rect 9680 5176 9732 5228
rect 9036 5040 9088 5092
rect 10416 5151 10468 5160
rect 10416 5117 10450 5151
rect 10450 5117 10468 5151
rect 10416 5108 10468 5117
rect 11980 5253 11989 5287
rect 11989 5253 12023 5287
rect 12023 5253 12032 5287
rect 11980 5244 12032 5253
rect 12440 5244 12492 5296
rect 14004 5244 14056 5296
rect 13636 5176 13688 5228
rect 14464 5176 14516 5228
rect 16396 5176 16448 5228
rect 17224 5219 17276 5228
rect 17224 5185 17233 5219
rect 17233 5185 17267 5219
rect 17267 5185 17276 5219
rect 17224 5176 17276 5185
rect 10324 5040 10376 5092
rect 12716 5108 12768 5160
rect 13268 5040 13320 5092
rect 16212 5108 16264 5160
rect 17040 5151 17092 5160
rect 17040 5117 17049 5151
rect 17049 5117 17083 5151
rect 17083 5117 17092 5151
rect 17040 5108 17092 5117
rect 4068 4972 4120 5024
rect 5632 4972 5684 5024
rect 8208 4972 8260 5024
rect 9220 4972 9272 5024
rect 9496 4972 9548 5024
rect 10692 4972 10744 5024
rect 11704 4972 11756 5024
rect 17408 5040 17460 5092
rect 14740 4972 14792 5024
rect 16028 4972 16080 5024
rect 6912 4870 6964 4922
rect 6976 4870 7028 4922
rect 7040 4870 7092 4922
rect 7104 4870 7156 4922
rect 12843 4870 12895 4922
rect 12907 4870 12959 4922
rect 12971 4870 13023 4922
rect 13035 4870 13087 4922
rect 1768 4768 1820 4820
rect 2780 4768 2832 4820
rect 2964 4768 3016 4820
rect 3148 4768 3200 4820
rect 4068 4768 4120 4820
rect 5264 4768 5316 4820
rect 5632 4811 5684 4820
rect 5632 4777 5641 4811
rect 5641 4777 5675 4811
rect 5675 4777 5684 4811
rect 5632 4768 5684 4777
rect 2320 4700 2372 4752
rect 2412 4675 2464 4684
rect 2412 4641 2421 4675
rect 2421 4641 2455 4675
rect 2455 4641 2464 4675
rect 2412 4632 2464 4641
rect 4804 4675 4856 4684
rect 4804 4641 4813 4675
rect 4813 4641 4847 4675
rect 4847 4641 4856 4675
rect 4804 4632 4856 4641
rect 4988 4632 5040 4684
rect 5540 4632 5592 4684
rect 6000 4675 6052 4684
rect 6000 4641 6009 4675
rect 6009 4641 6043 4675
rect 6043 4641 6052 4675
rect 6000 4632 6052 4641
rect 6460 4632 6512 4684
rect 8852 4768 8904 4820
rect 9036 4811 9088 4820
rect 9036 4777 9045 4811
rect 9045 4777 9079 4811
rect 9079 4777 9088 4811
rect 9036 4768 9088 4777
rect 9128 4768 9180 4820
rect 12440 4768 12492 4820
rect 13912 4768 13964 4820
rect 14464 4768 14516 4820
rect 16856 4811 16908 4820
rect 5080 4607 5132 4616
rect 5080 4573 5089 4607
rect 5089 4573 5123 4607
rect 5123 4573 5132 4607
rect 5080 4564 5132 4573
rect 5448 4564 5500 4616
rect 6368 4564 6420 4616
rect 6828 4564 6880 4616
rect 8024 4700 8076 4752
rect 11796 4743 11848 4752
rect 11796 4709 11805 4743
rect 11805 4709 11839 4743
rect 11839 4709 11848 4743
rect 11796 4700 11848 4709
rect 11980 4700 12032 4752
rect 13360 4700 13412 4752
rect 14096 4700 14148 4752
rect 15016 4700 15068 4752
rect 15384 4700 15436 4752
rect 16856 4777 16865 4811
rect 16865 4777 16899 4811
rect 16899 4777 16908 4811
rect 16856 4768 16908 4777
rect 8484 4632 8536 4684
rect 10692 4675 10744 4684
rect 10692 4641 10701 4675
rect 10701 4641 10735 4675
rect 10735 4641 10744 4675
rect 10692 4632 10744 4641
rect 16396 4632 16448 4684
rect 18236 4768 18288 4820
rect 8944 4564 8996 4616
rect 13820 4564 13872 4616
rect 15384 4607 15436 4616
rect 9496 4496 9548 4548
rect 14096 4496 14148 4548
rect 15384 4573 15393 4607
rect 15393 4573 15427 4607
rect 15427 4573 15436 4607
rect 15384 4564 15436 4573
rect 15568 4564 15620 4616
rect 16672 4564 16724 4616
rect 17316 4564 17368 4616
rect 17500 4607 17552 4616
rect 17500 4573 17509 4607
rect 17509 4573 17543 4607
rect 17543 4573 17552 4607
rect 17500 4564 17552 4573
rect 17684 4496 17736 4548
rect 3056 4428 3108 4480
rect 4436 4471 4488 4480
rect 4436 4437 4445 4471
rect 4445 4437 4479 4471
rect 4479 4437 4488 4471
rect 4436 4428 4488 4437
rect 9128 4428 9180 4480
rect 9772 4428 9824 4480
rect 16212 4428 16264 4480
rect 3947 4326 3999 4378
rect 4011 4326 4063 4378
rect 4075 4326 4127 4378
rect 4139 4326 4191 4378
rect 9878 4326 9930 4378
rect 9942 4326 9994 4378
rect 10006 4326 10058 4378
rect 10070 4326 10122 4378
rect 15808 4326 15860 4378
rect 15872 4326 15924 4378
rect 15936 4326 15988 4378
rect 16000 4326 16052 4378
rect 1860 4267 1912 4276
rect 1860 4233 1869 4267
rect 1869 4233 1903 4267
rect 1903 4233 1912 4267
rect 1860 4224 1912 4233
rect 4344 4224 4396 4276
rect 4528 4224 4580 4276
rect 204 4088 256 4140
rect 1952 4088 2004 4140
rect 4436 4131 4488 4140
rect 4436 4097 4445 4131
rect 4445 4097 4479 4131
rect 4479 4097 4488 4131
rect 4436 4088 4488 4097
rect 4712 4156 4764 4208
rect 6276 4156 6328 4208
rect 6368 4088 6420 4140
rect 6552 4224 6604 4276
rect 9496 4267 9548 4276
rect 9496 4233 9505 4267
rect 9505 4233 9539 4267
rect 9539 4233 9548 4267
rect 9496 4224 9548 4233
rect 8392 4156 8444 4208
rect 8944 4156 8996 4208
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 10048 4088 10100 4140
rect 2688 4020 2740 4072
rect 3148 4063 3200 4072
rect 3148 4029 3157 4063
rect 3157 4029 3191 4063
rect 3191 4029 3200 4063
rect 3148 4020 3200 4029
rect 3884 4020 3936 4072
rect 6000 4020 6052 4072
rect 6276 4020 6328 4072
rect 5540 3995 5592 4004
rect 2780 3884 2832 3936
rect 3332 3927 3384 3936
rect 3332 3893 3341 3927
rect 3341 3893 3375 3927
rect 3375 3893 3384 3927
rect 3332 3884 3384 3893
rect 5540 3961 5549 3995
rect 5549 3961 5583 3995
rect 5583 3961 5592 3995
rect 5540 3952 5592 3961
rect 5816 3952 5868 4004
rect 6552 3952 6604 4004
rect 6920 3952 6972 4004
rect 10416 4224 10468 4276
rect 13176 4088 13228 4140
rect 13268 4088 13320 4140
rect 13728 4131 13780 4140
rect 13728 4097 13737 4131
rect 13737 4097 13771 4131
rect 13771 4097 13780 4131
rect 13728 4088 13780 4097
rect 14924 4131 14976 4140
rect 14924 4097 14933 4131
rect 14933 4097 14967 4131
rect 14967 4097 14976 4131
rect 14924 4088 14976 4097
rect 17132 4131 17184 4140
rect 17132 4097 17141 4131
rect 17141 4097 17175 4131
rect 17175 4097 17184 4131
rect 17132 4088 17184 4097
rect 10324 4020 10376 4072
rect 7288 3952 7340 4004
rect 11888 4020 11940 4072
rect 10692 3952 10744 4004
rect 13544 3952 13596 4004
rect 14096 3952 14148 4004
rect 14556 3995 14608 4004
rect 14556 3961 14565 3995
rect 14565 3961 14599 3995
rect 14599 3961 14608 3995
rect 16212 3995 16264 4004
rect 14556 3952 14608 3961
rect 16212 3961 16221 3995
rect 16221 3961 16255 3995
rect 16255 3961 16264 3995
rect 16212 3952 16264 3961
rect 8484 3884 8536 3936
rect 8668 3884 8720 3936
rect 9312 3884 9364 3936
rect 9864 3884 9916 3936
rect 14280 3884 14332 3936
rect 15660 3884 15712 3936
rect 6912 3782 6964 3834
rect 6976 3782 7028 3834
rect 7040 3782 7092 3834
rect 7104 3782 7156 3834
rect 12843 3782 12895 3834
rect 12907 3782 12959 3834
rect 12971 3782 13023 3834
rect 13035 3782 13087 3834
rect 3884 3680 3936 3732
rect 7288 3723 7340 3732
rect 7288 3689 7297 3723
rect 7297 3689 7331 3723
rect 7331 3689 7340 3723
rect 7288 3680 7340 3689
rect 7748 3723 7800 3732
rect 7748 3689 7757 3723
rect 7757 3689 7791 3723
rect 7791 3689 7800 3723
rect 7748 3680 7800 3689
rect 8760 3680 8812 3732
rect 11980 3680 12032 3732
rect 12256 3680 12308 3732
rect 3608 3544 3660 3596
rect 4528 3612 4580 3664
rect 4620 3544 4672 3596
rect 3240 3476 3292 3528
rect 7380 3612 7432 3664
rect 7656 3612 7708 3664
rect 8024 3612 8076 3664
rect 9864 3612 9916 3664
rect 9036 3544 9088 3596
rect 10508 3612 10560 3664
rect 14648 3680 14700 3732
rect 15384 3680 15436 3732
rect 17776 3680 17828 3732
rect 15200 3612 15252 3664
rect 16304 3612 16356 3664
rect 17868 3612 17920 3664
rect 14464 3587 14516 3596
rect 14464 3553 14473 3587
rect 14473 3553 14507 3587
rect 14507 3553 14516 3587
rect 14464 3544 14516 3553
rect 7472 3476 7524 3528
rect 10784 3519 10836 3528
rect 10784 3485 10793 3519
rect 10793 3485 10827 3519
rect 10827 3485 10836 3519
rect 10784 3476 10836 3485
rect 11612 3476 11664 3528
rect 5448 3451 5500 3460
rect 5448 3417 5457 3451
rect 5457 3417 5491 3451
rect 5491 3417 5500 3451
rect 5448 3408 5500 3417
rect 8392 3451 8444 3460
rect 8392 3417 8401 3451
rect 8401 3417 8435 3451
rect 8435 3417 8444 3451
rect 8392 3408 8444 3417
rect 1860 3383 1912 3392
rect 1860 3349 1869 3383
rect 1869 3349 1903 3383
rect 1903 3349 1912 3383
rect 1860 3340 1912 3349
rect 2688 3340 2740 3392
rect 6276 3340 6328 3392
rect 6552 3340 6604 3392
rect 9772 3408 9824 3460
rect 10048 3451 10100 3460
rect 10048 3417 10057 3451
rect 10057 3417 10091 3451
rect 10091 3417 10100 3451
rect 10048 3408 10100 3417
rect 10416 3408 10468 3460
rect 11428 3408 11480 3460
rect 12164 3476 12216 3528
rect 13452 3519 13504 3528
rect 13452 3485 13461 3519
rect 13461 3485 13495 3519
rect 13495 3485 13504 3519
rect 13452 3476 13504 3485
rect 15108 3476 15160 3528
rect 17500 3519 17552 3528
rect 11796 3408 11848 3460
rect 17500 3485 17509 3519
rect 17509 3485 17543 3519
rect 17543 3485 17552 3519
rect 17500 3476 17552 3485
rect 8944 3340 8996 3392
rect 10784 3340 10836 3392
rect 15568 3340 15620 3392
rect 3947 3238 3999 3290
rect 4011 3238 4063 3290
rect 4075 3238 4127 3290
rect 4139 3238 4191 3290
rect 9878 3238 9930 3290
rect 9942 3238 9994 3290
rect 10006 3238 10058 3290
rect 10070 3238 10122 3290
rect 15808 3238 15860 3290
rect 15872 3238 15924 3290
rect 15936 3238 15988 3290
rect 16000 3238 16052 3290
rect 9680 3136 9732 3188
rect 17408 3179 17460 3188
rect 17408 3145 17417 3179
rect 17417 3145 17451 3179
rect 17451 3145 17460 3179
rect 17408 3136 17460 3145
rect 9772 3068 9824 3120
rect 1676 3000 1728 3052
rect 4528 3000 4580 3052
rect 6092 3000 6144 3052
rect 8208 3000 8260 3052
rect 10600 3000 10652 3052
rect 11152 3000 11204 3052
rect 12348 3000 12400 3052
rect 12532 3043 12584 3052
rect 12532 3009 12541 3043
rect 12541 3009 12575 3043
rect 12575 3009 12584 3043
rect 12532 3000 12584 3009
rect 12624 3000 12676 3052
rect 14924 3043 14976 3052
rect 14924 3009 14933 3043
rect 14933 3009 14967 3043
rect 14967 3009 14976 3043
rect 14924 3000 14976 3009
rect 16488 3043 16540 3052
rect 16488 3009 16497 3043
rect 16497 3009 16531 3043
rect 16531 3009 16540 3043
rect 16488 3000 16540 3009
rect 2044 2932 2096 2984
rect 1124 2864 1176 2916
rect 2136 2864 2188 2916
rect 3424 2932 3476 2984
rect 4252 2975 4304 2984
rect 4252 2941 4261 2975
rect 4261 2941 4295 2975
rect 4295 2941 4304 2975
rect 4252 2932 4304 2941
rect 5816 2932 5868 2984
rect 6552 2932 6604 2984
rect 6736 2932 6788 2984
rect 7288 2932 7340 2984
rect 7472 2932 7524 2984
rect 3148 2864 3200 2916
rect 7564 2864 7616 2916
rect 8576 2864 8628 2916
rect 8760 2907 8812 2916
rect 8760 2873 8769 2907
rect 8769 2873 8803 2907
rect 8803 2873 8812 2907
rect 8760 2864 8812 2873
rect 9588 2864 9640 2916
rect 10324 2907 10376 2916
rect 10324 2873 10333 2907
rect 10333 2873 10367 2907
rect 10367 2873 10376 2907
rect 10324 2864 10376 2873
rect 10416 2907 10468 2916
rect 10416 2873 10425 2907
rect 10425 2873 10459 2907
rect 10459 2873 10468 2907
rect 16580 2932 16632 2984
rect 10416 2864 10468 2873
rect 13544 2907 13596 2916
rect 13544 2873 13553 2907
rect 13553 2873 13587 2907
rect 13587 2873 13596 2907
rect 13544 2864 13596 2873
rect 9220 2796 9272 2848
rect 11152 2796 11204 2848
rect 12716 2796 12768 2848
rect 14556 2864 14608 2916
rect 15752 2907 15804 2916
rect 15752 2873 15761 2907
rect 15761 2873 15795 2907
rect 15795 2873 15804 2907
rect 15752 2864 15804 2873
rect 6912 2694 6964 2746
rect 6976 2694 7028 2746
rect 7040 2694 7092 2746
rect 7104 2694 7156 2746
rect 12843 2694 12895 2746
rect 12907 2694 12959 2746
rect 12971 2694 13023 2746
rect 13035 2694 13087 2746
rect 2964 2592 3016 2644
rect 3424 2635 3476 2644
rect 3424 2601 3433 2635
rect 3433 2601 3467 2635
rect 3467 2601 3476 2635
rect 3424 2592 3476 2601
rect 8208 2592 8260 2644
rect 8760 2592 8812 2644
rect 9220 2592 9272 2644
rect 16212 2635 16264 2644
rect 1584 2499 1636 2508
rect 1584 2465 1593 2499
rect 1593 2465 1627 2499
rect 1627 2465 1636 2499
rect 1584 2456 1636 2465
rect 2504 2499 2556 2508
rect 2504 2465 2513 2499
rect 2513 2465 2547 2499
rect 2547 2465 2556 2499
rect 2504 2456 2556 2465
rect 3056 2456 3108 2508
rect 5540 2524 5592 2576
rect 4804 2499 4856 2508
rect 4804 2465 4813 2499
rect 4813 2465 4847 2499
rect 4847 2465 4856 2499
rect 4804 2456 4856 2465
rect 8944 2524 8996 2576
rect 10232 2567 10284 2576
rect 10232 2533 10241 2567
rect 10241 2533 10275 2567
rect 10275 2533 10284 2567
rect 10232 2524 10284 2533
rect 10508 2524 10560 2576
rect 10692 2524 10744 2576
rect 11520 2524 11572 2576
rect 16212 2601 16221 2635
rect 16221 2601 16255 2635
rect 16255 2601 16264 2635
rect 16212 2592 16264 2601
rect 16948 2635 17000 2644
rect 16948 2601 16957 2635
rect 16957 2601 16991 2635
rect 16991 2601 17000 2635
rect 16948 2592 17000 2601
rect 17684 2635 17736 2644
rect 17684 2601 17693 2635
rect 17693 2601 17727 2635
rect 17727 2601 17736 2635
rect 17684 2592 17736 2601
rect 7380 2456 7432 2508
rect 8300 2456 8352 2508
rect 8484 2499 8536 2508
rect 8484 2465 8493 2499
rect 8493 2465 8527 2499
rect 8527 2465 8536 2499
rect 8484 2456 8536 2465
rect 11336 2456 11388 2508
rect 11796 2499 11848 2508
rect 11796 2465 11805 2499
rect 11805 2465 11839 2499
rect 11839 2465 11848 2499
rect 11796 2456 11848 2465
rect 14832 2567 14884 2576
rect 14832 2533 14841 2567
rect 14841 2533 14875 2567
rect 14875 2533 14884 2567
rect 14832 2524 14884 2533
rect 16028 2499 16080 2508
rect 16028 2465 16037 2499
rect 16037 2465 16071 2499
rect 16071 2465 16080 2499
rect 16028 2456 16080 2465
rect 16764 2499 16816 2508
rect 16764 2465 16773 2499
rect 16773 2465 16807 2499
rect 16807 2465 16816 2499
rect 16764 2456 16816 2465
rect 17500 2499 17552 2508
rect 17500 2465 17509 2499
rect 17509 2465 17543 2499
rect 17543 2465 17552 2499
rect 17500 2456 17552 2465
rect 664 2388 716 2440
rect 11060 2388 11112 2440
rect 6736 2320 6788 2372
rect 8392 2320 8444 2372
rect 3516 2252 3568 2304
rect 4988 2295 5040 2304
rect 4988 2261 4997 2295
rect 4997 2261 5031 2295
rect 5031 2261 5040 2295
rect 4988 2252 5040 2261
rect 10692 2252 10744 2304
rect 13084 2252 13136 2304
rect 16212 2252 16264 2304
rect 3947 2150 3999 2202
rect 4011 2150 4063 2202
rect 4075 2150 4127 2202
rect 4139 2150 4191 2202
rect 9878 2150 9930 2202
rect 9942 2150 9994 2202
rect 10006 2150 10058 2202
rect 10070 2150 10122 2202
rect 15808 2150 15860 2202
rect 15872 2150 15924 2202
rect 15936 2150 15988 2202
rect 16000 2150 16052 2202
rect 13084 2048 13136 2100
rect 15016 2048 15068 2100
rect 5172 1300 5224 1352
rect 8024 1300 8076 1352
rect 7104 1096 7156 1148
rect 7932 1096 7984 1148
rect 3700 688 3752 740
rect 4988 688 5040 740
<< metal2 >>
rect 294 16520 350 17000
rect 938 16520 994 17000
rect 1582 16520 1638 17000
rect 2226 16520 2282 17000
rect 2870 16520 2926 17000
rect 3514 16520 3570 17000
rect 3606 16688 3662 16697
rect 3606 16623 3662 16632
rect 308 13802 336 16520
rect 296 13796 348 13802
rect 296 13738 348 13744
rect 952 13530 980 16520
rect 1596 14618 1624 16520
rect 2240 14618 2268 16520
rect 2410 16280 2466 16289
rect 2410 16215 2466 16224
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 1676 14272 1728 14278
rect 1676 14214 1728 14220
rect 1492 13864 1544 13870
rect 1492 13806 1544 13812
rect 940 13524 992 13530
rect 940 13466 992 13472
rect 1504 11354 1532 13806
rect 1584 13456 1636 13462
rect 1584 13398 1636 13404
rect 1596 11694 1624 13398
rect 1584 11688 1636 11694
rect 1584 11630 1636 11636
rect 1492 11348 1544 11354
rect 1492 11290 1544 11296
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1596 10266 1624 11086
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1596 9042 1624 9454
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1584 8560 1636 8566
rect 1584 8502 1636 8508
rect 204 4140 256 4146
rect 204 4082 256 4088
rect 216 480 244 4082
rect 1124 2916 1176 2922
rect 1124 2858 1176 2864
rect 664 2440 716 2446
rect 664 2382 716 2388
rect 676 480 704 2382
rect 1136 480 1164 2858
rect 1596 2514 1624 8502
rect 1688 6798 1716 14214
rect 2044 14000 2096 14006
rect 2044 13942 2096 13948
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1872 12782 1900 13126
rect 1964 12986 1992 13670
rect 1952 12980 2004 12986
rect 1952 12922 2004 12928
rect 1860 12776 1912 12782
rect 1860 12718 1912 12724
rect 1952 12640 2004 12646
rect 1952 12582 2004 12588
rect 1964 12442 1992 12582
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1780 7993 1808 11494
rect 1872 11354 1900 11494
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1766 7984 1822 7993
rect 1766 7919 1822 7928
rect 1766 7304 1822 7313
rect 1766 7239 1822 7248
rect 1780 7002 1808 7239
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1688 6254 1716 6734
rect 1860 6384 1912 6390
rect 1858 6352 1860 6361
rect 1912 6352 1914 6361
rect 1858 6287 1914 6296
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1858 5944 1914 5953
rect 1858 5879 1914 5888
rect 1766 5536 1822 5545
rect 1766 5471 1822 5480
rect 1780 4826 1808 5471
rect 1872 5370 1900 5879
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 1860 5364 1912 5370
rect 1860 5306 1912 5312
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 1858 4720 1914 4729
rect 1858 4655 1914 4664
rect 1872 4282 1900 4655
rect 1860 4276 1912 4282
rect 1860 4218 1912 4224
rect 1964 4146 1992 5646
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 1860 3392 1912 3398
rect 1860 3334 1912 3340
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 1688 480 1716 2994
rect 1872 2281 1900 3334
rect 2056 2990 2084 13942
rect 2226 13832 2282 13841
rect 2226 13767 2282 13776
rect 2136 12844 2188 12850
rect 2136 12786 2188 12792
rect 2148 11150 2176 12786
rect 2240 11626 2268 13767
rect 2424 12306 2452 16215
rect 2884 14074 2912 16520
rect 3146 15872 3202 15881
rect 3146 15807 3202 15816
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2792 12714 2820 13262
rect 2780 12708 2832 12714
rect 3056 12708 3108 12714
rect 2780 12650 2832 12656
rect 2976 12668 3056 12696
rect 2412 12300 2464 12306
rect 2412 12242 2464 12248
rect 2792 12238 2820 12650
rect 2976 12442 3004 12668
rect 3056 12650 3108 12656
rect 3054 12608 3110 12617
rect 3054 12543 3110 12552
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 2780 12232 2832 12238
rect 2780 12174 2832 12180
rect 2228 11620 2280 11626
rect 2228 11562 2280 11568
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 2332 11014 2360 12174
rect 2688 11824 2740 11830
rect 2688 11766 2740 11772
rect 2320 11008 2372 11014
rect 2320 10950 2372 10956
rect 2136 8560 2188 8566
rect 2136 8502 2188 8508
rect 2148 7585 2176 8502
rect 2228 8288 2280 8294
rect 2228 8230 2280 8236
rect 2134 7576 2190 7585
rect 2240 7546 2268 8230
rect 2134 7511 2190 7520
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 2240 6458 2268 6734
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2332 4758 2360 10950
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2424 10198 2452 10542
rect 2700 10441 2728 11766
rect 2792 11762 2820 12174
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2976 11694 3004 12378
rect 3068 12238 3096 12543
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 3056 12096 3108 12102
rect 3056 12038 3108 12044
rect 2964 11688 3016 11694
rect 2964 11630 3016 11636
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2792 11354 2820 11494
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2780 10532 2832 10538
rect 2780 10474 2832 10480
rect 2872 10532 2924 10538
rect 2872 10474 2924 10480
rect 2686 10432 2742 10441
rect 2686 10367 2742 10376
rect 2412 10192 2464 10198
rect 2412 10134 2464 10140
rect 2596 10056 2648 10062
rect 2594 10024 2596 10033
rect 2648 10024 2650 10033
rect 2594 9959 2650 9968
rect 2608 9761 2636 9959
rect 2594 9752 2650 9761
rect 2594 9687 2650 9696
rect 2700 9382 2728 10367
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2688 9104 2740 9110
rect 2688 9046 2740 9052
rect 2700 8838 2728 9046
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2412 8356 2464 8362
rect 2412 8298 2464 8304
rect 2320 4752 2372 4758
rect 2320 4694 2372 4700
rect 2424 4690 2452 8298
rect 2700 7834 2728 8774
rect 2516 7806 2728 7834
rect 2516 7410 2544 7806
rect 2596 7744 2648 7750
rect 2596 7686 2648 7692
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2608 7342 2636 7686
rect 2596 7336 2648 7342
rect 2596 7278 2648 7284
rect 2792 7177 2820 10474
rect 2884 10441 2912 10474
rect 2870 10432 2926 10441
rect 2870 10367 2926 10376
rect 2976 10198 3004 11630
rect 3068 10248 3096 12038
rect 3160 11830 3188 15807
rect 3528 14822 3556 16520
rect 3620 15298 3648 16623
rect 4158 16520 4214 17000
rect 4802 16520 4858 17000
rect 5446 16520 5502 17000
rect 6090 16520 6146 17000
rect 6734 16520 6790 17000
rect 7378 16520 7434 17000
rect 8022 16520 8078 17000
rect 8666 16520 8722 17000
rect 9310 16520 9366 17000
rect 9954 16520 10010 17000
rect 10598 16520 10654 17000
rect 11242 16520 11298 17000
rect 11886 16520 11942 17000
rect 12530 16520 12586 17000
rect 13174 16520 13230 17000
rect 13818 16520 13874 17000
rect 14462 16520 14518 17000
rect 15106 16520 15162 17000
rect 15198 16688 15254 16697
rect 15198 16623 15254 16632
rect 3608 15292 3660 15298
rect 3608 15234 3660 15240
rect 3790 15056 3846 15065
rect 3790 14991 3846 15000
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 3698 14648 3754 14657
rect 3698 14583 3754 14592
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3514 14240 3570 14249
rect 3436 13802 3464 14214
rect 3514 14175 3570 14184
rect 3528 14074 3556 14175
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3424 13796 3476 13802
rect 3424 13738 3476 13744
rect 3514 13424 3570 13433
rect 3514 13359 3570 13368
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3148 11824 3200 11830
rect 3148 11766 3200 11772
rect 3146 11384 3202 11393
rect 3146 11319 3202 11328
rect 3160 11286 3188 11319
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3160 10606 3188 11086
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3068 10220 3188 10248
rect 2964 10192 3016 10198
rect 2964 10134 3016 10140
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2884 8430 2912 9862
rect 2976 9586 3004 10134
rect 3056 10124 3108 10130
rect 3056 10066 3108 10072
rect 3068 9722 3096 10066
rect 3056 9716 3108 9722
rect 3056 9658 3108 9664
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2976 9178 3004 9386
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 2976 8498 3004 9114
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 3068 8430 3096 9318
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 3056 8424 3108 8430
rect 3160 8401 3188 10220
rect 3056 8366 3108 8372
rect 3146 8392 3202 8401
rect 3146 8327 3202 8336
rect 3056 8288 3108 8294
rect 2870 8256 2926 8265
rect 3056 8230 3108 8236
rect 2870 8191 2926 8200
rect 2778 7168 2834 7177
rect 2778 7103 2834 7112
rect 2502 7032 2558 7041
rect 2502 6967 2558 6976
rect 2516 5273 2544 6967
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2700 5914 2728 6598
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2688 5908 2740 5914
rect 2688 5850 2740 5856
rect 2792 5846 2820 6394
rect 2780 5840 2832 5846
rect 2780 5782 2832 5788
rect 2502 5264 2558 5273
rect 2884 5234 2912 8191
rect 2964 7540 3016 7546
rect 2964 7482 3016 7488
rect 2976 7188 3004 7482
rect 3068 7342 3096 8230
rect 3252 8090 3280 13262
rect 3330 13016 3386 13025
rect 3330 12951 3386 12960
rect 3344 12345 3372 12951
rect 3528 12782 3556 13359
rect 3516 12776 3568 12782
rect 3516 12718 3568 12724
rect 3330 12336 3386 12345
rect 3330 12271 3386 12280
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3712 12186 3740 14583
rect 3804 12968 3832 14991
rect 4172 14362 4200 16520
rect 4172 14334 4292 14362
rect 3921 14172 4217 14192
rect 3977 14170 4001 14172
rect 4057 14170 4081 14172
rect 4137 14170 4161 14172
rect 3999 14118 4001 14170
rect 4063 14118 4075 14170
rect 4137 14118 4139 14170
rect 3977 14116 4001 14118
rect 4057 14116 4081 14118
rect 4137 14116 4161 14118
rect 3921 14096 4217 14116
rect 4264 13462 4292 14334
rect 4620 14000 4672 14006
rect 4620 13942 4672 13948
rect 4252 13456 4304 13462
rect 4252 13398 4304 13404
rect 4528 13252 4580 13258
rect 4528 13194 4580 13200
rect 3921 13084 4217 13104
rect 3977 13082 4001 13084
rect 4057 13082 4081 13084
rect 4137 13082 4161 13084
rect 3999 13030 4001 13082
rect 4063 13030 4075 13082
rect 4137 13030 4139 13082
rect 3977 13028 4001 13030
rect 4057 13028 4081 13030
rect 4137 13028 4161 13030
rect 3921 13008 4217 13028
rect 3804 12940 3924 12968
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 3344 11801 3372 12038
rect 3330 11792 3386 11801
rect 3330 11727 3386 11736
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 3344 10470 3372 11086
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3344 10062 3372 10406
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3344 9654 3372 9998
rect 3332 9648 3384 9654
rect 3332 9590 3384 9596
rect 3436 8401 3464 12174
rect 3608 12164 3660 12170
rect 3712 12158 3832 12186
rect 3896 12170 3924 12940
rect 4540 12850 4568 13194
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 4344 12640 4396 12646
rect 4344 12582 4396 12588
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4068 12232 4120 12238
rect 4066 12200 4068 12209
rect 4264 12209 4292 12242
rect 4120 12200 4122 12209
rect 3608 12106 3660 12112
rect 3516 11824 3568 11830
rect 3516 11766 3568 11772
rect 3528 10470 3556 11766
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3528 9994 3556 10406
rect 3516 9988 3568 9994
rect 3516 9930 3568 9936
rect 3514 9888 3570 9897
rect 3514 9823 3570 9832
rect 3422 8392 3478 8401
rect 3422 8327 3478 8336
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 2976 7160 3096 7188
rect 3068 6934 3096 7160
rect 3056 6928 3108 6934
rect 3054 6896 3056 6905
rect 3108 6896 3110 6905
rect 2964 6860 3016 6866
rect 3054 6831 3110 6840
rect 2964 6802 3016 6808
rect 2502 5199 2558 5208
rect 2872 5228 2924 5234
rect 2412 4684 2464 4690
rect 2412 4626 2464 4632
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 2136 2916 2188 2922
rect 2136 2858 2188 2864
rect 1858 2272 1914 2281
rect 1858 2207 1914 2216
rect 2148 480 2176 2858
rect 2516 2514 2544 5199
rect 2872 5170 2924 5176
rect 2778 5128 2834 5137
rect 2778 5063 2834 5072
rect 2872 5092 2924 5098
rect 2792 4826 2820 5063
rect 2872 5034 2924 5040
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2778 4312 2834 4321
rect 2778 4247 2834 4256
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2700 3398 2728 4014
rect 2792 3942 2820 4247
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2688 3392 2740 3398
rect 2688 3334 2740 3340
rect 2884 2938 2912 5034
rect 2976 4826 3004 6802
rect 3160 6338 3188 7686
rect 3240 7472 3292 7478
rect 3240 7414 3292 7420
rect 3068 6310 3188 6338
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 3068 4570 3096 6310
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 2976 4542 3096 4570
rect 2976 3380 3004 4542
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 3068 3505 3096 4422
rect 3160 4078 3188 4762
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 3252 3754 3280 7414
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3344 5846 3372 6734
rect 3436 6118 3464 6802
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3332 5840 3384 5846
rect 3332 5782 3384 5788
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3332 3936 3384 3942
rect 3330 3904 3332 3913
rect 3384 3904 3386 3913
rect 3330 3839 3386 3848
rect 3252 3726 3372 3754
rect 3240 3528 3292 3534
rect 3054 3496 3110 3505
rect 3240 3470 3292 3476
rect 3054 3431 3110 3440
rect 2976 3352 3096 3380
rect 2962 3088 3018 3097
rect 2962 3023 3018 3032
rect 2700 2910 2912 2938
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 2700 480 2728 2910
rect 2976 2650 3004 3023
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3068 2514 3096 3352
rect 3148 2916 3200 2922
rect 3148 2858 3200 2864
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 3160 480 3188 2858
rect 202 0 258 480
rect 662 0 718 480
rect 1122 0 1178 480
rect 1674 0 1730 480
rect 2134 0 2190 480
rect 2686 0 2742 480
rect 3146 0 3202 480
rect 3252 241 3280 3470
rect 3344 1873 3372 3726
rect 3436 2990 3464 5510
rect 3528 3482 3556 9823
rect 3620 9081 3648 12106
rect 3804 10146 3832 12158
rect 3884 12164 3936 12170
rect 4066 12135 4122 12144
rect 4250 12200 4306 12209
rect 4250 12135 4306 12144
rect 3884 12106 3936 12112
rect 3921 11996 4217 12016
rect 3977 11994 4001 11996
rect 4057 11994 4081 11996
rect 4137 11994 4161 11996
rect 3999 11942 4001 11994
rect 4063 11942 4075 11994
rect 4137 11942 4139 11994
rect 3977 11940 4001 11942
rect 4057 11940 4081 11942
rect 4137 11940 4161 11942
rect 3921 11920 4217 11940
rect 4356 11694 4384 12582
rect 4632 12374 4660 13942
rect 4816 13530 4844 16520
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 5460 12986 5488 16520
rect 5632 15292 5684 15298
rect 5632 15234 5684 15240
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4620 12368 4672 12374
rect 4526 12336 4582 12345
rect 4620 12310 4672 12316
rect 4526 12271 4528 12280
rect 4580 12271 4582 12280
rect 4528 12242 4580 12248
rect 4632 11898 4660 12310
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4436 11552 4488 11558
rect 4436 11494 4488 11500
rect 4344 11008 4396 11014
rect 4344 10950 4396 10956
rect 3921 10908 4217 10928
rect 3977 10906 4001 10908
rect 4057 10906 4081 10908
rect 4137 10906 4161 10908
rect 3999 10854 4001 10906
rect 4063 10854 4075 10906
rect 4137 10854 4139 10906
rect 3977 10852 4001 10854
rect 4057 10852 4081 10854
rect 4137 10852 4161 10854
rect 3921 10832 4217 10852
rect 4356 10674 4384 10950
rect 4448 10810 4476 11494
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3712 10118 3832 10146
rect 3606 9072 3662 9081
rect 3606 9007 3662 9016
rect 3606 8528 3662 8537
rect 3606 8463 3608 8472
rect 3660 8463 3662 8472
rect 3608 8434 3660 8440
rect 3712 7936 3740 10118
rect 3896 10044 3924 10542
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 3620 7908 3740 7936
rect 3804 10016 3924 10044
rect 3620 7546 3648 7908
rect 3700 7812 3752 7818
rect 3700 7754 3752 7760
rect 3608 7540 3660 7546
rect 3608 7482 3660 7488
rect 3608 7200 3660 7206
rect 3608 7142 3660 7148
rect 3620 6769 3648 7142
rect 3606 6760 3662 6769
rect 3606 6695 3662 6704
rect 3606 6352 3662 6361
rect 3606 6287 3662 6296
rect 3620 3602 3648 6287
rect 3608 3596 3660 3602
rect 3608 3538 3660 3544
rect 3528 3454 3648 3482
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 3422 2680 3478 2689
rect 3422 2615 3424 2624
rect 3476 2615 3478 2624
rect 3424 2586 3476 2592
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 3330 1864 3386 1873
rect 3330 1799 3386 1808
rect 3528 1465 3556 2246
rect 3514 1456 3570 1465
rect 3514 1391 3570 1400
rect 3620 480 3648 3454
rect 3712 1057 3740 7754
rect 3804 7041 3832 10016
rect 3921 9820 4217 9840
rect 3977 9818 4001 9820
rect 4057 9818 4081 9820
rect 4137 9818 4161 9820
rect 3999 9766 4001 9818
rect 4063 9766 4075 9818
rect 4137 9766 4139 9818
rect 3977 9764 4001 9766
rect 4057 9764 4081 9766
rect 4137 9764 4161 9766
rect 3921 9744 4217 9764
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 3974 9344 4030 9353
rect 3974 9279 4030 9288
rect 3988 9110 4016 9279
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 4080 9042 4108 9454
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 4172 9353 4200 9386
rect 4158 9344 4214 9353
rect 4158 9279 4214 9288
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 4172 8945 4200 9279
rect 4158 8936 4214 8945
rect 4158 8871 4214 8880
rect 3921 8732 4217 8752
rect 3977 8730 4001 8732
rect 4057 8730 4081 8732
rect 4137 8730 4161 8732
rect 3999 8678 4001 8730
rect 4063 8678 4075 8730
rect 4137 8678 4139 8730
rect 3977 8676 4001 8678
rect 4057 8676 4081 8678
rect 4137 8676 4161 8678
rect 3921 8656 4217 8676
rect 3921 7644 4217 7664
rect 3977 7642 4001 7644
rect 4057 7642 4081 7644
rect 4137 7642 4161 7644
rect 3999 7590 4001 7642
rect 4063 7590 4075 7642
rect 4137 7590 4139 7642
rect 3977 7588 4001 7590
rect 4057 7588 4081 7590
rect 4137 7588 4161 7590
rect 3921 7568 4217 7588
rect 4160 7268 4212 7274
rect 4160 7210 4212 7216
rect 3790 7032 3846 7041
rect 3790 6967 3846 6976
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 3804 6458 3832 6802
rect 4172 6746 4200 7210
rect 3988 6730 4200 6746
rect 3976 6724 4200 6730
rect 4028 6718 4200 6724
rect 3976 6666 4028 6672
rect 3921 6556 4217 6576
rect 3977 6554 4001 6556
rect 4057 6554 4081 6556
rect 4137 6554 4161 6556
rect 3999 6502 4001 6554
rect 4063 6502 4075 6554
rect 4137 6502 4139 6554
rect 3977 6500 4001 6502
rect 4057 6500 4081 6502
rect 4137 6500 4161 6502
rect 3921 6480 4217 6500
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 3804 5710 3832 6394
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3921 5468 4217 5488
rect 3977 5466 4001 5468
rect 4057 5466 4081 5468
rect 4137 5466 4161 5468
rect 3999 5414 4001 5466
rect 4063 5414 4075 5466
rect 4137 5414 4139 5466
rect 3977 5412 4001 5414
rect 4057 5412 4081 5414
rect 4137 5412 4161 5414
rect 3921 5392 4217 5412
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4080 4826 4108 4966
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 3921 4380 4217 4400
rect 3977 4378 4001 4380
rect 4057 4378 4081 4380
rect 4137 4378 4161 4380
rect 3999 4326 4001 4378
rect 4063 4326 4075 4378
rect 4137 4326 4139 4378
rect 3977 4324 4001 4326
rect 4057 4324 4081 4326
rect 4137 4324 4161 4326
rect 3921 4304 4217 4324
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 3896 3738 3924 4014
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3921 3292 4217 3312
rect 3977 3290 4001 3292
rect 4057 3290 4081 3292
rect 4137 3290 4161 3292
rect 3999 3238 4001 3290
rect 4063 3238 4075 3290
rect 4137 3238 4139 3290
rect 3977 3236 4001 3238
rect 4057 3236 4081 3238
rect 4137 3236 4161 3238
rect 3921 3216 4217 3236
rect 4264 2990 4292 10406
rect 4724 10146 4752 12718
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4816 10266 4844 11086
rect 5170 10704 5226 10713
rect 5170 10639 5226 10648
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4436 10124 4488 10130
rect 4436 10066 4488 10072
rect 4632 10118 4752 10146
rect 4344 8424 4396 8430
rect 4344 8366 4396 8372
rect 4356 8022 4384 8366
rect 4344 8016 4396 8022
rect 4344 7958 4396 7964
rect 4448 7546 4476 10066
rect 4528 10056 4580 10062
rect 4528 9998 4580 10004
rect 4540 8634 4568 9998
rect 4528 8628 4580 8634
rect 4528 8570 4580 8576
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4540 7886 4568 8434
rect 4632 8090 4660 10118
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4724 8838 4752 9998
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4986 9344 5042 9353
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4632 7206 4660 8026
rect 4712 7880 4764 7886
rect 4710 7848 4712 7857
rect 4764 7848 4766 7857
rect 4710 7783 4766 7792
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4724 7410 4752 7686
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4436 6248 4488 6254
rect 4436 6190 4488 6196
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4448 6118 4476 6190
rect 4620 6180 4672 6186
rect 4620 6122 4672 6128
rect 4436 6112 4488 6118
rect 4488 6072 4568 6100
rect 4436 6054 4488 6060
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 4356 4282 4384 5646
rect 4448 5370 4476 5714
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4540 5166 4568 6072
rect 4632 5710 4660 6122
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4724 5234 4752 6190
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4448 4146 4476 4422
rect 4540 4282 4568 5102
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4540 3670 4568 4218
rect 4724 4214 4752 5170
rect 4816 4690 4844 9318
rect 4986 9279 5042 9288
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 4908 8498 4936 8978
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4908 7750 4936 8434
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 4908 7410 4936 7686
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4896 5704 4948 5710
rect 4896 5646 4948 5652
rect 4908 5166 4936 5646
rect 4896 5160 4948 5166
rect 4896 5102 4948 5108
rect 5000 4690 5028 9279
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5092 7546 5120 8230
rect 5184 7857 5212 10639
rect 5276 9654 5304 11154
rect 5264 9648 5316 9654
rect 5264 9590 5316 9596
rect 5262 9480 5318 9489
rect 5262 9415 5318 9424
rect 5170 7848 5226 7857
rect 5170 7783 5226 7792
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5080 5092 5132 5098
rect 5080 5034 5132 5040
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 4528 3664 4580 3670
rect 4528 3606 4580 3612
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 4252 2984 4304 2990
rect 4252 2926 4304 2932
rect 3921 2204 4217 2224
rect 3977 2202 4001 2204
rect 4057 2202 4081 2204
rect 4137 2202 4161 2204
rect 3999 2150 4001 2202
rect 4063 2150 4075 2202
rect 4137 2150 4139 2202
rect 3977 2148 4001 2150
rect 4057 2148 4081 2150
rect 4137 2148 4161 2150
rect 3921 2128 4217 2148
rect 4540 1306 4568 2994
rect 4172 1278 4568 1306
rect 3698 1048 3754 1057
rect 3698 983 3754 992
rect 3700 740 3752 746
rect 3700 682 3752 688
rect 3712 649 3740 682
rect 3698 640 3754 649
rect 3698 575 3754 584
rect 4172 480 4200 1278
rect 4632 480 4660 3538
rect 4816 2514 4844 4626
rect 5092 4622 5120 5034
rect 5276 4826 5304 9415
rect 5368 8242 5396 11698
rect 5552 11642 5580 14010
rect 5460 11614 5580 11642
rect 5644 11626 5672 15234
rect 6104 13870 6132 16520
rect 6748 14090 6776 16520
rect 6886 14716 7182 14736
rect 6942 14714 6966 14716
rect 7022 14714 7046 14716
rect 7102 14714 7126 14716
rect 6964 14662 6966 14714
rect 7028 14662 7040 14714
rect 7102 14662 7104 14714
rect 6942 14660 6966 14662
rect 7022 14660 7046 14662
rect 7102 14660 7126 14662
rect 6886 14640 7182 14660
rect 6748 14074 6960 14090
rect 6748 14068 6972 14074
rect 6748 14062 6920 14068
rect 6920 14010 6972 14016
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 7392 13802 7420 16520
rect 5908 13796 5960 13802
rect 5908 13738 5960 13744
rect 7380 13796 7432 13802
rect 7380 13738 7432 13744
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 5632 11620 5684 11626
rect 5460 11234 5488 11614
rect 5632 11562 5684 11568
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5552 11354 5580 11494
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5460 11206 5672 11234
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5460 9722 5488 10746
rect 5552 10606 5580 10950
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5538 10160 5594 10169
rect 5538 10095 5594 10104
rect 5448 9716 5500 9722
rect 5448 9658 5500 9664
rect 5446 9616 5502 9625
rect 5446 9551 5502 9560
rect 5460 9382 5488 9551
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5552 8634 5580 10095
rect 5644 9450 5672 11206
rect 5736 9586 5764 12582
rect 5828 11898 5856 12582
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 5828 11762 5856 11834
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5920 11370 5948 13738
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6092 12844 6144 12850
rect 6092 12786 6144 12792
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 6012 12102 6040 12582
rect 6104 12442 6132 12786
rect 6092 12436 6144 12442
rect 6092 12378 6144 12384
rect 6090 12336 6146 12345
rect 6090 12271 6146 12280
rect 6104 12238 6132 12271
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 5828 11342 5948 11370
rect 5828 10690 5856 11342
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 5920 10810 5948 11154
rect 6012 11082 6040 12038
rect 6090 11792 6146 11801
rect 6090 11727 6092 11736
rect 6144 11727 6146 11736
rect 6092 11698 6144 11704
rect 6000 11076 6052 11082
rect 6000 11018 6052 11024
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 5828 10662 5948 10690
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5828 10266 5856 10542
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5632 9444 5684 9450
rect 5632 9386 5684 9392
rect 5828 9178 5856 9998
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5724 9104 5776 9110
rect 5724 9046 5776 9052
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5368 8214 5580 8242
rect 5446 7984 5502 7993
rect 5446 7919 5502 7928
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5368 5710 5396 7822
rect 5460 7818 5488 7919
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5460 7002 5488 7346
rect 5552 7188 5580 8214
rect 5644 7342 5672 8298
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5736 7206 5764 9046
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5724 7200 5776 7206
rect 5552 7160 5672 7188
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 5552 5778 5580 6326
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5356 5704 5408 5710
rect 5644 5658 5672 7160
rect 5724 7142 5776 7148
rect 5828 7018 5856 7482
rect 5356 5646 5408 5652
rect 5552 5630 5672 5658
rect 5736 6990 5856 7018
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5552 4690 5580 5630
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5644 4826 5672 4966
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5460 3466 5488 4558
rect 5540 4004 5592 4010
rect 5736 3992 5764 6990
rect 5592 3964 5764 3992
rect 5816 4004 5868 4010
rect 5540 3946 5592 3952
rect 5816 3946 5868 3952
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 5552 2582 5580 3946
rect 5828 2990 5856 3946
rect 5816 2984 5868 2990
rect 5816 2926 5868 2932
rect 5920 2802 5948 10662
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 6012 10062 6040 10610
rect 6092 10532 6144 10538
rect 6092 10474 6144 10480
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 6012 9586 6040 9998
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 6012 7954 6040 8434
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 6012 7410 6040 7890
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 6012 5778 6040 6054
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 6012 4690 6040 5170
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 6012 4078 6040 4626
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 6104 3058 6132 10474
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 5644 2774 5948 2802
rect 5540 2576 5592 2582
rect 5540 2518 5592 2524
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 4988 2304 5040 2310
rect 4988 2246 5040 2252
rect 5000 746 5028 2246
rect 5172 1352 5224 1358
rect 5172 1294 5224 1300
rect 4988 740 5040 746
rect 4988 682 5040 688
rect 5184 480 5212 1294
rect 5644 480 5672 2774
rect 6196 480 6224 13670
rect 6886 13628 7182 13648
rect 6942 13626 6966 13628
rect 7022 13626 7046 13628
rect 7102 13626 7126 13628
rect 6964 13574 6966 13626
rect 7028 13574 7040 13626
rect 7102 13574 7104 13626
rect 6942 13572 6966 13574
rect 7022 13572 7046 13574
rect 7102 13572 7126 13574
rect 6886 13552 7182 13572
rect 8036 12782 8064 16520
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8128 12782 8156 13126
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 8024 12776 8076 12782
rect 8024 12718 8076 12724
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 6886 12540 7182 12560
rect 6942 12538 6966 12540
rect 7022 12538 7046 12540
rect 7102 12538 7126 12540
rect 6964 12486 6966 12538
rect 7028 12486 7040 12538
rect 7102 12486 7104 12538
rect 6942 12484 6966 12486
rect 7022 12484 7046 12486
rect 7102 12484 7126 12486
rect 6886 12464 7182 12484
rect 6552 12436 6604 12442
rect 6552 12378 6604 12384
rect 6276 12368 6328 12374
rect 6274 12336 6276 12345
rect 6328 12336 6330 12345
rect 6274 12271 6330 12280
rect 6564 12288 6592 12378
rect 6644 12300 6696 12306
rect 6288 10470 6316 12271
rect 6564 12260 6644 12288
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6380 11694 6408 12174
rect 6458 11792 6514 11801
rect 6458 11727 6514 11736
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 6368 11076 6420 11082
rect 6368 11018 6420 11024
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6288 9897 6316 10066
rect 6274 9888 6330 9897
rect 6274 9823 6330 9832
rect 6276 9512 6328 9518
rect 6276 9454 6328 9460
rect 6288 9382 6316 9454
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6276 9104 6328 9110
rect 6276 9046 6328 9052
rect 6288 8022 6316 9046
rect 6380 8537 6408 11018
rect 6472 9489 6500 11727
rect 6458 9480 6514 9489
rect 6458 9415 6514 9424
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6366 8528 6422 8537
rect 6366 8463 6422 8472
rect 6276 8016 6328 8022
rect 6276 7958 6328 7964
rect 6288 7342 6316 7958
rect 6276 7336 6328 7342
rect 6368 7336 6420 7342
rect 6276 7278 6328 7284
rect 6366 7304 6368 7313
rect 6420 7304 6422 7313
rect 6366 7239 6422 7248
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6288 6458 6316 6802
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6288 5302 6316 6258
rect 6276 5296 6328 5302
rect 6276 5238 6328 5244
rect 6380 4706 6408 7142
rect 6472 6254 6500 9318
rect 6564 8974 6592 12260
rect 6644 12242 6696 12248
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6748 11762 6776 12038
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6748 11626 6776 11698
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 6644 11076 6696 11082
rect 6644 11018 6696 11024
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6460 6248 6512 6254
rect 6460 6190 6512 6196
rect 6564 6186 6592 6734
rect 6552 6180 6604 6186
rect 6552 6122 6604 6128
rect 6288 4678 6408 4706
rect 6460 4684 6512 4690
rect 6288 4214 6316 4678
rect 6460 4626 6512 4632
rect 6368 4616 6420 4622
rect 6472 4593 6500 4626
rect 6368 4558 6420 4564
rect 6458 4584 6514 4593
rect 6276 4208 6328 4214
rect 6276 4150 6328 4156
rect 6380 4146 6408 4558
rect 6458 4519 6514 4528
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 6288 3398 6316 4014
rect 6564 4010 6592 4218
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6564 2990 6592 3334
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 6656 480 6684 11018
rect 6748 10674 6776 11562
rect 6886 11452 7182 11472
rect 6942 11450 6966 11452
rect 7022 11450 7046 11452
rect 7102 11450 7126 11452
rect 6964 11398 6966 11450
rect 7028 11398 7040 11450
rect 7102 11398 7104 11450
rect 6942 11396 6966 11398
rect 7022 11396 7046 11398
rect 7102 11396 7126 11398
rect 6886 11376 7182 11396
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 7116 10606 7144 10746
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7208 10452 7236 11154
rect 7300 10606 7328 12582
rect 7656 12300 7708 12306
rect 7656 12242 7708 12248
rect 7470 12200 7526 12209
rect 7470 12135 7526 12144
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7208 10424 7328 10452
rect 6886 10364 7182 10384
rect 6942 10362 6966 10364
rect 7022 10362 7046 10364
rect 7102 10362 7126 10364
rect 6964 10310 6966 10362
rect 7028 10310 7040 10362
rect 7102 10310 7104 10362
rect 6942 10308 6966 10310
rect 7022 10308 7046 10310
rect 7102 10308 7126 10310
rect 6734 10296 6790 10305
rect 6886 10288 7182 10308
rect 7300 10282 7328 10424
rect 7300 10254 7420 10282
rect 6734 10231 6790 10240
rect 6748 10062 6776 10231
rect 7288 10192 7340 10198
rect 7288 10134 7340 10140
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6748 8498 6776 9862
rect 6932 9586 6960 9930
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6886 9276 7182 9296
rect 6942 9274 6966 9276
rect 7022 9274 7046 9276
rect 7102 9274 7126 9276
rect 6964 9222 6966 9274
rect 7028 9222 7040 9274
rect 7102 9222 7104 9274
rect 6942 9220 6966 9222
rect 7022 9220 7046 9222
rect 7102 9220 7126 9222
rect 6886 9200 7182 9220
rect 7300 9178 7328 10134
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7194 8936 7250 8945
rect 7194 8871 7250 8880
rect 7208 8634 7236 8871
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 6748 7546 6776 8434
rect 6886 8188 7182 8208
rect 6942 8186 6966 8188
rect 7022 8186 7046 8188
rect 7102 8186 7126 8188
rect 6964 8134 6966 8186
rect 7028 8134 7040 8186
rect 7102 8134 7104 8186
rect 6942 8132 6966 8134
rect 7022 8132 7046 8134
rect 7102 8132 7126 8134
rect 6886 8112 7182 8132
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 7208 7546 7236 7890
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7300 7206 7328 8434
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 6886 7100 7182 7120
rect 6942 7098 6966 7100
rect 7022 7098 7046 7100
rect 7102 7098 7126 7100
rect 6964 7046 6966 7098
rect 7028 7046 7040 7098
rect 7102 7046 7104 7098
rect 6942 7044 6966 7046
rect 7022 7044 7046 7046
rect 7102 7044 7126 7046
rect 6886 7024 7182 7044
rect 7392 6202 7420 10254
rect 7484 10130 7512 12135
rect 7571 11212 7623 11218
rect 7571 11154 7623 11160
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 7576 10062 7604 11154
rect 7564 10056 7616 10062
rect 7470 10024 7526 10033
rect 7564 9998 7616 10004
rect 7470 9959 7526 9968
rect 7484 9874 7512 9959
rect 7484 9846 7604 9874
rect 7470 9344 7526 9353
rect 7576 9330 7604 9846
rect 7526 9302 7604 9330
rect 7470 9279 7526 9288
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7484 8294 7512 9114
rect 7576 8498 7604 9302
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7472 8288 7524 8294
rect 7576 8265 7604 8298
rect 7472 8230 7524 8236
rect 7562 8256 7618 8265
rect 7484 8090 7512 8230
rect 7562 8191 7618 8200
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7472 6724 7524 6730
rect 7472 6666 7524 6672
rect 7300 6174 7420 6202
rect 6886 6012 7182 6032
rect 6942 6010 6966 6012
rect 7022 6010 7046 6012
rect 7102 6010 7126 6012
rect 6964 5958 6966 6010
rect 7028 5958 7040 6010
rect 7102 5958 7104 6010
rect 6942 5956 6966 5958
rect 7022 5956 7046 5958
rect 7102 5956 7126 5958
rect 6886 5936 7182 5956
rect 7300 5302 7328 6174
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7392 5846 7420 6054
rect 7380 5840 7432 5846
rect 7380 5782 7432 5788
rect 7288 5296 7340 5302
rect 7288 5238 7340 5244
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6748 2990 6776 5102
rect 6886 4924 7182 4944
rect 6942 4922 6966 4924
rect 7022 4922 7046 4924
rect 7102 4922 7126 4924
rect 6964 4870 6966 4922
rect 7028 4870 7040 4922
rect 7102 4870 7104 4922
rect 6942 4868 6966 4870
rect 7022 4868 7046 4870
rect 7102 4868 7126 4870
rect 6886 4848 7182 4868
rect 6918 4720 6974 4729
rect 6918 4655 6974 4664
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6840 4146 6868 4558
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6932 4010 6960 4655
rect 7300 4298 7328 5238
rect 7392 5166 7420 5782
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 7484 4729 7512 6666
rect 7470 4720 7526 4729
rect 7470 4655 7526 4664
rect 7300 4270 7512 4298
rect 6920 4004 6972 4010
rect 6920 3946 6972 3952
rect 7288 4004 7340 4010
rect 7288 3946 7340 3952
rect 6886 3836 7182 3856
rect 6942 3834 6966 3836
rect 7022 3834 7046 3836
rect 7102 3834 7126 3836
rect 6964 3782 6966 3834
rect 7028 3782 7040 3834
rect 7102 3782 7104 3834
rect 6942 3780 6966 3782
rect 7022 3780 7046 3782
rect 7102 3780 7126 3782
rect 6886 3760 7182 3780
rect 7300 3738 7328 3946
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7300 2990 7328 3674
rect 7380 3664 7432 3670
rect 7380 3606 7432 3612
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 6748 2378 6776 2926
rect 6886 2748 7182 2768
rect 6942 2746 6966 2748
rect 7022 2746 7046 2748
rect 7102 2746 7126 2748
rect 6964 2694 6966 2746
rect 7028 2694 7040 2746
rect 7102 2694 7104 2746
rect 6942 2692 6966 2694
rect 7022 2692 7046 2694
rect 7102 2692 7126 2694
rect 6886 2672 7182 2692
rect 7392 2514 7420 3606
rect 7484 3534 7512 4270
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7484 2990 7512 3470
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7576 2922 7604 7686
rect 7668 7002 7696 12242
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7760 7857 7788 10746
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7746 7848 7802 7857
rect 7746 7783 7802 7792
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7668 6322 7696 6734
rect 7760 6322 7788 7783
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7748 6180 7800 6186
rect 7748 6122 7800 6128
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7668 3670 7696 5510
rect 7760 3738 7788 6122
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7852 3516 7880 10406
rect 7932 9376 7984 9382
rect 7930 9344 7932 9353
rect 7984 9344 7986 9353
rect 7930 9279 7986 9288
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 7944 8945 7972 9114
rect 7930 8936 7986 8945
rect 7930 8871 7986 8880
rect 7932 8832 7984 8838
rect 7932 8774 7984 8780
rect 7944 8362 7972 8774
rect 7932 8356 7984 8362
rect 7932 8298 7984 8304
rect 7930 8120 7986 8129
rect 7930 8055 7986 8064
rect 7668 3488 7880 3516
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 7380 2508 7432 2514
rect 7380 2450 7432 2456
rect 6736 2372 6788 2378
rect 6736 2314 6788 2320
rect 7104 1148 7156 1154
rect 7104 1090 7156 1096
rect 7116 480 7144 1090
rect 7668 480 7696 3488
rect 7944 1154 7972 8055
rect 8036 6361 8064 12718
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 8128 7868 8156 12038
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8220 11286 8248 11494
rect 8208 11280 8260 11286
rect 8208 11222 8260 11228
rect 8300 11280 8352 11286
rect 8300 11222 8352 11228
rect 8312 10577 8340 11222
rect 8392 10736 8444 10742
rect 8392 10678 8444 10684
rect 8298 10568 8354 10577
rect 8298 10503 8354 10512
rect 8404 10198 8432 10678
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8220 8498 8248 9454
rect 8496 8838 8524 12786
rect 8680 12481 8708 16520
rect 8760 14816 8812 14822
rect 8760 14758 8812 14764
rect 8772 12850 8800 14758
rect 9324 13802 9352 16520
rect 9402 15464 9458 15473
rect 9402 15399 9458 15408
rect 9036 13796 9088 13802
rect 9036 13738 9088 13744
rect 9312 13796 9364 13802
rect 9312 13738 9364 13744
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8666 12472 8722 12481
rect 8666 12407 8722 12416
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 8680 11898 8708 12174
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8666 11112 8722 11121
rect 8666 11047 8722 11056
rect 8680 10606 8708 11047
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 8772 9654 8800 12174
rect 8852 11892 8904 11898
rect 8852 11834 8904 11840
rect 8864 11801 8892 11834
rect 8850 11792 8906 11801
rect 8850 11727 8906 11736
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8864 10577 8892 11494
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8850 10568 8906 10577
rect 8850 10503 8906 10512
rect 8864 10044 8892 10503
rect 8956 10198 8984 10950
rect 8944 10192 8996 10198
rect 8944 10134 8996 10140
rect 8864 10016 8984 10044
rect 8760 9648 8812 9654
rect 8680 9608 8760 9636
rect 8680 8922 8708 9608
rect 8760 9590 8812 9596
rect 8850 9616 8906 9625
rect 8850 9551 8906 9560
rect 8864 9382 8892 9551
rect 8760 9376 8812 9382
rect 8758 9344 8760 9353
rect 8852 9376 8904 9382
rect 8812 9344 8814 9353
rect 8852 9318 8904 9324
rect 8758 9279 8814 9288
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 8864 8945 8892 9114
rect 8588 8894 8708 8922
rect 8850 8936 8906 8945
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8588 8786 8616 8894
rect 8850 8871 8906 8880
rect 8852 8832 8904 8838
rect 8758 8800 8814 8809
rect 8588 8758 8708 8786
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8312 8072 8340 8570
rect 8312 8044 8432 8072
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8208 7880 8260 7886
rect 8128 7840 8208 7868
rect 8208 7822 8260 7828
rect 8206 7576 8262 7585
rect 8206 7511 8262 7520
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8128 6458 8156 6734
rect 8220 6730 8248 7511
rect 8312 7002 8340 7890
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8022 6352 8078 6361
rect 8022 6287 8078 6296
rect 8404 6254 8432 8044
rect 8484 7880 8536 7886
rect 8680 7834 8708 8758
rect 8852 8774 8904 8780
rect 8758 8735 8814 8744
rect 8484 7822 8536 7828
rect 8496 7002 8524 7822
rect 8588 7806 8708 7834
rect 8588 7274 8616 7806
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8680 7449 8708 7686
rect 8666 7440 8722 7449
rect 8666 7375 8722 7384
rect 8576 7268 8628 7274
rect 8576 7210 8628 7216
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8588 6390 8616 7210
rect 8484 6384 8536 6390
rect 8484 6326 8536 6332
rect 8576 6384 8628 6390
rect 8576 6326 8628 6332
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 8116 5636 8168 5642
rect 8116 5578 8168 5584
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 8036 5302 8064 5510
rect 8024 5296 8076 5302
rect 8024 5238 8076 5244
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 8036 4758 8064 5102
rect 8024 4752 8076 4758
rect 8024 4694 8076 4700
rect 8024 3664 8076 3670
rect 8024 3606 8076 3612
rect 8036 1358 8064 3606
rect 8024 1352 8076 1358
rect 8024 1294 8076 1300
rect 7932 1148 7984 1154
rect 7932 1090 7984 1096
rect 8128 480 8156 5578
rect 8312 5370 8340 6122
rect 8496 5574 8524 6326
rect 8588 5914 8616 6326
rect 8772 6254 8800 8735
rect 8864 8294 8892 8774
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 8864 6100 8892 7890
rect 8772 6072 8892 6100
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 8220 4593 8248 4966
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8206 4584 8262 4593
rect 8206 4519 8262 4528
rect 8392 4208 8444 4214
rect 8392 4150 8444 4156
rect 8404 3466 8432 4150
rect 8496 3942 8524 4626
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 8392 3460 8444 3466
rect 8392 3402 8444 3408
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8220 2650 8248 2994
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 8298 2544 8354 2553
rect 8298 2479 8300 2488
rect 8352 2479 8354 2488
rect 8300 2450 8352 2456
rect 8404 2378 8432 3402
rect 8496 2514 8524 3878
rect 8576 2916 8628 2922
rect 8576 2858 8628 2864
rect 8588 2825 8616 2858
rect 8574 2816 8630 2825
rect 8574 2751 8630 2760
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 8680 480 8708 3878
rect 8772 3738 8800 6072
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 8864 4826 8892 5850
rect 8956 5642 8984 10016
rect 9048 5710 9076 13738
rect 9128 12368 9180 12374
rect 9128 12310 9180 12316
rect 9310 12336 9366 12345
rect 9140 10169 9168 12310
rect 9416 12306 9444 15399
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9310 12271 9366 12280
rect 9404 12300 9456 12306
rect 9324 12238 9352 12271
rect 9404 12242 9456 12248
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9416 12170 9444 12242
rect 9404 12164 9456 12170
rect 9404 12106 9456 12112
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9232 11286 9260 11494
rect 9220 11280 9272 11286
rect 9220 11222 9272 11228
rect 9126 10160 9182 10169
rect 9126 10095 9182 10104
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 9140 8673 9168 9590
rect 9126 8664 9182 8673
rect 9126 8599 9182 8608
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9140 7041 9168 7822
rect 9126 7032 9182 7041
rect 9126 6967 9182 6976
rect 9128 6928 9180 6934
rect 9128 6870 9180 6876
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 8944 5636 8996 5642
rect 8944 5578 8996 5584
rect 9048 5216 9076 5646
rect 8956 5188 9076 5216
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8956 4622 8984 5188
rect 9036 5092 9088 5098
rect 9036 5034 9088 5040
rect 9048 4826 9076 5034
rect 9140 4826 9168 6870
rect 9232 5030 9260 11222
rect 9324 9994 9352 11698
rect 9312 9988 9364 9994
rect 9312 9930 9364 9936
rect 9404 9988 9456 9994
rect 9404 9930 9456 9936
rect 9324 9586 9352 9930
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9416 9364 9444 9930
rect 9496 9920 9548 9926
rect 9494 9888 9496 9897
rect 9548 9888 9550 9897
rect 9494 9823 9550 9832
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9324 9336 9444 9364
rect 9324 7993 9352 9336
rect 9404 8968 9456 8974
rect 9508 8945 9536 9522
rect 9404 8910 9456 8916
rect 9494 8936 9550 8945
rect 9416 8673 9444 8910
rect 9494 8871 9550 8880
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9402 8664 9458 8673
rect 9402 8599 9458 8608
rect 9508 8129 9536 8774
rect 9494 8120 9550 8129
rect 9404 8084 9456 8090
rect 9494 8055 9550 8064
rect 9404 8026 9456 8032
rect 9310 7984 9366 7993
rect 9310 7919 9366 7928
rect 9312 7812 9364 7818
rect 9312 7754 9364 7760
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 8956 4214 8984 4558
rect 8944 4208 8996 4214
rect 8944 4150 8996 4156
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 9048 3602 9076 4762
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 8772 2650 8800 2858
rect 8760 2644 8812 2650
rect 8760 2586 8812 2592
rect 8956 2582 8984 3334
rect 8944 2576 8996 2582
rect 8944 2518 8996 2524
rect 9140 480 9168 4422
rect 9324 3942 9352 7754
rect 9416 7410 9444 8026
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9508 7478 9536 7686
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9416 7002 9444 7346
rect 9508 7342 9536 7414
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9404 6996 9456 7002
rect 9404 6938 9456 6944
rect 9508 6798 9536 7278
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9508 5370 9536 5714
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9496 5024 9548 5030
rect 9494 4992 9496 5001
rect 9548 4992 9550 5001
rect 9494 4927 9550 4936
rect 9496 4548 9548 4554
rect 9496 4490 9548 4496
rect 9508 4282 9536 4490
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9600 2922 9628 14418
rect 9968 14362 9996 16520
rect 9968 14334 10272 14362
rect 9852 14172 10148 14192
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 9930 14118 9932 14170
rect 9994 14118 10006 14170
rect 10068 14118 10070 14170
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 9852 14096 10148 14116
rect 10244 13190 10272 14334
rect 10324 13796 10376 13802
rect 10324 13738 10376 13744
rect 10232 13184 10284 13190
rect 10232 13126 10284 13132
rect 9852 13084 10148 13104
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 9930 13030 9932 13082
rect 9994 13030 10006 13082
rect 10068 13030 10070 13082
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 9852 13008 10148 13028
rect 9852 11996 10148 12016
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 9930 11942 9932 11994
rect 9994 11942 10006 11994
rect 10068 11942 10070 11994
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 9852 11920 10148 11940
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 9852 10908 10148 10928
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 9930 10854 9932 10906
rect 9994 10854 10006 10906
rect 10068 10854 10070 10906
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 9852 10832 10148 10852
rect 10244 10810 10272 11086
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 9770 10704 9826 10713
rect 9770 10639 9826 10648
rect 9784 9994 9812 10639
rect 10138 10296 10194 10305
rect 10138 10231 10194 10240
rect 10152 10130 10180 10231
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9680 9376 9732 9382
rect 9678 9344 9680 9353
rect 9732 9344 9734 9353
rect 9678 9279 9734 9288
rect 9784 9110 9812 9930
rect 9852 9820 10148 9840
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 9930 9766 9932 9818
rect 9994 9766 10006 9818
rect 10068 9766 10070 9818
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 9852 9744 10148 9764
rect 10244 9704 10272 10066
rect 9876 9676 10272 9704
rect 9680 9104 9732 9110
rect 9680 9046 9732 9052
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 9692 8945 9720 9046
rect 9678 8936 9734 8945
rect 9876 8888 9904 9676
rect 10336 9602 10364 13738
rect 10612 13138 10640 16520
rect 11256 13734 11284 16520
rect 11900 13802 11928 16520
rect 12072 15224 12124 15230
rect 12072 15166 12124 15172
rect 11336 13796 11388 13802
rect 11336 13738 11388 13744
rect 11888 13796 11940 13802
rect 11888 13738 11940 13744
rect 11980 13796 12032 13802
rect 11980 13738 12032 13744
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 10612 13110 11008 13138
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10508 11076 10560 11082
rect 10508 11018 10560 11024
rect 10416 11008 10468 11014
rect 10416 10950 10468 10956
rect 10428 10674 10456 10950
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10428 10062 10456 10406
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10244 9574 10364 9602
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 10060 9382 10088 9454
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 9678 8871 9734 8880
rect 9784 8860 9904 8888
rect 9784 8616 9812 8860
rect 9852 8732 10148 8752
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 9930 8678 9932 8730
rect 9994 8678 10006 8730
rect 10068 8678 10070 8730
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 9852 8656 10148 8676
rect 9784 8588 10088 8616
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9968 8129 9996 8366
rect 9954 8120 10010 8129
rect 9954 8055 10010 8064
rect 10060 8022 10088 8588
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9692 7342 9720 7686
rect 9852 7644 10148 7664
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 9930 7590 9932 7642
rect 9994 7590 10006 7642
rect 10068 7590 10070 7642
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 9852 7568 10148 7588
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 9692 7206 9720 7278
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9692 6458 9720 7142
rect 9876 6934 9904 7142
rect 9864 6928 9916 6934
rect 9864 6870 9916 6876
rect 9956 6928 10008 6934
rect 9956 6870 10008 6876
rect 9968 6730 9996 6870
rect 10060 6730 10088 7278
rect 10138 7168 10194 7177
rect 10138 7103 10194 7112
rect 10152 6866 10180 7103
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 9956 6724 10008 6730
rect 9956 6666 10008 6672
rect 10048 6724 10100 6730
rect 10048 6666 10100 6672
rect 9852 6556 10148 6576
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 9930 6502 9932 6554
rect 9994 6502 10006 6554
rect 10068 6502 10070 6554
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 9852 6480 10148 6500
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9692 5710 9720 6394
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9692 5234 9720 5646
rect 9852 5468 10148 5488
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 9930 5414 9932 5466
rect 9994 5414 10006 5466
rect 10068 5414 10070 5466
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 9852 5392 10148 5412
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9784 3466 9812 4422
rect 9852 4380 10148 4400
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 9930 4326 9932 4378
rect 9994 4326 10006 4378
rect 10068 4326 10070 4378
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 9852 4304 10148 4324
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9876 3670 9904 3878
rect 9864 3664 9916 3670
rect 9864 3606 9916 3612
rect 10060 3466 10088 4082
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 9852 3292 10148 3312
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 9930 3238 9932 3290
rect 9994 3238 10006 3290
rect 10068 3238 10070 3290
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 9852 3216 10148 3236
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9588 2916 9640 2922
rect 9588 2858 9640 2864
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 9232 2650 9260 2790
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 9692 480 9720 3130
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 9784 1442 9812 3062
rect 10244 2582 10272 9574
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10336 6730 10364 9318
rect 10324 6724 10376 6730
rect 10324 6666 10376 6672
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10336 5778 10364 6394
rect 10428 6254 10456 9998
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 10336 5574 10364 5714
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10428 5166 10456 5510
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10324 5092 10376 5098
rect 10324 5034 10376 5040
rect 10336 4078 10364 5034
rect 10428 4282 10456 5102
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10324 4072 10376 4078
rect 10324 4014 10376 4020
rect 10520 3670 10548 11018
rect 10612 10130 10640 12718
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10612 9178 10640 9522
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10612 7274 10640 9114
rect 10704 9042 10732 11154
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10796 10810 10824 10950
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10796 10554 10824 10746
rect 10888 10742 10916 11154
rect 10876 10736 10928 10742
rect 10876 10678 10928 10684
rect 10796 10526 10916 10554
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10796 10198 10824 10406
rect 10784 10192 10836 10198
rect 10784 10134 10836 10140
rect 10888 9042 10916 10526
rect 10692 9036 10744 9042
rect 10876 9036 10928 9042
rect 10744 8996 10824 9024
rect 10692 8978 10744 8984
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10704 7750 10732 8298
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10704 7449 10732 7686
rect 10690 7440 10746 7449
rect 10690 7375 10746 7384
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10612 6390 10640 6734
rect 10692 6724 10744 6730
rect 10692 6666 10744 6672
rect 10600 6384 10652 6390
rect 10600 6326 10652 6332
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 10416 3460 10468 3466
rect 10416 3402 10468 3408
rect 10322 2952 10378 2961
rect 10428 2922 10456 3402
rect 10612 3176 10640 6190
rect 10704 5846 10732 6666
rect 10796 6254 10824 8996
rect 10876 8978 10928 8984
rect 10888 8129 10916 8978
rect 10874 8120 10930 8129
rect 10874 8055 10930 8064
rect 10876 8016 10928 8022
rect 10876 7958 10928 7964
rect 10888 6798 10916 7958
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 10692 5704 10744 5710
rect 10692 5646 10744 5652
rect 10704 5114 10732 5646
rect 10784 5636 10836 5642
rect 10784 5578 10836 5584
rect 10796 5370 10824 5578
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10704 5086 10824 5114
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10704 4690 10732 4966
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 10704 4010 10732 4626
rect 10692 4004 10744 4010
rect 10692 3946 10744 3952
rect 10796 3618 10824 5086
rect 10520 3148 10640 3176
rect 10704 3590 10824 3618
rect 10322 2887 10324 2896
rect 10376 2887 10378 2896
rect 10416 2916 10468 2922
rect 10324 2858 10376 2864
rect 10416 2858 10468 2864
rect 10520 2582 10548 3148
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10232 2576 10284 2582
rect 10508 2576 10560 2582
rect 10232 2518 10284 2524
rect 10506 2544 10508 2553
rect 10560 2544 10562 2553
rect 10506 2479 10562 2488
rect 9852 2204 10148 2224
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 9930 2150 9932 2202
rect 9994 2150 10006 2202
rect 10068 2150 10070 2202
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 9852 2128 10148 2148
rect 9784 1414 10180 1442
rect 10152 480 10180 1414
rect 10612 480 10640 2994
rect 10704 2582 10732 3590
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 10796 3398 10824 3470
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10796 2961 10824 3334
rect 10782 2952 10838 2961
rect 10782 2887 10838 2896
rect 10692 2576 10744 2582
rect 10692 2518 10744 2524
rect 10980 2530 11008 13110
rect 11242 12200 11298 12209
rect 11242 12135 11298 12144
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 11072 10305 11100 10406
rect 11058 10296 11114 10305
rect 11058 10231 11114 10240
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 11072 9654 11100 10066
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 11164 9518 11192 11494
rect 11256 10674 11284 12135
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11152 9512 11204 9518
rect 11152 9454 11204 9460
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11150 8936 11206 8945
rect 11150 8871 11206 8880
rect 11058 8664 11114 8673
rect 11058 8599 11114 8608
rect 11072 7002 11100 8599
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 11164 3058 11192 8871
rect 11256 8430 11284 9318
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11256 7818 11284 8230
rect 11244 7812 11296 7818
rect 11244 7754 11296 7760
rect 11242 7304 11298 7313
rect 11242 7239 11298 7248
rect 11152 3052 11204 3058
rect 11072 3012 11152 3040
rect 11072 2825 11100 3012
rect 11152 2994 11204 3000
rect 11152 2848 11204 2854
rect 11058 2816 11114 2825
rect 11152 2790 11204 2796
rect 11058 2751 11114 2760
rect 10704 2310 10732 2518
rect 10980 2502 11100 2530
rect 11072 2446 11100 2502
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 10692 2304 10744 2310
rect 10692 2246 10744 2252
rect 11164 480 11192 2790
rect 11256 2496 11284 7239
rect 11348 5846 11376 13738
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11428 13252 11480 13258
rect 11428 13194 11480 13200
rect 11440 12714 11468 13194
rect 11428 12708 11480 12714
rect 11428 12650 11480 12656
rect 11704 12708 11756 12714
rect 11704 12650 11756 12656
rect 11336 5840 11388 5846
rect 11336 5782 11388 5788
rect 11440 3466 11468 12650
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 11428 3460 11480 3466
rect 11428 3402 11480 3408
rect 11532 2582 11560 12378
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11624 11121 11652 12242
rect 11716 11150 11744 12650
rect 11704 11144 11756 11150
rect 11610 11112 11666 11121
rect 11704 11086 11756 11092
rect 11610 11047 11666 11056
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11624 10538 11652 10950
rect 11612 10532 11664 10538
rect 11612 10474 11664 10480
rect 11704 10532 11756 10538
rect 11704 10474 11756 10480
rect 11624 10062 11652 10474
rect 11612 10056 11664 10062
rect 11610 10024 11612 10033
rect 11664 10024 11666 10033
rect 11610 9959 11666 9968
rect 11716 9722 11744 10474
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11610 9616 11666 9625
rect 11610 9551 11666 9560
rect 11624 6458 11652 9551
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11716 8294 11744 8978
rect 11704 8288 11756 8294
rect 11704 8230 11756 8236
rect 11716 8022 11744 8230
rect 11704 8016 11756 8022
rect 11704 7958 11756 7964
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11716 6322 11744 7686
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11704 5024 11756 5030
rect 11702 4992 11704 5001
rect 11756 4992 11758 5001
rect 11702 4927 11758 4936
rect 11808 4758 11836 13670
rect 11992 13530 12020 13738
rect 11980 13524 12032 13530
rect 11980 13466 12032 13472
rect 12084 13410 12112 15166
rect 11992 13382 12112 13410
rect 11992 13326 12020 13382
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11900 8378 11928 11086
rect 11992 9518 12020 13262
rect 12544 13138 12572 16520
rect 12817 14716 13113 14736
rect 12873 14714 12897 14716
rect 12953 14714 12977 14716
rect 13033 14714 13057 14716
rect 12895 14662 12897 14714
rect 12959 14662 12971 14714
rect 13033 14662 13035 14714
rect 12873 14660 12897 14662
rect 12953 14660 12977 14662
rect 13033 14660 13057 14662
rect 12817 14640 13113 14660
rect 12817 13628 13113 13648
rect 12873 13626 12897 13628
rect 12953 13626 12977 13628
rect 13033 13626 13057 13628
rect 12895 13574 12897 13626
rect 12959 13574 12971 13626
rect 13033 13574 13035 13626
rect 12873 13572 12897 13574
rect 12953 13572 12977 13574
rect 13033 13572 13057 13574
rect 12817 13552 13113 13572
rect 12360 13110 12572 13138
rect 12624 13184 12676 13190
rect 13188 13161 13216 16520
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13544 14000 13596 14006
rect 13544 13942 13596 13948
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 12624 13126 12676 13132
rect 13174 13152 13230 13161
rect 12360 12220 12388 13110
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12360 12192 12480 12220
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12164 11552 12216 11558
rect 12164 11494 12216 11500
rect 12072 11280 12124 11286
rect 12072 11222 12124 11228
rect 12084 10742 12112 11222
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 12072 10464 12124 10470
rect 12072 10406 12124 10412
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 11978 9208 12034 9217
rect 11978 9143 12034 9152
rect 11992 8945 12020 9143
rect 11978 8936 12034 8945
rect 11978 8871 12034 8880
rect 12084 8566 12112 10406
rect 12176 9625 12204 11494
rect 12162 9616 12218 9625
rect 12162 9551 12218 9560
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 12072 8560 12124 8566
rect 12072 8502 12124 8508
rect 11900 8350 12020 8378
rect 11886 7304 11942 7313
rect 11886 7239 11942 7248
rect 11796 4752 11848 4758
rect 11796 4694 11848 4700
rect 11900 4078 11928 7239
rect 11992 5846 12020 8350
rect 12176 8022 12204 9386
rect 12164 8016 12216 8022
rect 12164 7958 12216 7964
rect 12072 7812 12124 7818
rect 12072 7754 12124 7760
rect 12084 7206 12112 7754
rect 12164 7472 12216 7478
rect 12164 7414 12216 7420
rect 12176 7342 12204 7414
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 12084 6866 12112 7142
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 12084 6186 12112 6802
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12176 6390 12204 6598
rect 12164 6384 12216 6390
rect 12164 6326 12216 6332
rect 12072 6180 12124 6186
rect 12072 6122 12124 6128
rect 12072 5908 12124 5914
rect 12072 5850 12124 5856
rect 11980 5840 12032 5846
rect 11980 5782 12032 5788
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11992 5302 12020 5646
rect 12084 5642 12112 5850
rect 12072 5636 12124 5642
rect 12072 5578 12124 5584
rect 11980 5296 12032 5302
rect 11980 5238 12032 5244
rect 11980 4752 12032 4758
rect 11980 4694 12032 4700
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 11992 3738 12020 4694
rect 12268 3738 12296 12038
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12360 10849 12388 11698
rect 12346 10840 12402 10849
rect 12346 10775 12402 10784
rect 12348 10736 12400 10742
rect 12348 10678 12400 10684
rect 12360 9489 12388 10678
rect 12346 9480 12402 9489
rect 12346 9415 12402 9424
rect 12452 9217 12480 12192
rect 12544 11558 12572 12242
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12636 11234 12664 13126
rect 13174 13087 13230 13096
rect 13372 12850 13400 13874
rect 13556 13530 13584 13942
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13268 12776 13320 12782
rect 13268 12718 13320 12724
rect 12817 12540 13113 12560
rect 12873 12538 12897 12540
rect 12953 12538 12977 12540
rect 13033 12538 13057 12540
rect 12895 12486 12897 12538
rect 12959 12486 12971 12538
rect 13033 12486 13035 12538
rect 12873 12484 12897 12486
rect 12953 12484 12977 12486
rect 13033 12484 13057 12486
rect 12817 12464 13113 12484
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12544 11206 12664 11234
rect 12438 9208 12494 9217
rect 12438 9143 12494 9152
rect 12438 9072 12494 9081
rect 12348 9036 12400 9042
rect 12438 9007 12494 9016
rect 12348 8978 12400 8984
rect 12360 8634 12388 8978
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 12452 8378 12480 9007
rect 12360 8350 12480 8378
rect 12360 7970 12388 8350
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12452 8090 12480 8230
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12360 7942 12480 7970
rect 12452 7886 12480 7942
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12360 7177 12388 7822
rect 12440 7200 12492 7206
rect 12346 7168 12402 7177
rect 12440 7142 12492 7148
rect 12346 7103 12402 7112
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 11520 2576 11572 2582
rect 11520 2518 11572 2524
rect 11336 2508 11388 2514
rect 11256 2468 11336 2496
rect 11336 2450 11388 2456
rect 11624 480 11652 3470
rect 11796 3460 11848 3466
rect 11796 3402 11848 3408
rect 11808 2553 11836 3402
rect 11794 2544 11850 2553
rect 11794 2479 11796 2488
rect 11848 2479 11850 2488
rect 11796 2450 11848 2456
rect 12176 480 12204 3470
rect 12360 3058 12388 6938
rect 12452 6254 12480 7142
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12440 5296 12492 5302
rect 12440 5238 12492 5244
rect 12452 4826 12480 5238
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12544 3058 12572 11206
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12636 10606 12664 10950
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12636 10266 12664 10406
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12728 10146 12756 12038
rect 13280 11898 13308 12718
rect 13360 12640 13412 12646
rect 13360 12582 13412 12588
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13372 11642 13400 12582
rect 13556 12050 13584 13262
rect 13648 12918 13676 13670
rect 13740 13326 13768 14350
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13832 13190 13860 16520
rect 14372 13864 14424 13870
rect 14476 13818 14504 16520
rect 14924 14544 14976 14550
rect 14924 14486 14976 14492
rect 14424 13812 14504 13818
rect 14372 13806 14504 13812
rect 14384 13790 14504 13806
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13636 12912 13688 12918
rect 13636 12854 13688 12860
rect 13728 12912 13780 12918
rect 13728 12854 13780 12860
rect 13280 11614 13400 11642
rect 13464 12022 13584 12050
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 12817 11452 13113 11472
rect 12873 11450 12897 11452
rect 12953 11450 12977 11452
rect 13033 11450 13057 11452
rect 12895 11398 12897 11450
rect 12959 11398 12971 11450
rect 13033 11398 13035 11450
rect 12873 11396 12897 11398
rect 12953 11396 12977 11398
rect 13033 11396 13057 11398
rect 12817 11376 13113 11396
rect 12817 10364 13113 10384
rect 12873 10362 12897 10364
rect 12953 10362 12977 10364
rect 13033 10362 13057 10364
rect 12895 10310 12897 10362
rect 12959 10310 12971 10362
rect 13033 10310 13035 10362
rect 12873 10308 12897 10310
rect 12953 10308 12977 10310
rect 13033 10308 13057 10310
rect 12817 10288 13113 10308
rect 12808 10192 12860 10198
rect 12636 10118 12756 10146
rect 12806 10160 12808 10169
rect 12860 10160 12862 10169
rect 12636 3210 12664 10118
rect 12806 10095 12862 10104
rect 12716 10056 12768 10062
rect 12808 10056 12860 10062
rect 12716 9998 12768 10004
rect 12806 10024 12808 10033
rect 12860 10024 12862 10033
rect 12728 9722 12756 9998
rect 12806 9959 12862 9968
rect 13082 10024 13138 10033
rect 13082 9959 13138 9968
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 13096 9364 13124 9959
rect 13188 9518 13216 11494
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 12728 9336 13124 9364
rect 13176 9376 13228 9382
rect 12728 7834 12756 9336
rect 13176 9318 13228 9324
rect 12817 9276 13113 9296
rect 12873 9274 12897 9276
rect 12953 9274 12977 9276
rect 13033 9274 13057 9276
rect 12895 9222 12897 9274
rect 12959 9222 12971 9274
rect 13033 9222 13035 9274
rect 12873 9220 12897 9222
rect 12953 9220 12977 9222
rect 13033 9220 13057 9222
rect 12817 9200 13113 9220
rect 13188 9178 13216 9318
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13084 9104 13136 9110
rect 13084 9046 13136 9052
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12912 8498 12940 8774
rect 13096 8498 13124 9046
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 13084 8492 13136 8498
rect 13136 8452 13216 8480
rect 13084 8434 13136 8440
rect 12806 8392 12862 8401
rect 12806 8327 12808 8336
rect 12860 8327 12862 8336
rect 12808 8298 12860 8304
rect 12817 8188 13113 8208
rect 12873 8186 12897 8188
rect 12953 8186 12977 8188
rect 13033 8186 13057 8188
rect 12895 8134 12897 8186
rect 12959 8134 12971 8186
rect 13033 8134 13035 8186
rect 12873 8132 12897 8134
rect 12953 8132 12977 8134
rect 13033 8132 13057 8134
rect 12817 8112 13113 8132
rect 12728 7806 12848 7834
rect 13188 7818 13216 8452
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12728 6322 12756 7686
rect 12820 7290 12848 7806
rect 13176 7812 13228 7818
rect 13176 7754 13228 7760
rect 13188 7410 13216 7754
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 12820 7262 13216 7290
rect 12817 7100 13113 7120
rect 12873 7098 12897 7100
rect 12953 7098 12977 7100
rect 13033 7098 13057 7100
rect 12895 7046 12897 7098
rect 12959 7046 12971 7098
rect 13033 7046 13035 7098
rect 12873 7044 12897 7046
rect 12953 7044 12977 7046
rect 13033 7044 13057 7046
rect 12817 7024 13113 7044
rect 13188 6984 13216 7262
rect 13096 6956 13216 6984
rect 13096 6644 13124 6956
rect 13176 6792 13228 6798
rect 13174 6760 13176 6769
rect 13228 6760 13230 6769
rect 13174 6695 13230 6704
rect 13096 6616 13216 6644
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12817 6012 13113 6032
rect 12873 6010 12897 6012
rect 12953 6010 12977 6012
rect 13033 6010 13057 6012
rect 12895 5958 12897 6010
rect 12959 5958 12971 6010
rect 13033 5958 13035 6010
rect 12873 5956 12897 5958
rect 12953 5956 12977 5958
rect 13033 5956 13057 5958
rect 12817 5936 13113 5956
rect 13188 5846 13216 6616
rect 13176 5840 13228 5846
rect 13176 5782 13228 5788
rect 12714 5672 12770 5681
rect 12714 5607 12770 5616
rect 13174 5672 13230 5681
rect 13174 5607 13230 5616
rect 12728 5574 12756 5607
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12728 5166 12756 5510
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 12817 4924 13113 4944
rect 12873 4922 12897 4924
rect 12953 4922 12977 4924
rect 13033 4922 13057 4924
rect 12895 4870 12897 4922
rect 12959 4870 12971 4922
rect 13033 4870 13035 4922
rect 12873 4868 12897 4870
rect 12953 4868 12977 4870
rect 13033 4868 13057 4870
rect 12817 4848 13113 4868
rect 13188 4298 13216 5607
rect 13280 5098 13308 11614
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13372 11286 13400 11494
rect 13360 11280 13412 11286
rect 13360 11222 13412 11228
rect 13464 11098 13492 12022
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13372 11070 13492 11098
rect 13372 10146 13400 11070
rect 13452 10668 13504 10674
rect 13452 10610 13504 10616
rect 13464 10577 13492 10610
rect 13450 10568 13506 10577
rect 13450 10503 13506 10512
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13464 10266 13492 10406
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13372 10118 13492 10146
rect 13360 9512 13412 9518
rect 13360 9454 13412 9460
rect 13372 9081 13400 9454
rect 13358 9072 13414 9081
rect 13358 9007 13414 9016
rect 13360 8968 13412 8974
rect 13358 8936 13360 8945
rect 13412 8936 13414 8945
rect 13358 8871 13414 8880
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13372 7002 13400 8570
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13372 5846 13400 6598
rect 13360 5840 13412 5846
rect 13360 5782 13412 5788
rect 13358 5128 13414 5137
rect 13268 5092 13320 5098
rect 13358 5063 13414 5072
rect 13268 5034 13320 5040
rect 13372 4758 13400 5063
rect 13360 4752 13412 4758
rect 13360 4694 13412 4700
rect 13188 4270 13308 4298
rect 13280 4146 13308 4270
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 12817 3836 13113 3856
rect 12873 3834 12897 3836
rect 12953 3834 12977 3836
rect 13033 3834 13057 3836
rect 12895 3782 12897 3834
rect 12959 3782 12971 3834
rect 13033 3782 13035 3834
rect 12873 3780 12897 3782
rect 12953 3780 12977 3782
rect 13033 3780 13057 3782
rect 12817 3760 13113 3780
rect 12636 3182 12756 3210
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 12636 480 12664 2994
rect 12728 2854 12756 3182
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 12817 2748 13113 2768
rect 12873 2746 12897 2748
rect 12953 2746 12977 2748
rect 13033 2746 13057 2748
rect 12895 2694 12897 2746
rect 12959 2694 12971 2746
rect 13033 2694 13035 2746
rect 12873 2692 12897 2694
rect 12953 2692 12977 2694
rect 13033 2692 13057 2694
rect 12817 2672 13113 2692
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 13096 2106 13124 2246
rect 13084 2100 13136 2106
rect 13084 2042 13136 2048
rect 13188 480 13216 4082
rect 13464 3534 13492 10118
rect 13556 4010 13584 11834
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 13648 11218 13676 11698
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13648 10470 13676 11154
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13648 9994 13676 10406
rect 13636 9988 13688 9994
rect 13636 9930 13688 9936
rect 13648 8974 13676 9930
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13634 7984 13690 7993
rect 13634 7919 13636 7928
rect 13688 7919 13690 7928
rect 13636 7890 13688 7896
rect 13636 7200 13688 7206
rect 13634 7168 13636 7177
rect 13688 7168 13690 7177
rect 13634 7103 13690 7112
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13544 4004 13596 4010
rect 13544 3946 13596 3952
rect 13542 3904 13598 3913
rect 13542 3839 13598 3848
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13556 2922 13584 3839
rect 13544 2916 13596 2922
rect 13544 2858 13596 2864
rect 13648 480 13676 5170
rect 13740 4146 13768 12854
rect 13912 12164 13964 12170
rect 13912 12106 13964 12112
rect 14004 12164 14056 12170
rect 14004 12106 14056 12112
rect 13924 11898 13952 12106
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 13912 11620 13964 11626
rect 13912 11562 13964 11568
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13832 10577 13860 10950
rect 13818 10568 13874 10577
rect 13818 10503 13874 10512
rect 13832 9586 13860 10503
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13818 9480 13874 9489
rect 13818 9415 13874 9424
rect 13832 9382 13860 9415
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13924 9110 13952 11562
rect 13912 9104 13964 9110
rect 13912 9046 13964 9052
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13832 6866 13860 8026
rect 13924 7750 13952 8910
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13818 6760 13874 6769
rect 13818 6695 13874 6704
rect 13832 4622 13860 6695
rect 13924 4826 13952 7686
rect 14016 6769 14044 12106
rect 14096 11620 14148 11626
rect 14096 11562 14148 11568
rect 14108 8566 14136 11562
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14200 10266 14228 10746
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 14200 9586 14228 10202
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 14200 9178 14228 9522
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14200 8974 14228 9114
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 14096 8560 14148 8566
rect 14096 8502 14148 8508
rect 14200 8498 14228 8910
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14096 8356 14148 8362
rect 14096 8298 14148 8304
rect 14108 7954 14136 8298
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 14096 7540 14148 7546
rect 14200 7528 14228 8434
rect 14148 7500 14228 7528
rect 14096 7482 14148 7488
rect 14096 6792 14148 6798
rect 14002 6760 14058 6769
rect 14096 6734 14148 6740
rect 14002 6695 14058 6704
rect 14004 6656 14056 6662
rect 14004 6598 14056 6604
rect 14016 5914 14044 6598
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 14108 5574 14136 6734
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 14200 5778 14228 6190
rect 14188 5772 14240 5778
rect 14188 5714 14240 5720
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 14004 5296 14056 5302
rect 14004 5238 14056 5244
rect 13912 4820 13964 4826
rect 13912 4762 13964 4768
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 3238 232 3294 241
rect 3238 167 3294 176
rect 3606 0 3662 480
rect 4158 0 4214 480
rect 4618 0 4674 480
rect 5170 0 5226 480
rect 5630 0 5686 480
rect 6182 0 6238 480
rect 6642 0 6698 480
rect 7102 0 7158 480
rect 7654 0 7710 480
rect 8114 0 8170 480
rect 8666 0 8722 480
rect 9126 0 9182 480
rect 9678 0 9734 480
rect 10138 0 10194 480
rect 10598 0 10654 480
rect 11150 0 11206 480
rect 11610 0 11666 480
rect 12162 0 12218 480
rect 12622 0 12678 480
rect 13174 0 13230 480
rect 13634 0 13690 480
rect 14016 241 14044 5238
rect 14096 4752 14148 4758
rect 14096 4694 14148 4700
rect 14108 4554 14136 4694
rect 14096 4548 14148 4554
rect 14096 4490 14148 4496
rect 14096 4004 14148 4010
rect 14096 3946 14148 3952
rect 14108 480 14136 3946
rect 14292 3942 14320 11494
rect 14372 11348 14424 11354
rect 14372 11290 14424 11296
rect 14384 9489 14412 11290
rect 14370 9480 14426 9489
rect 14370 9415 14426 9424
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14384 7002 14412 9318
rect 14372 6996 14424 7002
rect 14372 6938 14424 6944
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14384 6186 14412 6598
rect 14372 6180 14424 6186
rect 14372 6122 14424 6128
rect 14384 5642 14412 6122
rect 14372 5636 14424 5642
rect 14372 5578 14424 5584
rect 14476 5234 14504 13790
rect 14936 13530 14964 14486
rect 15120 13870 15148 16520
rect 15108 13864 15160 13870
rect 15028 13824 15108 13852
rect 14924 13524 14976 13530
rect 14924 13466 14976 13472
rect 14936 13433 14964 13466
rect 14922 13424 14978 13433
rect 14922 13359 14978 13368
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 14464 4820 14516 4826
rect 14464 4762 14516 4768
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 14476 3641 14504 4762
rect 14568 4010 14596 12038
rect 14556 4004 14608 4010
rect 14556 3946 14608 3952
rect 14660 3890 14688 13126
rect 15028 12458 15056 13824
rect 15108 13806 15160 13812
rect 15106 13424 15162 13433
rect 15106 13359 15108 13368
rect 15160 13359 15162 13368
rect 15108 13330 15160 13336
rect 15212 13274 15240 16623
rect 15750 16520 15806 17000
rect 16394 16520 16450 17000
rect 17038 16520 17094 17000
rect 17682 16520 17738 17000
rect 18326 16520 18382 17000
rect 18970 16520 19026 17000
rect 19614 16520 19670 17000
rect 15382 15056 15438 15065
rect 15382 14991 15438 15000
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15120 13246 15240 13274
rect 15120 12617 15148 13246
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15106 12608 15162 12617
rect 15106 12543 15162 12552
rect 14936 12430 15056 12458
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 14752 8129 14780 12242
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 14738 8120 14794 8129
rect 14738 8055 14794 8064
rect 14738 6896 14794 6905
rect 14738 6831 14794 6840
rect 14752 5778 14780 6831
rect 14740 5772 14792 5778
rect 14740 5714 14792 5720
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 14568 3862 14688 3890
rect 14462 3632 14518 3641
rect 14462 3567 14464 3576
rect 14516 3567 14518 3576
rect 14464 3538 14516 3544
rect 14568 2922 14596 3862
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14556 2916 14608 2922
rect 14556 2858 14608 2864
rect 14660 480 14688 3674
rect 14752 1873 14780 4966
rect 14844 2582 14872 11154
rect 14936 4146 14964 12430
rect 15014 11792 15070 11801
rect 15014 11727 15070 11736
rect 15028 10130 15056 11727
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15016 10124 15068 10130
rect 15016 10066 15068 10072
rect 15028 8673 15056 10066
rect 15120 9926 15148 11494
rect 15108 9920 15160 9926
rect 15108 9862 15160 9868
rect 15212 8922 15240 13126
rect 15304 12986 15332 13670
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15396 12753 15424 14991
rect 15566 14648 15622 14657
rect 15566 14583 15622 14592
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15488 13705 15516 14418
rect 15580 14278 15608 14583
rect 15764 14482 15792 16520
rect 15934 16280 15990 16289
rect 15934 16215 15990 16224
rect 15948 15230 15976 16215
rect 15936 15224 15988 15230
rect 15936 15166 15988 15172
rect 15752 14476 15804 14482
rect 15752 14418 15804 14424
rect 15568 14272 15620 14278
rect 15568 14214 15620 14220
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 16302 14240 16358 14249
rect 15566 13832 15622 13841
rect 15672 13802 15700 14214
rect 15782 14172 16078 14192
rect 16302 14175 16358 14184
rect 15838 14170 15862 14172
rect 15918 14170 15942 14172
rect 15998 14170 16022 14172
rect 15860 14118 15862 14170
rect 15924 14118 15936 14170
rect 15998 14118 16000 14170
rect 15838 14116 15862 14118
rect 15918 14116 15942 14118
rect 15998 14116 16022 14118
rect 15782 14096 16078 14116
rect 15566 13767 15622 13776
rect 15660 13796 15712 13802
rect 15474 13696 15530 13705
rect 15474 13631 15530 13640
rect 15476 12776 15528 12782
rect 15382 12744 15438 12753
rect 15476 12718 15528 12724
rect 15382 12679 15438 12688
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 15290 12472 15346 12481
rect 15290 12407 15346 12416
rect 15304 12238 15332 12407
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15292 10192 15344 10198
rect 15290 10160 15292 10169
rect 15344 10160 15346 10169
rect 15290 10095 15346 10104
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 15304 9722 15332 9930
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15304 8945 15332 9318
rect 15120 8894 15240 8922
rect 15290 8936 15346 8945
rect 15014 8664 15070 8673
rect 15014 8599 15070 8608
rect 15120 8548 15148 8894
rect 15290 8871 15346 8880
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 15028 8520 15148 8548
rect 15028 8106 15056 8520
rect 15212 8362 15240 8774
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 15200 8356 15252 8362
rect 15200 8298 15252 8304
rect 15028 8078 15240 8106
rect 15014 7984 15070 7993
rect 15014 7919 15070 7928
rect 15028 4758 15056 7919
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 15120 7546 15148 7822
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15120 6730 15148 7482
rect 15108 6724 15160 6730
rect 15108 6666 15160 6672
rect 15016 4752 15068 4758
rect 15016 4694 15068 4700
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 14922 4040 14978 4049
rect 14922 3975 14978 3984
rect 14936 3058 14964 3975
rect 15212 3670 15240 8078
rect 15304 7857 15332 8570
rect 15290 7848 15346 7857
rect 15290 7783 15346 7792
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15304 7546 15332 7686
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15290 6352 15346 6361
rect 15290 6287 15346 6296
rect 15304 5273 15332 6287
rect 15290 5264 15346 5273
rect 15290 5199 15346 5208
rect 15396 4758 15424 12582
rect 15488 10577 15516 12718
rect 15580 12209 15608 13767
rect 15660 13738 15712 13744
rect 15658 13696 15714 13705
rect 15658 13631 15714 13640
rect 15566 12200 15622 12209
rect 15566 12135 15622 12144
rect 15672 12084 15700 13631
rect 15782 13084 16078 13104
rect 15838 13082 15862 13084
rect 15918 13082 15942 13084
rect 15998 13082 16022 13084
rect 15860 13030 15862 13082
rect 15924 13030 15936 13082
rect 15998 13030 16000 13082
rect 15838 13028 15862 13030
rect 15918 13028 15942 13030
rect 15998 13028 16022 13030
rect 15782 13008 16078 13028
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 16224 12617 16252 12718
rect 16210 12608 16266 12617
rect 16210 12543 16266 12552
rect 15580 12056 15700 12084
rect 16120 12096 16172 12102
rect 15474 10568 15530 10577
rect 15474 10503 15530 10512
rect 15476 10464 15528 10470
rect 15476 10406 15528 10412
rect 15488 6905 15516 10406
rect 15580 10033 15608 12056
rect 16120 12038 16172 12044
rect 15782 11996 16078 12016
rect 15838 11994 15862 11996
rect 15918 11994 15942 11996
rect 15998 11994 16022 11996
rect 15860 11942 15862 11994
rect 15924 11942 15936 11994
rect 15998 11942 16000 11994
rect 15838 11940 15862 11942
rect 15918 11940 15942 11942
rect 15998 11940 16022 11942
rect 15782 11920 16078 11940
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15672 10538 15700 11698
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15764 11354 15792 11494
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 15782 10908 16078 10928
rect 15838 10906 15862 10908
rect 15918 10906 15942 10908
rect 15998 10906 16022 10908
rect 15860 10854 15862 10906
rect 15924 10854 15936 10906
rect 15998 10854 16000 10906
rect 15838 10852 15862 10854
rect 15918 10852 15942 10854
rect 15998 10852 16022 10854
rect 15782 10832 16078 10852
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15844 10532 15896 10538
rect 15844 10474 15896 10480
rect 15566 10024 15622 10033
rect 15566 9959 15622 9968
rect 15672 9908 15700 10474
rect 15856 10198 15884 10474
rect 15844 10192 15896 10198
rect 15844 10134 15896 10140
rect 15663 9880 15700 9908
rect 15566 9752 15622 9761
rect 15663 9738 15691 9880
rect 15782 9820 16078 9840
rect 15838 9818 15862 9820
rect 15918 9818 15942 9820
rect 15998 9818 16022 9820
rect 15860 9766 15862 9818
rect 15924 9766 15936 9818
rect 15998 9766 16000 9818
rect 15838 9764 15862 9766
rect 15918 9764 15942 9766
rect 15998 9764 16022 9766
rect 15782 9744 16078 9764
rect 15663 9710 15700 9738
rect 15566 9687 15622 9696
rect 15474 6896 15530 6905
rect 15474 6831 15530 6840
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15488 5370 15516 6734
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 15384 4752 15436 4758
rect 15384 4694 15436 4700
rect 15580 4622 15608 9687
rect 15672 9654 15700 9710
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 15658 9072 15714 9081
rect 15658 9007 15714 9016
rect 15672 7002 15700 9007
rect 15782 8732 16078 8752
rect 15838 8730 15862 8732
rect 15918 8730 15942 8732
rect 15998 8730 16022 8732
rect 15860 8678 15862 8730
rect 15924 8678 15936 8730
rect 15998 8678 16000 8730
rect 15838 8676 15862 8678
rect 15918 8676 15942 8678
rect 15998 8676 16022 8678
rect 15782 8656 16078 8676
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 15752 8356 15804 8362
rect 15752 8298 15804 8304
rect 15764 8265 15792 8298
rect 15750 8256 15806 8265
rect 15750 8191 15806 8200
rect 15856 7886 15884 8366
rect 16026 8120 16082 8129
rect 16026 8055 16028 8064
rect 16080 8055 16082 8064
rect 16028 8026 16080 8032
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 15782 7644 16078 7664
rect 15838 7642 15862 7644
rect 15918 7642 15942 7644
rect 15998 7642 16022 7644
rect 15860 7590 15862 7642
rect 15924 7590 15936 7642
rect 15998 7590 16000 7642
rect 15838 7588 15862 7590
rect 15918 7588 15942 7590
rect 15998 7588 16022 7590
rect 15782 7568 16078 7588
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 15672 6458 15700 6802
rect 15782 6556 16078 6576
rect 15838 6554 15862 6556
rect 15918 6554 15942 6556
rect 15998 6554 16022 6556
rect 15860 6502 15862 6554
rect 15924 6502 15936 6554
rect 15998 6502 16000 6554
rect 15838 6500 15862 6502
rect 15918 6500 15942 6502
rect 15998 6500 16022 6502
rect 15782 6480 16078 6500
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15752 6384 15804 6390
rect 15752 6326 15804 6332
rect 15660 6112 15712 6118
rect 15660 6054 15712 6060
rect 15672 5778 15700 6054
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15764 5710 15792 6326
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 15672 4865 15700 5510
rect 15782 5468 16078 5488
rect 15838 5466 15862 5468
rect 15918 5466 15942 5468
rect 15998 5466 16022 5468
rect 15860 5414 15862 5466
rect 15924 5414 15936 5466
rect 15998 5414 16000 5466
rect 15838 5412 15862 5414
rect 15918 5412 15942 5414
rect 15998 5412 16022 5414
rect 15782 5392 16078 5412
rect 16026 5128 16082 5137
rect 16026 5063 16082 5072
rect 16040 5030 16068 5063
rect 16028 5024 16080 5030
rect 16028 4966 16080 4972
rect 15658 4856 15714 4865
rect 15658 4791 15714 4800
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 15568 4616 15620 4622
rect 15568 4558 15620 4564
rect 15396 3738 15424 4558
rect 15782 4380 16078 4400
rect 15838 4378 15862 4380
rect 15918 4378 15942 4380
rect 15998 4378 16022 4380
rect 15860 4326 15862 4378
rect 15924 4326 15936 4378
rect 15998 4326 16000 4378
rect 15838 4324 15862 4326
rect 15918 4324 15942 4326
rect 15998 4324 16022 4326
rect 15782 4304 16078 4324
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15200 3664 15252 3670
rect 15200 3606 15252 3612
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 14832 2576 14884 2582
rect 14832 2518 14884 2524
rect 15016 2100 15068 2106
rect 15016 2042 15068 2048
rect 14738 1864 14794 1873
rect 14738 1799 14794 1808
rect 15028 1057 15056 2042
rect 15014 1048 15070 1057
rect 15014 983 15070 992
rect 15120 480 15148 3470
rect 15568 3392 15620 3398
rect 15568 3334 15620 3340
rect 15580 2553 15608 3334
rect 15566 2544 15622 2553
rect 15566 2479 15622 2488
rect 15672 480 15700 3878
rect 15782 3292 16078 3312
rect 15838 3290 15862 3292
rect 15918 3290 15942 3292
rect 15998 3290 16022 3292
rect 15860 3238 15862 3290
rect 15924 3238 15936 3290
rect 15998 3238 16000 3290
rect 15838 3236 15862 3238
rect 15918 3236 15942 3238
rect 15998 3236 16022 3238
rect 15782 3216 16078 3236
rect 15750 2952 15806 2961
rect 15750 2887 15752 2896
rect 15804 2887 15806 2896
rect 15752 2858 15804 2864
rect 16026 2680 16082 2689
rect 16026 2615 16082 2624
rect 16040 2514 16068 2615
rect 16028 2508 16080 2514
rect 16028 2450 16080 2456
rect 15782 2204 16078 2224
rect 15838 2202 15862 2204
rect 15918 2202 15942 2204
rect 15998 2202 16022 2204
rect 15860 2150 15862 2202
rect 15924 2150 15936 2202
rect 15998 2150 16000 2202
rect 15838 2148 15862 2150
rect 15918 2148 15942 2150
rect 15998 2148 16022 2150
rect 15782 2128 16078 2148
rect 16132 480 16160 12038
rect 16316 11830 16344 14175
rect 16408 13870 16436 16520
rect 17052 14550 17080 16520
rect 17040 14544 17092 14550
rect 17040 14486 17092 14492
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 16304 11824 16356 11830
rect 16304 11766 16356 11772
rect 16408 11370 16436 13806
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16316 11342 16436 11370
rect 16212 9376 16264 9382
rect 16212 9318 16264 9324
rect 16224 9110 16252 9318
rect 16212 9104 16264 9110
rect 16212 9046 16264 9052
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 16224 7342 16252 7890
rect 16212 7336 16264 7342
rect 16212 7278 16264 7284
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16224 6322 16252 7142
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 16224 5710 16252 6258
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16212 5568 16264 5574
rect 16212 5510 16264 5516
rect 16224 5166 16252 5510
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 16224 4049 16252 4422
rect 16210 4040 16266 4049
rect 16210 3975 16212 3984
rect 16264 3975 16266 3984
rect 16212 3946 16264 3952
rect 16316 3670 16344 11342
rect 16396 11212 16448 11218
rect 16396 11154 16448 11160
rect 16408 8634 16436 11154
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16396 7744 16448 7750
rect 16396 7686 16448 7692
rect 16408 6186 16436 7686
rect 16396 6180 16448 6186
rect 16396 6122 16448 6128
rect 16396 5704 16448 5710
rect 16396 5646 16448 5652
rect 16408 5234 16436 5646
rect 16396 5228 16448 5234
rect 16396 5170 16448 5176
rect 16394 4992 16450 5001
rect 16394 4927 16450 4936
rect 16408 4690 16436 4927
rect 16396 4684 16448 4690
rect 16396 4626 16448 4632
rect 16304 3664 16356 3670
rect 16304 3606 16356 3612
rect 16210 3088 16266 3097
rect 16500 3058 16528 11630
rect 16592 10305 16620 12718
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16776 11694 16804 11834
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16764 11688 16816 11694
rect 16868 11665 16896 11698
rect 16764 11630 16816 11636
rect 16854 11656 16910 11665
rect 16854 11591 16910 11600
rect 16948 11620 17000 11626
rect 16764 11348 16816 11354
rect 16764 11290 16816 11296
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16578 10296 16634 10305
rect 16578 10231 16634 10240
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16592 9178 16620 10066
rect 16684 9926 16712 11086
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 16684 9450 16712 9862
rect 16776 9466 16804 11290
rect 16868 9586 16896 11591
rect 16948 11562 17000 11568
rect 16960 11354 16988 11562
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 17040 11280 17092 11286
rect 17040 11222 17092 11228
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16960 10606 16988 10950
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16856 9580 16908 9586
rect 16856 9522 16908 9528
rect 16672 9444 16724 9450
rect 16776 9438 16988 9466
rect 16672 9386 16724 9392
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16776 9178 16804 9318
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 16764 9172 16816 9178
rect 16764 9114 16816 9120
rect 16592 8974 16620 9114
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16592 8498 16620 8910
rect 16684 8566 16712 8978
rect 16762 8800 16818 8809
rect 16762 8735 16818 8744
rect 16672 8560 16724 8566
rect 16672 8502 16724 8508
rect 16580 8492 16632 8498
rect 16580 8434 16632 8440
rect 16776 8412 16804 8735
rect 16868 8537 16896 9318
rect 16854 8528 16910 8537
rect 16854 8463 16910 8472
rect 16776 8384 16896 8412
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16592 7274 16620 7822
rect 16580 7268 16632 7274
rect 16580 7210 16632 7216
rect 16592 6458 16620 7210
rect 16684 6730 16712 8298
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16776 8090 16804 8230
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16868 7970 16896 8384
rect 16776 7942 16896 7970
rect 16672 6724 16724 6730
rect 16672 6666 16724 6672
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16580 5840 16632 5846
rect 16580 5782 16632 5788
rect 16210 3023 16266 3032
rect 16488 3052 16540 3058
rect 16224 2650 16252 3023
rect 16488 2994 16540 3000
rect 16592 2990 16620 5782
rect 16684 5370 16712 6054
rect 16672 5364 16724 5370
rect 16672 5306 16724 5312
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16580 2984 16632 2990
rect 16580 2926 16632 2932
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 16212 2304 16264 2310
rect 16210 2272 16212 2281
rect 16264 2272 16266 2281
rect 16210 2207 16266 2216
rect 16684 480 16712 4558
rect 16776 2514 16804 7942
rect 16856 7812 16908 7818
rect 16856 7754 16908 7760
rect 16868 6934 16896 7754
rect 16856 6928 16908 6934
rect 16856 6870 16908 6876
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16868 4826 16896 5714
rect 16856 4820 16908 4826
rect 16856 4762 16908 4768
rect 16960 3890 16988 9438
rect 17052 8906 17080 11222
rect 17040 8900 17092 8906
rect 17040 8842 17092 8848
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 17052 5166 17080 8570
rect 17040 5160 17092 5166
rect 17040 5102 17092 5108
rect 17144 4146 17172 12242
rect 17236 10146 17264 12582
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 17328 10266 17356 11154
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 17420 10810 17448 11086
rect 17408 10804 17460 10810
rect 17408 10746 17460 10752
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17236 10118 17356 10146
rect 17420 10130 17448 10610
rect 17224 9580 17276 9586
rect 17224 9522 17276 9528
rect 17236 8566 17264 9522
rect 17224 8560 17276 8566
rect 17224 8502 17276 8508
rect 17236 7886 17264 8502
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17236 6798 17264 7822
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17224 6452 17276 6458
rect 17224 6394 17276 6400
rect 17236 5710 17264 6394
rect 17224 5704 17276 5710
rect 17224 5646 17276 5652
rect 17236 5234 17264 5646
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 17328 4622 17356 10118
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 17406 9888 17462 9897
rect 17406 9823 17462 9832
rect 17420 7818 17448 9823
rect 17408 7812 17460 7818
rect 17408 7754 17460 7760
rect 17512 7041 17540 11494
rect 17604 10266 17632 13262
rect 17696 13258 17724 16520
rect 18340 13462 18368 16520
rect 18418 15872 18474 15881
rect 18418 15807 18474 15816
rect 18328 13456 18380 13462
rect 18328 13398 18380 13404
rect 17776 13388 17828 13394
rect 17776 13330 17828 13336
rect 17684 13252 17736 13258
rect 17684 13194 17736 13200
rect 17788 12186 17816 13330
rect 18326 13288 18382 13297
rect 18326 13223 18382 13232
rect 18144 12640 18196 12646
rect 18144 12582 18196 12588
rect 17868 12300 17920 12306
rect 17868 12242 17920 12248
rect 17696 12158 17816 12186
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17604 9625 17632 9998
rect 17590 9616 17646 9625
rect 17590 9551 17646 9560
rect 17498 7032 17554 7041
rect 17498 6967 17554 6976
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 17592 6112 17644 6118
rect 17592 6054 17644 6060
rect 17420 5681 17448 6054
rect 17406 5672 17462 5681
rect 17406 5607 17462 5616
rect 17500 5636 17552 5642
rect 17500 5578 17552 5584
rect 17408 5568 17460 5574
rect 17408 5510 17460 5516
rect 17420 5098 17448 5510
rect 17408 5092 17460 5098
rect 17408 5034 17460 5040
rect 17512 4622 17540 5578
rect 17316 4616 17368 4622
rect 17316 4558 17368 4564
rect 17500 4616 17552 4622
rect 17500 4558 17552 4564
rect 17406 4448 17462 4457
rect 17406 4383 17462 4392
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 16960 3862 17172 3890
rect 16946 3632 17002 3641
rect 16946 3567 17002 3576
rect 16960 2650 16988 3567
rect 16948 2644 17000 2650
rect 16948 2586 17000 2592
rect 16764 2508 16816 2514
rect 16764 2450 16816 2456
rect 17144 480 17172 3862
rect 17420 3194 17448 4383
rect 17512 3534 17540 4558
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17498 2680 17554 2689
rect 17498 2615 17554 2624
rect 17512 2514 17540 2615
rect 17500 2508 17552 2514
rect 17500 2450 17552 2456
rect 17604 480 17632 6054
rect 17696 4554 17724 12158
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17788 6118 17816 12038
rect 17880 11014 17908 12242
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 17868 11008 17920 11014
rect 17868 10950 17920 10956
rect 17972 10826 18000 11630
rect 17880 10798 18000 10826
rect 17880 9602 17908 10798
rect 17880 9574 18000 9602
rect 17866 9480 17922 9489
rect 17866 9415 17922 9424
rect 17880 8838 17908 9415
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 17776 5772 17828 5778
rect 17776 5714 17828 5720
rect 17684 4548 17736 4554
rect 17684 4490 17736 4496
rect 17682 4040 17738 4049
rect 17682 3975 17738 3984
rect 17696 2650 17724 3975
rect 17788 3738 17816 5714
rect 17776 3732 17828 3738
rect 17776 3674 17828 3680
rect 17880 3670 17908 8774
rect 17972 8634 18000 9574
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 18064 7449 18092 12038
rect 18050 7440 18106 7449
rect 18050 7375 18106 7384
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 18064 6089 18092 6598
rect 18050 6080 18106 6089
rect 18050 6015 18106 6024
rect 17868 3664 17920 3670
rect 17868 3606 17920 3612
rect 17684 2644 17736 2650
rect 17684 2586 17736 2592
rect 18156 480 18184 12582
rect 18234 11248 18290 11257
rect 18234 11183 18290 11192
rect 18248 4826 18276 11183
rect 18340 10606 18368 13223
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 18432 10266 18460 15807
rect 18984 13530 19012 16520
rect 18972 13524 19024 13530
rect 18972 13466 19024 13472
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18512 9104 18564 9110
rect 18512 9046 18564 9052
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 18340 6390 18368 8978
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18328 6384 18380 6390
rect 18328 6326 18380 6332
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 18432 649 18460 7482
rect 18524 6497 18552 9046
rect 18510 6488 18566 6497
rect 18510 6423 18566 6432
rect 18418 640 18474 649
rect 18418 575 18474 584
rect 18616 480 18644 13126
rect 19628 12918 19656 16520
rect 19616 12912 19668 12918
rect 19616 12854 19668 12860
rect 19156 12164 19208 12170
rect 19156 12106 19208 12112
rect 18880 7744 18932 7750
rect 18880 7686 18932 7692
rect 18892 1465 18920 7686
rect 18878 1456 18934 1465
rect 18878 1391 18934 1400
rect 19168 480 19196 12106
rect 19616 11824 19668 11830
rect 19616 11766 19668 11772
rect 19628 480 19656 11766
rect 14002 232 14058 241
rect 14002 167 14058 176
rect 14094 0 14150 480
rect 14646 0 14702 480
rect 15106 0 15162 480
rect 15658 0 15714 480
rect 16118 0 16174 480
rect 16670 0 16726 480
rect 17130 0 17186 480
rect 17590 0 17646 480
rect 18142 0 18198 480
rect 18602 0 18658 480
rect 19154 0 19210 480
rect 19614 0 19670 480
<< via2 >>
rect 3606 16632 3662 16688
rect 2410 16224 2466 16280
rect 1766 7928 1822 7984
rect 1766 7248 1822 7304
rect 1858 6332 1860 6352
rect 1860 6332 1912 6352
rect 1912 6332 1914 6352
rect 1858 6296 1914 6332
rect 1858 5888 1914 5944
rect 1766 5480 1822 5536
rect 1858 4664 1914 4720
rect 2226 13776 2282 13832
rect 3146 15816 3202 15872
rect 3054 12552 3110 12608
rect 2134 7520 2190 7576
rect 2686 10376 2742 10432
rect 2594 10004 2596 10024
rect 2596 10004 2648 10024
rect 2648 10004 2650 10024
rect 2594 9968 2650 10004
rect 2594 9696 2650 9752
rect 2870 10376 2926 10432
rect 15198 16632 15254 16688
rect 3790 15000 3846 15056
rect 3698 14592 3754 14648
rect 3514 14184 3570 14240
rect 3514 13368 3570 13424
rect 3146 11328 3202 11384
rect 3146 8336 3202 8392
rect 2870 8200 2926 8256
rect 2778 7112 2834 7168
rect 2502 6976 2558 7032
rect 2502 5208 2558 5264
rect 3330 12960 3386 13016
rect 3330 12280 3386 12336
rect 3921 14170 3977 14172
rect 4001 14170 4057 14172
rect 4081 14170 4137 14172
rect 4161 14170 4217 14172
rect 3921 14118 3947 14170
rect 3947 14118 3977 14170
rect 4001 14118 4011 14170
rect 4011 14118 4057 14170
rect 4081 14118 4127 14170
rect 4127 14118 4137 14170
rect 4161 14118 4191 14170
rect 4191 14118 4217 14170
rect 3921 14116 3977 14118
rect 4001 14116 4057 14118
rect 4081 14116 4137 14118
rect 4161 14116 4217 14118
rect 3921 13082 3977 13084
rect 4001 13082 4057 13084
rect 4081 13082 4137 13084
rect 4161 13082 4217 13084
rect 3921 13030 3947 13082
rect 3947 13030 3977 13082
rect 4001 13030 4011 13082
rect 4011 13030 4057 13082
rect 4081 13030 4127 13082
rect 4127 13030 4137 13082
rect 4161 13030 4191 13082
rect 4191 13030 4217 13082
rect 3921 13028 3977 13030
rect 4001 13028 4057 13030
rect 4081 13028 4137 13030
rect 4161 13028 4217 13030
rect 3330 11736 3386 11792
rect 4066 12180 4068 12200
rect 4068 12180 4120 12200
rect 4120 12180 4122 12200
rect 3514 9832 3570 9888
rect 3422 8336 3478 8392
rect 3054 6876 3056 6896
rect 3056 6876 3108 6896
rect 3108 6876 3110 6896
rect 3054 6840 3110 6876
rect 1858 2216 1914 2272
rect 2778 5072 2834 5128
rect 2778 4256 2834 4312
rect 3330 3884 3332 3904
rect 3332 3884 3384 3904
rect 3384 3884 3386 3904
rect 3330 3848 3386 3884
rect 3054 3440 3110 3496
rect 2962 3032 3018 3088
rect 4066 12144 4122 12180
rect 4250 12144 4306 12200
rect 3921 11994 3977 11996
rect 4001 11994 4057 11996
rect 4081 11994 4137 11996
rect 4161 11994 4217 11996
rect 3921 11942 3947 11994
rect 3947 11942 3977 11994
rect 4001 11942 4011 11994
rect 4011 11942 4057 11994
rect 4081 11942 4127 11994
rect 4127 11942 4137 11994
rect 4161 11942 4191 11994
rect 4191 11942 4217 11994
rect 3921 11940 3977 11942
rect 4001 11940 4057 11942
rect 4081 11940 4137 11942
rect 4161 11940 4217 11942
rect 4526 12300 4582 12336
rect 4526 12280 4528 12300
rect 4528 12280 4580 12300
rect 4580 12280 4582 12300
rect 3921 10906 3977 10908
rect 4001 10906 4057 10908
rect 4081 10906 4137 10908
rect 4161 10906 4217 10908
rect 3921 10854 3947 10906
rect 3947 10854 3977 10906
rect 4001 10854 4011 10906
rect 4011 10854 4057 10906
rect 4081 10854 4127 10906
rect 4127 10854 4137 10906
rect 4161 10854 4191 10906
rect 4191 10854 4217 10906
rect 3921 10852 3977 10854
rect 4001 10852 4057 10854
rect 4081 10852 4137 10854
rect 4161 10852 4217 10854
rect 3606 9016 3662 9072
rect 3606 8492 3662 8528
rect 3606 8472 3608 8492
rect 3608 8472 3660 8492
rect 3660 8472 3662 8492
rect 3606 6704 3662 6760
rect 3606 6296 3662 6352
rect 3422 2644 3478 2680
rect 3422 2624 3424 2644
rect 3424 2624 3476 2644
rect 3476 2624 3478 2644
rect 3330 1808 3386 1864
rect 3514 1400 3570 1456
rect 3921 9818 3977 9820
rect 4001 9818 4057 9820
rect 4081 9818 4137 9820
rect 4161 9818 4217 9820
rect 3921 9766 3947 9818
rect 3947 9766 3977 9818
rect 4001 9766 4011 9818
rect 4011 9766 4057 9818
rect 4081 9766 4127 9818
rect 4127 9766 4137 9818
rect 4161 9766 4191 9818
rect 4191 9766 4217 9818
rect 3921 9764 3977 9766
rect 4001 9764 4057 9766
rect 4081 9764 4137 9766
rect 4161 9764 4217 9766
rect 3974 9288 4030 9344
rect 4158 9288 4214 9344
rect 4158 8880 4214 8936
rect 3921 8730 3977 8732
rect 4001 8730 4057 8732
rect 4081 8730 4137 8732
rect 4161 8730 4217 8732
rect 3921 8678 3947 8730
rect 3947 8678 3977 8730
rect 4001 8678 4011 8730
rect 4011 8678 4057 8730
rect 4081 8678 4127 8730
rect 4127 8678 4137 8730
rect 4161 8678 4191 8730
rect 4191 8678 4217 8730
rect 3921 8676 3977 8678
rect 4001 8676 4057 8678
rect 4081 8676 4137 8678
rect 4161 8676 4217 8678
rect 3921 7642 3977 7644
rect 4001 7642 4057 7644
rect 4081 7642 4137 7644
rect 4161 7642 4217 7644
rect 3921 7590 3947 7642
rect 3947 7590 3977 7642
rect 4001 7590 4011 7642
rect 4011 7590 4057 7642
rect 4081 7590 4127 7642
rect 4127 7590 4137 7642
rect 4161 7590 4191 7642
rect 4191 7590 4217 7642
rect 3921 7588 3977 7590
rect 4001 7588 4057 7590
rect 4081 7588 4137 7590
rect 4161 7588 4217 7590
rect 3790 6976 3846 7032
rect 3921 6554 3977 6556
rect 4001 6554 4057 6556
rect 4081 6554 4137 6556
rect 4161 6554 4217 6556
rect 3921 6502 3947 6554
rect 3947 6502 3977 6554
rect 4001 6502 4011 6554
rect 4011 6502 4057 6554
rect 4081 6502 4127 6554
rect 4127 6502 4137 6554
rect 4161 6502 4191 6554
rect 4191 6502 4217 6554
rect 3921 6500 3977 6502
rect 4001 6500 4057 6502
rect 4081 6500 4137 6502
rect 4161 6500 4217 6502
rect 3921 5466 3977 5468
rect 4001 5466 4057 5468
rect 4081 5466 4137 5468
rect 4161 5466 4217 5468
rect 3921 5414 3947 5466
rect 3947 5414 3977 5466
rect 4001 5414 4011 5466
rect 4011 5414 4057 5466
rect 4081 5414 4127 5466
rect 4127 5414 4137 5466
rect 4161 5414 4191 5466
rect 4191 5414 4217 5466
rect 3921 5412 3977 5414
rect 4001 5412 4057 5414
rect 4081 5412 4137 5414
rect 4161 5412 4217 5414
rect 3921 4378 3977 4380
rect 4001 4378 4057 4380
rect 4081 4378 4137 4380
rect 4161 4378 4217 4380
rect 3921 4326 3947 4378
rect 3947 4326 3977 4378
rect 4001 4326 4011 4378
rect 4011 4326 4057 4378
rect 4081 4326 4127 4378
rect 4127 4326 4137 4378
rect 4161 4326 4191 4378
rect 4191 4326 4217 4378
rect 3921 4324 3977 4326
rect 4001 4324 4057 4326
rect 4081 4324 4137 4326
rect 4161 4324 4217 4326
rect 3921 3290 3977 3292
rect 4001 3290 4057 3292
rect 4081 3290 4137 3292
rect 4161 3290 4217 3292
rect 3921 3238 3947 3290
rect 3947 3238 3977 3290
rect 4001 3238 4011 3290
rect 4011 3238 4057 3290
rect 4081 3238 4127 3290
rect 4127 3238 4137 3290
rect 4161 3238 4191 3290
rect 4191 3238 4217 3290
rect 3921 3236 3977 3238
rect 4001 3236 4057 3238
rect 4081 3236 4137 3238
rect 4161 3236 4217 3238
rect 5170 10648 5226 10704
rect 4710 7828 4712 7848
rect 4712 7828 4764 7848
rect 4764 7828 4766 7848
rect 4710 7792 4766 7828
rect 4986 9288 5042 9344
rect 5262 9424 5318 9480
rect 5170 7792 5226 7848
rect 3921 2202 3977 2204
rect 4001 2202 4057 2204
rect 4081 2202 4137 2204
rect 4161 2202 4217 2204
rect 3921 2150 3947 2202
rect 3947 2150 3977 2202
rect 4001 2150 4011 2202
rect 4011 2150 4057 2202
rect 4081 2150 4127 2202
rect 4127 2150 4137 2202
rect 4161 2150 4191 2202
rect 4191 2150 4217 2202
rect 3921 2148 3977 2150
rect 4001 2148 4057 2150
rect 4081 2148 4137 2150
rect 4161 2148 4217 2150
rect 3698 992 3754 1048
rect 3698 584 3754 640
rect 6886 14714 6942 14716
rect 6966 14714 7022 14716
rect 7046 14714 7102 14716
rect 7126 14714 7182 14716
rect 6886 14662 6912 14714
rect 6912 14662 6942 14714
rect 6966 14662 6976 14714
rect 6976 14662 7022 14714
rect 7046 14662 7092 14714
rect 7092 14662 7102 14714
rect 7126 14662 7156 14714
rect 7156 14662 7182 14714
rect 6886 14660 6942 14662
rect 6966 14660 7022 14662
rect 7046 14660 7102 14662
rect 7126 14660 7182 14662
rect 5538 10104 5594 10160
rect 5446 9560 5502 9616
rect 6090 12280 6146 12336
rect 6090 11756 6146 11792
rect 6090 11736 6092 11756
rect 6092 11736 6144 11756
rect 6144 11736 6146 11756
rect 5446 7928 5502 7984
rect 6886 13626 6942 13628
rect 6966 13626 7022 13628
rect 7046 13626 7102 13628
rect 7126 13626 7182 13628
rect 6886 13574 6912 13626
rect 6912 13574 6942 13626
rect 6966 13574 6976 13626
rect 6976 13574 7022 13626
rect 7046 13574 7092 13626
rect 7092 13574 7102 13626
rect 7126 13574 7156 13626
rect 7156 13574 7182 13626
rect 6886 13572 6942 13574
rect 6966 13572 7022 13574
rect 7046 13572 7102 13574
rect 7126 13572 7182 13574
rect 6886 12538 6942 12540
rect 6966 12538 7022 12540
rect 7046 12538 7102 12540
rect 7126 12538 7182 12540
rect 6886 12486 6912 12538
rect 6912 12486 6942 12538
rect 6966 12486 6976 12538
rect 6976 12486 7022 12538
rect 7046 12486 7092 12538
rect 7092 12486 7102 12538
rect 7126 12486 7156 12538
rect 7156 12486 7182 12538
rect 6886 12484 6942 12486
rect 6966 12484 7022 12486
rect 7046 12484 7102 12486
rect 7126 12484 7182 12486
rect 6274 12316 6276 12336
rect 6276 12316 6328 12336
rect 6328 12316 6330 12336
rect 6274 12280 6330 12316
rect 6458 11736 6514 11792
rect 6274 9832 6330 9888
rect 6458 9424 6514 9480
rect 6366 8472 6422 8528
rect 6366 7284 6368 7304
rect 6368 7284 6420 7304
rect 6420 7284 6422 7304
rect 6366 7248 6422 7284
rect 6458 4528 6514 4584
rect 6886 11450 6942 11452
rect 6966 11450 7022 11452
rect 7046 11450 7102 11452
rect 7126 11450 7182 11452
rect 6886 11398 6912 11450
rect 6912 11398 6942 11450
rect 6966 11398 6976 11450
rect 6976 11398 7022 11450
rect 7046 11398 7092 11450
rect 7092 11398 7102 11450
rect 7126 11398 7156 11450
rect 7156 11398 7182 11450
rect 6886 11396 6942 11398
rect 6966 11396 7022 11398
rect 7046 11396 7102 11398
rect 7126 11396 7182 11398
rect 7470 12144 7526 12200
rect 6886 10362 6942 10364
rect 6966 10362 7022 10364
rect 7046 10362 7102 10364
rect 7126 10362 7182 10364
rect 6886 10310 6912 10362
rect 6912 10310 6942 10362
rect 6966 10310 6976 10362
rect 6976 10310 7022 10362
rect 7046 10310 7092 10362
rect 7092 10310 7102 10362
rect 7126 10310 7156 10362
rect 7156 10310 7182 10362
rect 6886 10308 6942 10310
rect 6966 10308 7022 10310
rect 7046 10308 7102 10310
rect 7126 10308 7182 10310
rect 6734 10240 6790 10296
rect 6886 9274 6942 9276
rect 6966 9274 7022 9276
rect 7046 9274 7102 9276
rect 7126 9274 7182 9276
rect 6886 9222 6912 9274
rect 6912 9222 6942 9274
rect 6966 9222 6976 9274
rect 6976 9222 7022 9274
rect 7046 9222 7092 9274
rect 7092 9222 7102 9274
rect 7126 9222 7156 9274
rect 7156 9222 7182 9274
rect 6886 9220 6942 9222
rect 6966 9220 7022 9222
rect 7046 9220 7102 9222
rect 7126 9220 7182 9222
rect 7194 8880 7250 8936
rect 6886 8186 6942 8188
rect 6966 8186 7022 8188
rect 7046 8186 7102 8188
rect 7126 8186 7182 8188
rect 6886 8134 6912 8186
rect 6912 8134 6942 8186
rect 6966 8134 6976 8186
rect 6976 8134 7022 8186
rect 7046 8134 7092 8186
rect 7092 8134 7102 8186
rect 7126 8134 7156 8186
rect 7156 8134 7182 8186
rect 6886 8132 6942 8134
rect 6966 8132 7022 8134
rect 7046 8132 7102 8134
rect 7126 8132 7182 8134
rect 6886 7098 6942 7100
rect 6966 7098 7022 7100
rect 7046 7098 7102 7100
rect 7126 7098 7182 7100
rect 6886 7046 6912 7098
rect 6912 7046 6942 7098
rect 6966 7046 6976 7098
rect 6976 7046 7022 7098
rect 7046 7046 7092 7098
rect 7092 7046 7102 7098
rect 7126 7046 7156 7098
rect 7156 7046 7182 7098
rect 6886 7044 6942 7046
rect 6966 7044 7022 7046
rect 7046 7044 7102 7046
rect 7126 7044 7182 7046
rect 7470 9968 7526 10024
rect 7470 9288 7526 9344
rect 7562 8200 7618 8256
rect 6886 6010 6942 6012
rect 6966 6010 7022 6012
rect 7046 6010 7102 6012
rect 7126 6010 7182 6012
rect 6886 5958 6912 6010
rect 6912 5958 6942 6010
rect 6966 5958 6976 6010
rect 6976 5958 7022 6010
rect 7046 5958 7092 6010
rect 7092 5958 7102 6010
rect 7126 5958 7156 6010
rect 7156 5958 7182 6010
rect 6886 5956 6942 5958
rect 6966 5956 7022 5958
rect 7046 5956 7102 5958
rect 7126 5956 7182 5958
rect 6886 4922 6942 4924
rect 6966 4922 7022 4924
rect 7046 4922 7102 4924
rect 7126 4922 7182 4924
rect 6886 4870 6912 4922
rect 6912 4870 6942 4922
rect 6966 4870 6976 4922
rect 6976 4870 7022 4922
rect 7046 4870 7092 4922
rect 7092 4870 7102 4922
rect 7126 4870 7156 4922
rect 7156 4870 7182 4922
rect 6886 4868 6942 4870
rect 6966 4868 7022 4870
rect 7046 4868 7102 4870
rect 7126 4868 7182 4870
rect 6918 4664 6974 4720
rect 7470 4664 7526 4720
rect 6886 3834 6942 3836
rect 6966 3834 7022 3836
rect 7046 3834 7102 3836
rect 7126 3834 7182 3836
rect 6886 3782 6912 3834
rect 6912 3782 6942 3834
rect 6966 3782 6976 3834
rect 6976 3782 7022 3834
rect 7046 3782 7092 3834
rect 7092 3782 7102 3834
rect 7126 3782 7156 3834
rect 7156 3782 7182 3834
rect 6886 3780 6942 3782
rect 6966 3780 7022 3782
rect 7046 3780 7102 3782
rect 7126 3780 7182 3782
rect 6886 2746 6942 2748
rect 6966 2746 7022 2748
rect 7046 2746 7102 2748
rect 7126 2746 7182 2748
rect 6886 2694 6912 2746
rect 6912 2694 6942 2746
rect 6966 2694 6976 2746
rect 6976 2694 7022 2746
rect 7046 2694 7092 2746
rect 7092 2694 7102 2746
rect 7126 2694 7156 2746
rect 7156 2694 7182 2746
rect 6886 2692 6942 2694
rect 6966 2692 7022 2694
rect 7046 2692 7102 2694
rect 7126 2692 7182 2694
rect 7746 7792 7802 7848
rect 7930 9324 7932 9344
rect 7932 9324 7984 9344
rect 7984 9324 7986 9344
rect 7930 9288 7986 9324
rect 7930 8880 7986 8936
rect 7930 8064 7986 8120
rect 8298 10512 8354 10568
rect 9402 15408 9458 15464
rect 8666 12416 8722 12472
rect 8666 11056 8722 11112
rect 8850 11736 8906 11792
rect 8850 10512 8906 10568
rect 8850 9560 8906 9616
rect 8758 9324 8760 9344
rect 8760 9324 8812 9344
rect 8812 9324 8814 9344
rect 8758 9288 8814 9324
rect 8850 8880 8906 8936
rect 8206 7520 8262 7576
rect 8022 6296 8078 6352
rect 8758 8744 8814 8800
rect 8666 7384 8722 7440
rect 8206 4528 8262 4584
rect 8298 2508 8354 2544
rect 8298 2488 8300 2508
rect 8300 2488 8352 2508
rect 8352 2488 8354 2508
rect 8574 2760 8630 2816
rect 9310 12280 9366 12336
rect 9126 10104 9182 10160
rect 9126 8608 9182 8664
rect 9126 6976 9182 7032
rect 9494 9868 9496 9888
rect 9496 9868 9548 9888
rect 9548 9868 9550 9888
rect 9494 9832 9550 9868
rect 9494 8880 9550 8936
rect 9402 8608 9458 8664
rect 9494 8064 9550 8120
rect 9310 7928 9366 7984
rect 9494 4972 9496 4992
rect 9496 4972 9548 4992
rect 9548 4972 9550 4992
rect 9494 4936 9550 4972
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9878 14170
rect 9878 14118 9908 14170
rect 9932 14118 9942 14170
rect 9942 14118 9988 14170
rect 10012 14118 10058 14170
rect 10058 14118 10068 14170
rect 10092 14118 10122 14170
rect 10122 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9878 13082
rect 9878 13030 9908 13082
rect 9932 13030 9942 13082
rect 9942 13030 9988 13082
rect 10012 13030 10058 13082
rect 10058 13030 10068 13082
rect 10092 13030 10122 13082
rect 10122 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9878 11994
rect 9878 11942 9908 11994
rect 9932 11942 9942 11994
rect 9942 11942 9988 11994
rect 10012 11942 10058 11994
rect 10058 11942 10068 11994
rect 10092 11942 10122 11994
rect 10122 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9878 10906
rect 9878 10854 9908 10906
rect 9932 10854 9942 10906
rect 9942 10854 9988 10906
rect 10012 10854 10058 10906
rect 10058 10854 10068 10906
rect 10092 10854 10122 10906
rect 10122 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 9770 10648 9826 10704
rect 10138 10240 10194 10296
rect 9678 9324 9680 9344
rect 9680 9324 9732 9344
rect 9732 9324 9734 9344
rect 9678 9288 9734 9324
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9878 9818
rect 9878 9766 9908 9818
rect 9932 9766 9942 9818
rect 9942 9766 9988 9818
rect 10012 9766 10058 9818
rect 10058 9766 10068 9818
rect 10092 9766 10122 9818
rect 10122 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 9678 8880 9734 8936
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9878 8730
rect 9878 8678 9908 8730
rect 9932 8678 9942 8730
rect 9942 8678 9988 8730
rect 10012 8678 10058 8730
rect 10058 8678 10068 8730
rect 10092 8678 10122 8730
rect 10122 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 9954 8064 10010 8120
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9878 7642
rect 9878 7590 9908 7642
rect 9932 7590 9942 7642
rect 9942 7590 9988 7642
rect 10012 7590 10058 7642
rect 10058 7590 10068 7642
rect 10092 7590 10122 7642
rect 10122 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 10138 7112 10194 7168
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9878 6554
rect 9878 6502 9908 6554
rect 9932 6502 9942 6554
rect 9942 6502 9988 6554
rect 10012 6502 10058 6554
rect 10058 6502 10068 6554
rect 10092 6502 10122 6554
rect 10122 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9878 5466
rect 9878 5414 9908 5466
rect 9932 5414 9942 5466
rect 9942 5414 9988 5466
rect 10012 5414 10058 5466
rect 10058 5414 10068 5466
rect 10092 5414 10122 5466
rect 10122 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9878 4378
rect 9878 4326 9908 4378
rect 9932 4326 9942 4378
rect 9942 4326 9988 4378
rect 10012 4326 10058 4378
rect 10058 4326 10068 4378
rect 10092 4326 10122 4378
rect 10122 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9878 3290
rect 9878 3238 9908 3290
rect 9932 3238 9942 3290
rect 9942 3238 9988 3290
rect 10012 3238 10058 3290
rect 10058 3238 10068 3290
rect 10092 3238 10122 3290
rect 10122 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 10690 7384 10746 7440
rect 10322 2916 10378 2952
rect 10874 8064 10930 8120
rect 10322 2896 10324 2916
rect 10324 2896 10376 2916
rect 10376 2896 10378 2916
rect 10506 2524 10508 2544
rect 10508 2524 10560 2544
rect 10560 2524 10562 2544
rect 10506 2488 10562 2524
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9878 2202
rect 9878 2150 9908 2202
rect 9932 2150 9942 2202
rect 9942 2150 9988 2202
rect 10012 2150 10058 2202
rect 10058 2150 10068 2202
rect 10092 2150 10122 2202
rect 10122 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 10782 2896 10838 2952
rect 11242 12144 11298 12200
rect 11058 10240 11114 10296
rect 11150 8880 11206 8936
rect 11058 8608 11114 8664
rect 11242 7248 11298 7304
rect 11058 2760 11114 2816
rect 11610 11056 11666 11112
rect 11610 10004 11612 10024
rect 11612 10004 11664 10024
rect 11664 10004 11666 10024
rect 11610 9968 11666 10004
rect 11610 9560 11666 9616
rect 11702 4972 11704 4992
rect 11704 4972 11756 4992
rect 11756 4972 11758 4992
rect 11702 4936 11758 4972
rect 12817 14714 12873 14716
rect 12897 14714 12953 14716
rect 12977 14714 13033 14716
rect 13057 14714 13113 14716
rect 12817 14662 12843 14714
rect 12843 14662 12873 14714
rect 12897 14662 12907 14714
rect 12907 14662 12953 14714
rect 12977 14662 13023 14714
rect 13023 14662 13033 14714
rect 13057 14662 13087 14714
rect 13087 14662 13113 14714
rect 12817 14660 12873 14662
rect 12897 14660 12953 14662
rect 12977 14660 13033 14662
rect 13057 14660 13113 14662
rect 12817 13626 12873 13628
rect 12897 13626 12953 13628
rect 12977 13626 13033 13628
rect 13057 13626 13113 13628
rect 12817 13574 12843 13626
rect 12843 13574 12873 13626
rect 12897 13574 12907 13626
rect 12907 13574 12953 13626
rect 12977 13574 13023 13626
rect 13023 13574 13033 13626
rect 13057 13574 13087 13626
rect 13087 13574 13113 13626
rect 12817 13572 12873 13574
rect 12897 13572 12953 13574
rect 12977 13572 13033 13574
rect 13057 13572 13113 13574
rect 11978 9152 12034 9208
rect 11978 8880 12034 8936
rect 12162 9560 12218 9616
rect 11886 7248 11942 7304
rect 12346 10784 12402 10840
rect 12346 9424 12402 9480
rect 13174 13096 13230 13152
rect 12817 12538 12873 12540
rect 12897 12538 12953 12540
rect 12977 12538 13033 12540
rect 13057 12538 13113 12540
rect 12817 12486 12843 12538
rect 12843 12486 12873 12538
rect 12897 12486 12907 12538
rect 12907 12486 12953 12538
rect 12977 12486 13023 12538
rect 13023 12486 13033 12538
rect 13057 12486 13087 12538
rect 13087 12486 13113 12538
rect 12817 12484 12873 12486
rect 12897 12484 12953 12486
rect 12977 12484 13033 12486
rect 13057 12484 13113 12486
rect 12438 9152 12494 9208
rect 12438 9016 12494 9072
rect 12346 7112 12402 7168
rect 11794 2508 11850 2544
rect 11794 2488 11796 2508
rect 11796 2488 11848 2508
rect 11848 2488 11850 2508
rect 12817 11450 12873 11452
rect 12897 11450 12953 11452
rect 12977 11450 13033 11452
rect 13057 11450 13113 11452
rect 12817 11398 12843 11450
rect 12843 11398 12873 11450
rect 12897 11398 12907 11450
rect 12907 11398 12953 11450
rect 12977 11398 13023 11450
rect 13023 11398 13033 11450
rect 13057 11398 13087 11450
rect 13087 11398 13113 11450
rect 12817 11396 12873 11398
rect 12897 11396 12953 11398
rect 12977 11396 13033 11398
rect 13057 11396 13113 11398
rect 12817 10362 12873 10364
rect 12897 10362 12953 10364
rect 12977 10362 13033 10364
rect 13057 10362 13113 10364
rect 12817 10310 12843 10362
rect 12843 10310 12873 10362
rect 12897 10310 12907 10362
rect 12907 10310 12953 10362
rect 12977 10310 13023 10362
rect 13023 10310 13033 10362
rect 13057 10310 13087 10362
rect 13087 10310 13113 10362
rect 12817 10308 12873 10310
rect 12897 10308 12953 10310
rect 12977 10308 13033 10310
rect 13057 10308 13113 10310
rect 12806 10140 12808 10160
rect 12808 10140 12860 10160
rect 12860 10140 12862 10160
rect 12806 10104 12862 10140
rect 12806 10004 12808 10024
rect 12808 10004 12860 10024
rect 12860 10004 12862 10024
rect 12806 9968 12862 10004
rect 13082 9968 13138 10024
rect 12817 9274 12873 9276
rect 12897 9274 12953 9276
rect 12977 9274 13033 9276
rect 13057 9274 13113 9276
rect 12817 9222 12843 9274
rect 12843 9222 12873 9274
rect 12897 9222 12907 9274
rect 12907 9222 12953 9274
rect 12977 9222 13023 9274
rect 13023 9222 13033 9274
rect 13057 9222 13087 9274
rect 13087 9222 13113 9274
rect 12817 9220 12873 9222
rect 12897 9220 12953 9222
rect 12977 9220 13033 9222
rect 13057 9220 13113 9222
rect 12806 8356 12862 8392
rect 12806 8336 12808 8356
rect 12808 8336 12860 8356
rect 12860 8336 12862 8356
rect 12817 8186 12873 8188
rect 12897 8186 12953 8188
rect 12977 8186 13033 8188
rect 13057 8186 13113 8188
rect 12817 8134 12843 8186
rect 12843 8134 12873 8186
rect 12897 8134 12907 8186
rect 12907 8134 12953 8186
rect 12977 8134 13023 8186
rect 13023 8134 13033 8186
rect 13057 8134 13087 8186
rect 13087 8134 13113 8186
rect 12817 8132 12873 8134
rect 12897 8132 12953 8134
rect 12977 8132 13033 8134
rect 13057 8132 13113 8134
rect 12817 7098 12873 7100
rect 12897 7098 12953 7100
rect 12977 7098 13033 7100
rect 13057 7098 13113 7100
rect 12817 7046 12843 7098
rect 12843 7046 12873 7098
rect 12897 7046 12907 7098
rect 12907 7046 12953 7098
rect 12977 7046 13023 7098
rect 13023 7046 13033 7098
rect 13057 7046 13087 7098
rect 13087 7046 13113 7098
rect 12817 7044 12873 7046
rect 12897 7044 12953 7046
rect 12977 7044 13033 7046
rect 13057 7044 13113 7046
rect 13174 6740 13176 6760
rect 13176 6740 13228 6760
rect 13228 6740 13230 6760
rect 13174 6704 13230 6740
rect 12817 6010 12873 6012
rect 12897 6010 12953 6012
rect 12977 6010 13033 6012
rect 13057 6010 13113 6012
rect 12817 5958 12843 6010
rect 12843 5958 12873 6010
rect 12897 5958 12907 6010
rect 12907 5958 12953 6010
rect 12977 5958 13023 6010
rect 13023 5958 13033 6010
rect 13057 5958 13087 6010
rect 13087 5958 13113 6010
rect 12817 5956 12873 5958
rect 12897 5956 12953 5958
rect 12977 5956 13033 5958
rect 13057 5956 13113 5958
rect 12714 5616 12770 5672
rect 13174 5616 13230 5672
rect 12817 4922 12873 4924
rect 12897 4922 12953 4924
rect 12977 4922 13033 4924
rect 13057 4922 13113 4924
rect 12817 4870 12843 4922
rect 12843 4870 12873 4922
rect 12897 4870 12907 4922
rect 12907 4870 12953 4922
rect 12977 4870 13023 4922
rect 13023 4870 13033 4922
rect 13057 4870 13087 4922
rect 13087 4870 13113 4922
rect 12817 4868 12873 4870
rect 12897 4868 12953 4870
rect 12977 4868 13033 4870
rect 13057 4868 13113 4870
rect 13450 10512 13506 10568
rect 13358 9016 13414 9072
rect 13358 8916 13360 8936
rect 13360 8916 13412 8936
rect 13412 8916 13414 8936
rect 13358 8880 13414 8916
rect 13358 5072 13414 5128
rect 12817 3834 12873 3836
rect 12897 3834 12953 3836
rect 12977 3834 13033 3836
rect 13057 3834 13113 3836
rect 12817 3782 12843 3834
rect 12843 3782 12873 3834
rect 12897 3782 12907 3834
rect 12907 3782 12953 3834
rect 12977 3782 13023 3834
rect 13023 3782 13033 3834
rect 13057 3782 13087 3834
rect 13087 3782 13113 3834
rect 12817 3780 12873 3782
rect 12897 3780 12953 3782
rect 12977 3780 13033 3782
rect 13057 3780 13113 3782
rect 12817 2746 12873 2748
rect 12897 2746 12953 2748
rect 12977 2746 13033 2748
rect 13057 2746 13113 2748
rect 12817 2694 12843 2746
rect 12843 2694 12873 2746
rect 12897 2694 12907 2746
rect 12907 2694 12953 2746
rect 12977 2694 13023 2746
rect 13023 2694 13033 2746
rect 13057 2694 13087 2746
rect 13087 2694 13113 2746
rect 12817 2692 12873 2694
rect 12897 2692 12953 2694
rect 12977 2692 13033 2694
rect 13057 2692 13113 2694
rect 13634 7948 13690 7984
rect 13634 7928 13636 7948
rect 13636 7928 13688 7948
rect 13688 7928 13690 7948
rect 13634 7148 13636 7168
rect 13636 7148 13688 7168
rect 13688 7148 13690 7168
rect 13634 7112 13690 7148
rect 13542 3848 13598 3904
rect 13818 10512 13874 10568
rect 13818 9424 13874 9480
rect 13818 6704 13874 6760
rect 14002 6704 14058 6760
rect 3238 176 3294 232
rect 14370 9424 14426 9480
rect 14922 13368 14978 13424
rect 15106 13388 15162 13424
rect 15106 13368 15108 13388
rect 15108 13368 15160 13388
rect 15160 13368 15162 13388
rect 15382 15000 15438 15056
rect 15106 12552 15162 12608
rect 14738 8064 14794 8120
rect 14738 6840 14794 6896
rect 14462 3596 14518 3632
rect 14462 3576 14464 3596
rect 14464 3576 14516 3596
rect 14516 3576 14518 3596
rect 15014 11736 15070 11792
rect 15566 14592 15622 14648
rect 15934 16224 15990 16280
rect 15566 13776 15622 13832
rect 16302 14184 16358 14240
rect 15782 14170 15838 14172
rect 15862 14170 15918 14172
rect 15942 14170 15998 14172
rect 16022 14170 16078 14172
rect 15782 14118 15808 14170
rect 15808 14118 15838 14170
rect 15862 14118 15872 14170
rect 15872 14118 15918 14170
rect 15942 14118 15988 14170
rect 15988 14118 15998 14170
rect 16022 14118 16052 14170
rect 16052 14118 16078 14170
rect 15782 14116 15838 14118
rect 15862 14116 15918 14118
rect 15942 14116 15998 14118
rect 16022 14116 16078 14118
rect 15474 13640 15530 13696
rect 15382 12688 15438 12744
rect 15290 12416 15346 12472
rect 15290 10140 15292 10160
rect 15292 10140 15344 10160
rect 15344 10140 15346 10160
rect 15290 10104 15346 10140
rect 15014 8608 15070 8664
rect 15290 8880 15346 8936
rect 15014 7928 15070 7984
rect 14922 3984 14978 4040
rect 15290 7792 15346 7848
rect 15290 6296 15346 6352
rect 15290 5208 15346 5264
rect 15658 13640 15714 13696
rect 15566 12144 15622 12200
rect 15782 13082 15838 13084
rect 15862 13082 15918 13084
rect 15942 13082 15998 13084
rect 16022 13082 16078 13084
rect 15782 13030 15808 13082
rect 15808 13030 15838 13082
rect 15862 13030 15872 13082
rect 15872 13030 15918 13082
rect 15942 13030 15988 13082
rect 15988 13030 15998 13082
rect 16022 13030 16052 13082
rect 16052 13030 16078 13082
rect 15782 13028 15838 13030
rect 15862 13028 15918 13030
rect 15942 13028 15998 13030
rect 16022 13028 16078 13030
rect 16210 12552 16266 12608
rect 15474 10512 15530 10568
rect 15782 11994 15838 11996
rect 15862 11994 15918 11996
rect 15942 11994 15998 11996
rect 16022 11994 16078 11996
rect 15782 11942 15808 11994
rect 15808 11942 15838 11994
rect 15862 11942 15872 11994
rect 15872 11942 15918 11994
rect 15942 11942 15988 11994
rect 15988 11942 15998 11994
rect 16022 11942 16052 11994
rect 16052 11942 16078 11994
rect 15782 11940 15838 11942
rect 15862 11940 15918 11942
rect 15942 11940 15998 11942
rect 16022 11940 16078 11942
rect 15782 10906 15838 10908
rect 15862 10906 15918 10908
rect 15942 10906 15998 10908
rect 16022 10906 16078 10908
rect 15782 10854 15808 10906
rect 15808 10854 15838 10906
rect 15862 10854 15872 10906
rect 15872 10854 15918 10906
rect 15942 10854 15988 10906
rect 15988 10854 15998 10906
rect 16022 10854 16052 10906
rect 16052 10854 16078 10906
rect 15782 10852 15838 10854
rect 15862 10852 15918 10854
rect 15942 10852 15998 10854
rect 16022 10852 16078 10854
rect 15566 9968 15622 10024
rect 15566 9696 15622 9752
rect 15782 9818 15838 9820
rect 15862 9818 15918 9820
rect 15942 9818 15998 9820
rect 16022 9818 16078 9820
rect 15782 9766 15808 9818
rect 15808 9766 15838 9818
rect 15862 9766 15872 9818
rect 15872 9766 15918 9818
rect 15942 9766 15988 9818
rect 15988 9766 15998 9818
rect 16022 9766 16052 9818
rect 16052 9766 16078 9818
rect 15782 9764 15838 9766
rect 15862 9764 15918 9766
rect 15942 9764 15998 9766
rect 16022 9764 16078 9766
rect 15474 6840 15530 6896
rect 15658 9016 15714 9072
rect 15782 8730 15838 8732
rect 15862 8730 15918 8732
rect 15942 8730 15998 8732
rect 16022 8730 16078 8732
rect 15782 8678 15808 8730
rect 15808 8678 15838 8730
rect 15862 8678 15872 8730
rect 15872 8678 15918 8730
rect 15942 8678 15988 8730
rect 15988 8678 15998 8730
rect 16022 8678 16052 8730
rect 16052 8678 16078 8730
rect 15782 8676 15838 8678
rect 15862 8676 15918 8678
rect 15942 8676 15998 8678
rect 16022 8676 16078 8678
rect 15750 8200 15806 8256
rect 16026 8084 16082 8120
rect 16026 8064 16028 8084
rect 16028 8064 16080 8084
rect 16080 8064 16082 8084
rect 15782 7642 15838 7644
rect 15862 7642 15918 7644
rect 15942 7642 15998 7644
rect 16022 7642 16078 7644
rect 15782 7590 15808 7642
rect 15808 7590 15838 7642
rect 15862 7590 15872 7642
rect 15872 7590 15918 7642
rect 15942 7590 15988 7642
rect 15988 7590 15998 7642
rect 16022 7590 16052 7642
rect 16052 7590 16078 7642
rect 15782 7588 15838 7590
rect 15862 7588 15918 7590
rect 15942 7588 15998 7590
rect 16022 7588 16078 7590
rect 15782 6554 15838 6556
rect 15862 6554 15918 6556
rect 15942 6554 15998 6556
rect 16022 6554 16078 6556
rect 15782 6502 15808 6554
rect 15808 6502 15838 6554
rect 15862 6502 15872 6554
rect 15872 6502 15918 6554
rect 15942 6502 15988 6554
rect 15988 6502 15998 6554
rect 16022 6502 16052 6554
rect 16052 6502 16078 6554
rect 15782 6500 15838 6502
rect 15862 6500 15918 6502
rect 15942 6500 15998 6502
rect 16022 6500 16078 6502
rect 15782 5466 15838 5468
rect 15862 5466 15918 5468
rect 15942 5466 15998 5468
rect 16022 5466 16078 5468
rect 15782 5414 15808 5466
rect 15808 5414 15838 5466
rect 15862 5414 15872 5466
rect 15872 5414 15918 5466
rect 15942 5414 15988 5466
rect 15988 5414 15998 5466
rect 16022 5414 16052 5466
rect 16052 5414 16078 5466
rect 15782 5412 15838 5414
rect 15862 5412 15918 5414
rect 15942 5412 15998 5414
rect 16022 5412 16078 5414
rect 16026 5072 16082 5128
rect 15658 4800 15714 4856
rect 15782 4378 15838 4380
rect 15862 4378 15918 4380
rect 15942 4378 15998 4380
rect 16022 4378 16078 4380
rect 15782 4326 15808 4378
rect 15808 4326 15838 4378
rect 15862 4326 15872 4378
rect 15872 4326 15918 4378
rect 15942 4326 15988 4378
rect 15988 4326 15998 4378
rect 16022 4326 16052 4378
rect 16052 4326 16078 4378
rect 15782 4324 15838 4326
rect 15862 4324 15918 4326
rect 15942 4324 15998 4326
rect 16022 4324 16078 4326
rect 14738 1808 14794 1864
rect 15014 992 15070 1048
rect 15566 2488 15622 2544
rect 15782 3290 15838 3292
rect 15862 3290 15918 3292
rect 15942 3290 15998 3292
rect 16022 3290 16078 3292
rect 15782 3238 15808 3290
rect 15808 3238 15838 3290
rect 15862 3238 15872 3290
rect 15872 3238 15918 3290
rect 15942 3238 15988 3290
rect 15988 3238 15998 3290
rect 16022 3238 16052 3290
rect 16052 3238 16078 3290
rect 15782 3236 15838 3238
rect 15862 3236 15918 3238
rect 15942 3236 15998 3238
rect 16022 3236 16078 3238
rect 15750 2916 15806 2952
rect 15750 2896 15752 2916
rect 15752 2896 15804 2916
rect 15804 2896 15806 2916
rect 16026 2624 16082 2680
rect 15782 2202 15838 2204
rect 15862 2202 15918 2204
rect 15942 2202 15998 2204
rect 16022 2202 16078 2204
rect 15782 2150 15808 2202
rect 15808 2150 15838 2202
rect 15862 2150 15872 2202
rect 15872 2150 15918 2202
rect 15942 2150 15988 2202
rect 15988 2150 15998 2202
rect 16022 2150 16052 2202
rect 16052 2150 16078 2202
rect 15782 2148 15838 2150
rect 15862 2148 15918 2150
rect 15942 2148 15998 2150
rect 16022 2148 16078 2150
rect 16210 4004 16266 4040
rect 16210 3984 16212 4004
rect 16212 3984 16264 4004
rect 16264 3984 16266 4004
rect 16394 4936 16450 4992
rect 16210 3032 16266 3088
rect 16854 11600 16910 11656
rect 16578 10240 16634 10296
rect 16762 8744 16818 8800
rect 16854 8472 16910 8528
rect 16210 2252 16212 2272
rect 16212 2252 16264 2272
rect 16264 2252 16266 2272
rect 16210 2216 16266 2252
rect 17406 9832 17462 9888
rect 18418 15816 18474 15872
rect 18326 13232 18382 13288
rect 17590 9560 17646 9616
rect 17498 6976 17554 7032
rect 17406 5616 17462 5672
rect 17406 4392 17462 4448
rect 16946 3576 17002 3632
rect 17498 2624 17554 2680
rect 17866 9424 17922 9480
rect 17682 3984 17738 4040
rect 18050 7384 18106 7440
rect 18050 6024 18106 6080
rect 18234 11192 18290 11248
rect 18510 6432 18566 6488
rect 18418 584 18474 640
rect 18878 1400 18934 1456
rect 14002 176 14058 232
<< metal3 >>
rect 0 16690 480 16720
rect 3601 16690 3667 16693
rect 0 16688 3667 16690
rect 0 16632 3606 16688
rect 3662 16632 3667 16688
rect 0 16630 3667 16632
rect 0 16600 480 16630
rect 3601 16627 3667 16630
rect 15193 16690 15259 16693
rect 19520 16690 20000 16720
rect 15193 16688 20000 16690
rect 15193 16632 15198 16688
rect 15254 16632 20000 16688
rect 15193 16630 20000 16632
rect 15193 16627 15259 16630
rect 19520 16600 20000 16630
rect 0 16282 480 16312
rect 2405 16282 2471 16285
rect 0 16280 2471 16282
rect 0 16224 2410 16280
rect 2466 16224 2471 16280
rect 0 16222 2471 16224
rect 0 16192 480 16222
rect 2405 16219 2471 16222
rect 15929 16282 15995 16285
rect 19520 16282 20000 16312
rect 15929 16280 20000 16282
rect 15929 16224 15934 16280
rect 15990 16224 20000 16280
rect 15929 16222 20000 16224
rect 15929 16219 15995 16222
rect 19520 16192 20000 16222
rect 0 15874 480 15904
rect 3141 15874 3207 15877
rect 0 15872 3207 15874
rect 0 15816 3146 15872
rect 3202 15816 3207 15872
rect 0 15814 3207 15816
rect 0 15784 480 15814
rect 3141 15811 3207 15814
rect 18413 15874 18479 15877
rect 19520 15874 20000 15904
rect 18413 15872 20000 15874
rect 18413 15816 18418 15872
rect 18474 15816 20000 15872
rect 18413 15814 20000 15816
rect 18413 15811 18479 15814
rect 19520 15784 20000 15814
rect 0 15466 480 15496
rect 9397 15466 9463 15469
rect 0 15464 9463 15466
rect 0 15408 9402 15464
rect 9458 15408 9463 15464
rect 0 15406 9463 15408
rect 0 15376 480 15406
rect 9397 15403 9463 15406
rect 16246 15404 16252 15468
rect 16316 15466 16322 15468
rect 19520 15466 20000 15496
rect 16316 15406 20000 15466
rect 16316 15404 16322 15406
rect 19520 15376 20000 15406
rect 0 15058 480 15088
rect 3785 15058 3851 15061
rect 0 15056 3851 15058
rect 0 15000 3790 15056
rect 3846 15000 3851 15056
rect 0 14998 3851 15000
rect 0 14968 480 14998
rect 3785 14995 3851 14998
rect 15377 15058 15443 15061
rect 19520 15058 20000 15088
rect 15377 15056 20000 15058
rect 15377 15000 15382 15056
rect 15438 15000 20000 15056
rect 15377 14998 20000 15000
rect 15377 14995 15443 14998
rect 19520 14968 20000 14998
rect 6874 14720 7194 14721
rect 0 14650 480 14680
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7194 14720
rect 6874 14655 7194 14656
rect 12805 14720 13125 14721
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 14655 13125 14656
rect 3693 14650 3759 14653
rect 0 14648 3759 14650
rect 0 14592 3698 14648
rect 3754 14592 3759 14648
rect 0 14590 3759 14592
rect 0 14560 480 14590
rect 3693 14587 3759 14590
rect 15561 14650 15627 14653
rect 19520 14650 20000 14680
rect 15561 14648 20000 14650
rect 15561 14592 15566 14648
rect 15622 14592 20000 14648
rect 15561 14590 20000 14592
rect 15561 14587 15627 14590
rect 19520 14560 20000 14590
rect 0 14242 480 14272
rect 3509 14242 3575 14245
rect 0 14240 3575 14242
rect 0 14184 3514 14240
rect 3570 14184 3575 14240
rect 0 14182 3575 14184
rect 0 14152 480 14182
rect 3509 14179 3575 14182
rect 16297 14242 16363 14245
rect 19520 14242 20000 14272
rect 16297 14240 20000 14242
rect 16297 14184 16302 14240
rect 16358 14184 20000 14240
rect 16297 14182 20000 14184
rect 16297 14179 16363 14182
rect 3909 14176 4229 14177
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 14111 4229 14112
rect 9840 14176 10160 14177
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 14111 10160 14112
rect 15770 14176 16090 14177
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 19520 14152 20000 14182
rect 15770 14111 16090 14112
rect 0 13834 480 13864
rect 2221 13834 2287 13837
rect 0 13832 2287 13834
rect 0 13776 2226 13832
rect 2282 13776 2287 13832
rect 0 13774 2287 13776
rect 0 13744 480 13774
rect 2221 13771 2287 13774
rect 15561 13834 15627 13837
rect 19520 13834 20000 13864
rect 15561 13832 20000 13834
rect 15561 13776 15566 13832
rect 15622 13776 20000 13832
rect 15561 13774 20000 13776
rect 15561 13771 15627 13774
rect 19520 13744 20000 13774
rect 15469 13698 15535 13701
rect 15653 13698 15719 13701
rect 15469 13696 15719 13698
rect 15469 13640 15474 13696
rect 15530 13640 15658 13696
rect 15714 13640 15719 13696
rect 15469 13638 15719 13640
rect 15469 13635 15535 13638
rect 15653 13635 15719 13638
rect 6874 13632 7194 13633
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7194 13632
rect 6874 13567 7194 13568
rect 12805 13632 13125 13633
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 13567 13125 13568
rect 0 13426 480 13456
rect 3509 13426 3575 13429
rect 0 13424 3575 13426
rect 0 13368 3514 13424
rect 3570 13368 3575 13424
rect 0 13366 3575 13368
rect 0 13336 480 13366
rect 3509 13363 3575 13366
rect 14774 13364 14780 13428
rect 14844 13426 14850 13428
rect 14917 13426 14983 13429
rect 14844 13424 14983 13426
rect 14844 13368 14922 13424
rect 14978 13368 14983 13424
rect 14844 13366 14983 13368
rect 14844 13364 14850 13366
rect 14917 13363 14983 13366
rect 15101 13428 15167 13429
rect 15101 13424 15148 13428
rect 15212 13426 15218 13428
rect 15101 13368 15106 13424
rect 15101 13364 15148 13368
rect 15212 13366 15258 13426
rect 15212 13364 15218 13366
rect 15101 13363 15167 13364
rect 18321 13290 18387 13293
rect 19520 13290 20000 13320
rect 18321 13288 20000 13290
rect 18321 13232 18326 13288
rect 18382 13232 20000 13288
rect 18321 13230 20000 13232
rect 18321 13227 18387 13230
rect 19520 13200 20000 13230
rect 13169 13154 13235 13157
rect 13302 13154 13308 13156
rect 13169 13152 13308 13154
rect 13169 13096 13174 13152
rect 13230 13096 13308 13152
rect 13169 13094 13308 13096
rect 13169 13091 13235 13094
rect 13302 13092 13308 13094
rect 13372 13092 13378 13156
rect 3909 13088 4229 13089
rect 0 13018 480 13048
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 13023 4229 13024
rect 9840 13088 10160 13089
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 13023 10160 13024
rect 15770 13088 16090 13089
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 15770 13023 16090 13024
rect 3325 13018 3391 13021
rect 0 13016 3391 13018
rect 0 12960 3330 13016
rect 3386 12960 3391 13016
rect 0 12958 3391 12960
rect 0 12928 480 12958
rect 3325 12955 3391 12958
rect 14958 12820 14964 12884
rect 15028 12882 15034 12884
rect 19520 12882 20000 12912
rect 15028 12822 20000 12882
rect 15028 12820 15034 12822
rect 19520 12792 20000 12822
rect 13854 12684 13860 12748
rect 13924 12746 13930 12748
rect 15377 12746 15443 12749
rect 13924 12744 15443 12746
rect 13924 12688 15382 12744
rect 15438 12688 15443 12744
rect 13924 12686 15443 12688
rect 13924 12684 13930 12686
rect 15377 12683 15443 12686
rect 0 12610 480 12640
rect 3049 12610 3115 12613
rect 0 12608 3115 12610
rect 0 12552 3054 12608
rect 3110 12552 3115 12608
rect 0 12550 3115 12552
rect 0 12520 480 12550
rect 3049 12547 3115 12550
rect 15101 12610 15167 12613
rect 16205 12610 16271 12613
rect 16430 12610 16436 12612
rect 15101 12608 15210 12610
rect 15101 12552 15106 12608
rect 15162 12552 15210 12608
rect 15101 12547 15210 12552
rect 16205 12608 16436 12610
rect 16205 12552 16210 12608
rect 16266 12552 16436 12608
rect 16205 12550 16436 12552
rect 16205 12547 16271 12550
rect 16430 12548 16436 12550
rect 16500 12548 16506 12612
rect 6874 12544 7194 12545
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7194 12544
rect 6874 12479 7194 12480
rect 12805 12544 13125 12545
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 12479 13125 12480
rect 8661 12474 8727 12477
rect 10358 12474 10364 12476
rect 8661 12472 10364 12474
rect 8661 12416 8666 12472
rect 8722 12416 10364 12472
rect 8661 12414 10364 12416
rect 8661 12411 8727 12414
rect 10358 12412 10364 12414
rect 10428 12412 10434 12476
rect 15150 12474 15210 12547
rect 15285 12474 15351 12477
rect 15150 12472 15351 12474
rect 15150 12416 15290 12472
rect 15346 12416 15351 12472
rect 15150 12414 15351 12416
rect 15285 12411 15351 12414
rect 15510 12412 15516 12476
rect 15580 12474 15586 12476
rect 19520 12474 20000 12504
rect 15580 12414 20000 12474
rect 15580 12412 15586 12414
rect 19520 12384 20000 12414
rect 2998 12276 3004 12340
rect 3068 12338 3074 12340
rect 3325 12338 3391 12341
rect 3068 12336 3391 12338
rect 3068 12280 3330 12336
rect 3386 12280 3391 12336
rect 3068 12278 3391 12280
rect 3068 12276 3074 12278
rect 3325 12275 3391 12278
rect 4521 12338 4587 12341
rect 6085 12338 6151 12341
rect 4521 12336 6151 12338
rect 4521 12280 4526 12336
rect 4582 12280 6090 12336
rect 6146 12280 6151 12336
rect 4521 12278 6151 12280
rect 4521 12275 4587 12278
rect 6085 12275 6151 12278
rect 6269 12338 6335 12341
rect 9305 12338 9371 12341
rect 6269 12336 9371 12338
rect 6269 12280 6274 12336
rect 6330 12280 9310 12336
rect 9366 12280 9371 12336
rect 6269 12278 9371 12280
rect 6269 12275 6335 12278
rect 9305 12275 9371 12278
rect 0 12202 480 12232
rect 4061 12202 4127 12205
rect 0 12200 4127 12202
rect 0 12144 4066 12200
rect 4122 12144 4127 12200
rect 0 12142 4127 12144
rect 0 12112 480 12142
rect 4061 12139 4127 12142
rect 4245 12202 4311 12205
rect 7465 12202 7531 12205
rect 4245 12200 7531 12202
rect 4245 12144 4250 12200
rect 4306 12144 7470 12200
rect 7526 12144 7531 12200
rect 4245 12142 7531 12144
rect 4245 12139 4311 12142
rect 7465 12139 7531 12142
rect 11237 12202 11303 12205
rect 15561 12202 15627 12205
rect 11237 12200 15627 12202
rect 11237 12144 11242 12200
rect 11298 12144 15566 12200
rect 15622 12144 15627 12200
rect 11237 12142 15627 12144
rect 11237 12139 11303 12142
rect 15561 12139 15627 12142
rect 19520 12066 20000 12096
rect 16208 12006 20000 12066
rect 3909 12000 4229 12001
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 11935 4229 11936
rect 9840 12000 10160 12001
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 11935 10160 11936
rect 15770 12000 16090 12001
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 15770 11935 16090 11936
rect 0 11794 480 11824
rect 3325 11794 3391 11797
rect 0 11792 3391 11794
rect 0 11736 3330 11792
rect 3386 11736 3391 11792
rect 0 11734 3391 11736
rect 0 11704 480 11734
rect 3325 11731 3391 11734
rect 6085 11794 6151 11797
rect 6453 11794 6519 11797
rect 8845 11794 8911 11797
rect 6085 11792 8911 11794
rect 6085 11736 6090 11792
rect 6146 11736 6458 11792
rect 6514 11736 8850 11792
rect 8906 11736 8911 11792
rect 6085 11734 8911 11736
rect 6085 11731 6151 11734
rect 6453 11731 6519 11734
rect 8845 11731 8911 11734
rect 15009 11794 15075 11797
rect 16208 11794 16268 12006
rect 19520 11976 20000 12006
rect 15009 11792 16268 11794
rect 15009 11736 15014 11792
rect 15070 11736 16268 11792
rect 15009 11734 16268 11736
rect 15009 11731 15075 11734
rect 16849 11658 16915 11661
rect 19520 11658 20000 11688
rect 16849 11656 20000 11658
rect 16849 11600 16854 11656
rect 16910 11600 20000 11656
rect 16849 11598 20000 11600
rect 16849 11595 16915 11598
rect 19520 11568 20000 11598
rect 6874 11456 7194 11457
rect 0 11386 480 11416
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7194 11456
rect 6874 11391 7194 11392
rect 12805 11456 13125 11457
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 11391 13125 11392
rect 3141 11386 3207 11389
rect 0 11384 3207 11386
rect 0 11328 3146 11384
rect 3202 11328 3207 11384
rect 0 11326 3207 11328
rect 0 11296 480 11326
rect 3141 11323 3207 11326
rect 18229 11250 18295 11253
rect 19520 11250 20000 11280
rect 18229 11248 20000 11250
rect 18229 11192 18234 11248
rect 18290 11192 20000 11248
rect 18229 11190 20000 11192
rect 18229 11187 18295 11190
rect 19520 11160 20000 11190
rect 8661 11114 8727 11117
rect 11278 11114 11284 11116
rect 8661 11112 11284 11114
rect 8661 11056 8666 11112
rect 8722 11056 11284 11112
rect 8661 11054 11284 11056
rect 8661 11051 8727 11054
rect 11278 11052 11284 11054
rect 11348 11114 11354 11116
rect 11605 11114 11671 11117
rect 11348 11112 11671 11114
rect 11348 11056 11610 11112
rect 11666 11056 11671 11112
rect 11348 11054 11671 11056
rect 11348 11052 11354 11054
rect 11605 11051 11671 11054
rect 0 10978 480 11008
rect 0 10918 3848 10978
rect 0 10888 480 10918
rect 3788 10706 3848 10918
rect 3909 10912 4229 10913
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 10847 4229 10848
rect 9840 10912 10160 10913
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 10847 10160 10848
rect 15770 10912 16090 10913
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15770 10847 16090 10848
rect 12014 10780 12020 10844
rect 12084 10842 12090 10844
rect 12341 10842 12407 10845
rect 19520 10842 20000 10872
rect 12084 10840 12407 10842
rect 12084 10784 12346 10840
rect 12402 10784 12407 10840
rect 12084 10782 12407 10784
rect 12084 10780 12090 10782
rect 12341 10779 12407 10782
rect 16208 10782 20000 10842
rect 5165 10706 5231 10709
rect 3788 10704 5231 10706
rect 3788 10648 5170 10704
rect 5226 10648 5231 10704
rect 3788 10646 5231 10648
rect 5165 10643 5231 10646
rect 9765 10706 9831 10709
rect 16208 10706 16268 10782
rect 19520 10752 20000 10782
rect 9765 10704 16268 10706
rect 9765 10648 9770 10704
rect 9826 10648 16268 10704
rect 9765 10646 16268 10648
rect 9765 10643 9831 10646
rect 0 10570 480 10600
rect 8293 10570 8359 10573
rect 0 10568 8359 10570
rect 0 10512 8298 10568
rect 8354 10512 8359 10568
rect 0 10510 8359 10512
rect 0 10480 480 10510
rect 8293 10507 8359 10510
rect 8845 10570 8911 10573
rect 13445 10570 13511 10573
rect 13813 10570 13879 10573
rect 8845 10568 13370 10570
rect 8845 10512 8850 10568
rect 8906 10512 13370 10568
rect 8845 10510 13370 10512
rect 8845 10507 8911 10510
rect 2681 10434 2747 10437
rect 2865 10434 2931 10437
rect 2681 10432 2931 10434
rect 2681 10376 2686 10432
rect 2742 10376 2870 10432
rect 2926 10376 2931 10432
rect 2681 10374 2931 10376
rect 13310 10434 13370 10510
rect 13445 10568 13879 10570
rect 13445 10512 13450 10568
rect 13506 10512 13818 10568
rect 13874 10512 13879 10568
rect 13445 10510 13879 10512
rect 13445 10507 13511 10510
rect 13813 10507 13879 10510
rect 15469 10570 15535 10573
rect 16798 10570 16804 10572
rect 15469 10568 16804 10570
rect 15469 10512 15474 10568
rect 15530 10512 16804 10568
rect 15469 10510 16804 10512
rect 15469 10507 15535 10510
rect 16798 10508 16804 10510
rect 16868 10508 16874 10572
rect 19520 10434 20000 10464
rect 13310 10374 20000 10434
rect 2681 10371 2747 10374
rect 2865 10371 2931 10374
rect 6874 10368 7194 10369
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7194 10368
rect 6874 10303 7194 10304
rect 12805 10368 13125 10369
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 19520 10344 20000 10374
rect 12805 10303 13125 10304
rect 3550 10236 3556 10300
rect 3620 10298 3626 10300
rect 6729 10298 6795 10301
rect 3620 10296 6795 10298
rect 3620 10240 6734 10296
rect 6790 10240 6795 10296
rect 3620 10238 6795 10240
rect 3620 10236 3626 10238
rect 6729 10235 6795 10238
rect 10133 10298 10199 10301
rect 11053 10298 11119 10301
rect 16573 10298 16639 10301
rect 10133 10296 11119 10298
rect 10133 10240 10138 10296
rect 10194 10240 11058 10296
rect 11114 10240 11119 10296
rect 10133 10238 11119 10240
rect 10133 10235 10199 10238
rect 11053 10235 11119 10238
rect 14598 10296 16639 10298
rect 14598 10240 16578 10296
rect 16634 10240 16639 10296
rect 14598 10238 16639 10240
rect 0 10162 480 10192
rect 5533 10162 5599 10165
rect 0 10160 5599 10162
rect 0 10104 5538 10160
rect 5594 10104 5599 10160
rect 0 10102 5599 10104
rect 0 10072 480 10102
rect 5533 10099 5599 10102
rect 9121 10162 9187 10165
rect 12801 10162 12867 10165
rect 9121 10160 12867 10162
rect 9121 10104 9126 10160
rect 9182 10104 12806 10160
rect 12862 10104 12867 10160
rect 9121 10102 12867 10104
rect 9121 10099 9187 10102
rect 12801 10099 12867 10102
rect 2589 10026 2655 10029
rect 7465 10026 7531 10029
rect 2589 10024 7531 10026
rect 2589 9968 2594 10024
rect 2650 9968 7470 10024
rect 7526 9968 7531 10024
rect 2589 9966 7531 9968
rect 2589 9963 2655 9966
rect 7465 9963 7531 9966
rect 11605 10026 11671 10029
rect 12801 10026 12867 10029
rect 11605 10024 12867 10026
rect 11605 9968 11610 10024
rect 11666 9968 12806 10024
rect 12862 9968 12867 10024
rect 11605 9966 12867 9968
rect 11605 9963 11671 9966
rect 12801 9963 12867 9966
rect 13077 10026 13143 10029
rect 14598 10026 14658 10238
rect 16573 10235 16639 10238
rect 15285 10162 15351 10165
rect 16614 10162 16620 10164
rect 15285 10160 16620 10162
rect 15285 10104 15290 10160
rect 15346 10104 16620 10160
rect 15285 10102 16620 10104
rect 15285 10099 15351 10102
rect 16614 10100 16620 10102
rect 16684 10100 16690 10164
rect 13077 10024 14658 10026
rect 13077 9968 13082 10024
rect 13138 9968 14658 10024
rect 13077 9966 14658 9968
rect 15561 10024 15627 10029
rect 15561 9968 15566 10024
rect 15622 9968 15627 10024
rect 13077 9963 13143 9966
rect 15561 9963 15627 9968
rect 3509 9892 3575 9893
rect 3509 9890 3556 9892
rect 3464 9888 3556 9890
rect 3464 9832 3514 9888
rect 3464 9830 3556 9832
rect 3509 9828 3556 9830
rect 3620 9828 3626 9892
rect 6269 9890 6335 9893
rect 9489 9890 9555 9893
rect 6269 9888 9555 9890
rect 6269 9832 6274 9888
rect 6330 9832 9494 9888
rect 9550 9832 9555 9888
rect 6269 9830 9555 9832
rect 3509 9827 3575 9828
rect 6269 9827 6335 9830
rect 9489 9827 9555 9830
rect 3909 9824 4229 9825
rect 0 9754 480 9784
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 9759 4229 9760
rect 9840 9824 10160 9825
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 9759 10160 9760
rect 15564 9757 15624 9963
rect 17401 9890 17467 9893
rect 19520 9890 20000 9920
rect 17401 9888 20000 9890
rect 17401 9832 17406 9888
rect 17462 9832 20000 9888
rect 17401 9830 20000 9832
rect 17401 9827 17467 9830
rect 15770 9824 16090 9825
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 19520 9800 20000 9830
rect 15770 9759 16090 9760
rect 2589 9754 2655 9757
rect 0 9752 2655 9754
rect 0 9696 2594 9752
rect 2650 9696 2655 9752
rect 0 9694 2655 9696
rect 0 9664 480 9694
rect 2589 9691 2655 9694
rect 15561 9752 15627 9757
rect 15561 9696 15566 9752
rect 15622 9696 15627 9752
rect 15561 9691 15627 9696
rect 5441 9618 5507 9621
rect 8845 9618 8911 9621
rect 11605 9618 11671 9621
rect 12157 9618 12223 9621
rect 5441 9616 11530 9618
rect 5441 9560 5446 9616
rect 5502 9560 8850 9616
rect 8906 9560 11530 9616
rect 5441 9558 11530 9560
rect 5441 9555 5507 9558
rect 8845 9555 8911 9558
rect 5257 9482 5323 9485
rect 6453 9482 6519 9485
rect 11470 9482 11530 9558
rect 11605 9616 12223 9618
rect 11605 9560 11610 9616
rect 11666 9560 12162 9616
rect 12218 9560 12223 9616
rect 11605 9558 12223 9560
rect 11605 9555 11671 9558
rect 12157 9555 12223 9558
rect 12382 9556 12388 9620
rect 12452 9618 12458 9620
rect 17585 9618 17651 9621
rect 12452 9616 17651 9618
rect 12452 9560 17590 9616
rect 17646 9560 17651 9616
rect 12452 9558 17651 9560
rect 12452 9556 12458 9558
rect 17585 9555 17651 9558
rect 12341 9482 12407 9485
rect 13813 9482 13879 9485
rect 5257 9480 6519 9482
rect 5257 9424 5262 9480
rect 5318 9424 6458 9480
rect 6514 9424 6519 9480
rect 5257 9422 6519 9424
rect 5257 9419 5323 9422
rect 6453 9419 6519 9422
rect 6686 9422 9690 9482
rect 0 9346 480 9376
rect 3969 9346 4035 9349
rect 0 9344 4035 9346
rect 0 9288 3974 9344
rect 4030 9288 4035 9344
rect 0 9286 4035 9288
rect 0 9256 480 9286
rect 3969 9283 4035 9286
rect 4153 9346 4219 9349
rect 4981 9346 5047 9349
rect 6686 9346 6746 9422
rect 9630 9380 9690 9422
rect 10550 9422 10932 9482
rect 11470 9480 13879 9482
rect 11470 9424 12346 9480
rect 12402 9424 13818 9480
rect 13874 9424 13879 9480
rect 11470 9422 13879 9424
rect 4153 9344 6746 9346
rect 4153 9288 4158 9344
rect 4214 9288 4986 9344
rect 5042 9288 6746 9344
rect 4153 9286 6746 9288
rect 7465 9344 7531 9349
rect 7465 9288 7470 9344
rect 7526 9288 7531 9344
rect 4153 9283 4219 9286
rect 4981 9283 5047 9286
rect 7465 9283 7531 9288
rect 7925 9346 7991 9349
rect 8753 9348 8819 9349
rect 8150 9346 8156 9348
rect 7925 9344 8156 9346
rect 7925 9288 7930 9344
rect 7986 9288 8156 9344
rect 7925 9286 8156 9288
rect 7925 9283 7991 9286
rect 8150 9284 8156 9286
rect 8220 9284 8226 9348
rect 8702 9346 8708 9348
rect 8662 9286 8708 9346
rect 8772 9344 8819 9348
rect 8814 9288 8819 9344
rect 9630 9346 9874 9380
rect 10550 9346 10610 9422
rect 9630 9344 10610 9346
rect 9630 9320 9678 9344
rect 8702 9284 8708 9286
rect 8772 9284 8819 9288
rect 8753 9283 8819 9284
rect 9673 9288 9678 9320
rect 9734 9320 10610 9344
rect 9734 9288 9739 9320
rect 9673 9283 9739 9288
rect 9814 9286 10610 9320
rect 10872 9346 10932 9422
rect 12341 9419 12407 9422
rect 13813 9419 13879 9422
rect 14365 9484 14431 9485
rect 14365 9480 14412 9484
rect 14476 9482 14482 9484
rect 17861 9482 17927 9485
rect 19520 9482 20000 9512
rect 14365 9424 14370 9480
rect 14365 9420 14412 9424
rect 14476 9422 14522 9482
rect 17861 9480 20000 9482
rect 17861 9424 17866 9480
rect 17922 9424 20000 9480
rect 17861 9422 20000 9424
rect 14476 9420 14482 9422
rect 14365 9419 14431 9420
rect 17861 9419 17927 9422
rect 19520 9392 20000 9422
rect 12014 9346 12020 9348
rect 10872 9286 12020 9346
rect 12014 9284 12020 9286
rect 12084 9284 12090 9348
rect 6874 9280 7194 9281
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7194 9280
rect 6874 9215 7194 9216
rect 7468 9210 7528 9283
rect 12805 9280 13125 9281
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 9215 13125 9216
rect 11973 9210 12039 9213
rect 7468 9208 12039 9210
rect 7468 9152 11978 9208
rect 12034 9152 12039 9208
rect 7468 9150 12039 9152
rect 11973 9147 12039 9150
rect 12433 9210 12499 9213
rect 12566 9210 12572 9212
rect 12433 9208 12572 9210
rect 12433 9152 12438 9208
rect 12494 9152 12572 9208
rect 12433 9150 12572 9152
rect 12433 9147 12499 9150
rect 12566 9148 12572 9150
rect 12636 9148 12642 9212
rect 3601 9074 3667 9077
rect 12433 9074 12499 9077
rect 13353 9074 13419 9077
rect 15653 9074 15719 9077
rect 19520 9074 20000 9104
rect 3601 9072 13419 9074
rect 3601 9016 3606 9072
rect 3662 9016 12438 9072
rect 12494 9016 13358 9072
rect 13414 9016 13419 9072
rect 3601 9014 13419 9016
rect 3601 9011 3667 9014
rect 12433 9011 12499 9014
rect 13353 9011 13419 9014
rect 13494 9072 20000 9074
rect 13494 9016 15658 9072
rect 15714 9016 20000 9072
rect 13494 9014 20000 9016
rect 0 8938 480 8968
rect 4153 8938 4219 8941
rect 0 8936 4219 8938
rect 0 8880 4158 8936
rect 4214 8880 4219 8936
rect 0 8878 4219 8880
rect 0 8848 480 8878
rect 4153 8875 4219 8878
rect 7189 8938 7255 8941
rect 7925 8940 7991 8941
rect 7925 8938 7972 8940
rect 7189 8936 7972 8938
rect 7189 8880 7194 8936
rect 7250 8880 7930 8936
rect 7189 8878 7972 8880
rect 7189 8875 7255 8878
rect 7925 8876 7972 8878
rect 8036 8876 8042 8940
rect 8845 8938 8911 8941
rect 9489 8938 9555 8941
rect 8845 8936 9555 8938
rect 8845 8880 8850 8936
rect 8906 8880 9494 8936
rect 9550 8880 9555 8936
rect 8845 8878 9555 8880
rect 7925 8875 7991 8876
rect 8845 8875 8911 8878
rect 9489 8875 9555 8878
rect 9673 8938 9739 8941
rect 11145 8938 11211 8941
rect 11278 8938 11284 8940
rect 9673 8936 10426 8938
rect 9673 8880 9678 8936
rect 9734 8880 10426 8936
rect 9673 8878 10426 8880
rect 9673 8875 9739 8878
rect 8753 8804 8819 8805
rect 8702 8740 8708 8804
rect 8772 8802 8819 8804
rect 10366 8802 10426 8878
rect 11145 8936 11284 8938
rect 11145 8880 11150 8936
rect 11206 8880 11284 8936
rect 11145 8878 11284 8880
rect 11145 8875 11211 8878
rect 11278 8876 11284 8878
rect 11348 8876 11354 8940
rect 11830 8876 11836 8940
rect 11900 8938 11906 8940
rect 11973 8938 12039 8941
rect 13353 8938 13419 8941
rect 11900 8936 13419 8938
rect 11900 8880 11978 8936
rect 12034 8880 13358 8936
rect 13414 8880 13419 8936
rect 11900 8878 13419 8880
rect 11900 8876 11906 8878
rect 11973 8875 12039 8878
rect 13353 8875 13419 8878
rect 13494 8802 13554 9014
rect 15653 9011 15719 9014
rect 19520 8984 20000 9014
rect 15285 8938 15351 8941
rect 15285 8936 16268 8938
rect 15285 8880 15290 8936
rect 15346 8880 16268 8936
rect 15285 8878 16268 8880
rect 15285 8875 15351 8878
rect 8772 8800 8864 8802
rect 8814 8744 8864 8800
rect 8772 8742 8864 8744
rect 10366 8742 13554 8802
rect 8772 8740 8819 8742
rect 8753 8739 8819 8740
rect 3909 8736 4229 8737
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 8671 4229 8672
rect 9840 8736 10160 8737
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 8671 10160 8672
rect 15770 8736 16090 8737
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 15770 8671 16090 8672
rect 9121 8666 9187 8669
rect 4294 8664 9187 8666
rect 4294 8608 9126 8664
rect 9182 8608 9187 8664
rect 4294 8606 9187 8608
rect 3601 8530 3667 8533
rect 4294 8530 4354 8606
rect 9121 8603 9187 8606
rect 9254 8604 9260 8668
rect 9324 8666 9330 8668
rect 9397 8666 9463 8669
rect 9324 8664 9463 8666
rect 9324 8608 9402 8664
rect 9458 8608 9463 8664
rect 9324 8606 9463 8608
rect 9324 8604 9330 8606
rect 9397 8603 9463 8606
rect 11053 8666 11119 8669
rect 15009 8666 15075 8669
rect 11053 8664 15075 8666
rect 11053 8608 11058 8664
rect 11114 8608 15014 8664
rect 15070 8608 15075 8664
rect 11053 8606 15075 8608
rect 16208 8666 16268 8878
rect 16614 8740 16620 8804
rect 16684 8802 16690 8804
rect 16757 8802 16823 8805
rect 16684 8800 16823 8802
rect 16684 8744 16762 8800
rect 16818 8744 16823 8800
rect 16684 8742 16823 8744
rect 16684 8740 16690 8742
rect 16757 8739 16823 8742
rect 19520 8666 20000 8696
rect 16208 8606 20000 8666
rect 11053 8603 11119 8606
rect 15009 8603 15075 8606
rect 19520 8576 20000 8606
rect 3601 8528 4354 8530
rect 3601 8472 3606 8528
rect 3662 8472 4354 8528
rect 3601 8470 4354 8472
rect 6361 8530 6427 8533
rect 15326 8530 15332 8532
rect 6361 8528 15332 8530
rect 6361 8472 6366 8528
rect 6422 8472 15332 8528
rect 6361 8470 15332 8472
rect 3601 8467 3667 8470
rect 6361 8467 6427 8470
rect 15326 8468 15332 8470
rect 15396 8530 15402 8532
rect 16849 8530 16915 8533
rect 15396 8528 16915 8530
rect 15396 8472 16854 8528
rect 16910 8472 16915 8528
rect 15396 8470 16915 8472
rect 15396 8468 15402 8470
rect 16849 8467 16915 8470
rect 0 8394 480 8424
rect 3141 8394 3207 8397
rect 0 8392 3207 8394
rect 0 8336 3146 8392
rect 3202 8336 3207 8392
rect 0 8334 3207 8336
rect 0 8304 480 8334
rect 3141 8331 3207 8334
rect 3417 8394 3483 8397
rect 12801 8394 12867 8397
rect 16614 8394 16620 8396
rect 3417 8392 16620 8394
rect 3417 8336 3422 8392
rect 3478 8336 12806 8392
rect 12862 8336 16620 8392
rect 3417 8334 16620 8336
rect 3417 8331 3483 8334
rect 12801 8331 12867 8334
rect 16614 8332 16620 8334
rect 16684 8332 16690 8396
rect 2865 8258 2931 8261
rect 2998 8258 3004 8260
rect 2865 8256 3004 8258
rect 2865 8200 2870 8256
rect 2926 8200 3004 8256
rect 2865 8198 3004 8200
rect 2865 8195 2931 8198
rect 2998 8196 3004 8198
rect 3068 8196 3074 8260
rect 7557 8258 7623 8261
rect 12382 8258 12388 8260
rect 7557 8256 12388 8258
rect 7557 8200 7562 8256
rect 7618 8200 12388 8256
rect 7557 8198 12388 8200
rect 7557 8195 7623 8198
rect 12382 8196 12388 8198
rect 12452 8196 12458 8260
rect 15745 8258 15811 8261
rect 19520 8258 20000 8288
rect 13494 8198 15164 8258
rect 6874 8192 7194 8193
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7194 8192
rect 6874 8127 7194 8128
rect 12805 8192 13125 8193
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 12805 8127 13125 8128
rect 7925 8122 7991 8125
rect 9489 8122 9555 8125
rect 7925 8120 9555 8122
rect 7925 8064 7930 8120
rect 7986 8064 9494 8120
rect 9550 8064 9555 8120
rect 7925 8062 9555 8064
rect 7925 8059 7991 8062
rect 9489 8059 9555 8062
rect 9949 8122 10015 8125
rect 10869 8122 10935 8125
rect 9949 8120 10935 8122
rect 9949 8064 9954 8120
rect 10010 8064 10874 8120
rect 10930 8064 10935 8120
rect 9949 8062 10935 8064
rect 9949 8059 10015 8062
rect 10869 8059 10935 8062
rect 0 7986 480 8016
rect 1761 7986 1827 7989
rect 0 7984 1827 7986
rect 0 7928 1766 7984
rect 1822 7928 1827 7984
rect 0 7926 1827 7928
rect 0 7896 480 7926
rect 1761 7923 1827 7926
rect 5441 7986 5507 7989
rect 9305 7986 9371 7989
rect 5441 7984 9371 7986
rect 5441 7928 5446 7984
rect 5502 7928 9310 7984
rect 9366 7928 9371 7984
rect 5441 7926 9371 7928
rect 5441 7923 5507 7926
rect 9305 7923 9371 7926
rect 4705 7850 4771 7853
rect 5165 7850 5231 7853
rect 7741 7850 7807 7853
rect 13494 7850 13554 8198
rect 14733 8122 14799 8125
rect 15104 8122 15164 8198
rect 15745 8256 20000 8258
rect 15745 8200 15750 8256
rect 15806 8200 20000 8256
rect 15745 8198 20000 8200
rect 15745 8195 15811 8198
rect 19520 8168 20000 8198
rect 16021 8122 16087 8125
rect 16246 8122 16252 8124
rect 14733 8120 15026 8122
rect 14733 8064 14738 8120
rect 14794 8064 15026 8120
rect 14733 8062 15026 8064
rect 15104 8120 16252 8122
rect 15104 8064 16026 8120
rect 16082 8064 16252 8120
rect 15104 8062 16252 8064
rect 14733 8059 14799 8062
rect 14966 7989 15026 8062
rect 16021 8059 16087 8062
rect 16246 8060 16252 8062
rect 16316 8060 16322 8124
rect 13629 7986 13695 7989
rect 13629 7984 13738 7986
rect 13629 7928 13634 7984
rect 13690 7928 13738 7984
rect 13629 7923 13738 7928
rect 14966 7984 15075 7989
rect 15510 7986 15516 7988
rect 14966 7928 15014 7984
rect 15070 7928 15075 7984
rect 14966 7926 15075 7928
rect 15009 7923 15075 7926
rect 15150 7926 15516 7986
rect 4705 7848 7666 7850
rect 4705 7792 4710 7848
rect 4766 7792 5170 7848
rect 5226 7792 7666 7848
rect 4705 7790 7666 7792
rect 4705 7787 4771 7790
rect 5165 7787 5231 7790
rect 7606 7714 7666 7790
rect 7741 7848 13554 7850
rect 7741 7792 7746 7848
rect 7802 7792 13554 7848
rect 7741 7790 13554 7792
rect 13678 7850 13738 7923
rect 15150 7850 15210 7926
rect 15510 7924 15516 7926
rect 15580 7924 15586 7988
rect 13678 7790 15210 7850
rect 15285 7850 15351 7853
rect 19520 7850 20000 7880
rect 15285 7848 20000 7850
rect 15285 7792 15290 7848
rect 15346 7792 20000 7848
rect 15285 7790 20000 7792
rect 7741 7787 7807 7790
rect 9254 7714 9260 7716
rect 7606 7654 9260 7714
rect 9254 7652 9260 7654
rect 9324 7652 9330 7716
rect 3909 7648 4229 7649
rect 0 7578 480 7608
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 7583 4229 7584
rect 9840 7648 10160 7649
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 7583 10160 7584
rect 2129 7578 2195 7581
rect 8201 7580 8267 7581
rect 8150 7578 8156 7580
rect 0 7576 2195 7578
rect 0 7520 2134 7576
rect 2190 7520 2195 7576
rect 0 7518 2195 7520
rect 8110 7518 8156 7578
rect 8220 7576 8267 7580
rect 8262 7520 8267 7576
rect 0 7488 480 7518
rect 2129 7515 2195 7518
rect 8150 7516 8156 7518
rect 8220 7516 8267 7520
rect 8201 7515 8267 7516
rect 8661 7442 8727 7445
rect 10685 7442 10751 7445
rect 8661 7440 10751 7442
rect 8661 7384 8666 7440
rect 8722 7384 10690 7440
rect 10746 7384 10751 7440
rect 8661 7382 10751 7384
rect 8661 7379 8727 7382
rect 10685 7379 10751 7382
rect 1761 7306 1827 7309
rect 6361 7306 6427 7309
rect 1761 7304 6427 7306
rect 1761 7248 1766 7304
rect 1822 7248 6366 7304
rect 6422 7248 6427 7304
rect 1761 7246 6427 7248
rect 1761 7243 1827 7246
rect 6361 7243 6427 7246
rect 9254 7244 9260 7308
rect 9324 7306 9330 7308
rect 11237 7306 11303 7309
rect 9324 7304 11303 7306
rect 9324 7248 11242 7304
rect 11298 7248 11303 7304
rect 9324 7246 11303 7248
rect 9324 7244 9330 7246
rect 11237 7243 11303 7246
rect 11881 7306 11947 7309
rect 13678 7306 13738 7790
rect 15285 7787 15351 7790
rect 19520 7760 20000 7790
rect 14958 7652 14964 7716
rect 15028 7714 15034 7716
rect 15510 7714 15516 7716
rect 15028 7654 15516 7714
rect 15028 7652 15034 7654
rect 15510 7652 15516 7654
rect 15580 7652 15586 7716
rect 15770 7648 16090 7649
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 7583 16090 7584
rect 18045 7442 18111 7445
rect 19520 7442 20000 7472
rect 18045 7440 20000 7442
rect 18045 7384 18050 7440
rect 18106 7384 20000 7440
rect 18045 7382 20000 7384
rect 18045 7379 18111 7382
rect 19520 7352 20000 7382
rect 11881 7304 13738 7306
rect 11881 7248 11886 7304
rect 11942 7248 13738 7304
rect 11881 7246 13738 7248
rect 11881 7243 11947 7246
rect 0 7170 480 7200
rect 2773 7170 2839 7173
rect 0 7168 2839 7170
rect 0 7112 2778 7168
rect 2834 7112 2839 7168
rect 0 7110 2839 7112
rect 0 7080 480 7110
rect 2773 7107 2839 7110
rect 7966 7108 7972 7172
rect 8036 7170 8042 7172
rect 10133 7170 10199 7173
rect 12341 7170 12407 7173
rect 8036 7168 12407 7170
rect 8036 7112 10138 7168
rect 10194 7112 12346 7168
rect 12402 7112 12407 7168
rect 8036 7110 12407 7112
rect 8036 7108 8042 7110
rect 10133 7107 10199 7110
rect 12341 7107 12407 7110
rect 13629 7170 13695 7173
rect 13854 7170 13860 7172
rect 13629 7168 13860 7170
rect 13629 7112 13634 7168
rect 13690 7112 13860 7168
rect 13629 7110 13860 7112
rect 13629 7107 13695 7110
rect 13854 7108 13860 7110
rect 13924 7108 13930 7172
rect 6874 7104 7194 7105
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7194 7104
rect 6874 7039 7194 7040
rect 12805 7104 13125 7105
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 7039 13125 7040
rect 2497 7034 2563 7037
rect 3785 7034 3851 7037
rect 2497 7032 3851 7034
rect 2497 6976 2502 7032
rect 2558 6976 3790 7032
rect 3846 6976 3851 7032
rect 2497 6974 3851 6976
rect 2497 6971 2563 6974
rect 3785 6971 3851 6974
rect 9121 7032 9187 7037
rect 9121 6976 9126 7032
rect 9182 6976 9187 7032
rect 9121 6971 9187 6976
rect 17493 7034 17559 7037
rect 19520 7034 20000 7064
rect 17493 7032 20000 7034
rect 17493 6976 17498 7032
rect 17554 6976 20000 7032
rect 17493 6974 20000 6976
rect 17493 6971 17559 6974
rect 3049 6898 3115 6901
rect 9124 6898 9184 6971
rect 19520 6944 20000 6974
rect 14733 6898 14799 6901
rect 15469 6898 15535 6901
rect 3049 6896 4032 6898
rect 3049 6840 3054 6896
rect 3110 6840 4032 6896
rect 3049 6838 4032 6840
rect 9124 6896 14799 6898
rect 9124 6840 14738 6896
rect 14794 6840 14799 6896
rect 9124 6838 14799 6840
rect 3049 6835 3115 6838
rect 0 6762 480 6792
rect 3601 6762 3667 6765
rect 0 6760 3667 6762
rect 0 6704 3606 6760
rect 3662 6704 3667 6760
rect 0 6702 3667 6704
rect 3972 6762 4032 6838
rect 14733 6835 14799 6838
rect 15288 6896 15535 6898
rect 15288 6840 15474 6896
rect 15530 6840 15535 6896
rect 15288 6838 15535 6840
rect 13169 6762 13235 6765
rect 3972 6760 13235 6762
rect 3972 6704 13174 6760
rect 13230 6704 13235 6760
rect 3972 6702 13235 6704
rect 0 6672 480 6702
rect 3601 6699 3667 6702
rect 13169 6699 13235 6702
rect 13813 6762 13879 6765
rect 13997 6762 14063 6765
rect 13813 6760 14063 6762
rect 13813 6704 13818 6760
rect 13874 6704 14002 6760
rect 14058 6704 14063 6760
rect 13813 6702 14063 6704
rect 13813 6699 13879 6702
rect 13997 6699 14063 6702
rect 3909 6560 4229 6561
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 6495 4229 6496
rect 9840 6560 10160 6561
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 6495 10160 6496
rect 0 6354 480 6384
rect 15288 6357 15348 6838
rect 15469 6835 15535 6838
rect 15770 6560 16090 6561
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 15770 6495 16090 6496
rect 18505 6490 18571 6493
rect 19520 6490 20000 6520
rect 18505 6488 20000 6490
rect 18505 6432 18510 6488
rect 18566 6432 20000 6488
rect 18505 6430 20000 6432
rect 18505 6427 18571 6430
rect 19520 6400 20000 6430
rect 1853 6354 1919 6357
rect 0 6352 1919 6354
rect 0 6296 1858 6352
rect 1914 6296 1919 6352
rect 0 6294 1919 6296
rect 0 6264 480 6294
rect 1853 6291 1919 6294
rect 3601 6354 3667 6357
rect 8017 6354 8083 6357
rect 3601 6352 8083 6354
rect 3601 6296 3606 6352
rect 3662 6296 8022 6352
rect 8078 6296 8083 6352
rect 3601 6294 8083 6296
rect 3601 6291 3667 6294
rect 8017 6291 8083 6294
rect 15285 6352 15351 6357
rect 15285 6296 15290 6352
rect 15346 6296 15351 6352
rect 15285 6291 15351 6296
rect 18045 6082 18111 6085
rect 19520 6082 20000 6112
rect 18045 6080 20000 6082
rect 18045 6024 18050 6080
rect 18106 6024 20000 6080
rect 18045 6022 20000 6024
rect 18045 6019 18111 6022
rect 6874 6016 7194 6017
rect 0 5946 480 5976
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7194 6016
rect 6874 5951 7194 5952
rect 12805 6016 13125 6017
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 19520 5992 20000 6022
rect 12805 5951 13125 5952
rect 1853 5946 1919 5949
rect 0 5944 1919 5946
rect 0 5888 1858 5944
rect 1914 5888 1919 5944
rect 0 5886 1919 5888
rect 0 5856 480 5886
rect 1853 5883 1919 5886
rect 12014 5612 12020 5676
rect 12084 5674 12090 5676
rect 12709 5674 12775 5677
rect 12084 5672 12775 5674
rect 12084 5616 12714 5672
rect 12770 5616 12775 5672
rect 12084 5614 12775 5616
rect 12084 5612 12090 5614
rect 12709 5611 12775 5614
rect 13169 5674 13235 5677
rect 13302 5674 13308 5676
rect 13169 5672 13308 5674
rect 13169 5616 13174 5672
rect 13230 5616 13308 5672
rect 13169 5614 13308 5616
rect 13169 5611 13235 5614
rect 13302 5612 13308 5614
rect 13372 5612 13378 5676
rect 17401 5674 17467 5677
rect 19520 5674 20000 5704
rect 17401 5672 20000 5674
rect 17401 5616 17406 5672
rect 17462 5616 20000 5672
rect 17401 5614 20000 5616
rect 17401 5611 17467 5614
rect 19520 5584 20000 5614
rect 0 5538 480 5568
rect 1761 5538 1827 5541
rect 0 5536 1827 5538
rect 0 5480 1766 5536
rect 1822 5480 1827 5536
rect 0 5478 1827 5480
rect 0 5448 480 5478
rect 1761 5475 1827 5478
rect 3909 5472 4229 5473
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 5407 4229 5408
rect 9840 5472 10160 5473
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 5407 10160 5408
rect 15770 5472 16090 5473
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 15770 5407 16090 5408
rect 2497 5266 2563 5269
rect 15285 5266 15351 5269
rect 19520 5266 20000 5296
rect 2497 5264 15026 5266
rect 2497 5208 2502 5264
rect 2558 5208 15026 5264
rect 2497 5206 15026 5208
rect 2497 5203 2563 5206
rect 0 5130 480 5160
rect 2773 5130 2839 5133
rect 0 5128 2839 5130
rect 0 5072 2778 5128
rect 2834 5072 2839 5128
rect 0 5070 2839 5072
rect 0 5040 480 5070
rect 2773 5067 2839 5070
rect 12566 5068 12572 5132
rect 12636 5130 12642 5132
rect 13353 5130 13419 5133
rect 12636 5128 13419 5130
rect 12636 5072 13358 5128
rect 13414 5072 13419 5128
rect 12636 5070 13419 5072
rect 12636 5068 12642 5070
rect 13353 5067 13419 5070
rect 9489 4994 9555 4997
rect 11697 4994 11763 4997
rect 9489 4992 11763 4994
rect 9489 4936 9494 4992
rect 9550 4936 11702 4992
rect 11758 4936 11763 4992
rect 9489 4934 11763 4936
rect 14966 4994 15026 5206
rect 15285 5264 20000 5266
rect 15285 5208 15290 5264
rect 15346 5208 20000 5264
rect 15285 5206 20000 5208
rect 15285 5203 15351 5206
rect 19520 5176 20000 5206
rect 15510 5068 15516 5132
rect 15580 5130 15586 5132
rect 16021 5130 16087 5133
rect 15580 5128 16087 5130
rect 15580 5072 16026 5128
rect 16082 5072 16087 5128
rect 15580 5070 16087 5072
rect 15580 5068 15586 5070
rect 16021 5067 16087 5070
rect 16389 4994 16455 4997
rect 14966 4992 16455 4994
rect 14966 4936 16394 4992
rect 16450 4936 16455 4992
rect 14966 4934 16455 4936
rect 9489 4931 9555 4934
rect 11697 4931 11763 4934
rect 16389 4931 16455 4934
rect 6874 4928 7194 4929
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7194 4928
rect 6874 4863 7194 4864
rect 12805 4928 13125 4929
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 4863 13125 4864
rect 15653 4858 15719 4861
rect 19520 4858 20000 4888
rect 15653 4856 20000 4858
rect 15653 4800 15658 4856
rect 15714 4800 20000 4856
rect 15653 4798 20000 4800
rect 15653 4795 15719 4798
rect 19520 4768 20000 4798
rect 0 4722 480 4752
rect 1853 4722 1919 4725
rect 0 4720 1919 4722
rect 0 4664 1858 4720
rect 1914 4664 1919 4720
rect 0 4662 1919 4664
rect 0 4632 480 4662
rect 1853 4659 1919 4662
rect 6913 4722 6979 4725
rect 7465 4722 7531 4725
rect 15510 4722 15516 4724
rect 6913 4720 15516 4722
rect 6913 4664 6918 4720
rect 6974 4664 7470 4720
rect 7526 4664 15516 4720
rect 6913 4662 15516 4664
rect 6913 4659 6979 4662
rect 7465 4659 7531 4662
rect 15510 4660 15516 4662
rect 15580 4660 15586 4724
rect 6453 4586 6519 4589
rect 8201 4586 8267 4589
rect 6453 4584 8267 4586
rect 6453 4528 6458 4584
rect 6514 4528 8206 4584
rect 8262 4528 8267 4584
rect 6453 4526 8267 4528
rect 6453 4523 6519 4526
rect 8201 4523 8267 4526
rect 17401 4450 17467 4453
rect 19520 4450 20000 4480
rect 17401 4448 20000 4450
rect 17401 4392 17406 4448
rect 17462 4392 20000 4448
rect 17401 4390 20000 4392
rect 17401 4387 17467 4390
rect 3909 4384 4229 4385
rect 0 4314 480 4344
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 4319 4229 4320
rect 9840 4384 10160 4385
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 4319 10160 4320
rect 15770 4384 16090 4385
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 19520 4360 20000 4390
rect 15770 4319 16090 4320
rect 2773 4314 2839 4317
rect 0 4312 2839 4314
rect 0 4256 2778 4312
rect 2834 4256 2839 4312
rect 0 4254 2839 4256
rect 0 4224 480 4254
rect 2773 4251 2839 4254
rect 14774 3980 14780 4044
rect 14844 4042 14850 4044
rect 14917 4042 14983 4045
rect 14844 4040 14983 4042
rect 14844 3984 14922 4040
rect 14978 3984 14983 4040
rect 14844 3982 14983 3984
rect 14844 3980 14850 3982
rect 14917 3979 14983 3982
rect 16205 4042 16271 4045
rect 16798 4042 16804 4044
rect 16205 4040 16804 4042
rect 16205 3984 16210 4040
rect 16266 3984 16804 4040
rect 16205 3982 16804 3984
rect 16205 3979 16271 3982
rect 16798 3980 16804 3982
rect 16868 3980 16874 4044
rect 17677 4042 17743 4045
rect 19520 4042 20000 4072
rect 17677 4040 20000 4042
rect 17677 3984 17682 4040
rect 17738 3984 20000 4040
rect 17677 3982 20000 3984
rect 17677 3979 17743 3982
rect 19520 3952 20000 3982
rect 0 3906 480 3936
rect 3325 3906 3391 3909
rect 0 3904 3391 3906
rect 0 3848 3330 3904
rect 3386 3848 3391 3904
rect 0 3846 3391 3848
rect 0 3816 480 3846
rect 3325 3843 3391 3846
rect 13537 3906 13603 3909
rect 16430 3906 16436 3908
rect 13537 3904 16436 3906
rect 13537 3848 13542 3904
rect 13598 3848 16436 3904
rect 13537 3846 16436 3848
rect 13537 3843 13603 3846
rect 16430 3844 16436 3846
rect 16500 3844 16506 3908
rect 6874 3840 7194 3841
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7194 3840
rect 6874 3775 7194 3776
rect 12805 3840 13125 3841
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 3775 13125 3776
rect 14457 3636 14523 3637
rect 14406 3572 14412 3636
rect 14476 3634 14523 3636
rect 16941 3634 17007 3637
rect 19520 3634 20000 3664
rect 14476 3632 14568 3634
rect 14518 3576 14568 3632
rect 14476 3574 14568 3576
rect 16941 3632 20000 3634
rect 16941 3576 16946 3632
rect 17002 3576 20000 3632
rect 16941 3574 20000 3576
rect 14476 3572 14523 3574
rect 14457 3571 14523 3572
rect 16941 3571 17007 3574
rect 19520 3544 20000 3574
rect 0 3498 480 3528
rect 3049 3498 3115 3501
rect 0 3496 3115 3498
rect 0 3440 3054 3496
rect 3110 3440 3115 3496
rect 0 3438 3115 3440
rect 0 3408 480 3438
rect 3049 3435 3115 3438
rect 3909 3296 4229 3297
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 3231 4229 3232
rect 9840 3296 10160 3297
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 3231 10160 3232
rect 15770 3296 16090 3297
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15770 3231 16090 3232
rect 0 3090 480 3120
rect 2957 3090 3023 3093
rect 0 3088 3023 3090
rect 0 3032 2962 3088
rect 3018 3032 3023 3088
rect 0 3030 3023 3032
rect 0 3000 480 3030
rect 2957 3027 3023 3030
rect 16205 3090 16271 3093
rect 19520 3090 20000 3120
rect 16205 3088 20000 3090
rect 16205 3032 16210 3088
rect 16266 3032 20000 3088
rect 16205 3030 20000 3032
rect 16205 3027 16271 3030
rect 19520 3000 20000 3030
rect 10317 2956 10383 2957
rect 10317 2954 10364 2956
rect 10272 2952 10364 2954
rect 10272 2896 10322 2952
rect 10272 2894 10364 2896
rect 10317 2892 10364 2894
rect 10428 2892 10434 2956
rect 10777 2954 10843 2957
rect 15142 2954 15148 2956
rect 10777 2952 15148 2954
rect 10777 2896 10782 2952
rect 10838 2896 15148 2952
rect 10777 2894 15148 2896
rect 10317 2891 10383 2892
rect 10777 2891 10843 2894
rect 15142 2892 15148 2894
rect 15212 2954 15218 2956
rect 15745 2954 15811 2957
rect 15212 2952 15811 2954
rect 15212 2896 15750 2952
rect 15806 2896 15811 2952
rect 15212 2894 15811 2896
rect 15212 2892 15218 2894
rect 15745 2891 15811 2894
rect 8569 2818 8635 2821
rect 11053 2818 11119 2821
rect 8569 2816 11119 2818
rect 8569 2760 8574 2816
rect 8630 2760 11058 2816
rect 11114 2760 11119 2816
rect 8569 2758 11119 2760
rect 8569 2755 8635 2758
rect 11053 2755 11119 2758
rect 6874 2752 7194 2753
rect 0 2682 480 2712
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7194 2752
rect 6874 2687 7194 2688
rect 12805 2752 13125 2753
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 12805 2687 13125 2688
rect 3417 2682 3483 2685
rect 0 2680 3483 2682
rect 0 2624 3422 2680
rect 3478 2624 3483 2680
rect 0 2622 3483 2624
rect 0 2592 480 2622
rect 3417 2619 3483 2622
rect 15326 2620 15332 2684
rect 15396 2682 15402 2684
rect 16021 2682 16087 2685
rect 15396 2680 16087 2682
rect 15396 2624 16026 2680
rect 16082 2624 16087 2680
rect 15396 2622 16087 2624
rect 15396 2620 15402 2622
rect 16021 2619 16087 2622
rect 16614 2620 16620 2684
rect 16684 2682 16690 2684
rect 17493 2682 17559 2685
rect 19520 2682 20000 2712
rect 16684 2680 17559 2682
rect 16684 2624 17498 2680
rect 17554 2624 17559 2680
rect 16684 2622 17559 2624
rect 16684 2620 16690 2622
rect 17493 2619 17559 2622
rect 17726 2622 20000 2682
rect 8293 2546 8359 2549
rect 10501 2546 10567 2549
rect 11789 2548 11855 2549
rect 11789 2546 11836 2548
rect 8293 2544 10567 2546
rect 8293 2488 8298 2544
rect 8354 2488 10506 2544
rect 10562 2488 10567 2544
rect 8293 2486 10567 2488
rect 11744 2544 11836 2546
rect 11744 2488 11794 2544
rect 11744 2486 11836 2488
rect 8293 2483 8359 2486
rect 10501 2483 10567 2486
rect 11789 2484 11836 2486
rect 11900 2484 11906 2548
rect 15561 2546 15627 2549
rect 17726 2546 17786 2622
rect 19520 2592 20000 2622
rect 15561 2544 17786 2546
rect 15561 2488 15566 2544
rect 15622 2488 17786 2544
rect 15561 2486 17786 2488
rect 11789 2483 11855 2484
rect 15561 2483 15627 2486
rect 0 2274 480 2304
rect 1853 2274 1919 2277
rect 0 2272 1919 2274
rect 0 2216 1858 2272
rect 1914 2216 1919 2272
rect 0 2214 1919 2216
rect 0 2184 480 2214
rect 1853 2211 1919 2214
rect 16205 2274 16271 2277
rect 19520 2274 20000 2304
rect 16205 2272 20000 2274
rect 16205 2216 16210 2272
rect 16266 2216 20000 2272
rect 16205 2214 20000 2216
rect 16205 2211 16271 2214
rect 3909 2208 4229 2209
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2143 4229 2144
rect 9840 2208 10160 2209
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2143 10160 2144
rect 15770 2208 16090 2209
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 19520 2184 20000 2214
rect 15770 2143 16090 2144
rect 0 1866 480 1896
rect 3325 1866 3391 1869
rect 0 1864 3391 1866
rect 0 1808 3330 1864
rect 3386 1808 3391 1864
rect 0 1806 3391 1808
rect 0 1776 480 1806
rect 3325 1803 3391 1806
rect 14733 1866 14799 1869
rect 19520 1866 20000 1896
rect 14733 1864 20000 1866
rect 14733 1808 14738 1864
rect 14794 1808 20000 1864
rect 14733 1806 20000 1808
rect 14733 1803 14799 1806
rect 19520 1776 20000 1806
rect 0 1458 480 1488
rect 3509 1458 3575 1461
rect 0 1456 3575 1458
rect 0 1400 3514 1456
rect 3570 1400 3575 1456
rect 0 1398 3575 1400
rect 0 1368 480 1398
rect 3509 1395 3575 1398
rect 18873 1458 18939 1461
rect 19520 1458 20000 1488
rect 18873 1456 20000 1458
rect 18873 1400 18878 1456
rect 18934 1400 20000 1456
rect 18873 1398 20000 1400
rect 18873 1395 18939 1398
rect 19520 1368 20000 1398
rect 0 1050 480 1080
rect 3693 1050 3759 1053
rect 0 1048 3759 1050
rect 0 992 3698 1048
rect 3754 992 3759 1048
rect 0 990 3759 992
rect 0 960 480 990
rect 3693 987 3759 990
rect 15009 1050 15075 1053
rect 19520 1050 20000 1080
rect 15009 1048 20000 1050
rect 15009 992 15014 1048
rect 15070 992 20000 1048
rect 15009 990 20000 992
rect 15009 987 15075 990
rect 19520 960 20000 990
rect 0 642 480 672
rect 3693 642 3759 645
rect 0 640 3759 642
rect 0 584 3698 640
rect 3754 584 3759 640
rect 0 582 3759 584
rect 0 552 480 582
rect 3693 579 3759 582
rect 18413 642 18479 645
rect 19520 642 20000 672
rect 18413 640 20000 642
rect 18413 584 18418 640
rect 18474 584 20000 640
rect 18413 582 20000 584
rect 18413 579 18479 582
rect 19520 552 20000 582
rect 0 234 480 264
rect 3233 234 3299 237
rect 0 232 3299 234
rect 0 176 3238 232
rect 3294 176 3299 232
rect 0 174 3299 176
rect 0 144 480 174
rect 3233 171 3299 174
rect 13997 234 14063 237
rect 19520 234 20000 264
rect 13997 232 20000 234
rect 13997 176 14002 232
rect 14058 176 20000 232
rect 13997 174 20000 176
rect 13997 171 14063 174
rect 19520 144 20000 174
<< via3 >>
rect 16252 15404 16316 15468
rect 6882 14716 6946 14720
rect 6882 14660 6886 14716
rect 6886 14660 6942 14716
rect 6942 14660 6946 14716
rect 6882 14656 6946 14660
rect 6962 14716 7026 14720
rect 6962 14660 6966 14716
rect 6966 14660 7022 14716
rect 7022 14660 7026 14716
rect 6962 14656 7026 14660
rect 7042 14716 7106 14720
rect 7042 14660 7046 14716
rect 7046 14660 7102 14716
rect 7102 14660 7106 14716
rect 7042 14656 7106 14660
rect 7122 14716 7186 14720
rect 7122 14660 7126 14716
rect 7126 14660 7182 14716
rect 7182 14660 7186 14716
rect 7122 14656 7186 14660
rect 12813 14716 12877 14720
rect 12813 14660 12817 14716
rect 12817 14660 12873 14716
rect 12873 14660 12877 14716
rect 12813 14656 12877 14660
rect 12893 14716 12957 14720
rect 12893 14660 12897 14716
rect 12897 14660 12953 14716
rect 12953 14660 12957 14716
rect 12893 14656 12957 14660
rect 12973 14716 13037 14720
rect 12973 14660 12977 14716
rect 12977 14660 13033 14716
rect 13033 14660 13037 14716
rect 12973 14656 13037 14660
rect 13053 14716 13117 14720
rect 13053 14660 13057 14716
rect 13057 14660 13113 14716
rect 13113 14660 13117 14716
rect 13053 14656 13117 14660
rect 3917 14172 3981 14176
rect 3917 14116 3921 14172
rect 3921 14116 3977 14172
rect 3977 14116 3981 14172
rect 3917 14112 3981 14116
rect 3997 14172 4061 14176
rect 3997 14116 4001 14172
rect 4001 14116 4057 14172
rect 4057 14116 4061 14172
rect 3997 14112 4061 14116
rect 4077 14172 4141 14176
rect 4077 14116 4081 14172
rect 4081 14116 4137 14172
rect 4137 14116 4141 14172
rect 4077 14112 4141 14116
rect 4157 14172 4221 14176
rect 4157 14116 4161 14172
rect 4161 14116 4217 14172
rect 4217 14116 4221 14172
rect 4157 14112 4221 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 15778 14172 15842 14176
rect 15778 14116 15782 14172
rect 15782 14116 15838 14172
rect 15838 14116 15842 14172
rect 15778 14112 15842 14116
rect 15858 14172 15922 14176
rect 15858 14116 15862 14172
rect 15862 14116 15918 14172
rect 15918 14116 15922 14172
rect 15858 14112 15922 14116
rect 15938 14172 16002 14176
rect 15938 14116 15942 14172
rect 15942 14116 15998 14172
rect 15998 14116 16002 14172
rect 15938 14112 16002 14116
rect 16018 14172 16082 14176
rect 16018 14116 16022 14172
rect 16022 14116 16078 14172
rect 16078 14116 16082 14172
rect 16018 14112 16082 14116
rect 6882 13628 6946 13632
rect 6882 13572 6886 13628
rect 6886 13572 6942 13628
rect 6942 13572 6946 13628
rect 6882 13568 6946 13572
rect 6962 13628 7026 13632
rect 6962 13572 6966 13628
rect 6966 13572 7022 13628
rect 7022 13572 7026 13628
rect 6962 13568 7026 13572
rect 7042 13628 7106 13632
rect 7042 13572 7046 13628
rect 7046 13572 7102 13628
rect 7102 13572 7106 13628
rect 7042 13568 7106 13572
rect 7122 13628 7186 13632
rect 7122 13572 7126 13628
rect 7126 13572 7182 13628
rect 7182 13572 7186 13628
rect 7122 13568 7186 13572
rect 12813 13628 12877 13632
rect 12813 13572 12817 13628
rect 12817 13572 12873 13628
rect 12873 13572 12877 13628
rect 12813 13568 12877 13572
rect 12893 13628 12957 13632
rect 12893 13572 12897 13628
rect 12897 13572 12953 13628
rect 12953 13572 12957 13628
rect 12893 13568 12957 13572
rect 12973 13628 13037 13632
rect 12973 13572 12977 13628
rect 12977 13572 13033 13628
rect 13033 13572 13037 13628
rect 12973 13568 13037 13572
rect 13053 13628 13117 13632
rect 13053 13572 13057 13628
rect 13057 13572 13113 13628
rect 13113 13572 13117 13628
rect 13053 13568 13117 13572
rect 14780 13364 14844 13428
rect 15148 13424 15212 13428
rect 15148 13368 15162 13424
rect 15162 13368 15212 13424
rect 15148 13364 15212 13368
rect 13308 13092 13372 13156
rect 3917 13084 3981 13088
rect 3917 13028 3921 13084
rect 3921 13028 3977 13084
rect 3977 13028 3981 13084
rect 3917 13024 3981 13028
rect 3997 13084 4061 13088
rect 3997 13028 4001 13084
rect 4001 13028 4057 13084
rect 4057 13028 4061 13084
rect 3997 13024 4061 13028
rect 4077 13084 4141 13088
rect 4077 13028 4081 13084
rect 4081 13028 4137 13084
rect 4137 13028 4141 13084
rect 4077 13024 4141 13028
rect 4157 13084 4221 13088
rect 4157 13028 4161 13084
rect 4161 13028 4217 13084
rect 4217 13028 4221 13084
rect 4157 13024 4221 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 15778 13084 15842 13088
rect 15778 13028 15782 13084
rect 15782 13028 15838 13084
rect 15838 13028 15842 13084
rect 15778 13024 15842 13028
rect 15858 13084 15922 13088
rect 15858 13028 15862 13084
rect 15862 13028 15918 13084
rect 15918 13028 15922 13084
rect 15858 13024 15922 13028
rect 15938 13084 16002 13088
rect 15938 13028 15942 13084
rect 15942 13028 15998 13084
rect 15998 13028 16002 13084
rect 15938 13024 16002 13028
rect 16018 13084 16082 13088
rect 16018 13028 16022 13084
rect 16022 13028 16078 13084
rect 16078 13028 16082 13084
rect 16018 13024 16082 13028
rect 14964 12820 15028 12884
rect 13860 12684 13924 12748
rect 16436 12548 16500 12612
rect 6882 12540 6946 12544
rect 6882 12484 6886 12540
rect 6886 12484 6942 12540
rect 6942 12484 6946 12540
rect 6882 12480 6946 12484
rect 6962 12540 7026 12544
rect 6962 12484 6966 12540
rect 6966 12484 7022 12540
rect 7022 12484 7026 12540
rect 6962 12480 7026 12484
rect 7042 12540 7106 12544
rect 7042 12484 7046 12540
rect 7046 12484 7102 12540
rect 7102 12484 7106 12540
rect 7042 12480 7106 12484
rect 7122 12540 7186 12544
rect 7122 12484 7126 12540
rect 7126 12484 7182 12540
rect 7182 12484 7186 12540
rect 7122 12480 7186 12484
rect 12813 12540 12877 12544
rect 12813 12484 12817 12540
rect 12817 12484 12873 12540
rect 12873 12484 12877 12540
rect 12813 12480 12877 12484
rect 12893 12540 12957 12544
rect 12893 12484 12897 12540
rect 12897 12484 12953 12540
rect 12953 12484 12957 12540
rect 12893 12480 12957 12484
rect 12973 12540 13037 12544
rect 12973 12484 12977 12540
rect 12977 12484 13033 12540
rect 13033 12484 13037 12540
rect 12973 12480 13037 12484
rect 13053 12540 13117 12544
rect 13053 12484 13057 12540
rect 13057 12484 13113 12540
rect 13113 12484 13117 12540
rect 13053 12480 13117 12484
rect 10364 12412 10428 12476
rect 15516 12412 15580 12476
rect 3004 12276 3068 12340
rect 3917 11996 3981 12000
rect 3917 11940 3921 11996
rect 3921 11940 3977 11996
rect 3977 11940 3981 11996
rect 3917 11936 3981 11940
rect 3997 11996 4061 12000
rect 3997 11940 4001 11996
rect 4001 11940 4057 11996
rect 4057 11940 4061 11996
rect 3997 11936 4061 11940
rect 4077 11996 4141 12000
rect 4077 11940 4081 11996
rect 4081 11940 4137 11996
rect 4137 11940 4141 11996
rect 4077 11936 4141 11940
rect 4157 11996 4221 12000
rect 4157 11940 4161 11996
rect 4161 11940 4217 11996
rect 4217 11940 4221 11996
rect 4157 11936 4221 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 15778 11996 15842 12000
rect 15778 11940 15782 11996
rect 15782 11940 15838 11996
rect 15838 11940 15842 11996
rect 15778 11936 15842 11940
rect 15858 11996 15922 12000
rect 15858 11940 15862 11996
rect 15862 11940 15918 11996
rect 15918 11940 15922 11996
rect 15858 11936 15922 11940
rect 15938 11996 16002 12000
rect 15938 11940 15942 11996
rect 15942 11940 15998 11996
rect 15998 11940 16002 11996
rect 15938 11936 16002 11940
rect 16018 11996 16082 12000
rect 16018 11940 16022 11996
rect 16022 11940 16078 11996
rect 16078 11940 16082 11996
rect 16018 11936 16082 11940
rect 6882 11452 6946 11456
rect 6882 11396 6886 11452
rect 6886 11396 6942 11452
rect 6942 11396 6946 11452
rect 6882 11392 6946 11396
rect 6962 11452 7026 11456
rect 6962 11396 6966 11452
rect 6966 11396 7022 11452
rect 7022 11396 7026 11452
rect 6962 11392 7026 11396
rect 7042 11452 7106 11456
rect 7042 11396 7046 11452
rect 7046 11396 7102 11452
rect 7102 11396 7106 11452
rect 7042 11392 7106 11396
rect 7122 11452 7186 11456
rect 7122 11396 7126 11452
rect 7126 11396 7182 11452
rect 7182 11396 7186 11452
rect 7122 11392 7186 11396
rect 12813 11452 12877 11456
rect 12813 11396 12817 11452
rect 12817 11396 12873 11452
rect 12873 11396 12877 11452
rect 12813 11392 12877 11396
rect 12893 11452 12957 11456
rect 12893 11396 12897 11452
rect 12897 11396 12953 11452
rect 12953 11396 12957 11452
rect 12893 11392 12957 11396
rect 12973 11452 13037 11456
rect 12973 11396 12977 11452
rect 12977 11396 13033 11452
rect 13033 11396 13037 11452
rect 12973 11392 13037 11396
rect 13053 11452 13117 11456
rect 13053 11396 13057 11452
rect 13057 11396 13113 11452
rect 13113 11396 13117 11452
rect 13053 11392 13117 11396
rect 11284 11052 11348 11116
rect 3917 10908 3981 10912
rect 3917 10852 3921 10908
rect 3921 10852 3977 10908
rect 3977 10852 3981 10908
rect 3917 10848 3981 10852
rect 3997 10908 4061 10912
rect 3997 10852 4001 10908
rect 4001 10852 4057 10908
rect 4057 10852 4061 10908
rect 3997 10848 4061 10852
rect 4077 10908 4141 10912
rect 4077 10852 4081 10908
rect 4081 10852 4137 10908
rect 4137 10852 4141 10908
rect 4077 10848 4141 10852
rect 4157 10908 4221 10912
rect 4157 10852 4161 10908
rect 4161 10852 4217 10908
rect 4217 10852 4221 10908
rect 4157 10848 4221 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 15778 10908 15842 10912
rect 15778 10852 15782 10908
rect 15782 10852 15838 10908
rect 15838 10852 15842 10908
rect 15778 10848 15842 10852
rect 15858 10908 15922 10912
rect 15858 10852 15862 10908
rect 15862 10852 15918 10908
rect 15918 10852 15922 10908
rect 15858 10848 15922 10852
rect 15938 10908 16002 10912
rect 15938 10852 15942 10908
rect 15942 10852 15998 10908
rect 15998 10852 16002 10908
rect 15938 10848 16002 10852
rect 16018 10908 16082 10912
rect 16018 10852 16022 10908
rect 16022 10852 16078 10908
rect 16078 10852 16082 10908
rect 16018 10848 16082 10852
rect 12020 10780 12084 10844
rect 16804 10508 16868 10572
rect 6882 10364 6946 10368
rect 6882 10308 6886 10364
rect 6886 10308 6942 10364
rect 6942 10308 6946 10364
rect 6882 10304 6946 10308
rect 6962 10364 7026 10368
rect 6962 10308 6966 10364
rect 6966 10308 7022 10364
rect 7022 10308 7026 10364
rect 6962 10304 7026 10308
rect 7042 10364 7106 10368
rect 7042 10308 7046 10364
rect 7046 10308 7102 10364
rect 7102 10308 7106 10364
rect 7042 10304 7106 10308
rect 7122 10364 7186 10368
rect 7122 10308 7126 10364
rect 7126 10308 7182 10364
rect 7182 10308 7186 10364
rect 7122 10304 7186 10308
rect 12813 10364 12877 10368
rect 12813 10308 12817 10364
rect 12817 10308 12873 10364
rect 12873 10308 12877 10364
rect 12813 10304 12877 10308
rect 12893 10364 12957 10368
rect 12893 10308 12897 10364
rect 12897 10308 12953 10364
rect 12953 10308 12957 10364
rect 12893 10304 12957 10308
rect 12973 10364 13037 10368
rect 12973 10308 12977 10364
rect 12977 10308 13033 10364
rect 13033 10308 13037 10364
rect 12973 10304 13037 10308
rect 13053 10364 13117 10368
rect 13053 10308 13057 10364
rect 13057 10308 13113 10364
rect 13113 10308 13117 10364
rect 13053 10304 13117 10308
rect 3556 10236 3620 10300
rect 16620 10100 16684 10164
rect 3556 9888 3620 9892
rect 3556 9832 3570 9888
rect 3570 9832 3620 9888
rect 3556 9828 3620 9832
rect 3917 9820 3981 9824
rect 3917 9764 3921 9820
rect 3921 9764 3977 9820
rect 3977 9764 3981 9820
rect 3917 9760 3981 9764
rect 3997 9820 4061 9824
rect 3997 9764 4001 9820
rect 4001 9764 4057 9820
rect 4057 9764 4061 9820
rect 3997 9760 4061 9764
rect 4077 9820 4141 9824
rect 4077 9764 4081 9820
rect 4081 9764 4137 9820
rect 4137 9764 4141 9820
rect 4077 9760 4141 9764
rect 4157 9820 4221 9824
rect 4157 9764 4161 9820
rect 4161 9764 4217 9820
rect 4217 9764 4221 9820
rect 4157 9760 4221 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 15778 9820 15842 9824
rect 15778 9764 15782 9820
rect 15782 9764 15838 9820
rect 15838 9764 15842 9820
rect 15778 9760 15842 9764
rect 15858 9820 15922 9824
rect 15858 9764 15862 9820
rect 15862 9764 15918 9820
rect 15918 9764 15922 9820
rect 15858 9760 15922 9764
rect 15938 9820 16002 9824
rect 15938 9764 15942 9820
rect 15942 9764 15998 9820
rect 15998 9764 16002 9820
rect 15938 9760 16002 9764
rect 16018 9820 16082 9824
rect 16018 9764 16022 9820
rect 16022 9764 16078 9820
rect 16078 9764 16082 9820
rect 16018 9760 16082 9764
rect 12388 9556 12452 9620
rect 8156 9284 8220 9348
rect 8708 9344 8772 9348
rect 8708 9288 8758 9344
rect 8758 9288 8772 9344
rect 8708 9284 8772 9288
rect 14412 9480 14476 9484
rect 14412 9424 14426 9480
rect 14426 9424 14476 9480
rect 14412 9420 14476 9424
rect 12020 9284 12084 9348
rect 6882 9276 6946 9280
rect 6882 9220 6886 9276
rect 6886 9220 6942 9276
rect 6942 9220 6946 9276
rect 6882 9216 6946 9220
rect 6962 9276 7026 9280
rect 6962 9220 6966 9276
rect 6966 9220 7022 9276
rect 7022 9220 7026 9276
rect 6962 9216 7026 9220
rect 7042 9276 7106 9280
rect 7042 9220 7046 9276
rect 7046 9220 7102 9276
rect 7102 9220 7106 9276
rect 7042 9216 7106 9220
rect 7122 9276 7186 9280
rect 7122 9220 7126 9276
rect 7126 9220 7182 9276
rect 7182 9220 7186 9276
rect 7122 9216 7186 9220
rect 12813 9276 12877 9280
rect 12813 9220 12817 9276
rect 12817 9220 12873 9276
rect 12873 9220 12877 9276
rect 12813 9216 12877 9220
rect 12893 9276 12957 9280
rect 12893 9220 12897 9276
rect 12897 9220 12953 9276
rect 12953 9220 12957 9276
rect 12893 9216 12957 9220
rect 12973 9276 13037 9280
rect 12973 9220 12977 9276
rect 12977 9220 13033 9276
rect 13033 9220 13037 9276
rect 12973 9216 13037 9220
rect 13053 9276 13117 9280
rect 13053 9220 13057 9276
rect 13057 9220 13113 9276
rect 13113 9220 13117 9276
rect 13053 9216 13117 9220
rect 12572 9148 12636 9212
rect 7972 8936 8036 8940
rect 7972 8880 7986 8936
rect 7986 8880 8036 8936
rect 7972 8876 8036 8880
rect 8708 8800 8772 8804
rect 11284 8876 11348 8940
rect 11836 8876 11900 8940
rect 8708 8744 8758 8800
rect 8758 8744 8772 8800
rect 8708 8740 8772 8744
rect 3917 8732 3981 8736
rect 3917 8676 3921 8732
rect 3921 8676 3977 8732
rect 3977 8676 3981 8732
rect 3917 8672 3981 8676
rect 3997 8732 4061 8736
rect 3997 8676 4001 8732
rect 4001 8676 4057 8732
rect 4057 8676 4061 8732
rect 3997 8672 4061 8676
rect 4077 8732 4141 8736
rect 4077 8676 4081 8732
rect 4081 8676 4137 8732
rect 4137 8676 4141 8732
rect 4077 8672 4141 8676
rect 4157 8732 4221 8736
rect 4157 8676 4161 8732
rect 4161 8676 4217 8732
rect 4217 8676 4221 8732
rect 4157 8672 4221 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 15778 8732 15842 8736
rect 15778 8676 15782 8732
rect 15782 8676 15838 8732
rect 15838 8676 15842 8732
rect 15778 8672 15842 8676
rect 15858 8732 15922 8736
rect 15858 8676 15862 8732
rect 15862 8676 15918 8732
rect 15918 8676 15922 8732
rect 15858 8672 15922 8676
rect 15938 8732 16002 8736
rect 15938 8676 15942 8732
rect 15942 8676 15998 8732
rect 15998 8676 16002 8732
rect 15938 8672 16002 8676
rect 16018 8732 16082 8736
rect 16018 8676 16022 8732
rect 16022 8676 16078 8732
rect 16078 8676 16082 8732
rect 16018 8672 16082 8676
rect 9260 8604 9324 8668
rect 16620 8740 16684 8804
rect 15332 8468 15396 8532
rect 16620 8332 16684 8396
rect 3004 8196 3068 8260
rect 12388 8196 12452 8260
rect 6882 8188 6946 8192
rect 6882 8132 6886 8188
rect 6886 8132 6942 8188
rect 6942 8132 6946 8188
rect 6882 8128 6946 8132
rect 6962 8188 7026 8192
rect 6962 8132 6966 8188
rect 6966 8132 7022 8188
rect 7022 8132 7026 8188
rect 6962 8128 7026 8132
rect 7042 8188 7106 8192
rect 7042 8132 7046 8188
rect 7046 8132 7102 8188
rect 7102 8132 7106 8188
rect 7042 8128 7106 8132
rect 7122 8188 7186 8192
rect 7122 8132 7126 8188
rect 7126 8132 7182 8188
rect 7182 8132 7186 8188
rect 7122 8128 7186 8132
rect 12813 8188 12877 8192
rect 12813 8132 12817 8188
rect 12817 8132 12873 8188
rect 12873 8132 12877 8188
rect 12813 8128 12877 8132
rect 12893 8188 12957 8192
rect 12893 8132 12897 8188
rect 12897 8132 12953 8188
rect 12953 8132 12957 8188
rect 12893 8128 12957 8132
rect 12973 8188 13037 8192
rect 12973 8132 12977 8188
rect 12977 8132 13033 8188
rect 13033 8132 13037 8188
rect 12973 8128 13037 8132
rect 13053 8188 13117 8192
rect 13053 8132 13057 8188
rect 13057 8132 13113 8188
rect 13113 8132 13117 8188
rect 13053 8128 13117 8132
rect 16252 8060 16316 8124
rect 15516 7924 15580 7988
rect 9260 7652 9324 7716
rect 3917 7644 3981 7648
rect 3917 7588 3921 7644
rect 3921 7588 3977 7644
rect 3977 7588 3981 7644
rect 3917 7584 3981 7588
rect 3997 7644 4061 7648
rect 3997 7588 4001 7644
rect 4001 7588 4057 7644
rect 4057 7588 4061 7644
rect 3997 7584 4061 7588
rect 4077 7644 4141 7648
rect 4077 7588 4081 7644
rect 4081 7588 4137 7644
rect 4137 7588 4141 7644
rect 4077 7584 4141 7588
rect 4157 7644 4221 7648
rect 4157 7588 4161 7644
rect 4161 7588 4217 7644
rect 4217 7588 4221 7644
rect 4157 7584 4221 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 8156 7576 8220 7580
rect 8156 7520 8206 7576
rect 8206 7520 8220 7576
rect 8156 7516 8220 7520
rect 9260 7244 9324 7308
rect 14964 7652 15028 7716
rect 15516 7652 15580 7716
rect 15778 7644 15842 7648
rect 15778 7588 15782 7644
rect 15782 7588 15838 7644
rect 15838 7588 15842 7644
rect 15778 7584 15842 7588
rect 15858 7644 15922 7648
rect 15858 7588 15862 7644
rect 15862 7588 15918 7644
rect 15918 7588 15922 7644
rect 15858 7584 15922 7588
rect 15938 7644 16002 7648
rect 15938 7588 15942 7644
rect 15942 7588 15998 7644
rect 15998 7588 16002 7644
rect 15938 7584 16002 7588
rect 16018 7644 16082 7648
rect 16018 7588 16022 7644
rect 16022 7588 16078 7644
rect 16078 7588 16082 7644
rect 16018 7584 16082 7588
rect 7972 7108 8036 7172
rect 13860 7108 13924 7172
rect 6882 7100 6946 7104
rect 6882 7044 6886 7100
rect 6886 7044 6942 7100
rect 6942 7044 6946 7100
rect 6882 7040 6946 7044
rect 6962 7100 7026 7104
rect 6962 7044 6966 7100
rect 6966 7044 7022 7100
rect 7022 7044 7026 7100
rect 6962 7040 7026 7044
rect 7042 7100 7106 7104
rect 7042 7044 7046 7100
rect 7046 7044 7102 7100
rect 7102 7044 7106 7100
rect 7042 7040 7106 7044
rect 7122 7100 7186 7104
rect 7122 7044 7126 7100
rect 7126 7044 7182 7100
rect 7182 7044 7186 7100
rect 7122 7040 7186 7044
rect 12813 7100 12877 7104
rect 12813 7044 12817 7100
rect 12817 7044 12873 7100
rect 12873 7044 12877 7100
rect 12813 7040 12877 7044
rect 12893 7100 12957 7104
rect 12893 7044 12897 7100
rect 12897 7044 12953 7100
rect 12953 7044 12957 7100
rect 12893 7040 12957 7044
rect 12973 7100 13037 7104
rect 12973 7044 12977 7100
rect 12977 7044 13033 7100
rect 13033 7044 13037 7100
rect 12973 7040 13037 7044
rect 13053 7100 13117 7104
rect 13053 7044 13057 7100
rect 13057 7044 13113 7100
rect 13113 7044 13117 7100
rect 13053 7040 13117 7044
rect 3917 6556 3981 6560
rect 3917 6500 3921 6556
rect 3921 6500 3977 6556
rect 3977 6500 3981 6556
rect 3917 6496 3981 6500
rect 3997 6556 4061 6560
rect 3997 6500 4001 6556
rect 4001 6500 4057 6556
rect 4057 6500 4061 6556
rect 3997 6496 4061 6500
rect 4077 6556 4141 6560
rect 4077 6500 4081 6556
rect 4081 6500 4137 6556
rect 4137 6500 4141 6556
rect 4077 6496 4141 6500
rect 4157 6556 4221 6560
rect 4157 6500 4161 6556
rect 4161 6500 4217 6556
rect 4217 6500 4221 6556
rect 4157 6496 4221 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 15778 6556 15842 6560
rect 15778 6500 15782 6556
rect 15782 6500 15838 6556
rect 15838 6500 15842 6556
rect 15778 6496 15842 6500
rect 15858 6556 15922 6560
rect 15858 6500 15862 6556
rect 15862 6500 15918 6556
rect 15918 6500 15922 6556
rect 15858 6496 15922 6500
rect 15938 6556 16002 6560
rect 15938 6500 15942 6556
rect 15942 6500 15998 6556
rect 15998 6500 16002 6556
rect 15938 6496 16002 6500
rect 16018 6556 16082 6560
rect 16018 6500 16022 6556
rect 16022 6500 16078 6556
rect 16078 6500 16082 6556
rect 16018 6496 16082 6500
rect 6882 6012 6946 6016
rect 6882 5956 6886 6012
rect 6886 5956 6942 6012
rect 6942 5956 6946 6012
rect 6882 5952 6946 5956
rect 6962 6012 7026 6016
rect 6962 5956 6966 6012
rect 6966 5956 7022 6012
rect 7022 5956 7026 6012
rect 6962 5952 7026 5956
rect 7042 6012 7106 6016
rect 7042 5956 7046 6012
rect 7046 5956 7102 6012
rect 7102 5956 7106 6012
rect 7042 5952 7106 5956
rect 7122 6012 7186 6016
rect 7122 5956 7126 6012
rect 7126 5956 7182 6012
rect 7182 5956 7186 6012
rect 7122 5952 7186 5956
rect 12813 6012 12877 6016
rect 12813 5956 12817 6012
rect 12817 5956 12873 6012
rect 12873 5956 12877 6012
rect 12813 5952 12877 5956
rect 12893 6012 12957 6016
rect 12893 5956 12897 6012
rect 12897 5956 12953 6012
rect 12953 5956 12957 6012
rect 12893 5952 12957 5956
rect 12973 6012 13037 6016
rect 12973 5956 12977 6012
rect 12977 5956 13033 6012
rect 13033 5956 13037 6012
rect 12973 5952 13037 5956
rect 13053 6012 13117 6016
rect 13053 5956 13057 6012
rect 13057 5956 13113 6012
rect 13113 5956 13117 6012
rect 13053 5952 13117 5956
rect 12020 5612 12084 5676
rect 13308 5612 13372 5676
rect 3917 5468 3981 5472
rect 3917 5412 3921 5468
rect 3921 5412 3977 5468
rect 3977 5412 3981 5468
rect 3917 5408 3981 5412
rect 3997 5468 4061 5472
rect 3997 5412 4001 5468
rect 4001 5412 4057 5468
rect 4057 5412 4061 5468
rect 3997 5408 4061 5412
rect 4077 5468 4141 5472
rect 4077 5412 4081 5468
rect 4081 5412 4137 5468
rect 4137 5412 4141 5468
rect 4077 5408 4141 5412
rect 4157 5468 4221 5472
rect 4157 5412 4161 5468
rect 4161 5412 4217 5468
rect 4217 5412 4221 5468
rect 4157 5408 4221 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 15778 5468 15842 5472
rect 15778 5412 15782 5468
rect 15782 5412 15838 5468
rect 15838 5412 15842 5468
rect 15778 5408 15842 5412
rect 15858 5468 15922 5472
rect 15858 5412 15862 5468
rect 15862 5412 15918 5468
rect 15918 5412 15922 5468
rect 15858 5408 15922 5412
rect 15938 5468 16002 5472
rect 15938 5412 15942 5468
rect 15942 5412 15998 5468
rect 15998 5412 16002 5468
rect 15938 5408 16002 5412
rect 16018 5468 16082 5472
rect 16018 5412 16022 5468
rect 16022 5412 16078 5468
rect 16078 5412 16082 5468
rect 16018 5408 16082 5412
rect 12572 5068 12636 5132
rect 15516 5068 15580 5132
rect 6882 4924 6946 4928
rect 6882 4868 6886 4924
rect 6886 4868 6942 4924
rect 6942 4868 6946 4924
rect 6882 4864 6946 4868
rect 6962 4924 7026 4928
rect 6962 4868 6966 4924
rect 6966 4868 7022 4924
rect 7022 4868 7026 4924
rect 6962 4864 7026 4868
rect 7042 4924 7106 4928
rect 7042 4868 7046 4924
rect 7046 4868 7102 4924
rect 7102 4868 7106 4924
rect 7042 4864 7106 4868
rect 7122 4924 7186 4928
rect 7122 4868 7126 4924
rect 7126 4868 7182 4924
rect 7182 4868 7186 4924
rect 7122 4864 7186 4868
rect 12813 4924 12877 4928
rect 12813 4868 12817 4924
rect 12817 4868 12873 4924
rect 12873 4868 12877 4924
rect 12813 4864 12877 4868
rect 12893 4924 12957 4928
rect 12893 4868 12897 4924
rect 12897 4868 12953 4924
rect 12953 4868 12957 4924
rect 12893 4864 12957 4868
rect 12973 4924 13037 4928
rect 12973 4868 12977 4924
rect 12977 4868 13033 4924
rect 13033 4868 13037 4924
rect 12973 4864 13037 4868
rect 13053 4924 13117 4928
rect 13053 4868 13057 4924
rect 13057 4868 13113 4924
rect 13113 4868 13117 4924
rect 13053 4864 13117 4868
rect 15516 4660 15580 4724
rect 3917 4380 3981 4384
rect 3917 4324 3921 4380
rect 3921 4324 3977 4380
rect 3977 4324 3981 4380
rect 3917 4320 3981 4324
rect 3997 4380 4061 4384
rect 3997 4324 4001 4380
rect 4001 4324 4057 4380
rect 4057 4324 4061 4380
rect 3997 4320 4061 4324
rect 4077 4380 4141 4384
rect 4077 4324 4081 4380
rect 4081 4324 4137 4380
rect 4137 4324 4141 4380
rect 4077 4320 4141 4324
rect 4157 4380 4221 4384
rect 4157 4324 4161 4380
rect 4161 4324 4217 4380
rect 4217 4324 4221 4380
rect 4157 4320 4221 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 15778 4380 15842 4384
rect 15778 4324 15782 4380
rect 15782 4324 15838 4380
rect 15838 4324 15842 4380
rect 15778 4320 15842 4324
rect 15858 4380 15922 4384
rect 15858 4324 15862 4380
rect 15862 4324 15918 4380
rect 15918 4324 15922 4380
rect 15858 4320 15922 4324
rect 15938 4380 16002 4384
rect 15938 4324 15942 4380
rect 15942 4324 15998 4380
rect 15998 4324 16002 4380
rect 15938 4320 16002 4324
rect 16018 4380 16082 4384
rect 16018 4324 16022 4380
rect 16022 4324 16078 4380
rect 16078 4324 16082 4380
rect 16018 4320 16082 4324
rect 14780 3980 14844 4044
rect 16804 3980 16868 4044
rect 16436 3844 16500 3908
rect 6882 3836 6946 3840
rect 6882 3780 6886 3836
rect 6886 3780 6942 3836
rect 6942 3780 6946 3836
rect 6882 3776 6946 3780
rect 6962 3836 7026 3840
rect 6962 3780 6966 3836
rect 6966 3780 7022 3836
rect 7022 3780 7026 3836
rect 6962 3776 7026 3780
rect 7042 3836 7106 3840
rect 7042 3780 7046 3836
rect 7046 3780 7102 3836
rect 7102 3780 7106 3836
rect 7042 3776 7106 3780
rect 7122 3836 7186 3840
rect 7122 3780 7126 3836
rect 7126 3780 7182 3836
rect 7182 3780 7186 3836
rect 7122 3776 7186 3780
rect 12813 3836 12877 3840
rect 12813 3780 12817 3836
rect 12817 3780 12873 3836
rect 12873 3780 12877 3836
rect 12813 3776 12877 3780
rect 12893 3836 12957 3840
rect 12893 3780 12897 3836
rect 12897 3780 12953 3836
rect 12953 3780 12957 3836
rect 12893 3776 12957 3780
rect 12973 3836 13037 3840
rect 12973 3780 12977 3836
rect 12977 3780 13033 3836
rect 13033 3780 13037 3836
rect 12973 3776 13037 3780
rect 13053 3836 13117 3840
rect 13053 3780 13057 3836
rect 13057 3780 13113 3836
rect 13113 3780 13117 3836
rect 13053 3776 13117 3780
rect 14412 3632 14476 3636
rect 14412 3576 14462 3632
rect 14462 3576 14476 3632
rect 14412 3572 14476 3576
rect 3917 3292 3981 3296
rect 3917 3236 3921 3292
rect 3921 3236 3977 3292
rect 3977 3236 3981 3292
rect 3917 3232 3981 3236
rect 3997 3292 4061 3296
rect 3997 3236 4001 3292
rect 4001 3236 4057 3292
rect 4057 3236 4061 3292
rect 3997 3232 4061 3236
rect 4077 3292 4141 3296
rect 4077 3236 4081 3292
rect 4081 3236 4137 3292
rect 4137 3236 4141 3292
rect 4077 3232 4141 3236
rect 4157 3292 4221 3296
rect 4157 3236 4161 3292
rect 4161 3236 4217 3292
rect 4217 3236 4221 3292
rect 4157 3232 4221 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 15778 3292 15842 3296
rect 15778 3236 15782 3292
rect 15782 3236 15838 3292
rect 15838 3236 15842 3292
rect 15778 3232 15842 3236
rect 15858 3292 15922 3296
rect 15858 3236 15862 3292
rect 15862 3236 15918 3292
rect 15918 3236 15922 3292
rect 15858 3232 15922 3236
rect 15938 3292 16002 3296
rect 15938 3236 15942 3292
rect 15942 3236 15998 3292
rect 15998 3236 16002 3292
rect 15938 3232 16002 3236
rect 16018 3292 16082 3296
rect 16018 3236 16022 3292
rect 16022 3236 16078 3292
rect 16078 3236 16082 3292
rect 16018 3232 16082 3236
rect 10364 2952 10428 2956
rect 10364 2896 10378 2952
rect 10378 2896 10428 2952
rect 10364 2892 10428 2896
rect 15148 2892 15212 2956
rect 6882 2748 6946 2752
rect 6882 2692 6886 2748
rect 6886 2692 6942 2748
rect 6942 2692 6946 2748
rect 6882 2688 6946 2692
rect 6962 2748 7026 2752
rect 6962 2692 6966 2748
rect 6966 2692 7022 2748
rect 7022 2692 7026 2748
rect 6962 2688 7026 2692
rect 7042 2748 7106 2752
rect 7042 2692 7046 2748
rect 7046 2692 7102 2748
rect 7102 2692 7106 2748
rect 7042 2688 7106 2692
rect 7122 2748 7186 2752
rect 7122 2692 7126 2748
rect 7126 2692 7182 2748
rect 7182 2692 7186 2748
rect 7122 2688 7186 2692
rect 12813 2748 12877 2752
rect 12813 2692 12817 2748
rect 12817 2692 12873 2748
rect 12873 2692 12877 2748
rect 12813 2688 12877 2692
rect 12893 2748 12957 2752
rect 12893 2692 12897 2748
rect 12897 2692 12953 2748
rect 12953 2692 12957 2748
rect 12893 2688 12957 2692
rect 12973 2748 13037 2752
rect 12973 2692 12977 2748
rect 12977 2692 13033 2748
rect 13033 2692 13037 2748
rect 12973 2688 13037 2692
rect 13053 2748 13117 2752
rect 13053 2692 13057 2748
rect 13057 2692 13113 2748
rect 13113 2692 13117 2748
rect 13053 2688 13117 2692
rect 15332 2620 15396 2684
rect 16620 2620 16684 2684
rect 11836 2544 11900 2548
rect 11836 2488 11850 2544
rect 11850 2488 11900 2544
rect 11836 2484 11900 2488
rect 3917 2204 3981 2208
rect 3917 2148 3921 2204
rect 3921 2148 3977 2204
rect 3977 2148 3981 2204
rect 3917 2144 3981 2148
rect 3997 2204 4061 2208
rect 3997 2148 4001 2204
rect 4001 2148 4057 2204
rect 4057 2148 4061 2204
rect 3997 2144 4061 2148
rect 4077 2204 4141 2208
rect 4077 2148 4081 2204
rect 4081 2148 4137 2204
rect 4137 2148 4141 2204
rect 4077 2144 4141 2148
rect 4157 2204 4221 2208
rect 4157 2148 4161 2204
rect 4161 2148 4217 2204
rect 4217 2148 4221 2204
rect 4157 2144 4221 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 15778 2204 15842 2208
rect 15778 2148 15782 2204
rect 15782 2148 15838 2204
rect 15838 2148 15842 2204
rect 15778 2144 15842 2148
rect 15858 2204 15922 2208
rect 15858 2148 15862 2204
rect 15862 2148 15918 2204
rect 15918 2148 15922 2204
rect 15858 2144 15922 2148
rect 15938 2204 16002 2208
rect 15938 2148 15942 2204
rect 15942 2148 15998 2204
rect 15998 2148 16002 2204
rect 15938 2144 16002 2148
rect 16018 2204 16082 2208
rect 16018 2148 16022 2204
rect 16022 2148 16078 2204
rect 16078 2148 16082 2204
rect 16018 2144 16082 2148
<< metal4 >>
rect 16251 15468 16317 15469
rect 16251 15404 16252 15468
rect 16316 15404 16317 15468
rect 16251 15403 16317 15404
rect 3909 14176 4229 14736
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 13088 4229 14112
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3003 12340 3069 12341
rect 3003 12276 3004 12340
rect 3068 12276 3069 12340
rect 3003 12275 3069 12276
rect 3006 8261 3066 12275
rect 3909 12000 4229 13024
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 10912 4229 11936
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3555 10300 3621 10301
rect 3555 10236 3556 10300
rect 3620 10236 3621 10300
rect 3555 10235 3621 10236
rect 3558 9893 3618 10235
rect 3555 9892 3621 9893
rect 3555 9828 3556 9892
rect 3620 9828 3621 9892
rect 3555 9827 3621 9828
rect 3909 9824 4229 10848
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 8736 4229 9760
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3003 8260 3069 8261
rect 3003 8196 3004 8260
rect 3068 8196 3069 8260
rect 3003 8195 3069 8196
rect 3909 7648 4229 8672
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 6560 4229 7584
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 5472 4229 6496
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 4384 4229 5408
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 3296 4229 4320
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 2208 4229 3232
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2128 4229 2144
rect 6874 14720 7195 14736
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7195 14720
rect 6874 13632 7195 14656
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7195 13632
rect 6874 12544 7195 13568
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7195 12544
rect 6874 11456 7195 12480
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7195 11456
rect 6874 10368 7195 11392
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7195 10368
rect 6874 9280 7195 10304
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 12000 10160 13024
rect 12805 14720 13125 14736
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 13632 13125 14656
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 12544 13125 13568
rect 15770 14176 16090 14736
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 14779 13428 14845 13429
rect 14779 13364 14780 13428
rect 14844 13364 14845 13428
rect 14779 13363 14845 13364
rect 15147 13428 15213 13429
rect 15147 13364 15148 13428
rect 15212 13364 15213 13428
rect 15147 13363 15213 13364
rect 13307 13156 13373 13157
rect 13307 13092 13308 13156
rect 13372 13092 13373 13156
rect 13307 13091 13373 13092
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 10363 12476 10429 12477
rect 10363 12412 10364 12476
rect 10428 12412 10429 12476
rect 10363 12411 10429 12412
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 8155 9348 8221 9349
rect 8155 9284 8156 9348
rect 8220 9284 8221 9348
rect 8155 9283 8221 9284
rect 8707 9348 8773 9349
rect 8707 9284 8708 9348
rect 8772 9284 8773 9348
rect 8707 9283 8773 9284
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7195 9280
rect 6874 8192 7195 9216
rect 7971 8940 8037 8941
rect 7971 8876 7972 8940
rect 8036 8876 8037 8940
rect 7971 8875 8037 8876
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7195 8192
rect 6874 7104 7195 8128
rect 7974 7173 8034 8875
rect 8158 7581 8218 9283
rect 8710 8805 8770 9283
rect 8707 8804 8773 8805
rect 8707 8740 8708 8804
rect 8772 8740 8773 8804
rect 8707 8739 8773 8740
rect 9840 8736 10160 9760
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9259 8668 9325 8669
rect 9259 8604 9260 8668
rect 9324 8604 9325 8668
rect 9259 8603 9325 8604
rect 9262 7717 9322 8603
rect 9259 7716 9325 7717
rect 9259 7652 9260 7716
rect 9324 7652 9325 7716
rect 9259 7651 9325 7652
rect 8155 7580 8221 7581
rect 8155 7516 8156 7580
rect 8220 7516 8221 7580
rect 8155 7515 8221 7516
rect 9262 7309 9322 7651
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9259 7308 9325 7309
rect 9259 7244 9260 7308
rect 9324 7244 9325 7308
rect 9259 7243 9325 7244
rect 7971 7172 8037 7173
rect 7971 7108 7972 7172
rect 8036 7108 8037 7172
rect 7971 7107 8037 7108
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7195 7104
rect 6874 6016 7195 7040
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7195 6016
rect 6874 4928 7195 5952
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7195 4928
rect 6874 3840 7195 4864
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7195 3840
rect 6874 2752 7195 3776
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7195 2752
rect 6874 2128 7195 2688
rect 9840 6560 10160 7584
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 2208 10160 3232
rect 10366 2957 10426 12411
rect 12805 11456 13125 12480
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 11283 11116 11349 11117
rect 11283 11052 11284 11116
rect 11348 11052 11349 11116
rect 11283 11051 11349 11052
rect 11286 8941 11346 11051
rect 12019 10844 12085 10845
rect 12019 10780 12020 10844
rect 12084 10780 12085 10844
rect 12019 10779 12085 10780
rect 12022 9349 12082 10779
rect 12805 10368 13125 11392
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 12387 9620 12453 9621
rect 12387 9556 12388 9620
rect 12452 9556 12453 9620
rect 12387 9555 12453 9556
rect 12019 9348 12085 9349
rect 12019 9284 12020 9348
rect 12084 9284 12085 9348
rect 12019 9283 12085 9284
rect 11283 8940 11349 8941
rect 11283 8876 11284 8940
rect 11348 8876 11349 8940
rect 11283 8875 11349 8876
rect 11835 8940 11901 8941
rect 11835 8876 11836 8940
rect 11900 8876 11901 8940
rect 11835 8875 11901 8876
rect 10363 2956 10429 2957
rect 10363 2892 10364 2956
rect 10428 2892 10429 2956
rect 10363 2891 10429 2892
rect 11838 2549 11898 8875
rect 12022 5677 12082 9283
rect 12390 8261 12450 9555
rect 12805 9280 13125 10304
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12571 9212 12637 9213
rect 12571 9148 12572 9212
rect 12636 9148 12637 9212
rect 12571 9147 12637 9148
rect 12387 8260 12453 8261
rect 12387 8196 12388 8260
rect 12452 8196 12453 8260
rect 12387 8195 12453 8196
rect 12019 5676 12085 5677
rect 12019 5612 12020 5676
rect 12084 5612 12085 5676
rect 12019 5611 12085 5612
rect 12574 5133 12634 9147
rect 12805 8192 13125 9216
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 12805 7104 13125 8128
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 6016 13125 7040
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12571 5132 12637 5133
rect 12571 5068 12572 5132
rect 12636 5068 12637 5132
rect 12571 5067 12637 5068
rect 12805 4928 13125 5952
rect 13310 5677 13370 13091
rect 13859 12748 13925 12749
rect 13859 12684 13860 12748
rect 13924 12684 13925 12748
rect 13859 12683 13925 12684
rect 13862 7173 13922 12683
rect 14411 9484 14477 9485
rect 14411 9420 14412 9484
rect 14476 9420 14477 9484
rect 14411 9419 14477 9420
rect 13859 7172 13925 7173
rect 13859 7108 13860 7172
rect 13924 7108 13925 7172
rect 13859 7107 13925 7108
rect 13307 5676 13373 5677
rect 13307 5612 13308 5676
rect 13372 5612 13373 5676
rect 13307 5611 13373 5612
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 3840 13125 4864
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 2752 13125 3776
rect 14414 3637 14474 9419
rect 14782 4045 14842 13363
rect 14963 12884 15029 12885
rect 14963 12820 14964 12884
rect 15028 12820 15029 12884
rect 14963 12819 15029 12820
rect 14966 7717 15026 12819
rect 14963 7716 15029 7717
rect 14963 7652 14964 7716
rect 15028 7652 15029 7716
rect 14963 7651 15029 7652
rect 14779 4044 14845 4045
rect 14779 3980 14780 4044
rect 14844 3980 14845 4044
rect 14779 3979 14845 3980
rect 14411 3636 14477 3637
rect 14411 3572 14412 3636
rect 14476 3572 14477 3636
rect 14411 3571 14477 3572
rect 15150 2957 15210 13363
rect 15770 13088 16090 14112
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 15515 12476 15581 12477
rect 15515 12412 15516 12476
rect 15580 12412 15581 12476
rect 15515 12411 15581 12412
rect 15331 8532 15397 8533
rect 15331 8468 15332 8532
rect 15396 8468 15397 8532
rect 15331 8467 15397 8468
rect 15147 2956 15213 2957
rect 15147 2892 15148 2956
rect 15212 2892 15213 2956
rect 15147 2891 15213 2892
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 11835 2548 11901 2549
rect 11835 2484 11836 2548
rect 11900 2484 11901 2548
rect 11835 2483 11901 2484
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12805 2128 13125 2688
rect 15334 2685 15394 8467
rect 15518 7989 15578 12411
rect 15770 12000 16090 13024
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 15770 10912 16090 11936
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15770 9824 16090 10848
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 15770 8736 16090 9760
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 15515 7988 15581 7989
rect 15515 7924 15516 7988
rect 15580 7924 15581 7988
rect 15515 7923 15581 7924
rect 15515 7716 15581 7717
rect 15515 7652 15516 7716
rect 15580 7652 15581 7716
rect 15515 7651 15581 7652
rect 15518 5133 15578 7651
rect 15770 7648 16090 8672
rect 16254 8125 16314 15403
rect 16435 12612 16501 12613
rect 16435 12548 16436 12612
rect 16500 12548 16501 12612
rect 16435 12547 16501 12548
rect 16251 8124 16317 8125
rect 16251 8060 16252 8124
rect 16316 8060 16317 8124
rect 16251 8059 16317 8060
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 6560 16090 7584
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 15770 5472 16090 6496
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 15515 5132 15581 5133
rect 15515 5068 15516 5132
rect 15580 5068 15581 5132
rect 15515 5067 15581 5068
rect 15518 4725 15578 5067
rect 15515 4724 15581 4725
rect 15515 4660 15516 4724
rect 15580 4660 15581 4724
rect 15515 4659 15581 4660
rect 15770 4384 16090 5408
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 15770 3296 16090 4320
rect 16438 3909 16498 12547
rect 16803 10572 16869 10573
rect 16803 10508 16804 10572
rect 16868 10508 16869 10572
rect 16803 10507 16869 10508
rect 16619 10164 16685 10165
rect 16619 10100 16620 10164
rect 16684 10100 16685 10164
rect 16619 10099 16685 10100
rect 16622 8805 16682 10099
rect 16619 8804 16685 8805
rect 16619 8740 16620 8804
rect 16684 8740 16685 8804
rect 16619 8739 16685 8740
rect 16619 8396 16685 8397
rect 16619 8332 16620 8396
rect 16684 8332 16685 8396
rect 16619 8331 16685 8332
rect 16435 3908 16501 3909
rect 16435 3844 16436 3908
rect 16500 3844 16501 3908
rect 16435 3843 16501 3844
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15331 2684 15397 2685
rect 15331 2620 15332 2684
rect 15396 2620 15397 2684
rect 15331 2619 15397 2620
rect 15770 2208 16090 3232
rect 16622 2685 16682 8331
rect 16806 4045 16866 10507
rect 16803 4044 16869 4045
rect 16803 3980 16804 4044
rect 16868 3980 16869 4044
rect 16803 3979 16869 3980
rect 16619 2684 16685 2685
rect 16619 2620 16620 2684
rect 16684 2620 16685 2684
rect 16619 2619 16685 2620
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 15770 2128 16090 2144
use sky130_fd_sc_hd__fill_1  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1606821651
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1472 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1564 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_10 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2024 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11
timestamp 1606821651
transform 1 0 2116 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_20
timestamp 1606821651
transform 1 0 2944 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19
timestamp 1606821651
transform 1 0 2852 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2392 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _26_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2484 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1606821651
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 3312 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _27_
timestamp 1606821651
transform 1 0 3220 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1606821651
transform 1 0 3864 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 4232 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _30_
timestamp 1606821651
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_40
timestamp 1606821651
transform 1 0 4784 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36
timestamp 1606821651
transform 1 0 4416 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1606821651
transform 1 0 4784 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_49
timestamp 1606821651
transform 1 0 5612 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_44
timestamp 1606821651
transform 1 0 5152 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 5152 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1606821651
transform 1 0 5244 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1606821651
transform 1 0 6348 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58
timestamp 1606821651
transform 1 0 6440 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52
timestamp 1606821651
transform 1 0 5888 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1606821651
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1606821651
transform 1 0 5980 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1606821651
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1606821651
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 8004 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 8648 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1606821651
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1606821651
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72
timestamp 1606821651
transform 1 0 7728 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_71
timestamp 1606821651
transform 1 0 7636 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_78
timestamp 1606821651
transform 1 0 8280 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606821651
transform 1 0 10212 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606821651
transform 1 0 10120 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1606821651
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1606821651
transform 1 0 8924 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1606821651
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_95
timestamp 1606821651
transform 1 0 9844 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_112
timestamp 1606821651
transform 1 0 11408 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_111
timestamp 1606821651
transform 1 0 11316 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1606821651
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1606821651
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1606821651
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115
timestamp 1606821651
transform 1 0 11684 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1606821651
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1606821651
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1606821651
transform 1 0 11776 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606821651
transform 1 0 12420 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1606821651
transform 1 0 12972 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1606821651
transform 1 0 13984 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606821651
transform 1 0 13708 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_0_133
timestamp 1606821651
transform 1 0 13340 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_136
timestamp 1606821651
transform 1 0 13616 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1606821651
transform 1 0 16008 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606821651
transform 1 0 15548 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1606821651
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_150
timestamp 1606821651
transform 1 0 14904 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154
timestamp 1606821651
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_156 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 15456 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_166
timestamp 1606821651
transform 1 0 16376 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_153
timestamp 1606821651
transform 1 0 15180 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_170
timestamp 1606821651
transform 1 0 16744 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1606821651
transform 1 0 16744 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_179
timestamp 1606821651
transform 1 0 17572 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_174
timestamp 1606821651
transform 1 0 17112 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_174
timestamp 1606821651
transform 1 0 17112 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1606821651
transform 1 0 17480 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1606821651
transform 1 0 17204 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_184
timestamp 1606821651
transform 1 0 18032 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp 1606821651
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1606821651
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1606821651
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1606821651
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606821651
transform -1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606821651
transform -1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _28_
timestamp 1606821651
transform 1 0 1656 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01
timestamp 1606821651
transform 1 0 2668 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606821651
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1606821651
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_10
timestamp 1606821651
transform 1 0 2024 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_16
timestamp 1606821651
transform 1 0 2576 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 4048 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1606821651
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_23
timestamp 1606821651
transform 1 0 3220 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5888 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_48
timestamp 1606821651
transform 1 0 5520 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _09_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 7728 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1606821651
transform 1 0 8372 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_68
timestamp 1606821651
transform 1 0 7360 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_75
timestamp 1606821651
transform 1 0 8004 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1606821651
transform 1 0 10028 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1606821651
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_88
timestamp 1606821651
transform 1 0 9200 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_93
timestamp 1606821651
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1606821651
transform 1 0 11224 0 -1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_2_106
timestamp 1606821651
transform 1 0 10856 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_123
timestamp 1606821651
transform 1 0 12420 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1606821651
transform 1 0 14444 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1606821651
transform 1 0 12788 0 -1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_2_140
timestamp 1606821651
transform 1 0 13984 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_144
timestamp 1606821651
transform 1 0 14352 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1606821651
transform 1 0 15272 0 -1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1606821651
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1606821651
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 16836 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_167
timestamp 1606821651
transform 1 0 16468 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_180
timestamp 1606821651
transform 1 0 17664 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606821651
transform -1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_188
timestamp 1606821651
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _22_
timestamp 1606821651
transform 1 0 1656 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _23_
timestamp 1606821651
transform 1 0 2392 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606821651
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1606821651
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_10
timestamp 1606821651
transform 1 0 2024 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_18
timestamp 1606821651
transform 1 0 2760 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _24_
timestamp 1606821651
transform 1 0 3128 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 3956 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_26
timestamp 1606821651
transform 1 0 3496 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_30
timestamp 1606821651
transform 1 0 3864 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_40
timestamp 1606821651
transform 1 0 4784 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6808 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1606821651
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1606821651
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_53
timestamp 1606821651
transform 1 0 5980 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_78
timestamp 1606821651
transform 1 0 8280 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1606821651
transform 1 0 9016 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10212 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_95
timestamp 1606821651
transform 1 0 9844 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1606821651
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_115
timestamp 1606821651
transform 1 0 11684 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1606821651
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_123
timestamp 1606821651
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1606821651
transform 1 0 12788 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1606821651
transform 1 0 14352 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_3_140
timestamp 1606821651
transform 1 0 13984 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606821651
transform 1 0 16008 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_3_157
timestamp 1606821651
transform 1 0 15548 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_161
timestamp 1606821651
transform 1 0 15916 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1606821651
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_175
timestamp 1606821651
transform 1 0 17204 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_184
timestamp 1606821651
transform 1 0 18032 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606821651
transform -1 0 18860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _20_
timestamp 1606821651
transform 1 0 1656 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1606821651
transform 1 0 2392 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606821651
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1606821651
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_10
timestamp 1606821651
transform 1 0 2024 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_18
timestamp 1606821651
transform 1 0 2760 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _25_
timestamp 1606821651
transform 1 0 3128 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4416 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1606821651
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_26
timestamp 1606821651
transform 1 0 3496 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_30
timestamp 1606821651
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1606821651
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1606821651
transform 1 0 5612 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_45
timestamp 1606821651
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_58
timestamp 1606821651
transform 1 0 6440 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_62
timestamp 1606821651
transform 1 0 6808 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1606821651
transform 1 0 6900 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7636 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_67
timestamp 1606821651
transform 1 0 7268 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _13_
timestamp 1606821651
transform 1 0 9660 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1606821651
transform 1 0 10304 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1606821651
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_87
timestamp 1606821651
transform 1 0 9108 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1606821651
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_96
timestamp 1606821651
transform 1 0 9936 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606821651
transform 1 0 11684 0 -1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_4_109
timestamp 1606821651
transform 1 0 11132 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606821651
transform 1 0 13616 0 -1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_4_128
timestamp 1606821651
transform 1 0 12880 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1606821651
transform 1 0 15272 0 -1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1606821651
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1606821651
transform 1 0 14812 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_2_
timestamp 1606821651
transform 1 0 16836 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_167
timestamp 1606821651
transform 1 0 16468 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_180
timestamp 1606821651
transform 1 0 17664 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606821651
transform -1 0 18860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_188
timestamp 1606821651
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _19_
timestamp 1606821651
transform 1 0 1656 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2576 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606821651
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 1606821651
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_10
timestamp 1606821651
transform 1 0 2024 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4876 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1606821651
transform 1 0 3680 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_22
timestamp 1606821651
transform 1 0 3128 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_37
timestamp 1606821651
transform 1 0 4508 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1606821651
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1606821651
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1606821651
transform 1 0 6348 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 8096 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_71
timestamp 1606821651
transform 1 0 7636 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_75
timestamp 1606821651
transform 1 0 8004 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10120 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_5_92
timestamp 1606821651
transform 1 0 9568 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1606821651
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1606821651
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 11960 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_114
timestamp 1606821651
transform 1 0 11592 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1606821651
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1606821651
transform 1 0 13156 0 1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_5_127
timestamp 1606821651
transform 1 0 12788 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_144
timestamp 1606821651
transform 1 0 14352 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1606821651
transform 1 0 14720 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1606821651
transform 1 0 15456 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_152
timestamp 1606821651
transform 1 0 15088 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_165
timestamp 1606821651
transform 1 0 16284 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1606821651
transform 1 0 16652 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1606821651
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_178
timestamp 1606821651
transform 1 0 17480 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1606821651
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_184
timestamp 1606821651
transform 1 0 18032 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606821651
transform -1 0 18860 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_10
timestamp 1606821651
transform 1 0 2024 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1606821651
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1606821651
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606821651
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606821651
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1748 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _18_
timestamp 1606821651
transform 1 0 1656 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_17
timestamp 1606821651
transform 1 0 2668 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_13
timestamp 1606821651
transform 1 0 2300 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1606821651
transform 1 0 2760 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 2392 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 4416 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606821651
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606821651
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_41
timestamp 1606821651
transform 1 0 4876 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_30
timestamp 1606821651
transform 1 0 3864 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1606821651
transform 1 0 5520 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6256 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1606821651
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606821651
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 6256 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_47
timestamp 1606821651
transform 1 0 5428 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_52
timestamp 1606821651
transform 1 0 5888 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1606821651
transform 1 0 5888 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1606821651
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1606821651
transform 1 0 8372 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8096 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_6_72
timestamp 1606821651
transform 1 0 7728 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_78
timestamp 1606821651
transform 1 0 8280 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_71
timestamp 1606821651
transform 1 0 7636 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_75
timestamp 1606821651
transform 1 0 8004 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9292 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606821651
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_88
timestamp 1606821651
transform 1 0 9200 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_85
timestamp 1606821651
transform 1 0 8924 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606821651
transform 1 0 11500 0 -1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1606821651
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1606821651
transform 1 0 11132 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606821651
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_109
timestamp 1606821651
transform 1 0 11132 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_105
timestamp 1606821651
transform 1 0 10764 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1606821651
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13064 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 14168 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_126
timestamp 1606821651
transform 1 0 12696 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_132
timestamp 1606821651
transform 1 0 13248 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_140
timestamp 1606821651
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1606821651
transform 1 0 15456 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1606821651
transform 1 0 16192 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1606821651
transform 1 0 16008 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606821651
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_146
timestamp 1606821651
transform 1 0 14536 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1606821651
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_154
timestamp 1606821651
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_160
timestamp 1606821651
transform 1 0 15824 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_158
timestamp 1606821651
transform 1 0 15640 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1606821651
transform 1 0 17204 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1606821651
transform 1 0 17388 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606821651
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_173
timestamp 1606821651
transform 1 0 17020 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_186
timestamp 1606821651
transform 1 0 18216 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_171
timestamp 1606821651
transform 1 0 16836 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_179
timestamp 1606821651
transform 1 0 17572 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_184
timestamp 1606821651
transform 1 0 18032 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606821651
transform -1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606821651
transform -1 0 18860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1606821651
transform 1 0 2760 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1606821651
transform 1 0 1564 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606821651
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1606821651
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_14
timestamp 1606821651
transform 1 0 2392 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4048 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606821651
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606821651
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1606821651
transform 1 0 5888 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_48
timestamp 1606821651
transform 1 0 5520 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_61
timestamp 1606821651
transform 1 0 6716 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1606821651
transform 1 0 7084 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1606821651
transform 1 0 8280 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_74
timestamp 1606821651
transform 1 0 7912 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _14_
timestamp 1606821651
transform 1 0 9660 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_1_
timestamp 1606821651
transform 1 0 10304 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606821651
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_87
timestamp 1606821651
transform 1 0 9108 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1606821651
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_96
timestamp 1606821651
transform 1 0 9936 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 11500 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_109
timestamp 1606821651
transform 1 0 11132 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _15_
timestamp 1606821651
transform 1 0 13340 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13984 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_129
timestamp 1606821651
transform 1 0 12972 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1606821651
transform 1 0 13616 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1606821651
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606821651
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1606821651
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_163
timestamp 1606821651
transform 1 0 16100 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1606821651
transform 1 0 17848 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16652 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_178
timestamp 1606821651
transform 1 0 17480 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_186
timestamp 1606821651
transform 1 0 18216 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606821651
transform -1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _29_
timestamp 1606821651
transform 1 0 1472 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1606821651
transform 1 0 2208 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606821651
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1606821651
transform 1 0 1380 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_8
timestamp 1606821651
transform 1 0 1840 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1606821651
transform 1 0 3404 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1606821651
transform 1 0 4232 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_21
timestamp 1606821651
transform 1 0 3036 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_29
timestamp 1606821651
transform 1 0 3772 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_33
timestamp 1606821651
transform 1 0 4140 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5428 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606821651
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_43
timestamp 1606821651
transform 1 0 5060 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_56
timestamp 1606821651
transform 1 0 6256 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1606821651
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1606821651
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 8372 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1606821651
transform 1 0 7176 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_75
timestamp 1606821651
transform 1 0 8004 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 10396 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_9_95
timestamp 1606821651
transform 1 0 9844 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1606821651
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606821651
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_117
timestamp 1606821651
transform 1 0 11868 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1606821651
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 13708 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_132
timestamp 1606821651
transform 1 0 13248 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_136
timestamp 1606821651
transform 1 0 13616 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 15548 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_153
timestamp 1606821651
transform 1 0 15180 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606821651
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_173
timestamp 1606821651
transform 1 0 17020 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1606821651
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_184
timestamp 1606821651
transform 1 0 18032 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606821651
transform -1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _31_
timestamp 1606821651
transform 1 0 1656 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1606821651
transform 1 0 2668 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606821651
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1606821651
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_10
timestamp 1606821651
transform 1 0 2024 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_16
timestamp 1606821651
transform 1 0 2576 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_2_
timestamp 1606821651
transform 1 0 4508 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606821651
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_26
timestamp 1606821651
transform 1 0 3496 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_30
timestamp 1606821651
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_32
timestamp 1606821651
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_36
timestamp 1606821651
transform 1 0 4416 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 5704 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_46
timestamp 1606821651
transform 1 0 5336 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1606821651
transform 1 0 8740 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1606821651
transform 1 0 7544 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_66
timestamp 1606821651
transform 1 0 7176 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_79
timestamp 1606821651
transform 1 0 8372 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 9660 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606821651
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_87
timestamp 1606821651
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1606821651
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1606821651
transform 1 0 11684 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_10_109
timestamp 1606821651
transform 1 0 11132 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_124
timestamp 1606821651
transform 1 0 12512 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1606821651
transform 1 0 14444 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1606821651
transform 1 0 12880 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 14076 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_137
timestamp 1606821651
transform 1 0 13708 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_144
timestamp 1606821651
transform 1 0 14352 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1606821651
transform 1 0 15456 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606821651
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_149
timestamp 1606821651
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_154
timestamp 1606821651
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_165
timestamp 1606821651
transform 1 0 16284 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1606821651
transform 1 0 17848 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1606821651
transform 1 0 16652 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_178
timestamp 1606821651
transform 1 0 17480 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_186
timestamp 1606821651
transform 1 0 18216 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606821651
transform -1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1606821651
transform 1 0 1840 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606821651
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1606821651
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 1606821651
transform 1 0 1748 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_17
timestamp 1606821651
transform 1 0 2668 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4232 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1606821651
transform 1 0 3036 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_30
timestamp 1606821651
transform 1 0 3864 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1606821651
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_1_
timestamp 1606821651
transform 1 0 5428 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606821651
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_43
timestamp 1606821651
transform 1 0 5060 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_56
timestamp 1606821651
transform 1 0 6256 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1606821651
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1606821651
transform 1 0 7360 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 8556 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_11_66
timestamp 1606821651
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_77
timestamp 1606821651
transform 1 0 8188 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10396 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606821651
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_117
timestamp 1606821651
transform 1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1606821651
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1606821651
transform 1 0 13800 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_134
timestamp 1606821651
transform 1 0 13432 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_142
timestamp 1606821651
transform 1 0 14168 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 14536 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_162
timestamp 1606821651
transform 1 0 16008 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606821651
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_175
timestamp 1606821651
transform 1 0 17204 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_184
timestamp 1606821651
transform 1 0 18032 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606821651
transform -1 0 18860 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 1564 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606821651
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1606821651
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 4048 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606821651
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_21
timestamp 1606821651
transform 1 0 3036 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1606821651
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5888 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_48
timestamp 1606821651
transform 1 0 5520 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_61
timestamp 1606821651
transform 1 0 6716 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1606821651
transform 1 0 7084 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8372 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_74
timestamp 1606821651
transform 1 0 7912 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_78
timestamp 1606821651
transform 1 0 8280 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1606821651
transform 1 0 10488 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_2_
timestamp 1606821651
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606821651
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1606821651
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10948 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_12_106
timestamp 1606821651
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_123
timestamp 1606821651
transform 1 0 12420 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1606821651
transform 1 0 14444 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1606821651
transform 1 0 12972 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 14168 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_138
timestamp 1606821651
transform 1 0 13800 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15272 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606821651
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1606821651
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1606821651
transform 1 0 17112 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_170
timestamp 1606821651
transform 1 0 16744 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_183
timestamp 1606821651
transform 1 0 17940 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606821651
transform -1 0 18860 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_189
timestamp 1606821651
transform 1 0 18492 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 1840 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_1_
timestamp 1606821651
transform 1 0 2760 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1606821651
transform 1 0 1564 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606821651
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606821651
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1606821651
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1606821651
transform 1 0 1748 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1606821651
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_14
timestamp 1606821651
transform 1 0 2392 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1606821651
transform 1 0 3680 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606821651
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_24
timestamp 1606821651
transform 1 0 3312 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_37
timestamp 1606821651
transform 1 0 4508 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_41
timestamp 1606821651
transform 1 0 4876 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1606821651
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_41
timestamp 1606821651
transform 1 0 4876 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_45
timestamp 1606821651
transform 1 0 5244 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 4968 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1606821651
transform 1 0 5244 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5336 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_55
timestamp 1606821651
transform 1 0 6164 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_54
timestamp 1606821651
transform 1 0 6072 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 6440 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606821651
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 6532 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_62
timestamp 1606821651
transform 1 0 6808 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7544 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6900 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8740 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_79
timestamp 1606821651
transform 1 0 8372 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_65
timestamp 1606821651
transform 1 0 7084 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_69
timestamp 1606821651
transform 1 0 7452 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9752 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1606821651
transform 1 0 9844 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606821651
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_92
timestamp 1606821651
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_103
timestamp 1606821651
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_86
timestamp 1606821651
transform 1 0 9016 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1606821651
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_104
timestamp 1606821651
transform 1 0 10672 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1606821651
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1606821651
transform 1 0 12236 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1606821651
transform 1 0 11040 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606821651
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_114
timestamp 1606821651
transform 1 0 11592 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_117
timestamp 1606821651
transform 1 0 11868 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 14168 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1606821651
transform 1 0 13432 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_132
timestamp 1606821651
transform 1 0 13248 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_140
timestamp 1606821651
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_130
timestamp 1606821651
transform 1 0 13064 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_143
timestamp 1606821651
transform 1 0 14260 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1606821651
transform 1 0 16008 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 15364 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606821651
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_158
timestamp 1606821651
transform 1 0 15640 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_166
timestamp 1606821651
transform 1 0 16376 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1606821651
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_154
timestamp 1606821651
transform 1 0 15272 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1606821651
transform 1 0 16744 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1606821651
transform 1 0 17204 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606821651
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_179
timestamp 1606821651
transform 1 0 17572 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_184
timestamp 1606821651
transform 1 0 18032 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_171
timestamp 1606821651
transform 1 0 16836 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_184
timestamp 1606821651
transform 1 0 18032 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606821651
transform -1 0 18860 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606821651
transform -1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1606821651
transform 1 0 1656 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 2392 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606821651
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1606821651
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_10
timestamp 1606821651
transform 1 0 2024 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1606821651
transform 1 0 4600 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_30
timestamp 1606821651
transform 1 0 3864 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1606821651
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 5796 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606821651
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_47
timestamp 1606821651
transform 1 0 5428 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1606821651
transform 1 0 6348 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1606821651
transform 1 0 8004 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_71
timestamp 1606821651
transform 1 0 7636 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_79
timestamp 1606821651
transform 1 0 8372 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 8924 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_101
timestamp 1606821651
transform 1 0 10396 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1606821651
transform 1 0 10764 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606821651
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_114
timestamp 1606821651
transform 1 0 11592 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13800 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_15_132
timestamp 1606821651
transform 1 0 13248 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1606821651
transform 1 0 16008 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_154
timestamp 1606821651
transform 1 0 15272 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_166
timestamp 1606821651
transform 1 0 16376 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1606821651
transform 1 0 16744 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606821651
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_179
timestamp 1606821651
transform 1 0 17572 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_184
timestamp 1606821651
transform 1 0 18032 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606821651
transform -1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_2_
timestamp 1606821651
transform 1 0 2668 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1606821651
transform 1 0 1472 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606821651
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1606821651
transform 1 0 1380 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_13
timestamp 1606821651
transform 1 0 2300 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4324 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606821651
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_26
timestamp 1606821651
transform 1 0 3496 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1606821651
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_32
timestamp 1606821651
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1606821651
transform 1 0 6808 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1606821651
transform 1 0 5520 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_44
timestamp 1606821651
transform 1 0 5152 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_57
timestamp 1606821651
transform 1 0 6348 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_61
timestamp 1606821651
transform 1 0 6716 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 7544 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_66
timestamp 1606821651
transform 1 0 7176 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1606821651
transform 1 0 9936 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 10580 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606821651
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_86
timestamp 1606821651
transform 1 0 9016 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_16_93
timestamp 1606821651
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_99
timestamp 1606821651
transform 1 0 10212 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 12604 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_16_119
timestamp 1606821651
transform 1 0 12052 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1606821651
transform 1 0 14444 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1606821651
transform 1 0 14076 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1606821651
transform 1 0 15732 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606821651
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1606821651
transform 1 0 14812 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_154
timestamp 1606821651
transform 1 0 15272 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_158
timestamp 1606821651
transform 1 0 15640 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1606821651
transform 1 0 16928 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_168
timestamp 1606821651
transform 1 0 16560 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_181
timestamp 1606821651
transform 1 0 17756 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606821651
transform -1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_189
timestamp 1606821651
transform 1 0 18492 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1606821651
transform 1 0 1564 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1606821651
transform 1 0 2300 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606821651
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1606821651
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_9
timestamp 1606821651
transform 1 0 1932 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 3496 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_22
timestamp 1606821651
transform 1 0 3128 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 6808 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1606821651
transform 1 0 5520 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606821651
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_42
timestamp 1606821651
transform 1 0 4968 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1606821651
transform 1 0 6348 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1606821651
transform 1 0 8740 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_78
timestamp 1606821651
transform 1 0 8280 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_82
timestamp 1606821651
transform 1 0 8648 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_92 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 9568 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_104
timestamp 1606821651
transform 1 0 10672 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1606821651
transform 1 0 11132 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606821651
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_108
timestamp 1606821651
transform 1 0 11040 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_112
timestamp 1606821651
transform 1 0 11408 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1606821651
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_123
timestamp 1606821651
transform 1 0 12420 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1606821651
transform 1 0 14352 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12972 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_17_138
timestamp 1606821651
transform 1 0 13800 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1606821651
transform 1 0 15088 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_148
timestamp 1606821651
transform 1 0 14720 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1606821651
transform 1 0 15916 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1606821651
transform 1 0 17204 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1606821651
transform 1 0 16468 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606821651
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_171
timestamp 1606821651
transform 1 0 16836 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_179
timestamp 1606821651
transform 1 0 17572 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_184
timestamp 1606821651
transform 1 0 18032 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606821651
transform -1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1606821651
transform 1 0 1472 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1606821651
transform 1 0 2208 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606821651
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1606821651
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_8
timestamp 1606821651
transform 1 0 1840 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4508 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606821651
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_21
timestamp 1606821651
transform 1 0 3036 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1606821651
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_32
timestamp 1606821651
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_36
timestamp 1606821651
transform 1 0 4416 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6348 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_53
timestamp 1606821651
transform 1 0 5980 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1606821651
transform 1 0 8188 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_73
timestamp 1606821651
transform 1 0 7820 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606821651
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_86
timestamp 1606821651
transform 1 0 9016 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1606821651
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1606821651
transform 1 0 12236 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1606821651
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_117
timestamp 1606821651
transform 1 0 11868 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_124
timestamp 1606821651
transform 1 0 12512 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1606821651
transform 1 0 13248 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1606821651
transform 1 0 14168 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_135
timestamp 1606821651
transform 1 0 13524 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_141
timestamp 1606821651
transform 1 0 14076 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_145
timestamp 1606821651
transform 1 0 14444 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1606821651
transform 1 0 16376 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1606821651
transform 1 0 15548 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606821651
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_154
timestamp 1606821651
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_161
timestamp 1606821651
transform 1 0 15916 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_165
timestamp 1606821651
transform 1 0 16284 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1606821651
transform 1 0 17848 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1606821651
transform 1 0 17112 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_170
timestamp 1606821651
transform 1 0 16744 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_178
timestamp 1606821651
transform 1 0 17480 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_186
timestamp 1606821651
transform 1 0 18216 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606821651
transform -1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_8
timestamp 1606821651
transform 1 0 1840 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1606821651
transform 1 0 1380 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 1606821651
transform 1 0 1380 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606821651
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606821651
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1606821651
transform 1 0 1472 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1606821651
transform 1 0 1472 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_13
timestamp 1606821651
transform 1 0 2300 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1606821651
transform 1 0 2208 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 2668 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _10_
timestamp 1606821651
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _11_
timestamp 1606821651
transform 1 0 4508 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606821651
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_33
timestamp 1606821651
transform 1 0 4140 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_40
timestamp 1606821651
transform 1 0 4784 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_21
timestamp 1606821651
transform 1 0 3036 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1606821651
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_35
timestamp 1606821651
transform 1 0 4324 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _12_
timestamp 1606821651
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1606821651
transform 1 0 5520 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606821651
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1606821651
transform 1 0 6348 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_47
timestamp 1606821651
transform 1 0 5428 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_59
timestamp 1606821651
transform 1 0 6532 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 7820 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_65
timestamp 1606821651
transform 1 0 7084 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_71
timestamp 1606821651
transform 1 0 7636 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_83
timestamp 1606821651
transform 1 0 8740 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606821651
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_85
timestamp 1606821651
transform 1 0 8924 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_97
timestamp 1606821651
transform 1 0 10028 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1606821651
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1606821651
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1606821651
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606821651
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_109
timestamp 1606821651
transform 1 0 11132 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1606821651
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1606821651
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1606821651
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1606821651
transform 1 0 13064 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_126
timestamp 1606821651
transform 1 0 12696 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_133
timestamp 1606821651
transform 1 0 13340 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_145
timestamp 1606821651
transform 1 0 14444 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1606821651
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1606821651
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1606821651
transform 1 0 16192 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1606821651
transform 1 0 15180 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1606821651
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606821651
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_156
timestamp 1606821651
transform 1 0 15456 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_157
timestamp 1606821651
transform 1 0 15548 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_169
timestamp 1606821651
transform 1 0 16652 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_168
timestamp 1606821651
transform 1 0 16560 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_178
timestamp 1606821651
transform 1 0 17480 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_179
timestamp 1606821651
transform 1 0 17572 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_174
timestamp 1606821651
transform 1 0 17112 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1606821651
transform 1 0 17204 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1606821651
transform 1 0 17204 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_186
timestamp 1606821651
transform 1 0 18216 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_184
timestamp 1606821651
transform 1 0 18032 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606821651
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1606821651
transform 1 0 17848 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606821651
transform -1 0 18860 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606821651
transform -1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1606821651
transform 1 0 1564 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606821651
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1606821651
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_14
timestamp 1606821651
transform 1 0 2392 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1606821651
transform 1 0 3128 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_26
timestamp 1606821651
transform 1 0 3496 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_38
timestamp 1606821651
transform 1 0 4600 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1606821651
transform 1 0 5980 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1606821651
transform 1 0 6808 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606821651
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_50
timestamp 1606821651
transform 1 0 5704 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1606821651
transform 1 0 6348 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_66
timestamp 1606821651
transform 1 0 7176 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_78
timestamp 1606821651
transform 1 0 8280 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_90
timestamp 1606821651
transform 1 0 9384 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_102
timestamp 1606821651
transform 1 0 10488 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606821651
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_114
timestamp 1606821651
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_123
timestamp 1606821651
transform 1 0 12420 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1606821651
transform 1 0 13432 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1606821651
transform 1 0 14444 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_131
timestamp 1606821651
transform 1 0 13156 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_138
timestamp 1606821651
transform 1 0 13800 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_144
timestamp 1606821651
transform 1 0 14352 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1606821651
transform 1 0 15548 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_149
timestamp 1606821651
transform 1 0 14812 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_161
timestamp 1606821651
transform 1 0 15916 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606821651
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_173
timestamp 1606821651
transform 1 0 17020 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1606821651
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_184
timestamp 1606821651
transform 1 0 18032 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606821651
transform -1 0 18860 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1606821651
transform 1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1606821651
transform 1 0 2484 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606821651
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1606821651
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_11
timestamp 1606821651
transform 1 0 2116 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_19
timestamp 1606821651
transform 1 0 2852 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1606821651
transform 1 0 3220 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606821651
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1606821651
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1606821651
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606821651
transform 1 0 6808 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1606821651
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_56
timestamp 1606821651
transform 1 0 6256 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_63
timestamp 1606821651
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_75
timestamp 1606821651
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606821651
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_87
timestamp 1606821651
transform 1 0 9108 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_94
timestamp 1606821651
transform 1 0 9752 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606821651
transform 1 0 12512 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_106
timestamp 1606821651
transform 1 0 10856 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_118
timestamp 1606821651
transform 1 0 11960 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_125
timestamp 1606821651
transform 1 0 12604 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_137
timestamp 1606821651
transform 1 0 13708 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1606821651
transform 1 0 15456 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606821651
transform 1 0 15364 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_149
timestamp 1606821651
transform 1 0 14812 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_160
timestamp 1606821651
transform 1 0 15824 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606821651
transform 1 0 18216 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_172
timestamp 1606821651
transform 1 0 16928 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_184
timestamp 1606821651
transform 1 0 18032 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_187
timestamp 1606821651
transform 1 0 18308 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606821651
transform -1 0 18860 0 -1 14688
box -38 -48 314 592
<< labels >>
rlabel metal2 s 7378 16520 7434 17000 6 IO_ISOL_N
port 0 nsew default input
rlabel metal2 s 5630 0 5686 480 6 SC_IN_BOT
port 1 nsew default input
rlabel metal2 s 6090 16520 6146 17000 6 SC_IN_TOP
port 2 nsew default input
rlabel metal2 s 6182 0 6238 480 6 SC_OUT_BOT
port 3 nsew default tristate
rlabel metal2 s 6734 16520 6790 17000 6 SC_OUT_TOP
port 4 nsew default tristate
rlabel metal2 s 202 0 258 480 6 bottom_grid_pin_0_
port 5 nsew default tristate
rlabel metal2 s 2686 0 2742 480 6 bottom_grid_pin_10_
port 6 nsew default tristate
rlabel metal2 s 3146 0 3202 480 6 bottom_grid_pin_12_
port 7 nsew default tristate
rlabel metal2 s 3606 0 3662 480 6 bottom_grid_pin_14_
port 8 nsew default tristate
rlabel metal2 s 4158 0 4214 480 6 bottom_grid_pin_16_
port 9 nsew default tristate
rlabel metal2 s 662 0 718 480 6 bottom_grid_pin_2_
port 10 nsew default tristate
rlabel metal2 s 1122 0 1178 480 6 bottom_grid_pin_4_
port 11 nsew default tristate
rlabel metal2 s 1674 0 1730 480 6 bottom_grid_pin_6_
port 12 nsew default tristate
rlabel metal2 s 2134 0 2190 480 6 bottom_grid_pin_8_
port 13 nsew default tristate
rlabel metal2 s 4618 0 4674 480 6 ccff_head
port 14 nsew default input
rlabel metal2 s 5170 0 5226 480 6 ccff_tail
port 15 nsew default tristate
rlabel metal3 s 0 8848 480 8968 6 chanx_left_in[0]
port 16 nsew default input
rlabel metal3 s 0 12928 480 13048 6 chanx_left_in[10]
port 17 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_left_in[11]
port 18 nsew default input
rlabel metal3 s 0 13744 480 13864 6 chanx_left_in[12]
port 19 nsew default input
rlabel metal3 s 0 14152 480 14272 6 chanx_left_in[13]
port 20 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[14]
port 21 nsew default input
rlabel metal3 s 0 14968 480 15088 6 chanx_left_in[15]
port 22 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chanx_left_in[16]
port 23 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[17]
port 24 nsew default input
rlabel metal3 s 0 16192 480 16312 6 chanx_left_in[18]
port 25 nsew default input
rlabel metal3 s 0 16600 480 16720 6 chanx_left_in[19]
port 26 nsew default input
rlabel metal3 s 0 9256 480 9376 6 chanx_left_in[1]
port 27 nsew default input
rlabel metal3 s 0 9664 480 9784 6 chanx_left_in[2]
port 28 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[3]
port 29 nsew default input
rlabel metal3 s 0 10480 480 10600 6 chanx_left_in[4]
port 30 nsew default input
rlabel metal3 s 0 10888 480 11008 6 chanx_left_in[5]
port 31 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[6]
port 32 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[7]
port 33 nsew default input
rlabel metal3 s 0 12112 480 12232 6 chanx_left_in[8]
port 34 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[9]
port 35 nsew default input
rlabel metal3 s 0 552 480 672 6 chanx_left_out[0]
port 36 nsew default tristate
rlabel metal3 s 0 4632 480 4752 6 chanx_left_out[10]
port 37 nsew default tristate
rlabel metal3 s 0 5040 480 5160 6 chanx_left_out[11]
port 38 nsew default tristate
rlabel metal3 s 0 5448 480 5568 6 chanx_left_out[12]
port 39 nsew default tristate
rlabel metal3 s 0 5856 480 5976 6 chanx_left_out[13]
port 40 nsew default tristate
rlabel metal3 s 0 6264 480 6384 6 chanx_left_out[14]
port 41 nsew default tristate
rlabel metal3 s 0 6672 480 6792 6 chanx_left_out[15]
port 42 nsew default tristate
rlabel metal3 s 0 7080 480 7200 6 chanx_left_out[16]
port 43 nsew default tristate
rlabel metal3 s 0 7488 480 7608 6 chanx_left_out[17]
port 44 nsew default tristate
rlabel metal3 s 0 7896 480 8016 6 chanx_left_out[18]
port 45 nsew default tristate
rlabel metal3 s 0 8304 480 8424 6 chanx_left_out[19]
port 46 nsew default tristate
rlabel metal3 s 0 960 480 1080 6 chanx_left_out[1]
port 47 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[2]
port 48 nsew default tristate
rlabel metal3 s 0 1776 480 1896 6 chanx_left_out[3]
port 49 nsew default tristate
rlabel metal3 s 0 2184 480 2304 6 chanx_left_out[4]
port 50 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 chanx_left_out[5]
port 51 nsew default tristate
rlabel metal3 s 0 3000 480 3120 6 chanx_left_out[6]
port 52 nsew default tristate
rlabel metal3 s 0 3408 480 3528 6 chanx_left_out[7]
port 53 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_out[8]
port 54 nsew default tristate
rlabel metal3 s 0 4224 480 4344 6 chanx_left_out[9]
port 55 nsew default tristate
rlabel metal3 s 19520 8576 20000 8696 6 chanx_right_in[0]
port 56 nsew default input
rlabel metal3 s 19520 12792 20000 12912 6 chanx_right_in[10]
port 57 nsew default input
rlabel metal3 s 19520 13200 20000 13320 6 chanx_right_in[11]
port 58 nsew default input
rlabel metal3 s 19520 13744 20000 13864 6 chanx_right_in[12]
port 59 nsew default input
rlabel metal3 s 19520 14152 20000 14272 6 chanx_right_in[13]
port 60 nsew default input
rlabel metal3 s 19520 14560 20000 14680 6 chanx_right_in[14]
port 61 nsew default input
rlabel metal3 s 19520 14968 20000 15088 6 chanx_right_in[15]
port 62 nsew default input
rlabel metal3 s 19520 15376 20000 15496 6 chanx_right_in[16]
port 63 nsew default input
rlabel metal3 s 19520 15784 20000 15904 6 chanx_right_in[17]
port 64 nsew default input
rlabel metal3 s 19520 16192 20000 16312 6 chanx_right_in[18]
port 65 nsew default input
rlabel metal3 s 19520 16600 20000 16720 6 chanx_right_in[19]
port 66 nsew default input
rlabel metal3 s 19520 8984 20000 9104 6 chanx_right_in[1]
port 67 nsew default input
rlabel metal3 s 19520 9392 20000 9512 6 chanx_right_in[2]
port 68 nsew default input
rlabel metal3 s 19520 9800 20000 9920 6 chanx_right_in[3]
port 69 nsew default input
rlabel metal3 s 19520 10344 20000 10464 6 chanx_right_in[4]
port 70 nsew default input
rlabel metal3 s 19520 10752 20000 10872 6 chanx_right_in[5]
port 71 nsew default input
rlabel metal3 s 19520 11160 20000 11280 6 chanx_right_in[6]
port 72 nsew default input
rlabel metal3 s 19520 11568 20000 11688 6 chanx_right_in[7]
port 73 nsew default input
rlabel metal3 s 19520 11976 20000 12096 6 chanx_right_in[8]
port 74 nsew default input
rlabel metal3 s 19520 12384 20000 12504 6 chanx_right_in[9]
port 75 nsew default input
rlabel metal3 s 19520 144 20000 264 6 chanx_right_out[0]
port 76 nsew default tristate
rlabel metal3 s 19520 4360 20000 4480 6 chanx_right_out[10]
port 77 nsew default tristate
rlabel metal3 s 19520 4768 20000 4888 6 chanx_right_out[11]
port 78 nsew default tristate
rlabel metal3 s 19520 5176 20000 5296 6 chanx_right_out[12]
port 79 nsew default tristate
rlabel metal3 s 19520 5584 20000 5704 6 chanx_right_out[13]
port 80 nsew default tristate
rlabel metal3 s 19520 5992 20000 6112 6 chanx_right_out[14]
port 81 nsew default tristate
rlabel metal3 s 19520 6400 20000 6520 6 chanx_right_out[15]
port 82 nsew default tristate
rlabel metal3 s 19520 6944 20000 7064 6 chanx_right_out[16]
port 83 nsew default tristate
rlabel metal3 s 19520 7352 20000 7472 6 chanx_right_out[17]
port 84 nsew default tristate
rlabel metal3 s 19520 7760 20000 7880 6 chanx_right_out[18]
port 85 nsew default tristate
rlabel metal3 s 19520 8168 20000 8288 6 chanx_right_out[19]
port 86 nsew default tristate
rlabel metal3 s 19520 552 20000 672 6 chanx_right_out[1]
port 87 nsew default tristate
rlabel metal3 s 19520 960 20000 1080 6 chanx_right_out[2]
port 88 nsew default tristate
rlabel metal3 s 19520 1368 20000 1488 6 chanx_right_out[3]
port 89 nsew default tristate
rlabel metal3 s 19520 1776 20000 1896 6 chanx_right_out[4]
port 90 nsew default tristate
rlabel metal3 s 19520 2184 20000 2304 6 chanx_right_out[5]
port 91 nsew default tristate
rlabel metal3 s 19520 2592 20000 2712 6 chanx_right_out[6]
port 92 nsew default tristate
rlabel metal3 s 19520 3000 20000 3120 6 chanx_right_out[7]
port 93 nsew default tristate
rlabel metal3 s 19520 3544 20000 3664 6 chanx_right_out[8]
port 94 nsew default tristate
rlabel metal3 s 19520 3952 20000 4072 6 chanx_right_out[9]
port 95 nsew default tristate
rlabel metal2 s 6642 0 6698 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
port 96 nsew default tristate
rlabel metal2 s 7102 0 7158 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
port 97 nsew default tristate
rlabel metal2 s 7654 0 7710 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
port 98 nsew default tristate
rlabel metal2 s 8114 0 8170 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
port 99 nsew default tristate
rlabel metal2 s 8666 0 8722 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
port 100 nsew default tristate
rlabel metal2 s 9126 0 9182 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
port 101 nsew default tristate
rlabel metal2 s 9678 0 9734 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
port 102 nsew default tristate
rlabel metal2 s 10138 0 10194 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
port 103 nsew default tristate
rlabel metal2 s 10598 0 10654 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
port 104 nsew default tristate
rlabel metal2 s 11150 0 11206 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
port 105 nsew default input
rlabel metal2 s 11610 0 11666 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
port 106 nsew default input
rlabel metal2 s 12162 0 12218 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
port 107 nsew default input
rlabel metal2 s 12622 0 12678 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
port 108 nsew default input
rlabel metal2 s 13174 0 13230 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
port 109 nsew default input
rlabel metal2 s 13634 0 13690 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
port 110 nsew default input
rlabel metal2 s 14094 0 14150 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
port 111 nsew default input
rlabel metal2 s 14646 0 14702 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
port 112 nsew default input
rlabel metal2 s 15106 0 15162 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
port 113 nsew default input
rlabel metal2 s 15658 0 15714 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
port 114 nsew default tristate
rlabel metal2 s 16118 0 16174 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
port 115 nsew default tristate
rlabel metal2 s 16670 0 16726 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
port 116 nsew default tristate
rlabel metal2 s 17130 0 17186 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
port 117 nsew default tristate
rlabel metal2 s 17590 0 17646 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
port 118 nsew default tristate
rlabel metal2 s 18142 0 18198 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
port 119 nsew default tristate
rlabel metal2 s 18602 0 18658 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
port 120 nsew default tristate
rlabel metal2 s 19154 0 19210 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
port 121 nsew default tristate
rlabel metal2 s 19614 0 19670 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
port 122 nsew default tristate
rlabel metal2 s 8022 16520 8078 17000 6 prog_clk_0_N_in
port 123 nsew default input
rlabel metal3 s 0 144 480 264 6 prog_clk_0_W_out
port 124 nsew default tristate
rlabel metal2 s 8666 16520 8722 17000 6 top_width_0_height_0__pin_0_
port 125 nsew default input
rlabel metal2 s 11886 16520 11942 17000 6 top_width_0_height_0__pin_10_
port 126 nsew default input
rlabel metal2 s 14462 16520 14518 17000 6 top_width_0_height_0__pin_11_lower
port 127 nsew default tristate
rlabel metal2 s 3514 16520 3570 17000 6 top_width_0_height_0__pin_11_upper
port 128 nsew default tristate
rlabel metal2 s 12530 16520 12586 17000 6 top_width_0_height_0__pin_12_
port 129 nsew default input
rlabel metal2 s 15106 16520 15162 17000 6 top_width_0_height_0__pin_13_lower
port 130 nsew default tristate
rlabel metal2 s 4158 16520 4214 17000 6 top_width_0_height_0__pin_13_upper
port 131 nsew default tristate
rlabel metal2 s 13174 16520 13230 17000 6 top_width_0_height_0__pin_14_
port 132 nsew default input
rlabel metal2 s 15750 16520 15806 17000 6 top_width_0_height_0__pin_15_lower
port 133 nsew default tristate
rlabel metal2 s 4802 16520 4858 17000 6 top_width_0_height_0__pin_15_upper
port 134 nsew default tristate
rlabel metal2 s 13818 16520 13874 17000 6 top_width_0_height_0__pin_16_
port 135 nsew default input
rlabel metal2 s 16394 16520 16450 17000 6 top_width_0_height_0__pin_17_lower
port 136 nsew default tristate
rlabel metal2 s 5446 16520 5502 17000 6 top_width_0_height_0__pin_17_upper
port 137 nsew default tristate
rlabel metal2 s 17038 16520 17094 17000 6 top_width_0_height_0__pin_1_lower
port 138 nsew default tristate
rlabel metal2 s 294 16520 350 17000 6 top_width_0_height_0__pin_1_upper
port 139 nsew default tristate
rlabel metal2 s 9310 16520 9366 17000 6 top_width_0_height_0__pin_2_
port 140 nsew default input
rlabel metal2 s 17682 16520 17738 17000 6 top_width_0_height_0__pin_3_lower
port 141 nsew default tristate
rlabel metal2 s 938 16520 994 17000 6 top_width_0_height_0__pin_3_upper
port 142 nsew default tristate
rlabel metal2 s 9954 16520 10010 17000 6 top_width_0_height_0__pin_4_
port 143 nsew default input
rlabel metal2 s 18326 16520 18382 17000 6 top_width_0_height_0__pin_5_lower
port 144 nsew default tristate
rlabel metal2 s 1582 16520 1638 17000 6 top_width_0_height_0__pin_5_upper
port 145 nsew default tristate
rlabel metal2 s 10598 16520 10654 17000 6 top_width_0_height_0__pin_6_
port 146 nsew default input
rlabel metal2 s 18970 16520 19026 17000 6 top_width_0_height_0__pin_7_lower
port 147 nsew default tristate
rlabel metal2 s 2226 16520 2282 17000 6 top_width_0_height_0__pin_7_upper
port 148 nsew default tristate
rlabel metal2 s 11242 16520 11298 17000 6 top_width_0_height_0__pin_8_
port 149 nsew default input
rlabel metal2 s 19614 16520 19670 17000 6 top_width_0_height_0__pin_9_lower
port 150 nsew default tristate
rlabel metal2 s 2870 16520 2926 17000 6 top_width_0_height_0__pin_9_upper
port 151 nsew default tristate
rlabel metal4 s 3909 2128 4229 14736 6 VPWR
port 152 nsew default input
rlabel metal4 s 6875 2128 7195 14736 6 VGND
port 153 nsew default input
<< properties >>
string FIXED_BBOX 0 0 20000 17000
<< end >>
