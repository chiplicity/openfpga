VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_1__0_
  CLASS BLOCK ;
  FOREIGN sb_1__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 114.000 BY 114.000 ;
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.010 110.000 1.290 114.000 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_TOP
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.790 110.000 113.070 114.000 ;
    END
  END SC_OUT_TOP
  PIN Test_en_N_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 21.710 110.000 21.990 114.000 ;
    END
  END Test_en_N_out
  PIN Test_en_S_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END Test_en_S_in
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 4.000 103.320 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 21.120 114.000 21.720 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 44.920 114.000 45.520 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 46.960 114.000 47.560 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 49.680 114.000 50.280 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 51.720 114.000 52.320 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 53.760 114.000 54.360 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 56.480 114.000 57.080 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 58.520 114.000 59.120 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 61.240 114.000 61.840 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 63.280 114.000 63.880 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 66.000 114.000 66.600 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 23.840 114.000 24.440 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 25.880 114.000 26.480 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 28.600 114.000 29.200 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 30.640 114.000 31.240 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 33.360 114.000 33.960 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 35.400 114.000 36.000 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 37.440 114.000 38.040 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 40.160 114.000 40.760 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 42.200 114.000 42.800 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 68.040 114.000 68.640 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 91.160 114.000 91.760 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 93.880 114.000 94.480 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 95.920 114.000 96.520 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 98.640 114.000 99.240 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 100.680 114.000 101.280 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 102.720 114.000 103.320 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 105.440 114.000 106.040 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 107.480 114.000 108.080 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 110.200 114.000 110.800 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 112.240 114.000 112.840 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 70.080 114.000 70.680 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 72.800 114.000 73.400 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 74.840 114.000 75.440 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 77.560 114.000 78.160 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 79.600 114.000 80.200 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 82.320 114.000 82.920 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 84.360 114.000 84.960 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 86.400 114.000 87.000 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 89.120 114.000 89.720 ;
    END
  END chanx_right_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.150 110.000 28.430 114.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.310 110.000 49.590 114.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.610 110.000 51.890 114.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.450 110.000 53.730 114.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.750 110.000 56.030 114.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 110.000 58.330 114.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 110.000 60.170 114.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.190 110.000 62.470 114.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.030 110.000 64.310 114.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.330 110.000 66.610 114.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.170 110.000 68.450 114.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.450 110.000 30.730 114.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.290 110.000 32.570 114.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 110.000 34.870 114.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.890 110.000 37.170 114.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.730 110.000 39.010 114.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.030 110.000 41.310 114.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.870 110.000 43.150 114.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.170 110.000 45.450 114.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.470 110.000 47.750 114.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.470 110.000 70.750 114.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.630 110.000 91.910 114.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.930 110.000 94.210 114.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.770 110.000 96.050 114.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.070 110.000 98.350 114.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 99.910 110.000 100.190 114.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.210 110.000 102.490 114.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.510 110.000 104.790 114.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.350 110.000 106.630 114.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.650 110.000 108.930 114.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.490 110.000 110.770 114.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.770 110.000 73.050 114.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.610 110.000 74.890 114.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.910 110.000 77.190 114.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.750 110.000 79.030 114.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.050 110.000 81.330 114.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.350 110.000 83.630 114.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.190 110.000 85.470 114.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.490 110.000 87.770 114.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.330 110.000 89.610 114.000 ;
    END
  END chany_top_out[9]
  PIN clk_3_N_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.010 110.000 24.290 114.000 ;
    END
  END clk_3_N_out
  PIN clk_3_S_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END clk_3_S_in
  PIN left_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END left_bottom_grid_pin_11_
  PIN left_bottom_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END left_bottom_grid_pin_13_
  PIN left_bottom_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END left_bottom_grid_pin_15_
  PIN left_bottom_grid_pin_17_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END left_bottom_grid_pin_17_
  PIN left_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 4.000 1.320 ;
    END
  END left_bottom_grid_pin_1_
  PIN left_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END left_bottom_grid_pin_3_
  PIN left_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END left_bottom_grid_pin_5_
  PIN left_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END left_bottom_grid_pin_7_
  PIN left_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END left_bottom_grid_pin_9_
  PIN prog_clk_0_N_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.870 110.000 20.150 114.000 ;
    END
  END prog_clk_0_N_in
  PIN prog_clk_3_N_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.310 110.000 26.590 114.000 ;
    END
  END prog_clk_3_N_out
  PIN prog_clk_3_S_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END prog_clk_3_S_in
  PIN right_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 12.280 114.000 12.880 ;
    END
  END right_bottom_grid_pin_11_
  PIN right_bottom_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 14.320 114.000 14.920 ;
    END
  END right_bottom_grid_pin_13_
  PIN right_bottom_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 17.040 114.000 17.640 ;
    END
  END right_bottom_grid_pin_15_
  PIN right_bottom_grid_pin_17_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 19.080 114.000 19.680 ;
    END
  END right_bottom_grid_pin_17_
  PIN right_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 0.720 114.000 1.320 ;
    END
  END right_bottom_grid_pin_1_
  PIN right_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 2.760 114.000 3.360 ;
    END
  END right_bottom_grid_pin_3_
  PIN right_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 4.800 114.000 5.400 ;
    END
  END right_bottom_grid_pin_5_
  PIN right_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 7.520 114.000 8.120 ;
    END
  END right_bottom_grid_pin_7_
  PIN right_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 9.560 114.000 10.160 ;
    END
  END right_bottom_grid_pin_9_
  PIN top_left_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 110.000 3.130 114.000 ;
    END
  END top_left_grid_pin_42_
  PIN top_left_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.150 110.000 5.430 114.000 ;
    END
  END top_left_grid_pin_43_
  PIN top_left_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 110.000 7.270 114.000 ;
    END
  END top_left_grid_pin_44_
  PIN top_left_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.290 110.000 9.570 114.000 ;
    END
  END top_left_grid_pin_45_
  PIN top_left_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.130 110.000 11.410 114.000 ;
    END
  END top_left_grid_pin_46_
  PIN top_left_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.430 110.000 13.710 114.000 ;
    END
  END top_left_grid_pin_47_
  PIN top_left_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.730 110.000 16.010 114.000 ;
    END
  END top_left_grid_pin_48_
  PIN top_left_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 110.000 17.850 114.000 ;
    END
  END top_left_grid_pin_49_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.880 10.640 23.480 100.880 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.040 10.640 40.640 100.880 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 108.100 100.725 ;
      LAYER met1 ;
        RECT 0.990 5.820 110.790 105.020 ;
      LAYER met2 ;
        RECT 1.570 109.720 2.570 112.725 ;
        RECT 3.410 109.720 4.870 112.725 ;
        RECT 5.710 109.720 6.710 112.725 ;
        RECT 7.550 109.720 9.010 112.725 ;
        RECT 9.850 109.720 10.850 112.725 ;
        RECT 11.690 109.720 13.150 112.725 ;
        RECT 13.990 109.720 15.450 112.725 ;
        RECT 16.290 109.720 17.290 112.725 ;
        RECT 18.130 109.720 19.590 112.725 ;
        RECT 20.430 109.720 21.430 112.725 ;
        RECT 22.270 109.720 23.730 112.725 ;
        RECT 24.570 109.720 26.030 112.725 ;
        RECT 26.870 109.720 27.870 112.725 ;
        RECT 28.710 109.720 30.170 112.725 ;
        RECT 31.010 109.720 32.010 112.725 ;
        RECT 32.850 109.720 34.310 112.725 ;
        RECT 35.150 109.720 36.610 112.725 ;
        RECT 37.450 109.720 38.450 112.725 ;
        RECT 39.290 109.720 40.750 112.725 ;
        RECT 41.590 109.720 42.590 112.725 ;
        RECT 43.430 109.720 44.890 112.725 ;
        RECT 45.730 109.720 47.190 112.725 ;
        RECT 48.030 109.720 49.030 112.725 ;
        RECT 49.870 109.720 51.330 112.725 ;
        RECT 52.170 109.720 53.170 112.725 ;
        RECT 54.010 109.720 55.470 112.725 ;
        RECT 56.310 109.720 57.770 112.725 ;
        RECT 58.610 109.720 59.610 112.725 ;
        RECT 60.450 109.720 61.910 112.725 ;
        RECT 62.750 109.720 63.750 112.725 ;
        RECT 64.590 109.720 66.050 112.725 ;
        RECT 66.890 109.720 67.890 112.725 ;
        RECT 68.730 109.720 70.190 112.725 ;
        RECT 71.030 109.720 72.490 112.725 ;
        RECT 73.330 109.720 74.330 112.725 ;
        RECT 75.170 109.720 76.630 112.725 ;
        RECT 77.470 109.720 78.470 112.725 ;
        RECT 79.310 109.720 80.770 112.725 ;
        RECT 81.610 109.720 83.070 112.725 ;
        RECT 83.910 109.720 84.910 112.725 ;
        RECT 85.750 109.720 87.210 112.725 ;
        RECT 88.050 109.720 89.050 112.725 ;
        RECT 89.890 109.720 91.350 112.725 ;
        RECT 92.190 109.720 93.650 112.725 ;
        RECT 94.490 109.720 95.490 112.725 ;
        RECT 96.330 109.720 97.790 112.725 ;
        RECT 98.630 109.720 99.630 112.725 ;
        RECT 100.470 109.720 101.930 112.725 ;
        RECT 102.770 109.720 104.230 112.725 ;
        RECT 105.070 109.720 106.070 112.725 ;
        RECT 106.910 109.720 108.370 112.725 ;
        RECT 109.210 109.720 110.210 112.725 ;
        RECT 111.050 109.720 112.510 112.725 ;
        RECT 1.020 4.280 113.000 109.720 ;
        RECT 1.020 0.835 10.850 4.280 ;
        RECT 11.690 0.835 33.390 4.280 ;
        RECT 34.230 0.835 56.390 4.280 ;
        RECT 57.230 0.835 78.930 4.280 ;
        RECT 79.770 0.835 101.930 4.280 ;
        RECT 102.770 0.835 113.000 4.280 ;
      LAYER met3 ;
        RECT 4.400 111.840 109.600 112.705 ;
        RECT 4.000 111.200 110.090 111.840 ;
        RECT 4.400 109.800 109.600 111.200 ;
        RECT 4.000 108.480 110.090 109.800 ;
        RECT 4.400 107.080 109.600 108.480 ;
        RECT 4.000 106.440 110.090 107.080 ;
        RECT 4.400 105.040 109.600 106.440 ;
        RECT 4.000 103.720 110.090 105.040 ;
        RECT 4.400 102.320 109.600 103.720 ;
        RECT 4.000 101.680 110.090 102.320 ;
        RECT 4.400 100.280 109.600 101.680 ;
        RECT 4.000 99.640 110.090 100.280 ;
        RECT 4.400 98.240 109.600 99.640 ;
        RECT 4.000 96.920 110.090 98.240 ;
        RECT 4.400 95.520 109.600 96.920 ;
        RECT 4.000 94.880 110.090 95.520 ;
        RECT 4.400 93.480 109.600 94.880 ;
        RECT 4.000 92.160 110.090 93.480 ;
        RECT 4.400 90.760 109.600 92.160 ;
        RECT 4.000 90.120 110.090 90.760 ;
        RECT 4.400 88.720 109.600 90.120 ;
        RECT 4.000 87.400 110.090 88.720 ;
        RECT 4.400 86.000 109.600 87.400 ;
        RECT 4.000 85.360 110.090 86.000 ;
        RECT 4.400 83.960 109.600 85.360 ;
        RECT 4.000 83.320 110.090 83.960 ;
        RECT 4.400 81.920 109.600 83.320 ;
        RECT 4.000 80.600 110.090 81.920 ;
        RECT 4.400 79.200 109.600 80.600 ;
        RECT 4.000 78.560 110.090 79.200 ;
        RECT 4.400 77.160 109.600 78.560 ;
        RECT 4.000 75.840 110.090 77.160 ;
        RECT 4.400 74.440 109.600 75.840 ;
        RECT 4.000 73.800 110.090 74.440 ;
        RECT 4.400 72.400 109.600 73.800 ;
        RECT 4.000 71.080 110.090 72.400 ;
        RECT 4.400 69.680 109.600 71.080 ;
        RECT 4.000 69.040 110.090 69.680 ;
        RECT 4.400 67.640 109.600 69.040 ;
        RECT 4.000 67.000 110.090 67.640 ;
        RECT 4.400 65.600 109.600 67.000 ;
        RECT 4.000 64.280 110.090 65.600 ;
        RECT 4.400 62.880 109.600 64.280 ;
        RECT 4.000 62.240 110.090 62.880 ;
        RECT 4.400 60.840 109.600 62.240 ;
        RECT 4.000 59.520 110.090 60.840 ;
        RECT 4.400 58.120 109.600 59.520 ;
        RECT 4.000 57.480 110.090 58.120 ;
        RECT 4.400 56.080 109.600 57.480 ;
        RECT 4.000 54.760 110.090 56.080 ;
        RECT 4.400 53.360 109.600 54.760 ;
        RECT 4.000 52.720 110.090 53.360 ;
        RECT 4.400 51.320 109.600 52.720 ;
        RECT 4.000 50.680 110.090 51.320 ;
        RECT 4.400 49.280 109.600 50.680 ;
        RECT 4.000 47.960 110.090 49.280 ;
        RECT 4.400 46.560 109.600 47.960 ;
        RECT 4.000 45.920 110.090 46.560 ;
        RECT 4.400 44.520 109.600 45.920 ;
        RECT 4.000 43.200 110.090 44.520 ;
        RECT 4.400 41.800 109.600 43.200 ;
        RECT 4.000 41.160 110.090 41.800 ;
        RECT 4.400 39.760 109.600 41.160 ;
        RECT 4.000 38.440 110.090 39.760 ;
        RECT 4.400 37.040 109.600 38.440 ;
        RECT 4.000 36.400 110.090 37.040 ;
        RECT 4.400 35.000 109.600 36.400 ;
        RECT 4.000 34.360 110.090 35.000 ;
        RECT 4.400 32.960 109.600 34.360 ;
        RECT 4.000 31.640 110.090 32.960 ;
        RECT 4.400 30.240 109.600 31.640 ;
        RECT 4.000 29.600 110.090 30.240 ;
        RECT 4.400 28.200 109.600 29.600 ;
        RECT 4.000 26.880 110.090 28.200 ;
        RECT 4.400 25.480 109.600 26.880 ;
        RECT 4.000 24.840 110.090 25.480 ;
        RECT 4.400 23.440 109.600 24.840 ;
        RECT 4.000 22.120 110.090 23.440 ;
        RECT 4.400 20.720 109.600 22.120 ;
        RECT 4.000 20.080 110.090 20.720 ;
        RECT 4.400 18.680 109.600 20.080 ;
        RECT 4.000 18.040 110.090 18.680 ;
        RECT 4.400 16.640 109.600 18.040 ;
        RECT 4.000 15.320 110.090 16.640 ;
        RECT 4.400 13.920 109.600 15.320 ;
        RECT 4.000 13.280 110.090 13.920 ;
        RECT 4.400 11.880 109.600 13.280 ;
        RECT 4.000 10.560 110.090 11.880 ;
        RECT 4.400 9.160 109.600 10.560 ;
        RECT 4.000 8.520 110.090 9.160 ;
        RECT 4.400 7.120 109.600 8.520 ;
        RECT 4.000 5.800 110.090 7.120 ;
        RECT 4.400 4.400 109.600 5.800 ;
        RECT 4.000 3.760 110.090 4.400 ;
        RECT 4.400 2.360 109.600 3.760 ;
        RECT 4.000 1.720 110.090 2.360 ;
        RECT 4.400 0.855 109.600 1.720 ;
      LAYER met4 ;
        RECT 26.055 10.640 38.640 100.880 ;
        RECT 41.040 10.640 96.305 100.880 ;
  END
END sb_1__0_
END LIBRARY

