VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_io_top_top
  CLASS BLOCK ;
  FOREIGN grid_io_top_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 79.670 BY 45.000 ;
  PIN IO_ISOL_N
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.270 38.800 79.670 39.400 ;
    END
  END IO_ISOL_N
  PIN bottom_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.060 0.000 20.340 2.400 ;
    END
  END bottom_width_0_height_0__pin_0_
  PIN bottom_width_0_height_0__pin_1_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.080 0.000 37.360 2.400 ;
    END
  END bottom_width_0_height_0__pin_1_lower
  PIN bottom_width_0_height_0__pin_1_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 3.040 0.000 3.320 2.400 ;
    END
  END bottom_width_0_height_0__pin_1_upper
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.270 16.360 79.670 16.960 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.270 27.920 79.670 28.520 ;
    END
  END ccff_tail
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 54.100 0.000 54.380 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.120 0.000 71.400 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.080 42.600 37.360 45.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.270 5.480 79.670 6.080 ;
    END
  END prog_clk
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 11.715 10.640 13.315 32.880 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.045 10.640 25.645 32.880 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.190 10.795 73.790 32.725 ;
      LAYER met1 ;
        RECT 0.190 10.640 73.790 32.880 ;
      LAYER met2 ;
        RECT 3.050 42.320 36.800 42.600 ;
        RECT 37.640 42.320 71.390 42.600 ;
        RECT 3.050 2.680 71.390 42.320 ;
        RECT 3.600 2.400 19.780 2.680 ;
        RECT 20.620 2.400 36.800 2.680 ;
        RECT 37.640 2.400 53.820 2.680 ;
        RECT 54.660 2.400 70.840 2.680 ;
      LAYER met3 ;
        RECT 11.715 38.400 76.870 39.265 ;
        RECT 11.715 28.920 77.270 38.400 ;
        RECT 11.715 27.520 76.870 28.920 ;
        RECT 11.715 17.360 77.270 27.520 ;
        RECT 11.715 15.960 76.870 17.360 ;
        RECT 11.715 6.480 77.270 15.960 ;
        RECT 11.715 5.615 76.870 6.480 ;
      LAYER met4 ;
        RECT 26.045 10.640 62.620 32.880 ;
  END
END grid_io_top_top
END LIBRARY

