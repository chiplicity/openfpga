magic
tech EFS8A
magscale 1 2
timestamp 1602873447
<< locali >>
rect 9631 22049 9758 22083
rect 4847 20961 4974 20995
rect 12535 17833 12541 17867
rect 12535 17765 12569 17833
rect 4939 17697 5066 17731
rect 8585 17051 8619 17221
rect 10609 16983 10643 17085
rect 18647 15521 18682 15555
rect 13547 13719 13581 13787
rect 17693 13719 17727 13889
rect 18981 13787 19015 14025
rect 13547 13685 13553 13719
rect 24823 12665 24961 12699
rect 19579 12393 19717 12427
rect 7952 12325 8020 12359
rect 6929 12223 6963 12325
rect 15243 12257 15370 12291
rect 24087 11849 24225 11883
rect 10149 11679 10183 11781
rect 12535 11305 12541 11339
rect 12535 11237 12569 11305
rect 16899 10081 16934 10115
rect 15676 9401 15748 9435
rect 15939 9129 15945 9163
rect 22287 9129 22293 9163
rect 15939 9061 15973 9129
rect 22287 9061 22321 9129
rect 21051 8857 21189 8891
rect 25375 8789 25421 8823
rect 13553 7191 13587 7497
rect 9969 6885 10044 6919
rect 22143 6885 22188 6919
rect 19383 6817 19418 6851
rect 6101 6239 6135 6409
rect 23305 6239 23339 6409
rect 22195 6103 22229 6171
rect 22195 6069 22201 6103
rect 15663 5865 15669 5899
rect 21275 5865 21281 5899
rect 15663 5797 15697 5865
rect 21275 5797 21309 5865
rect 1547 5321 1685 5355
rect 3847 5321 3985 5355
rect 8769 5015 8803 5253
rect 12265 5151 12299 5253
rect 13553 5219 13587 5321
rect 12265 5117 12357 5151
rect 14473 4471 14507 4573
rect 9045 3927 9079 4233
rect 10885 4063 10919 4233
rect 14657 3995 14691 4233
rect 18699 3927 18733 3995
rect 18699 3893 18705 3927
rect 18607 3689 18613 3723
rect 22103 3689 22109 3723
rect 18607 3621 18641 3689
rect 22103 3621 22137 3689
rect 3007 3553 3042 3587
rect 7297 3383 7331 3553
<< viali >>
rect 24777 24905 24811 24939
rect 24593 24701 24627 24735
rect 25145 24701 25179 24735
rect 24777 24361 24811 24395
rect 23489 24225 23523 24259
rect 24593 24225 24627 24259
rect 23673 24089 23707 24123
rect 14013 23817 14047 23851
rect 16589 23817 16623 23851
rect 18337 23817 18371 23851
rect 19441 23817 19475 23851
rect 22201 23817 22235 23851
rect 24777 23817 24811 23851
rect 20637 23749 20671 23783
rect 23857 23749 23891 23783
rect 1460 23613 1494 23647
rect 1869 23613 1903 23647
rect 13829 23613 13863 23647
rect 14381 23613 14415 23647
rect 16405 23613 16439 23647
rect 16957 23613 16991 23647
rect 18153 23613 18187 23647
rect 18705 23613 18739 23647
rect 19257 23613 19291 23647
rect 19809 23613 19843 23647
rect 20453 23613 20487 23647
rect 22017 23613 22051 23647
rect 22569 23613 22603 23647
rect 1547 23545 1581 23579
rect 21005 23545 21039 23579
rect 25145 23545 25179 23579
rect 24777 23273 24811 23307
rect 24593 23137 24627 23171
rect 24593 22389 24627 22423
rect 24777 22185 24811 22219
rect 9597 22049 9631 22083
rect 24593 22049 24627 22083
rect 9827 21845 9861 21879
rect 14381 21641 14415 21675
rect 9388 21437 9422 21471
rect 9781 21437 9815 21471
rect 13896 21437 13930 21471
rect 10149 21369 10183 21403
rect 9459 21301 9493 21335
rect 13967 21301 14001 21335
rect 24593 21301 24627 21335
rect 4813 20961 4847 20995
rect 11412 20961 11446 20995
rect 12884 20961 12918 20995
rect 10333 20893 10367 20927
rect 14013 20893 14047 20927
rect 5043 20757 5077 20791
rect 10885 20757 10919 20791
rect 11483 20757 11517 20791
rect 12955 20757 12989 20791
rect 4905 20553 4939 20587
rect 11621 20553 11655 20587
rect 13277 20553 13311 20587
rect 10701 20417 10735 20451
rect 9632 20349 9666 20383
rect 10057 20349 10091 20383
rect 12852 20349 12886 20383
rect 13737 20349 13771 20383
rect 13921 20349 13955 20383
rect 15460 20349 15494 20383
rect 10793 20281 10827 20315
rect 11345 20281 11379 20315
rect 13829 20281 13863 20315
rect 9735 20213 9769 20247
rect 10517 20213 10551 20247
rect 12633 20213 12667 20247
rect 12955 20213 12989 20247
rect 15531 20213 15565 20247
rect 15853 20213 15887 20247
rect 13461 20009 13495 20043
rect 24777 20009 24811 20043
rect 10241 19941 10275 19975
rect 11805 19941 11839 19975
rect 13737 19941 13771 19975
rect 13829 19941 13863 19975
rect 15945 19873 15979 19907
rect 24593 19873 24627 19907
rect 10149 19805 10183 19839
rect 10793 19805 10827 19839
rect 11713 19805 11747 19839
rect 14381 19805 14415 19839
rect 15301 19805 15335 19839
rect 12265 19737 12299 19771
rect 9965 19669 9999 19703
rect 10241 19465 10275 19499
rect 12633 19465 12667 19499
rect 13277 19465 13311 19499
rect 14381 19465 14415 19499
rect 15945 19465 15979 19499
rect 9965 19329 9999 19363
rect 10609 19329 10643 19363
rect 10885 19329 10919 19363
rect 13461 19329 13495 19363
rect 16635 19329 16669 19363
rect 24593 19329 24627 19363
rect 9137 19261 9171 19295
rect 9321 19261 9355 19295
rect 16532 19261 16566 19295
rect 16957 19261 16991 19295
rect 10977 19193 11011 19227
rect 11529 19193 11563 19227
rect 13553 19193 13587 19227
rect 14105 19193 14139 19227
rect 15025 19193 15059 19227
rect 15117 19193 15151 19227
rect 15669 19193 15703 19227
rect 11805 19125 11839 19159
rect 12265 19125 12299 19159
rect 14841 19125 14875 19159
rect 13461 18921 13495 18955
rect 15025 18921 15059 18955
rect 10701 18853 10735 18887
rect 11621 18853 11655 18887
rect 11713 18853 11747 18887
rect 12265 18853 12299 18887
rect 13829 18853 13863 18887
rect 15485 18853 15519 18887
rect 10609 18785 10643 18819
rect 14381 18785 14415 18819
rect 10977 18717 11011 18751
rect 13737 18717 13771 18751
rect 15393 18717 15427 18751
rect 15669 18717 15703 18751
rect 9689 18377 9723 18411
rect 9919 18377 9953 18411
rect 10609 18377 10643 18411
rect 11805 18377 11839 18411
rect 13093 18377 13127 18411
rect 15301 18377 15335 18411
rect 14841 18309 14875 18343
rect 16773 18309 16807 18343
rect 7481 18241 7515 18275
rect 8953 18241 8987 18275
rect 10885 18241 10919 18275
rect 11529 18241 11563 18275
rect 12173 18241 12207 18275
rect 14289 18241 14323 18275
rect 6996 18173 7030 18207
rect 9816 18173 9850 18207
rect 10241 18173 10275 18207
rect 13236 18173 13270 18207
rect 13645 18173 13679 18207
rect 15669 18173 15703 18207
rect 15853 18173 15887 18207
rect 8309 18105 8343 18139
rect 8401 18105 8435 18139
rect 10977 18105 11011 18139
rect 13323 18105 13357 18139
rect 14381 18105 14415 18139
rect 7067 18037 7101 18071
rect 8033 18037 8067 18071
rect 14013 18037 14047 18071
rect 16037 18037 16071 18071
rect 7113 17833 7147 17867
rect 11345 17833 11379 17867
rect 12541 17833 12575 17867
rect 13093 17833 13127 17867
rect 14105 17833 14139 17867
rect 14473 17833 14507 17867
rect 7389 17765 7423 17799
rect 10746 17765 10780 17799
rect 13737 17765 13771 17799
rect 15393 17765 15427 17799
rect 15485 17765 15519 17799
rect 17049 17765 17083 17799
rect 4905 17697 4939 17731
rect 13921 17697 13955 17731
rect 7297 17629 7331 17663
rect 7665 17629 7699 17663
rect 8217 17629 8251 17663
rect 10425 17629 10459 17663
rect 12173 17629 12207 17663
rect 16037 17629 16071 17663
rect 16957 17629 16991 17663
rect 17601 17629 17635 17663
rect 16405 17561 16439 17595
rect 5135 17493 5169 17527
rect 8953 17493 8987 17527
rect 11989 17493 12023 17527
rect 5089 17289 5123 17323
rect 6653 17289 6687 17323
rect 13829 17289 13863 17323
rect 15577 17289 15611 17323
rect 16221 17289 16255 17323
rect 17417 17289 17451 17323
rect 24777 17289 24811 17323
rect 8585 17221 8619 17255
rect 8677 17221 8711 17255
rect 15945 17221 15979 17255
rect 7389 17153 7423 17187
rect 8033 17153 8067 17187
rect 8953 17153 8987 17187
rect 9229 17153 9263 17187
rect 16497 17153 16531 17187
rect 16773 17153 16807 17187
rect 10609 17085 10643 17119
rect 12173 17085 12207 17119
rect 12725 17085 12759 17119
rect 12909 17085 12943 17119
rect 14105 17085 14139 17119
rect 14657 17085 14691 17119
rect 24593 17085 24627 17119
rect 25145 17085 25179 17119
rect 7481 17017 7515 17051
rect 8585 17017 8619 17051
rect 9045 17017 9079 17051
rect 10149 17017 10183 17051
rect 13230 17017 13264 17051
rect 14565 17017 14599 17051
rect 14978 17017 15012 17051
rect 16589 17017 16623 17051
rect 7205 16949 7239 16983
rect 8401 16949 8435 16983
rect 10425 16949 10459 16983
rect 10609 16949 10643 16983
rect 10793 16949 10827 16983
rect 11253 16949 11287 16983
rect 11897 16949 11931 16983
rect 18061 16949 18095 16983
rect 11529 16745 11563 16779
rect 14657 16745 14691 16779
rect 15485 16745 15519 16779
rect 17141 16745 17175 16779
rect 6745 16677 6779 16711
rect 7757 16677 7791 16711
rect 8309 16677 8343 16711
rect 11161 16677 11195 16711
rect 13461 16677 13495 16711
rect 14105 16677 14139 16711
rect 16313 16677 16347 16711
rect 17877 16677 17911 16711
rect 6653 16609 6687 16643
rect 9137 16609 9171 16643
rect 9505 16609 9539 16643
rect 9965 16609 9999 16643
rect 10425 16609 10459 16643
rect 10517 16609 10551 16643
rect 11069 16609 11103 16643
rect 12265 16609 12299 16643
rect 12449 16609 12483 16643
rect 12817 16609 12851 16643
rect 13369 16609 13403 16643
rect 7665 16541 7699 16575
rect 16221 16541 16255 16575
rect 17785 16541 17819 16575
rect 16773 16473 16807 16507
rect 18337 16473 18371 16507
rect 7297 16405 7331 16439
rect 8677 16405 8711 16439
rect 11805 16405 11839 16439
rect 13737 16405 13771 16439
rect 6653 16201 6687 16235
rect 7665 16201 7699 16235
rect 9229 16201 9263 16235
rect 16221 16201 16255 16235
rect 17785 16201 17819 16235
rect 18521 16201 18555 16235
rect 24777 16201 24811 16235
rect 6285 16133 6319 16167
rect 11437 16133 11471 16167
rect 13829 16133 13863 16167
rect 15669 16133 15703 16167
rect 6837 16065 6871 16099
rect 5784 15997 5818 16031
rect 8309 15997 8343 16031
rect 10333 15997 10367 16031
rect 10517 15997 10551 16031
rect 10885 15997 10919 16031
rect 11253 15997 11287 16031
rect 12633 15997 12667 16031
rect 12909 15997 12943 16031
rect 13277 15997 13311 16031
rect 13645 15997 13679 16031
rect 14749 15997 14783 16031
rect 18096 15997 18130 16031
rect 18889 15997 18923 16031
rect 24593 15997 24627 16031
rect 25145 15997 25179 16031
rect 5871 15929 5905 15963
rect 8217 15929 8251 15963
rect 8671 15929 8705 15963
rect 14197 15929 14231 15963
rect 14657 15929 14691 15963
rect 15111 15929 15145 15963
rect 18199 15929 18233 15963
rect 9505 15861 9539 15895
rect 9873 15861 9907 15895
rect 11897 15861 11931 15895
rect 12173 15861 12207 15895
rect 16497 15861 16531 15895
rect 17049 15861 17083 15895
rect 7481 15657 7515 15691
rect 8585 15657 8619 15691
rect 10057 15657 10091 15691
rect 11713 15657 11747 15691
rect 14013 15657 14047 15691
rect 16221 15657 16255 15691
rect 18751 15657 18785 15691
rect 6837 15589 6871 15623
rect 8027 15589 8061 15623
rect 15663 15589 15697 15623
rect 17233 15589 17267 15623
rect 6745 15521 6779 15555
rect 9137 15521 9171 15555
rect 10149 15521 10183 15555
rect 10701 15521 10735 15555
rect 10793 15521 10827 15555
rect 11345 15521 11379 15555
rect 12173 15521 12207 15555
rect 12449 15521 12483 15555
rect 12725 15521 12759 15555
rect 13093 15521 13127 15555
rect 13461 15521 13495 15555
rect 18613 15521 18647 15555
rect 7665 15453 7699 15487
rect 13737 15453 13771 15487
rect 15301 15453 15335 15487
rect 17141 15453 17175 15487
rect 17601 15453 17635 15487
rect 9505 15317 9539 15351
rect 14749 15317 14783 15351
rect 18061 15317 18095 15351
rect 6193 15113 6227 15147
rect 6653 15113 6687 15147
rect 8125 15113 8159 15147
rect 9137 15113 9171 15147
rect 16129 15113 16163 15147
rect 17693 15113 17727 15147
rect 7665 15045 7699 15079
rect 14197 15045 14231 15079
rect 13921 14977 13955 15011
rect 15301 14977 15335 15011
rect 17049 14977 17083 15011
rect 17325 14977 17359 15011
rect 19073 14977 19107 15011
rect 8861 14909 8895 14943
rect 8953 14909 8987 14943
rect 10149 14909 10183 14943
rect 10701 14909 10735 14943
rect 10793 14909 10827 14943
rect 11161 14909 11195 14943
rect 12449 14909 12483 14943
rect 12909 14909 12943 14943
rect 13277 14909 13311 14943
rect 13645 14909 13679 14943
rect 16865 14909 16899 14943
rect 18096 14909 18130 14943
rect 7113 14841 7147 14875
rect 7205 14841 7239 14875
rect 8493 14841 8527 14875
rect 11713 14841 11747 14875
rect 12173 14841 12207 14875
rect 14841 14841 14875 14875
rect 14933 14841 14967 14875
rect 18199 14841 18233 14875
rect 9413 14773 9447 14807
rect 9781 14773 9815 14807
rect 10057 14773 10091 14807
rect 14657 14773 14691 14807
rect 15761 14773 15795 14807
rect 18705 14773 18739 14807
rect 9137 14569 9171 14603
rect 11253 14569 11287 14603
rect 11897 14569 11931 14603
rect 13093 14569 13127 14603
rect 14841 14569 14875 14603
rect 15439 14569 15473 14603
rect 16405 14569 16439 14603
rect 24777 14569 24811 14603
rect 9965 14501 9999 14535
rect 11621 14501 11655 14535
rect 16681 14501 16715 14535
rect 16773 14501 16807 14535
rect 6688 14433 6722 14467
rect 8192 14433 8226 14467
rect 10057 14433 10091 14467
rect 11069 14433 11103 14467
rect 12081 14433 12115 14467
rect 12633 14433 12667 14467
rect 14289 14433 14323 14467
rect 15368 14433 15402 14467
rect 18153 14433 18187 14467
rect 18613 14433 18647 14467
rect 19717 14433 19751 14467
rect 24593 14433 24627 14467
rect 10517 14365 10551 14399
rect 12817 14365 12851 14399
rect 14381 14365 14415 14399
rect 16957 14365 16991 14399
rect 18797 14365 18831 14399
rect 7113 14297 7147 14331
rect 9505 14297 9539 14331
rect 10241 14297 10275 14331
rect 13461 14297 13495 14331
rect 6791 14229 6825 14263
rect 7849 14229 7883 14263
rect 8263 14229 8297 14263
rect 16037 14229 16071 14263
rect 19901 14229 19935 14263
rect 14105 14025 14139 14059
rect 14381 14025 14415 14059
rect 14841 14025 14875 14059
rect 15393 14025 15427 14059
rect 18981 14025 19015 14059
rect 19073 14025 19107 14059
rect 24593 14025 24627 14059
rect 7849 13889 7883 13923
rect 8217 13889 8251 13923
rect 16129 13889 16163 13923
rect 16773 13889 16807 13923
rect 17693 13889 17727 13923
rect 1476 13821 1510 13855
rect 1869 13821 1903 13855
rect 9321 13821 9355 13855
rect 9689 13821 9723 13855
rect 11161 13821 11195 13855
rect 13185 13821 13219 13855
rect 15000 13821 15034 13855
rect 7021 13753 7055 13787
rect 7665 13753 7699 13787
rect 7941 13753 7975 13787
rect 10333 13753 10367 13787
rect 12173 13753 12207 13787
rect 15761 13753 15795 13787
rect 16221 13753 16255 13787
rect 18337 13821 18371 13855
rect 18613 13821 18647 13855
rect 24823 13957 24857 13991
rect 19717 13889 19751 13923
rect 20244 13821 20278 13855
rect 20637 13821 20671 13855
rect 21256 13821 21290 13855
rect 22636 13821 22670 13855
rect 24720 13821 24754 13855
rect 17785 13753 17819 13787
rect 18981 13753 19015 13787
rect 21649 13753 21683 13787
rect 23121 13753 23155 13787
rect 25237 13753 25271 13787
rect 1547 13685 1581 13719
rect 8861 13685 8895 13719
rect 9137 13685 9171 13719
rect 11345 13685 11379 13719
rect 12725 13685 12759 13719
rect 13093 13685 13127 13719
rect 13553 13685 13587 13719
rect 15071 13685 15105 13719
rect 17049 13685 17083 13719
rect 17509 13685 17543 13719
rect 17693 13685 17727 13719
rect 18337 13685 18371 13719
rect 20315 13685 20349 13719
rect 21327 13685 21361 13719
rect 22707 13685 22741 13719
rect 23673 13685 23707 13719
rect 13829 13481 13863 13515
rect 16589 13481 16623 13515
rect 18705 13481 18739 13515
rect 21005 13481 21039 13515
rect 22707 13481 22741 13515
rect 6377 13413 6411 13447
rect 6561 13413 6595 13447
rect 6653 13413 6687 13447
rect 8217 13413 8251 13447
rect 9873 13413 9907 13447
rect 11069 13413 11103 13447
rect 15622 13413 15656 13447
rect 17049 13413 17083 13447
rect 18245 13413 18279 13447
rect 12081 13345 12115 13379
rect 12541 13345 12575 13379
rect 13093 13345 13127 13379
rect 13461 13345 13495 13379
rect 16221 13345 16255 13379
rect 17417 13345 17451 13379
rect 18889 13345 18923 13379
rect 19073 13345 19107 13379
rect 20913 13345 20947 13379
rect 21373 13345 21407 13379
rect 22636 13345 22670 13379
rect 23648 13345 23682 13379
rect 24660 13345 24694 13379
rect 8125 13277 8159 13311
rect 9781 13277 9815 13311
rect 10057 13277 10091 13311
rect 13553 13277 13587 13311
rect 15301 13277 15335 13311
rect 7113 13209 7147 13243
rect 8677 13209 8711 13243
rect 10793 13209 10827 13243
rect 7941 13141 7975 13175
rect 9045 13141 9079 13175
rect 9505 13141 9539 13175
rect 11529 13141 11563 13175
rect 11897 13141 11931 13175
rect 23719 13141 23753 13175
rect 24731 13141 24765 13175
rect 7665 12937 7699 12971
rect 8033 12937 8067 12971
rect 9045 12937 9079 12971
rect 11805 12937 11839 12971
rect 12173 12937 12207 12971
rect 14657 12937 14691 12971
rect 16221 12937 16255 12971
rect 17417 12937 17451 12971
rect 19073 12937 19107 12971
rect 13829 12869 13863 12903
rect 15853 12869 15887 12903
rect 23811 12869 23845 12903
rect 24593 12869 24627 12903
rect 14197 12801 14231 12835
rect 14933 12801 14967 12835
rect 15301 12801 15335 12835
rect 16497 12801 16531 12835
rect 16773 12801 16807 12835
rect 18613 12801 18647 12835
rect 21281 12801 21315 12835
rect 25237 12801 25271 12835
rect 5089 12733 5123 12767
rect 5825 12733 5859 12767
rect 8125 12733 8159 12767
rect 9413 12733 9447 12767
rect 10149 12733 10183 12767
rect 10609 12733 10643 12767
rect 10793 12733 10827 12767
rect 11069 12733 11103 12767
rect 12449 12733 12483 12767
rect 12909 12733 12943 12767
rect 13277 12733 13311 12767
rect 13645 12733 13679 12767
rect 19809 12733 19843 12767
rect 19901 12733 19935 12767
rect 20361 12733 20395 12767
rect 21465 12733 21499 12767
rect 21925 12733 21959 12767
rect 23740 12733 23774 12767
rect 24752 12733 24786 12767
rect 5917 12665 5951 12699
rect 6469 12665 6503 12699
rect 8446 12665 8480 12699
rect 15025 12665 15059 12699
rect 16589 12665 16623 12699
rect 18153 12665 18187 12699
rect 18245 12665 18279 12699
rect 20637 12665 20671 12699
rect 24961 12665 24995 12699
rect 6837 12597 6871 12631
rect 9781 12597 9815 12631
rect 9965 12597 9999 12631
rect 17785 12597 17819 12631
rect 20913 12597 20947 12631
rect 21741 12597 21775 12631
rect 22477 12597 22511 12631
rect 22845 12597 22879 12631
rect 24225 12597 24259 12631
rect 25513 12597 25547 12631
rect 7113 12393 7147 12427
rect 7573 12393 7607 12427
rect 9873 12393 9907 12427
rect 14841 12393 14875 12427
rect 15439 12393 15473 12427
rect 17693 12393 17727 12427
rect 19717 12393 19751 12427
rect 21925 12393 21959 12427
rect 22569 12393 22603 12427
rect 6285 12325 6319 12359
rect 6929 12325 6963 12359
rect 7918 12325 7952 12359
rect 9137 12325 9171 12359
rect 13829 12325 13863 12359
rect 16497 12325 16531 12359
rect 17325 12325 17359 12359
rect 17969 12325 18003 12359
rect 18061 12325 18095 12359
rect 6837 12257 6871 12291
rect 7665 12257 7699 12291
rect 8585 12257 8619 12291
rect 10057 12257 10091 12291
rect 10241 12257 10275 12291
rect 10609 12257 10643 12291
rect 10977 12257 11011 12291
rect 12725 12257 12759 12291
rect 15209 12257 15243 12291
rect 15761 12257 15795 12291
rect 19476 12257 19510 12291
rect 20913 12257 20947 12291
rect 21373 12257 21407 12291
rect 22477 12257 22511 12291
rect 22937 12257 22971 12291
rect 24108 12257 24142 12291
rect 25120 12257 25154 12291
rect 6193 12189 6227 12223
rect 6929 12189 6963 12223
rect 13737 12189 13771 12223
rect 14381 12189 14415 12223
rect 16405 12189 16439 12223
rect 17049 12189 17083 12223
rect 19901 12189 19935 12223
rect 21649 12189 21683 12223
rect 11529 12121 11563 12155
rect 13093 12121 13127 12155
rect 18521 12121 18555 12155
rect 9505 12053 9539 12087
rect 11897 12053 11931 12087
rect 12357 12053 12391 12087
rect 16221 12053 16255 12087
rect 18889 12053 18923 12087
rect 19349 12053 19383 12087
rect 20637 12053 20671 12087
rect 24179 12053 24213 12087
rect 25191 12053 25225 12087
rect 5917 11849 5951 11883
rect 6653 11849 6687 11883
rect 7941 11849 7975 11883
rect 8769 11849 8803 11883
rect 12265 11849 12299 11883
rect 14289 11849 14323 11883
rect 16221 11849 16255 11883
rect 16497 11849 16531 11883
rect 17877 11849 17911 11883
rect 20913 11849 20947 11883
rect 22201 11849 22235 11883
rect 22569 11849 22603 11883
rect 24225 11849 24259 11883
rect 24501 11849 24535 11883
rect 9137 11781 9171 11815
rect 9321 11781 9355 11815
rect 10149 11781 10183 11815
rect 13461 11781 13495 11815
rect 18705 11781 18739 11815
rect 21833 11781 21867 11815
rect 6929 11713 6963 11747
rect 7573 11713 7607 11747
rect 12541 11713 12575 11747
rect 13185 11713 13219 11747
rect 15301 11713 15335 11747
rect 16865 11713 16899 11747
rect 18153 11713 18187 11747
rect 19993 11713 20027 11747
rect 5733 11645 5767 11679
rect 6193 11645 6227 11679
rect 9229 11645 9263 11679
rect 9505 11645 9539 11679
rect 10149 11645 10183 11679
rect 10793 11645 10827 11679
rect 10885 11645 10919 11679
rect 11069 11645 11103 11679
rect 11529 11645 11563 11679
rect 14105 11645 14139 11679
rect 14657 11645 14691 11679
rect 17417 11645 17451 11679
rect 22937 11645 22971 11679
rect 24016 11645 24050 11679
rect 24777 11645 24811 11679
rect 25028 11645 25062 11679
rect 7021 11577 7055 11611
rect 8401 11577 8435 11611
rect 9965 11577 9999 11611
rect 12633 11577 12667 11611
rect 15663 11577 15697 11611
rect 18245 11577 18279 11611
rect 19717 11577 19751 11611
rect 19809 11577 19843 11611
rect 21281 11577 21315 11611
rect 21373 11577 21407 11611
rect 25513 11577 25547 11611
rect 5549 11509 5583 11543
rect 10241 11509 10275 11543
rect 10701 11509 10735 11543
rect 11897 11509 11931 11543
rect 13829 11509 13863 11543
rect 15117 11509 15151 11543
rect 19073 11509 19107 11543
rect 19441 11509 19475 11543
rect 25099 11509 25133 11543
rect 25881 11509 25915 11543
rect 6193 11305 6227 11339
rect 7757 11305 7791 11339
rect 12541 11305 12575 11339
rect 13093 11305 13127 11339
rect 14013 11305 14047 11339
rect 16221 11305 16255 11339
rect 16589 11305 16623 11339
rect 17969 11305 18003 11339
rect 18705 11305 18739 11339
rect 21925 11305 21959 11339
rect 24225 11305 24259 11339
rect 8033 11237 8067 11271
rect 13737 11237 13771 11271
rect 15663 11237 15697 11271
rect 17370 11237 17404 11271
rect 18245 11237 18279 11271
rect 18981 11237 19015 11271
rect 19533 11237 19567 11271
rect 20177 11237 20211 11271
rect 22753 11237 22787 11271
rect 23305 11237 23339 11271
rect 1476 11169 1510 11203
rect 6888 11169 6922 11203
rect 10057 11169 10091 11203
rect 10333 11169 10367 11203
rect 10885 11169 10919 11203
rect 11161 11169 11195 11203
rect 14264 11169 14298 11203
rect 17049 11169 17083 11203
rect 21097 11169 21131 11203
rect 21373 11169 21407 11203
rect 24225 11169 24259 11203
rect 24593 11169 24627 11203
rect 6975 11101 7009 11135
rect 7941 11101 7975 11135
rect 8217 11101 8251 11135
rect 9321 11101 9355 11135
rect 11345 11101 11379 11135
rect 12173 11101 12207 11135
rect 15301 11101 15335 11135
rect 18889 11101 18923 11135
rect 21649 11101 21683 11135
rect 22661 11101 22695 11135
rect 20637 11033 20671 11067
rect 1547 10965 1581 10999
rect 7389 10965 7423 10999
rect 8861 10965 8895 10999
rect 14335 10965 14369 10999
rect 15025 10965 15059 10999
rect 19809 10965 19843 10999
rect 23765 10965 23799 10999
rect 1593 10761 1627 10795
rect 8769 10761 8803 10795
rect 9229 10761 9263 10795
rect 11437 10761 11471 10795
rect 11805 10761 11839 10795
rect 12265 10761 12299 10795
rect 15209 10761 15243 10795
rect 17003 10761 17037 10795
rect 18981 10761 19015 10795
rect 19257 10761 19291 10795
rect 19947 10761 19981 10795
rect 20729 10761 20763 10795
rect 22109 10761 22143 10795
rect 22661 10761 22695 10795
rect 24685 10761 24719 10795
rect 5917 10693 5951 10727
rect 13829 10693 13863 10727
rect 16681 10693 16715 10727
rect 17693 10693 17727 10727
rect 19717 10693 19751 10727
rect 20361 10693 20395 10727
rect 6285 10625 6319 10659
rect 12541 10625 12575 10659
rect 13185 10625 13219 10659
rect 16037 10625 16071 10659
rect 18061 10625 18095 10659
rect 21189 10625 21223 10659
rect 23765 10625 23799 10659
rect 24041 10625 24075 10659
rect 5733 10557 5767 10591
rect 7573 10557 7607 10591
rect 9597 10557 9631 10591
rect 9781 10557 9815 10591
rect 10333 10557 10367 10591
rect 10517 10557 10551 10591
rect 14013 10557 14047 10591
rect 16900 10557 16934 10591
rect 17325 10557 17359 10591
rect 19876 10557 19910 10591
rect 22937 10557 22971 10591
rect 25272 10557 25306 10591
rect 25697 10557 25731 10591
rect 7481 10489 7515 10523
rect 7935 10489 7969 10523
rect 12633 10489 12667 10523
rect 15393 10489 15427 10523
rect 15485 10489 15519 10523
rect 18382 10489 18416 10523
rect 21005 10489 21039 10523
rect 21510 10489 21544 10523
rect 23397 10489 23431 10523
rect 23857 10489 23891 10523
rect 7113 10421 7147 10455
rect 8493 10421 8527 10455
rect 9413 10421 9447 10455
rect 11069 10421 11103 10455
rect 14197 10421 14231 10455
rect 14565 10421 14599 10455
rect 16405 10421 16439 10455
rect 25375 10421 25409 10455
rect 7297 10217 7331 10251
rect 9045 10217 9079 10251
rect 9413 10217 9447 10251
rect 9965 10217 9999 10251
rect 10609 10217 10643 10251
rect 12541 10217 12575 10251
rect 12817 10217 12851 10251
rect 15577 10217 15611 10251
rect 17417 10217 17451 10251
rect 21097 10217 21131 10251
rect 22477 10217 22511 10251
rect 24317 10217 24351 10251
rect 7573 10149 7607 10183
rect 8125 10149 8159 10183
rect 18245 10149 18279 10183
rect 18797 10149 18831 10183
rect 21878 10149 21912 10183
rect 23489 10149 23523 10183
rect 24041 10149 24075 10183
rect 25053 10149 25087 10183
rect 4848 10081 4882 10115
rect 5825 10081 5859 10115
rect 6377 10081 6411 10115
rect 10149 10081 10183 10115
rect 11805 10081 11839 10115
rect 13921 10081 13955 10115
rect 14105 10081 14139 10115
rect 15485 10081 15519 10115
rect 15853 10081 15887 10115
rect 16865 10081 16899 10115
rect 19660 10081 19694 10115
rect 21557 10081 21591 10115
rect 6469 10013 6503 10047
rect 7481 10013 7515 10047
rect 11161 10013 11195 10047
rect 14381 10013 14415 10047
rect 18153 10013 18187 10047
rect 22845 10013 22879 10047
rect 23397 10013 23431 10047
rect 24961 10013 24995 10047
rect 25237 10013 25271 10047
rect 10333 9945 10367 9979
rect 4951 9877 4985 9911
rect 8401 9877 8435 9911
rect 13553 9877 13587 9911
rect 15117 9877 15151 9911
rect 17003 9877 17037 9911
rect 19763 9877 19797 9911
rect 23213 9877 23247 9911
rect 4813 9673 4847 9707
rect 6561 9673 6595 9707
rect 12587 9673 12621 9707
rect 15301 9673 15335 9707
rect 18337 9673 18371 9707
rect 19717 9673 19751 9707
rect 21557 9673 21591 9707
rect 25375 9673 25409 9707
rect 10609 9605 10643 9639
rect 19441 9605 19475 9639
rect 20177 9605 20211 9639
rect 24961 9605 24995 9639
rect 7849 9537 7883 9571
rect 8125 9537 8159 9571
rect 17877 9537 17911 9571
rect 18521 9537 18555 9571
rect 20361 9537 20395 9571
rect 20637 9537 20671 9571
rect 21833 9537 21867 9571
rect 23765 9537 23799 9571
rect 24133 9537 24167 9571
rect 5641 9469 5675 9503
rect 5733 9469 5767 9503
rect 7205 9469 7239 9503
rect 8677 9469 8711 9503
rect 9229 9469 9263 9503
rect 11069 9469 11103 9503
rect 11253 9469 11287 9503
rect 12516 9469 12550 9503
rect 12909 9469 12943 9503
rect 13461 9469 13495 9503
rect 13921 9469 13955 9503
rect 15393 9469 15427 9503
rect 16313 9469 16347 9503
rect 25272 9469 25306 9503
rect 25697 9469 25731 9503
rect 6193 9401 6227 9435
rect 10241 9401 10275 9435
rect 11529 9401 11563 9435
rect 14197 9401 14231 9435
rect 14565 9401 14599 9435
rect 14933 9401 14967 9435
rect 15642 9401 15676 9435
rect 16865 9401 16899 9435
rect 18883 9401 18917 9435
rect 20453 9401 20487 9435
rect 22154 9401 22188 9435
rect 23029 9401 23063 9435
rect 23857 9401 23891 9435
rect 5917 9333 5951 9367
rect 8493 9333 8527 9367
rect 8769 9333 8803 9367
rect 11897 9333 11931 9367
rect 13277 9333 13311 9367
rect 17509 9333 17543 9367
rect 22753 9333 22787 9367
rect 23397 9333 23431 9367
rect 5181 9129 5215 9163
rect 7205 9129 7239 9163
rect 9873 9129 9907 9163
rect 13921 9129 13955 9163
rect 15025 9129 15059 9163
rect 15945 9129 15979 9163
rect 16497 9129 16531 9163
rect 18153 9129 18187 9163
rect 20269 9129 20303 9163
rect 20729 9129 20763 9163
rect 21741 9129 21775 9163
rect 22293 9129 22327 9163
rect 22845 9129 22879 9163
rect 24777 9129 24811 9163
rect 6193 9061 6227 9095
rect 6285 9061 6319 9095
rect 7941 9061 7975 9095
rect 8217 9061 8251 9095
rect 12954 9061 12988 9095
rect 18883 9061 18917 9095
rect 23305 9061 23339 9095
rect 23765 9061 23799 9095
rect 23857 9061 23891 9095
rect 9689 8993 9723 9027
rect 11069 8993 11103 9027
rect 11529 8993 11563 9027
rect 15577 8993 15611 9027
rect 17576 8993 17610 9027
rect 20948 8993 20982 9027
rect 21925 8993 21959 9027
rect 25304 8993 25338 9027
rect 6469 8925 6503 8959
rect 8125 8925 8159 8959
rect 11805 8925 11839 8959
rect 12633 8925 12667 8959
rect 18521 8925 18555 8959
rect 24041 8925 24075 8959
rect 7481 8857 7515 8891
rect 8677 8857 8711 8891
rect 19717 8857 19751 8891
rect 21189 8857 21223 8891
rect 25145 8857 25179 8891
rect 9137 8789 9171 8823
rect 10149 8789 10183 8823
rect 10793 8789 10827 8823
rect 12541 8789 12575 8823
rect 13553 8789 13587 8823
rect 14289 8789 14323 8823
rect 17417 8789 17451 8823
rect 17647 8789 17681 8823
rect 19441 8789 19475 8823
rect 21465 8789 21499 8823
rect 25421 8789 25455 8823
rect 6561 8585 6595 8619
rect 8033 8585 8067 8619
rect 9045 8585 9079 8619
rect 11069 8585 11103 8619
rect 11805 8585 11839 8619
rect 14013 8585 14047 8619
rect 15301 8585 15335 8619
rect 15669 8585 15703 8619
rect 20913 8585 20947 8619
rect 22661 8585 22695 8619
rect 23489 8585 23523 8619
rect 23857 8585 23891 8619
rect 25421 8585 25455 8619
rect 9781 8517 9815 8551
rect 21925 8517 21959 8551
rect 24961 8517 24995 8551
rect 5273 8449 5307 8483
rect 5917 8449 5951 8483
rect 8125 8449 8159 8483
rect 10425 8449 10459 8483
rect 12449 8449 12483 8483
rect 14289 8449 14323 8483
rect 14565 8449 14599 8483
rect 18245 8449 18279 8483
rect 18889 8449 18923 8483
rect 19809 8449 19843 8483
rect 20453 8449 20487 8483
rect 21373 8449 21407 8483
rect 23029 8449 23063 8483
rect 24409 8449 24443 8483
rect 25697 8449 25731 8483
rect 1444 8381 1478 8415
rect 1869 8381 1903 8415
rect 7113 8381 7147 8415
rect 7573 8381 7607 8415
rect 9965 8381 9999 8415
rect 10333 8381 10367 8415
rect 16681 8381 16715 8415
rect 16957 8381 16991 8415
rect 22293 8381 22327 8415
rect 1547 8313 1581 8347
rect 5089 8313 5123 8347
rect 5365 8313 5399 8347
rect 6285 8313 6319 8347
rect 8446 8313 8480 8347
rect 12770 8313 12804 8347
rect 14381 8313 14415 8347
rect 16313 8313 16347 8347
rect 17141 8313 17175 8347
rect 18337 8313 18371 8347
rect 19625 8313 19659 8347
rect 19901 8313 19935 8347
rect 21465 8313 21499 8347
rect 24501 8313 24535 8347
rect 7297 8245 7331 8279
rect 9413 8245 9447 8279
rect 11437 8245 11471 8279
rect 12173 8245 12207 8279
rect 13369 8245 13403 8279
rect 17601 8245 17635 8279
rect 19165 8245 19199 8279
rect 7297 8041 7331 8075
rect 7757 8041 7791 8075
rect 9045 8041 9079 8075
rect 12449 8041 12483 8075
rect 12725 8041 12759 8075
rect 15393 8041 15427 8075
rect 16497 8041 16531 8075
rect 18061 8041 18095 8075
rect 18705 8041 18739 8075
rect 19165 8041 19199 8075
rect 23673 8041 23707 8075
rect 6469 7973 6503 8007
rect 8170 7973 8204 8007
rect 11891 7973 11925 8007
rect 13829 7973 13863 8007
rect 21281 7973 21315 8007
rect 22845 7973 22879 8007
rect 24409 7973 24443 8007
rect 24961 7973 24995 8007
rect 5308 7905 5342 7939
rect 7849 7905 7883 7939
rect 9965 7905 9999 7939
rect 10425 7905 10459 7939
rect 15301 7905 15335 7939
rect 15761 7905 15795 7939
rect 16957 7905 16991 7939
rect 17509 7905 17543 7939
rect 19257 7905 19291 7939
rect 19809 7905 19843 7939
rect 4261 7837 4295 7871
rect 6377 7837 6411 7871
rect 7021 7837 7055 7871
rect 10701 7837 10735 7871
rect 11529 7837 11563 7871
rect 13553 7837 13587 7871
rect 13737 7837 13771 7871
rect 17601 7837 17635 7871
rect 19993 7837 20027 7871
rect 21189 7837 21223 7871
rect 21465 7837 21499 7871
rect 22753 7837 22787 7871
rect 24317 7837 24351 7871
rect 14289 7769 14323 7803
rect 16773 7769 16807 7803
rect 23305 7769 23339 7803
rect 5411 7701 5445 7735
rect 6101 7701 6135 7735
rect 8769 7701 8803 7735
rect 9413 7701 9447 7735
rect 18429 7701 18463 7735
rect 22109 7701 22143 7735
rect 24133 7701 24167 7735
rect 5273 7497 5307 7531
rect 6561 7497 6595 7531
rect 7941 7497 7975 7531
rect 11897 7497 11931 7531
rect 13553 7497 13587 7531
rect 13645 7497 13679 7531
rect 15531 7497 15565 7531
rect 17417 7497 17451 7531
rect 17877 7497 17911 7531
rect 19809 7497 19843 7531
rect 23397 7497 23431 7531
rect 25375 7497 25409 7531
rect 4629 7429 4663 7463
rect 6929 7361 6963 7395
rect 8769 7361 8803 7395
rect 10977 7361 11011 7395
rect 4721 7293 4755 7327
rect 5800 7293 5834 7327
rect 6285 7293 6319 7327
rect 9965 7293 9999 7327
rect 10425 7293 10459 7327
rect 12868 7293 12902 7327
rect 7021 7225 7055 7259
rect 7573 7225 7607 7259
rect 8493 7225 8527 7259
rect 8585 7225 8619 7259
rect 10701 7225 10735 7259
rect 12955 7225 12989 7259
rect 14841 7429 14875 7463
rect 24685 7429 24719 7463
rect 25053 7429 25087 7463
rect 14289 7361 14323 7395
rect 16313 7361 16347 7395
rect 18429 7361 18463 7395
rect 20729 7361 20763 7395
rect 23765 7361 23799 7395
rect 24409 7361 24443 7395
rect 15460 7293 15494 7327
rect 15853 7293 15887 7327
rect 16681 7293 16715 7327
rect 16865 7293 16899 7327
rect 19073 7293 19107 7327
rect 25304 7293 25338 7327
rect 13921 7225 13955 7259
rect 14013 7225 14047 7259
rect 17141 7225 17175 7259
rect 18521 7225 18555 7259
rect 19349 7225 19383 7259
rect 20453 7225 20487 7259
rect 20545 7225 20579 7259
rect 22109 7225 22143 7259
rect 22201 7225 22235 7259
rect 22753 7225 22787 7259
rect 23857 7225 23891 7259
rect 4905 7157 4939 7191
rect 5871 7157 5905 7191
rect 8309 7157 8343 7191
rect 9413 7157 9447 7191
rect 9873 7157 9907 7191
rect 11621 7157 11655 7191
rect 13369 7157 13403 7191
rect 13553 7157 13587 7191
rect 15209 7157 15243 7191
rect 20269 7157 20303 7191
rect 21465 7157 21499 7191
rect 21833 7157 21867 7191
rect 23121 7157 23155 7191
rect 25789 7157 25823 7191
rect 6285 6953 6319 6987
rect 8217 6953 8251 6987
rect 10885 6953 10919 6987
rect 11989 6953 12023 6987
rect 13461 6953 13495 6987
rect 14657 6953 14691 6987
rect 15485 6953 15519 6987
rect 19487 6953 19521 6987
rect 21189 6953 21223 6987
rect 22753 6953 22787 6987
rect 4629 6885 4663 6919
rect 6745 6885 6779 6919
rect 6837 6885 6871 6919
rect 7389 6885 7423 6919
rect 7941 6885 7975 6919
rect 9935 6885 9969 6919
rect 13829 6885 13863 6919
rect 17922 6885 17956 6919
rect 18797 6885 18831 6919
rect 19809 6885 19843 6919
rect 22109 6885 22143 6919
rect 23857 6885 23891 6919
rect 4144 6817 4178 6851
rect 5089 6817 5123 6851
rect 5365 6817 5399 6851
rect 8585 6817 8619 6851
rect 11529 6817 11563 6851
rect 11621 6817 11655 6851
rect 11805 6817 11839 6851
rect 16313 6817 16347 6851
rect 16589 6817 16623 6851
rect 17601 6817 17635 6851
rect 19349 6817 19383 6851
rect 21833 6817 21867 6851
rect 25304 6817 25338 6851
rect 4997 6749 5031 6783
rect 5825 6749 5859 6783
rect 9689 6749 9723 6783
rect 13185 6749 13219 6783
rect 13737 6749 13771 6783
rect 16773 6749 16807 6783
rect 23765 6749 23799 6783
rect 24041 6749 24075 6783
rect 4215 6681 4249 6715
rect 5181 6681 5215 6715
rect 8769 6681 8803 6715
rect 14289 6681 14323 6715
rect 20453 6681 20487 6715
rect 9229 6613 9263 6647
rect 10609 6613 10643 6647
rect 18521 6613 18555 6647
rect 25375 6613 25409 6647
rect 4721 6409 4755 6443
rect 5089 6409 5123 6443
rect 6101 6409 6135 6443
rect 6653 6409 6687 6443
rect 8309 6409 8343 6443
rect 11805 6409 11839 6443
rect 12679 6409 12713 6443
rect 17049 6409 17083 6443
rect 23305 6409 23339 6443
rect 25467 6409 25501 6443
rect 26157 6409 26191 6443
rect 5273 6341 5307 6375
rect 6193 6341 6227 6375
rect 9321 6341 9355 6375
rect 16313 6341 16347 6375
rect 16773 6341 16807 6375
rect 19441 6341 19475 6375
rect 7205 6273 7239 6307
rect 7941 6273 7975 6307
rect 15393 6273 15427 6307
rect 18061 6273 18095 6307
rect 19809 6273 19843 6307
rect 24777 6341 24811 6375
rect 24133 6273 24167 6307
rect 4215 6205 4249 6239
rect 5181 6205 5215 6239
rect 5457 6205 5491 6239
rect 6101 6205 6135 6239
rect 9229 6205 9263 6239
rect 9505 6205 9539 6239
rect 10701 6205 10735 6239
rect 11437 6205 11471 6239
rect 11529 6205 11563 6239
rect 12173 6205 12207 6239
rect 12608 6205 12642 6239
rect 13553 6205 13587 6239
rect 14105 6205 14139 6239
rect 14565 6205 14599 6239
rect 16865 6205 16899 6239
rect 17325 6205 17359 6239
rect 21833 6205 21867 6239
rect 23305 6205 23339 6239
rect 23397 6205 23431 6239
rect 25396 6205 25430 6239
rect 6929 6137 6963 6171
rect 7021 6137 7055 6171
rect 9965 6137 9999 6171
rect 14289 6137 14323 6171
rect 15485 6137 15519 6171
rect 16037 6137 16071 6171
rect 18382 6137 18416 6171
rect 20130 6137 20164 6171
rect 23857 6137 23891 6171
rect 23949 6137 23983 6171
rect 3985 6069 4019 6103
rect 4307 6069 4341 6103
rect 5641 6069 5675 6103
rect 8677 6069 8711 6103
rect 9045 6069 9079 6103
rect 10333 6069 10367 6103
rect 13093 6069 13127 6103
rect 13369 6069 13403 6103
rect 15117 6069 15151 6103
rect 17693 6069 17727 6103
rect 18981 6069 19015 6103
rect 20729 6069 20763 6103
rect 21281 6069 21315 6103
rect 21649 6069 21683 6103
rect 22201 6069 22235 6103
rect 22753 6069 22787 6103
rect 23121 6069 23155 6103
rect 25789 6069 25823 6103
rect 8493 5865 8527 5899
rect 9045 5865 9079 5899
rect 10149 5865 10183 5899
rect 10701 5865 10735 5899
rect 11529 5865 11563 5899
rect 13553 5865 13587 5899
rect 15669 5865 15703 5899
rect 17601 5865 17635 5899
rect 18889 5865 18923 5899
rect 19349 5865 19383 5899
rect 19901 5865 19935 5899
rect 20269 5865 20303 5899
rect 21281 5865 21315 5899
rect 22109 5865 22143 5899
rect 22477 5865 22511 5899
rect 23121 5865 23155 5899
rect 23765 5865 23799 5899
rect 6285 5797 6319 5831
rect 7205 5797 7239 5831
rect 7573 5797 7607 5831
rect 7941 5797 7975 5831
rect 13829 5797 13863 5831
rect 17969 5797 18003 5831
rect 18061 5797 18095 5831
rect 18613 5797 18647 5831
rect 24225 5797 24259 5831
rect 24317 5797 24351 5831
rect 2973 5729 3007 5763
rect 4905 5729 4939 5763
rect 5181 5729 5215 5763
rect 6009 5729 6043 5763
rect 6469 5729 6503 5763
rect 6745 5729 6779 5763
rect 8033 5729 8067 5763
rect 8309 5729 8343 5763
rect 9689 5729 9723 5763
rect 9965 5729 9999 5763
rect 12081 5729 12115 5763
rect 12633 5729 12667 5763
rect 15301 5729 15335 5763
rect 19508 5729 19542 5763
rect 20913 5729 20947 5763
rect 21833 5729 21867 5763
rect 4813 5661 4847 5695
rect 5365 5661 5399 5695
rect 12817 5661 12851 5695
rect 13737 5661 13771 5695
rect 14381 5661 14415 5695
rect 24501 5661 24535 5695
rect 4997 5593 5031 5627
rect 6561 5593 6595 5627
rect 8125 5593 8159 5627
rect 9781 5593 9815 5627
rect 16497 5593 16531 5627
rect 3157 5525 3191 5559
rect 9413 5525 9447 5559
rect 13093 5525 13127 5559
rect 16221 5525 16255 5559
rect 19579 5525 19613 5559
rect 1685 5321 1719 5355
rect 3249 5321 3283 5355
rect 3985 5321 4019 5355
rect 4629 5321 4663 5355
rect 9321 5321 9355 5355
rect 12081 5321 12115 5355
rect 13553 5321 13587 5355
rect 13829 5321 13863 5355
rect 15209 5321 15243 5355
rect 17785 5321 17819 5355
rect 18245 5321 18279 5355
rect 19717 5321 19751 5355
rect 20085 5321 20119 5355
rect 21833 5321 21867 5355
rect 25375 5321 25409 5355
rect 25697 5321 25731 5355
rect 2881 5253 2915 5287
rect 3617 5253 3651 5287
rect 6561 5253 6595 5287
rect 8493 5253 8527 5287
rect 8769 5253 8803 5287
rect 5641 5185 5675 5219
rect 1444 5117 1478 5151
rect 1869 5117 1903 5151
rect 2697 5117 2731 5151
rect 3776 5117 3810 5151
rect 4721 5117 4755 5151
rect 5273 5117 5307 5151
rect 5768 5117 5802 5151
rect 7481 5117 7515 5151
rect 8125 5117 8159 5151
rect 4261 5049 4295 5083
rect 7389 5049 7423 5083
rect 12265 5253 12299 5287
rect 20913 5253 20947 5287
rect 24685 5253 24719 5287
rect 13553 5185 13587 5219
rect 14289 5185 14323 5219
rect 16129 5185 16163 5219
rect 18797 5185 18831 5219
rect 20361 5185 20395 5219
rect 22385 5185 22419 5219
rect 24041 5185 24075 5219
rect 8953 5117 8987 5151
rect 9597 5117 9631 5151
rect 10793 5117 10827 5151
rect 11345 5117 11379 5151
rect 12357 5117 12391 5151
rect 12725 5117 12759 5151
rect 13185 5117 13219 5151
rect 13461 5117 13495 5151
rect 25304 5117 25338 5151
rect 10149 5049 10183 5083
rect 11529 5049 11563 5083
rect 14610 5049 14644 5083
rect 15485 5049 15519 5083
rect 16221 5049 16255 5083
rect 16773 5049 16807 5083
rect 18889 5049 18923 5083
rect 19441 5049 19475 5083
rect 20453 5049 20487 5083
rect 22109 5049 22143 5083
rect 22201 5049 22235 5083
rect 23765 5049 23799 5083
rect 23857 5049 23891 5083
rect 4905 4981 4939 5015
rect 5871 4981 5905 5015
rect 8769 4981 8803 5015
rect 10701 4981 10735 5015
rect 14105 4981 14139 5015
rect 15853 4981 15887 5015
rect 21281 4981 21315 5015
rect 23397 4981 23431 5015
rect 3111 4777 3145 4811
rect 4445 4777 4479 4811
rect 4813 4777 4847 4811
rect 7941 4777 7975 4811
rect 10885 4777 10919 4811
rect 12173 4777 12207 4811
rect 12541 4777 12575 4811
rect 13553 4777 13587 4811
rect 13829 4777 13863 4811
rect 14289 4777 14323 4811
rect 15485 4777 15519 4811
rect 18337 4777 18371 4811
rect 20361 4777 20395 4811
rect 22477 4777 22511 4811
rect 24225 4777 24259 4811
rect 6285 4709 6319 4743
rect 6469 4709 6503 4743
rect 12954 4709 12988 4743
rect 16221 4709 16255 4743
rect 19165 4709 19199 4743
rect 21281 4709 21315 4743
rect 22845 4709 22879 4743
rect 24685 4709 24719 4743
rect 3008 4641 3042 4675
rect 4905 4641 4939 4675
rect 5457 4641 5491 4675
rect 7113 4641 7147 4675
rect 7573 4641 7607 4675
rect 8033 4641 8067 4675
rect 8585 4641 8619 4675
rect 9689 4641 9723 4675
rect 9965 4641 9999 4675
rect 11253 4641 11287 4675
rect 11805 4641 11839 4675
rect 14749 4641 14783 4675
rect 17693 4641 17727 4675
rect 22109 4641 22143 4675
rect 5641 4573 5675 4607
rect 8677 4573 8711 4607
rect 10425 4573 10459 4607
rect 12633 4573 12667 4607
rect 14473 4573 14507 4607
rect 16129 4573 16163 4607
rect 16405 4573 16439 4607
rect 19073 4573 19107 4607
rect 19441 4573 19475 4607
rect 21189 4573 21223 4607
rect 21465 4573 21499 4607
rect 22753 4573 22787 4607
rect 23029 4573 23063 4607
rect 24593 4573 24627 4607
rect 24869 4573 24903 4607
rect 9781 4505 9815 4539
rect 23765 4505 23799 4539
rect 9413 4437 9447 4471
rect 11437 4437 11471 4471
rect 14473 4437 14507 4471
rect 17877 4437 17911 4471
rect 18797 4437 18831 4471
rect 3617 4233 3651 4267
rect 4077 4233 4111 4267
rect 7573 4233 7607 4267
rect 9045 4233 9079 4267
rect 10701 4233 10735 4267
rect 10885 4233 10919 4267
rect 11161 4233 11195 4267
rect 11437 4233 11471 4267
rect 12909 4233 12943 4267
rect 14657 4233 14691 4267
rect 16405 4233 16439 4267
rect 17141 4233 17175 4267
rect 21189 4233 21223 4267
rect 22569 4233 22603 4267
rect 22845 4233 22879 4267
rect 25421 4233 25455 4267
rect 2973 4097 3007 4131
rect 7297 4097 7331 4131
rect 8769 4097 8803 4131
rect 3224 4029 3258 4063
rect 4236 4029 4270 4063
rect 5181 4029 5215 4063
rect 5733 4029 5767 4063
rect 7757 4029 7791 4063
rect 8217 4029 8251 4063
rect 5917 3961 5951 3995
rect 8493 3961 8527 3995
rect 9413 4165 9447 4199
rect 10333 4165 10367 4199
rect 11805 4165 11839 4199
rect 13369 4097 13403 4131
rect 9321 4029 9355 4063
rect 9597 4029 9631 4063
rect 10885 4029 10919 4063
rect 11253 4029 11287 4063
rect 12725 4029 12759 4063
rect 17785 4097 17819 4131
rect 18337 4097 18371 4131
rect 20453 4097 20487 4131
rect 21649 4097 21683 4131
rect 24777 4097 24811 4131
rect 16957 4029 16991 4063
rect 17417 4029 17451 4063
rect 19257 4029 19291 4063
rect 13921 3961 13955 3995
rect 14013 3961 14047 3995
rect 14565 3961 14599 3995
rect 14657 3961 14691 3995
rect 15485 3961 15519 3995
rect 15577 3961 15611 3995
rect 16129 3961 16163 3995
rect 20177 3961 20211 3995
rect 20269 3961 20303 3995
rect 21970 3961 22004 3995
rect 24225 3961 24259 3995
rect 24501 3961 24535 3995
rect 24593 3961 24627 3995
rect 3295 3893 3329 3927
rect 4307 3893 4341 3927
rect 4721 3893 4755 3927
rect 4997 3893 5031 3927
rect 6561 3893 6595 3927
rect 9045 3893 9079 3927
rect 9137 3893 9171 3927
rect 9781 3893 9815 3927
rect 12265 3893 12299 3927
rect 13645 3893 13679 3927
rect 14841 3893 14875 3927
rect 15301 3893 15335 3927
rect 16773 3893 16807 3927
rect 18705 3893 18739 3927
rect 19533 3893 19567 3927
rect 19993 3893 20027 3927
rect 21557 3893 21591 3927
rect 23213 3893 23247 3927
rect 23949 3893 23983 3927
rect 5917 3689 5951 3723
rect 9413 3689 9447 3723
rect 11437 3689 11471 3723
rect 12081 3689 12115 3723
rect 18613 3689 18647 3723
rect 19809 3689 19843 3723
rect 20729 3689 20763 3723
rect 22109 3689 22143 3723
rect 22661 3689 22695 3723
rect 24685 3689 24719 3723
rect 3111 3621 3145 3655
rect 8769 3621 8803 3655
rect 12627 3621 12661 3655
rect 13921 3621 13955 3655
rect 15485 3621 15519 3655
rect 20177 3621 20211 3655
rect 23857 3621 23891 3655
rect 24409 3621 24443 3655
rect 2028 3553 2062 3587
rect 2973 3553 3007 3587
rect 5181 3553 5215 3587
rect 5457 3553 5491 3587
rect 7021 3553 7055 3587
rect 7205 3553 7239 3587
rect 7297 3553 7331 3587
rect 8033 3553 8067 3587
rect 8309 3553 8343 3587
rect 9689 3553 9723 3587
rect 9965 3553 9999 3587
rect 11253 3553 11287 3587
rect 11713 3553 11747 3587
rect 14105 3553 14139 3587
rect 15025 3553 15059 3587
rect 17141 3553 17175 3587
rect 18245 3553 18279 3587
rect 19165 3553 19199 3587
rect 4813 3485 4847 3519
rect 5641 3485 5675 3519
rect 2099 3417 2133 3451
rect 10149 3485 10183 3519
rect 12265 3485 12299 3519
rect 13461 3485 13495 3519
rect 15393 3485 15427 3519
rect 15669 3485 15703 3519
rect 21741 3485 21775 3519
rect 23765 3485 23799 3519
rect 25237 3485 25271 3519
rect 7941 3417 7975 3451
rect 8125 3417 8159 3451
rect 9781 3417 9815 3451
rect 10885 3417 10919 3451
rect 17325 3417 17359 3451
rect 7297 3349 7331 3383
rect 7573 3349 7607 3383
rect 13185 3349 13219 3383
rect 14289 3349 14323 3383
rect 14657 3349 14691 3383
rect 16313 3349 16347 3383
rect 17693 3349 17727 3383
rect 19441 3349 19475 3383
rect 21281 3349 21315 3383
rect 2283 3145 2317 3179
rect 3985 3145 4019 3179
rect 4353 3145 4387 3179
rect 6285 3145 6319 3179
rect 6653 3145 6687 3179
rect 9137 3145 9171 3179
rect 14105 3145 14139 3179
rect 15393 3145 15427 3179
rect 17141 3145 17175 3179
rect 18797 3145 18831 3179
rect 20821 3145 20855 3179
rect 24685 3145 24719 3179
rect 25375 3145 25409 3179
rect 5273 3077 5307 3111
rect 7389 3077 7423 3111
rect 13369 3077 13403 3111
rect 15117 3077 15151 3111
rect 15761 3077 15795 3111
rect 18337 3077 18371 3111
rect 4721 3009 4755 3043
rect 10885 3009 10919 3043
rect 11529 3009 11563 3043
rect 12449 3009 12483 3043
rect 14197 3009 14231 3043
rect 16037 3009 16071 3043
rect 16313 3009 16347 3043
rect 23029 3009 23063 3043
rect 23489 3009 23523 3043
rect 23765 3009 23799 3043
rect 24225 3009 24259 3043
rect 2212 2941 2246 2975
rect 4169 2941 4203 2975
rect 5181 2941 5215 2975
rect 5457 2941 5491 2975
rect 7297 2941 7331 2975
rect 7573 2941 7607 2975
rect 8401 2941 8435 2975
rect 8953 2941 8987 2975
rect 10241 2941 10275 2975
rect 11897 2941 11931 2975
rect 12265 2941 12299 2975
rect 18153 2941 18187 2975
rect 19257 2941 19291 2975
rect 21281 2941 21315 2975
rect 22201 2941 22235 2975
rect 25304 2941 25338 2975
rect 3065 2873 3099 2907
rect 5089 2873 5123 2907
rect 7205 2873 7239 2907
rect 10609 2873 10643 2907
rect 10977 2873 11011 2907
rect 12811 2873 12845 2907
rect 14518 2873 14552 2907
rect 16129 2873 16163 2907
rect 19578 2873 19612 2907
rect 21097 2873 21131 2907
rect 21602 2873 21636 2907
rect 22477 2873 22511 2907
rect 23857 2873 23891 2907
rect 2053 2805 2087 2839
rect 2605 2805 2639 2839
rect 3157 2805 3191 2839
rect 5641 2805 5675 2839
rect 7757 2805 7791 2839
rect 8677 2805 8711 2839
rect 9873 2805 9907 2839
rect 13645 2805 13679 2839
rect 17785 2805 17819 2839
rect 19073 2805 19107 2839
rect 20177 2805 20211 2839
rect 25789 2805 25823 2839
rect 2099 2601 2133 2635
rect 4721 2601 4755 2635
rect 4997 2601 5031 2635
rect 5365 2601 5399 2635
rect 6009 2601 6043 2635
rect 6377 2601 6411 2635
rect 7665 2601 7699 2635
rect 9137 2601 9171 2635
rect 10057 2601 10091 2635
rect 12265 2601 12299 2635
rect 16865 2601 16899 2635
rect 18981 2601 19015 2635
rect 21327 2601 21361 2635
rect 21741 2601 21775 2635
rect 5733 2533 5767 2567
rect 8861 2533 8895 2567
rect 9597 2533 9631 2567
rect 11161 2533 11195 2567
rect 11713 2533 11747 2567
rect 13737 2533 13771 2567
rect 14013 2533 14047 2567
rect 14565 2533 14599 2567
rect 15209 2533 15243 2567
rect 15945 2533 15979 2567
rect 16497 2533 16531 2567
rect 19441 2533 19475 2567
rect 19717 2533 19751 2567
rect 22017 2533 22051 2567
rect 22293 2533 22327 2567
rect 22385 2533 22419 2567
rect 22937 2533 22971 2567
rect 23673 2533 23707 2567
rect 24501 2533 24535 2567
rect 25329 2533 25363 2567
rect 2028 2465 2062 2499
rect 3040 2465 3074 2499
rect 4353 2465 4387 2499
rect 4813 2465 4847 2499
rect 5825 2465 5859 2499
rect 7113 2465 7147 2499
rect 8033 2465 8067 2499
rect 8769 2465 8803 2499
rect 9873 2465 9907 2499
rect 10425 2465 10459 2499
rect 10885 2465 10919 2499
rect 12725 2465 12759 2499
rect 13277 2465 13311 2499
rect 18153 2465 18187 2499
rect 18429 2465 18463 2499
rect 21256 2465 21290 2499
rect 11069 2397 11103 2431
rect 13921 2397 13955 2431
rect 14933 2397 14967 2431
rect 15853 2397 15887 2431
rect 19625 2397 19659 2431
rect 20545 2397 20579 2431
rect 23213 2397 23247 2431
rect 24409 2397 24443 2431
rect 25697 2397 25731 2431
rect 7297 2329 7331 2363
rect 18613 2329 18647 2363
rect 20177 2329 20211 2363
rect 24961 2329 24995 2363
rect 2513 2261 2547 2295
rect 3111 2261 3145 2295
rect 3525 2261 3559 2295
rect 12909 2261 12943 2295
<< metal1 >>
rect 2222 27480 2228 27532
rect 2280 27520 2286 27532
rect 3418 27520 3424 27532
rect 2280 27492 3424 27520
rect 2280 27480 2286 27492
rect 3418 27480 3424 27492
rect 3476 27480 3482 27532
rect 14366 27480 14372 27532
rect 14424 27520 14430 27532
rect 16206 27520 16212 27532
rect 14424 27492 16212 27520
rect 14424 27480 14430 27492
rect 16206 27480 16212 27492
rect 16264 27480 16270 27532
rect 750 26732 756 26784
rect 808 26772 814 26784
rect 2774 26772 2780 26784
rect 808 26744 2780 26772
rect 808 26732 814 26744
rect 2774 26732 2780 26744
rect 2832 26732 2838 26784
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 24765 24939 24823 24945
rect 24765 24905 24777 24939
rect 24811 24936 24823 24939
rect 27154 24936 27160 24948
rect 24811 24908 27160 24936
rect 24811 24905 24823 24908
rect 24765 24899 24823 24905
rect 27154 24896 27160 24908
rect 27212 24896 27218 24948
rect 24118 24692 24124 24744
rect 24176 24732 24182 24744
rect 24581 24735 24639 24741
rect 24581 24732 24593 24735
rect 24176 24704 24593 24732
rect 24176 24692 24182 24704
rect 24581 24701 24593 24704
rect 24627 24732 24639 24735
rect 25133 24735 25191 24741
rect 25133 24732 25145 24735
rect 24627 24704 25145 24732
rect 24627 24701 24639 24704
rect 24581 24695 24639 24701
rect 25133 24701 25145 24704
rect 25179 24701 25191 24735
rect 25133 24695 25191 24701
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 24762 24392 24768 24404
rect 24723 24364 24768 24392
rect 24762 24352 24768 24364
rect 24820 24352 24826 24404
rect 23477 24259 23535 24265
rect 23477 24225 23489 24259
rect 23523 24256 23535 24259
rect 23842 24256 23848 24268
rect 23523 24228 23848 24256
rect 23523 24225 23535 24228
rect 23477 24219 23535 24225
rect 23842 24216 23848 24228
rect 23900 24216 23906 24268
rect 24581 24259 24639 24265
rect 24581 24225 24593 24259
rect 24627 24256 24639 24259
rect 24670 24256 24676 24268
rect 24627 24228 24676 24256
rect 24627 24225 24639 24228
rect 24581 24219 24639 24225
rect 24670 24216 24676 24228
rect 24728 24216 24734 24268
rect 23661 24123 23719 24129
rect 23661 24089 23673 24123
rect 23707 24120 23719 24123
rect 25590 24120 25596 24132
rect 23707 24092 25596 24120
rect 23707 24089 23719 24092
rect 23661 24083 23719 24089
rect 25590 24080 25596 24092
rect 25648 24080 25654 24132
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 14001 23851 14059 23857
rect 14001 23817 14013 23851
rect 14047 23848 14059 23851
rect 14734 23848 14740 23860
rect 14047 23820 14740 23848
rect 14047 23817 14059 23820
rect 14001 23811 14059 23817
rect 14734 23808 14740 23820
rect 14792 23808 14798 23860
rect 16577 23851 16635 23857
rect 16577 23817 16589 23851
rect 16623 23848 16635 23851
rect 17770 23848 17776 23860
rect 16623 23820 17776 23848
rect 16623 23817 16635 23820
rect 16577 23811 16635 23817
rect 17770 23808 17776 23820
rect 17828 23808 17834 23860
rect 18325 23851 18383 23857
rect 18325 23817 18337 23851
rect 18371 23848 18383 23851
rect 19334 23848 19340 23860
rect 18371 23820 19340 23848
rect 18371 23817 18383 23820
rect 18325 23811 18383 23817
rect 19334 23808 19340 23820
rect 19392 23808 19398 23860
rect 19429 23851 19487 23857
rect 19429 23817 19441 23851
rect 19475 23848 19487 23851
rect 20898 23848 20904 23860
rect 19475 23820 20904 23848
rect 19475 23817 19487 23820
rect 19429 23811 19487 23817
rect 20898 23808 20904 23820
rect 20956 23808 20962 23860
rect 22189 23851 22247 23857
rect 22189 23817 22201 23851
rect 22235 23848 22247 23851
rect 24026 23848 24032 23860
rect 22235 23820 24032 23848
rect 22235 23817 22247 23820
rect 22189 23811 22247 23817
rect 24026 23808 24032 23820
rect 24084 23808 24090 23860
rect 24765 23851 24823 23857
rect 24765 23817 24777 23851
rect 24811 23848 24823 23851
rect 24946 23848 24952 23860
rect 24811 23820 24952 23848
rect 24811 23817 24823 23820
rect 24765 23811 24823 23817
rect 24946 23808 24952 23820
rect 25004 23808 25010 23860
rect 20625 23783 20683 23789
rect 20625 23749 20637 23783
rect 20671 23780 20683 23783
rect 22462 23780 22468 23792
rect 20671 23752 22468 23780
rect 20671 23749 20683 23752
rect 20625 23743 20683 23749
rect 22462 23740 22468 23752
rect 22520 23740 22526 23792
rect 23842 23780 23848 23792
rect 23803 23752 23848 23780
rect 23842 23740 23848 23752
rect 23900 23740 23906 23792
rect 1448 23647 1506 23653
rect 1448 23613 1460 23647
rect 1494 23644 1506 23647
rect 1854 23644 1860 23656
rect 1494 23616 1860 23644
rect 1494 23613 1506 23616
rect 1448 23607 1506 23613
rect 1854 23604 1860 23616
rect 1912 23604 1918 23656
rect 12710 23604 12716 23656
rect 12768 23644 12774 23656
rect 13817 23647 13875 23653
rect 13817 23644 13829 23647
rect 12768 23616 13829 23644
rect 12768 23604 12774 23616
rect 13817 23613 13829 23616
rect 13863 23644 13875 23647
rect 14369 23647 14427 23653
rect 14369 23644 14381 23647
rect 13863 23616 14381 23644
rect 13863 23613 13875 23616
rect 13817 23607 13875 23613
rect 14369 23613 14381 23616
rect 14415 23613 14427 23647
rect 14369 23607 14427 23613
rect 15378 23604 15384 23656
rect 15436 23644 15442 23656
rect 16393 23647 16451 23653
rect 16393 23644 16405 23647
rect 15436 23616 16405 23644
rect 15436 23604 15442 23616
rect 16393 23613 16405 23616
rect 16439 23644 16451 23647
rect 16945 23647 17003 23653
rect 16945 23644 16957 23647
rect 16439 23616 16957 23644
rect 16439 23613 16451 23616
rect 16393 23607 16451 23613
rect 16945 23613 16957 23616
rect 16991 23613 17003 23647
rect 16945 23607 17003 23613
rect 17218 23604 17224 23656
rect 17276 23644 17282 23656
rect 18141 23647 18199 23653
rect 18141 23644 18153 23647
rect 17276 23616 18153 23644
rect 17276 23604 17282 23616
rect 18141 23613 18153 23616
rect 18187 23644 18199 23647
rect 18693 23647 18751 23653
rect 18693 23644 18705 23647
rect 18187 23616 18705 23644
rect 18187 23613 18199 23616
rect 18141 23607 18199 23613
rect 18693 23613 18705 23616
rect 18739 23613 18751 23647
rect 18693 23607 18751 23613
rect 19245 23647 19303 23653
rect 19245 23613 19257 23647
rect 19291 23644 19303 23647
rect 19518 23644 19524 23656
rect 19291 23616 19524 23644
rect 19291 23613 19303 23616
rect 19245 23607 19303 23613
rect 19518 23604 19524 23616
rect 19576 23644 19582 23656
rect 19797 23647 19855 23653
rect 19797 23644 19809 23647
rect 19576 23616 19809 23644
rect 19576 23604 19582 23616
rect 19797 23613 19809 23616
rect 19843 23613 19855 23647
rect 19797 23607 19855 23613
rect 20441 23647 20499 23653
rect 20441 23613 20453 23647
rect 20487 23613 20499 23647
rect 22002 23644 22008 23656
rect 21915 23616 22008 23644
rect 20441 23607 20499 23613
rect 1535 23579 1593 23585
rect 1535 23545 1547 23579
rect 1581 23576 1593 23579
rect 7098 23576 7104 23588
rect 1581 23548 7104 23576
rect 1581 23545 1593 23548
rect 1535 23539 1593 23545
rect 7098 23536 7104 23548
rect 7156 23536 7162 23588
rect 19334 23536 19340 23588
rect 19392 23576 19398 23588
rect 20456 23576 20484 23607
rect 22002 23604 22008 23616
rect 22060 23644 22066 23656
rect 22557 23647 22615 23653
rect 22557 23644 22569 23647
rect 22060 23616 22569 23644
rect 22060 23604 22066 23616
rect 22557 23613 22569 23616
rect 22603 23613 22615 23647
rect 22557 23607 22615 23613
rect 20993 23579 21051 23585
rect 20993 23576 21005 23579
rect 19392 23548 21005 23576
rect 19392 23536 19398 23548
rect 20993 23545 21005 23548
rect 21039 23545 21051 23579
rect 20993 23539 21051 23545
rect 22646 23536 22652 23588
rect 22704 23576 22710 23588
rect 24670 23576 24676 23588
rect 22704 23548 24676 23576
rect 22704 23536 22710 23548
rect 24670 23536 24676 23548
rect 24728 23576 24734 23588
rect 25133 23579 25191 23585
rect 25133 23576 25145 23579
rect 24728 23548 25145 23576
rect 24728 23536 24734 23548
rect 25133 23545 25145 23548
rect 25179 23545 25191 23579
rect 25133 23539 25191 23545
rect 22738 23468 22744 23520
rect 22796 23508 22802 23520
rect 23842 23508 23848 23520
rect 22796 23480 23848 23508
rect 22796 23468 22802 23480
rect 23842 23468 23848 23480
rect 23900 23468 23906 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 24762 23304 24768 23316
rect 24723 23276 24768 23304
rect 24762 23264 24768 23276
rect 24820 23264 24826 23316
rect 24026 23128 24032 23180
rect 24084 23168 24090 23180
rect 24581 23171 24639 23177
rect 24581 23168 24593 23171
rect 24084 23140 24593 23168
rect 24084 23128 24090 23140
rect 24581 23137 24593 23140
rect 24627 23137 24639 23171
rect 24581 23131 24639 23137
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 24026 22380 24032 22432
rect 24084 22420 24090 22432
rect 24581 22423 24639 22429
rect 24581 22420 24593 22423
rect 24084 22392 24593 22420
rect 24084 22380 24090 22392
rect 24581 22389 24593 22392
rect 24627 22389 24639 22423
rect 24581 22383 24639 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 24762 22216 24768 22228
rect 24723 22188 24768 22216
rect 24762 22176 24768 22188
rect 24820 22176 24826 22228
rect 7098 22108 7104 22160
rect 7156 22148 7162 22160
rect 11974 22148 11980 22160
rect 7156 22120 11980 22148
rect 7156 22108 7162 22120
rect 11974 22108 11980 22120
rect 12032 22108 12038 22160
rect 9582 22080 9588 22092
rect 9543 22052 9588 22080
rect 9582 22040 9588 22052
rect 9640 22040 9646 22092
rect 24210 22040 24216 22092
rect 24268 22080 24274 22092
rect 24581 22083 24639 22089
rect 24581 22080 24593 22083
rect 24268 22052 24593 22080
rect 24268 22040 24274 22052
rect 24581 22049 24593 22052
rect 24627 22049 24639 22083
rect 24581 22043 24639 22049
rect 9815 21879 9873 21885
rect 9815 21845 9827 21879
rect 9861 21876 9873 21879
rect 18598 21876 18604 21888
rect 9861 21848 18604 21876
rect 9861 21845 9873 21848
rect 9815 21839 9873 21845
rect 18598 21836 18604 21848
rect 18656 21836 18662 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 14369 21675 14427 21681
rect 14369 21641 14381 21675
rect 14415 21672 14427 21675
rect 14734 21672 14740 21684
rect 14415 21644 14740 21672
rect 14415 21641 14427 21644
rect 14369 21635 14427 21641
rect 8938 21428 8944 21480
rect 8996 21468 9002 21480
rect 9376 21471 9434 21477
rect 9376 21468 9388 21471
rect 8996 21440 9388 21468
rect 8996 21428 9002 21440
rect 9376 21437 9388 21440
rect 9422 21468 9434 21471
rect 9769 21471 9827 21477
rect 9769 21468 9781 21471
rect 9422 21440 9781 21468
rect 9422 21437 9434 21440
rect 9376 21431 9434 21437
rect 9769 21437 9781 21440
rect 9815 21437 9827 21471
rect 9769 21431 9827 21437
rect 13884 21471 13942 21477
rect 13884 21437 13896 21471
rect 13930 21468 13942 21471
rect 14384 21468 14412 21635
rect 14734 21632 14740 21644
rect 14792 21672 14798 21684
rect 22002 21672 22008 21684
rect 14792 21644 22008 21672
rect 14792 21632 14798 21644
rect 22002 21632 22008 21644
rect 22060 21632 22066 21684
rect 13930 21440 14412 21468
rect 13930 21437 13942 21440
rect 13884 21431 13942 21437
rect 8570 21360 8576 21412
rect 8628 21400 8634 21412
rect 9582 21400 9588 21412
rect 8628 21372 9588 21400
rect 8628 21360 8634 21372
rect 9582 21360 9588 21372
rect 9640 21400 9646 21412
rect 10137 21403 10195 21409
rect 10137 21400 10149 21403
rect 9640 21372 10149 21400
rect 9640 21360 9646 21372
rect 10137 21369 10149 21372
rect 10183 21369 10195 21403
rect 10137 21363 10195 21369
rect 9447 21335 9505 21341
rect 9447 21301 9459 21335
rect 9493 21332 9505 21335
rect 10042 21332 10048 21344
rect 9493 21304 10048 21332
rect 9493 21301 9505 21304
rect 9447 21295 9505 21301
rect 10042 21292 10048 21304
rect 10100 21292 10106 21344
rect 13955 21335 14013 21341
rect 13955 21301 13967 21335
rect 14001 21332 14013 21335
rect 14090 21332 14096 21344
rect 14001 21304 14096 21332
rect 14001 21301 14013 21304
rect 13955 21295 14013 21301
rect 14090 21292 14096 21304
rect 14148 21292 14154 21344
rect 24210 21292 24216 21344
rect 24268 21332 24274 21344
rect 24581 21335 24639 21341
rect 24581 21332 24593 21335
rect 24268 21304 24593 21332
rect 24268 21292 24274 21304
rect 24581 21301 24593 21304
rect 24627 21301 24639 21335
rect 24581 21295 24639 21301
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 4801 20995 4859 21001
rect 4801 20961 4813 20995
rect 4847 20992 4859 20995
rect 4890 20992 4896 21004
rect 4847 20964 4896 20992
rect 4847 20961 4859 20964
rect 4801 20955 4859 20961
rect 4890 20952 4896 20964
rect 4948 20952 4954 21004
rect 11400 20995 11458 21001
rect 11400 20961 11412 20995
rect 11446 20992 11458 20995
rect 11606 20992 11612 21004
rect 11446 20964 11612 20992
rect 11446 20961 11458 20964
rect 11400 20955 11458 20961
rect 11606 20952 11612 20964
rect 11664 20952 11670 21004
rect 12872 20995 12930 21001
rect 12872 20961 12884 20995
rect 12918 20992 12930 20995
rect 13170 20992 13176 21004
rect 12918 20964 13176 20992
rect 12918 20961 12930 20964
rect 12872 20955 12930 20961
rect 13170 20952 13176 20964
rect 13228 20952 13234 21004
rect 10134 20884 10140 20936
rect 10192 20924 10198 20936
rect 10321 20927 10379 20933
rect 10321 20924 10333 20927
rect 10192 20896 10333 20924
rect 10192 20884 10198 20896
rect 10321 20893 10333 20896
rect 10367 20893 10379 20927
rect 10321 20887 10379 20893
rect 13630 20884 13636 20936
rect 13688 20924 13694 20936
rect 14001 20927 14059 20933
rect 14001 20924 14013 20927
rect 13688 20896 14013 20924
rect 13688 20884 13694 20896
rect 14001 20893 14013 20896
rect 14047 20893 14059 20927
rect 14001 20887 14059 20893
rect 4706 20748 4712 20800
rect 4764 20788 4770 20800
rect 5031 20791 5089 20797
rect 5031 20788 5043 20791
rect 4764 20760 5043 20788
rect 4764 20748 4770 20760
rect 5031 20757 5043 20760
rect 5077 20757 5089 20791
rect 5031 20751 5089 20757
rect 10686 20748 10692 20800
rect 10744 20788 10750 20800
rect 10873 20791 10931 20797
rect 10873 20788 10885 20791
rect 10744 20760 10885 20788
rect 10744 20748 10750 20760
rect 10873 20757 10885 20760
rect 10919 20788 10931 20791
rect 11471 20791 11529 20797
rect 11471 20788 11483 20791
rect 10919 20760 11483 20788
rect 10919 20757 10931 20760
rect 10873 20751 10931 20757
rect 11471 20757 11483 20760
rect 11517 20757 11529 20791
rect 11471 20751 11529 20757
rect 12943 20791 13001 20797
rect 12943 20757 12955 20791
rect 12989 20788 13001 20791
rect 13446 20788 13452 20800
rect 12989 20760 13452 20788
rect 12989 20757 13001 20760
rect 12943 20751 13001 20757
rect 13446 20748 13452 20760
rect 13504 20748 13510 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 4890 20584 4896 20596
rect 4851 20556 4896 20584
rect 4890 20544 4896 20556
rect 4948 20544 4954 20596
rect 11606 20584 11612 20596
rect 11567 20556 11612 20584
rect 11606 20544 11612 20556
rect 11664 20544 11670 20596
rect 13170 20544 13176 20596
rect 13228 20584 13234 20596
rect 13265 20587 13323 20593
rect 13265 20584 13277 20587
rect 13228 20556 13277 20584
rect 13228 20544 13234 20556
rect 13265 20553 13277 20556
rect 13311 20553 13323 20587
rect 13265 20547 13323 20553
rect 10686 20448 10692 20460
rect 10647 20420 10692 20448
rect 10686 20408 10692 20420
rect 10744 20408 10750 20460
rect 4430 20340 4436 20392
rect 4488 20380 4494 20392
rect 9620 20383 9678 20389
rect 9620 20380 9632 20383
rect 4488 20352 9632 20380
rect 4488 20340 4494 20352
rect 9620 20349 9632 20352
rect 9666 20380 9678 20383
rect 10045 20383 10103 20389
rect 10045 20380 10057 20383
rect 9666 20352 10057 20380
rect 9666 20349 9678 20352
rect 9620 20343 9678 20349
rect 10045 20349 10057 20352
rect 10091 20380 10103 20383
rect 10226 20380 10232 20392
rect 10091 20352 10232 20380
rect 10091 20349 10103 20352
rect 10045 20343 10103 20349
rect 10226 20340 10232 20352
rect 10284 20340 10290 20392
rect 12840 20383 12898 20389
rect 12840 20380 12852 20383
rect 12636 20352 12852 20380
rect 10781 20315 10839 20321
rect 10781 20312 10793 20315
rect 10704 20284 10793 20312
rect 10704 20256 10732 20284
rect 10781 20281 10793 20284
rect 10827 20281 10839 20315
rect 10781 20275 10839 20281
rect 11333 20315 11391 20321
rect 11333 20281 11345 20315
rect 11379 20312 11391 20315
rect 11698 20312 11704 20324
rect 11379 20284 11704 20312
rect 11379 20281 11391 20284
rect 11333 20275 11391 20281
rect 11698 20272 11704 20284
rect 11756 20272 11762 20324
rect 9723 20247 9781 20253
rect 9723 20213 9735 20247
rect 9769 20244 9781 20247
rect 9950 20244 9956 20256
rect 9769 20216 9956 20244
rect 9769 20213 9781 20216
rect 9723 20207 9781 20213
rect 9950 20204 9956 20216
rect 10008 20204 10014 20256
rect 10505 20247 10563 20253
rect 10505 20213 10517 20247
rect 10551 20244 10563 20247
rect 10686 20244 10692 20256
rect 10551 20216 10692 20244
rect 10551 20213 10563 20216
rect 10505 20207 10563 20213
rect 10686 20204 10692 20216
rect 10744 20204 10750 20256
rect 12250 20204 12256 20256
rect 12308 20244 12314 20256
rect 12636 20253 12664 20352
rect 12840 20349 12852 20352
rect 12886 20349 12898 20383
rect 13722 20380 13728 20392
rect 13635 20352 13728 20380
rect 12840 20343 12898 20349
rect 13722 20340 13728 20352
rect 13780 20380 13786 20392
rect 13909 20383 13967 20389
rect 13909 20380 13921 20383
rect 13780 20352 13921 20380
rect 13780 20340 13786 20352
rect 13909 20349 13921 20352
rect 13955 20349 13967 20383
rect 13909 20343 13967 20349
rect 15286 20340 15292 20392
rect 15344 20380 15350 20392
rect 15448 20383 15506 20389
rect 15448 20380 15460 20383
rect 15344 20352 15460 20380
rect 15344 20340 15350 20352
rect 15448 20349 15460 20352
rect 15494 20380 15506 20383
rect 15494 20352 15884 20380
rect 15494 20349 15506 20352
rect 15448 20343 15506 20349
rect 13814 20272 13820 20324
rect 13872 20312 13878 20324
rect 13872 20284 13917 20312
rect 13872 20272 13878 20284
rect 15856 20256 15884 20352
rect 12621 20247 12679 20253
rect 12621 20244 12633 20247
rect 12308 20216 12633 20244
rect 12308 20204 12314 20216
rect 12621 20213 12633 20216
rect 12667 20213 12679 20247
rect 12621 20207 12679 20213
rect 12943 20247 13001 20253
rect 12943 20213 12955 20247
rect 12989 20244 13001 20247
rect 13354 20244 13360 20256
rect 12989 20216 13360 20244
rect 12989 20213 13001 20216
rect 12943 20207 13001 20213
rect 13354 20204 13360 20216
rect 13412 20204 13418 20256
rect 14642 20204 14648 20256
rect 14700 20244 14706 20256
rect 15519 20247 15577 20253
rect 15519 20244 15531 20247
rect 14700 20216 15531 20244
rect 14700 20204 14706 20216
rect 15519 20213 15531 20216
rect 15565 20213 15577 20247
rect 15838 20244 15844 20256
rect 15799 20216 15844 20244
rect 15519 20207 15577 20213
rect 15838 20204 15844 20216
rect 15896 20204 15902 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 13446 20040 13452 20052
rect 13407 20012 13452 20040
rect 13446 20000 13452 20012
rect 13504 20040 13510 20052
rect 24765 20043 24823 20049
rect 13504 20012 13768 20040
rect 13504 20000 13510 20012
rect 10226 19972 10232 19984
rect 10187 19944 10232 19972
rect 10226 19932 10232 19944
rect 10284 19932 10290 19984
rect 11793 19975 11851 19981
rect 11793 19941 11805 19975
rect 11839 19972 11851 19975
rect 11882 19972 11888 19984
rect 11839 19944 11888 19972
rect 11839 19941 11851 19944
rect 11793 19935 11851 19941
rect 11882 19932 11888 19944
rect 11940 19932 11946 19984
rect 13740 19981 13768 20012
rect 24765 20009 24777 20043
rect 24811 20040 24823 20043
rect 25222 20040 25228 20052
rect 24811 20012 25228 20040
rect 24811 20009 24823 20012
rect 24765 20003 24823 20009
rect 25222 20000 25228 20012
rect 25280 20000 25286 20052
rect 13725 19975 13783 19981
rect 13725 19941 13737 19975
rect 13771 19941 13783 19975
rect 13725 19935 13783 19941
rect 13814 19932 13820 19984
rect 13872 19972 13878 19984
rect 13872 19944 13917 19972
rect 13872 19932 13878 19944
rect 15930 19904 15936 19916
rect 15891 19876 15936 19904
rect 15930 19864 15936 19876
rect 15988 19864 15994 19916
rect 24581 19907 24639 19913
rect 24581 19873 24593 19907
rect 24627 19904 24639 19907
rect 24670 19904 24676 19916
rect 24627 19876 24676 19904
rect 24627 19873 24639 19876
rect 24581 19867 24639 19873
rect 24670 19864 24676 19876
rect 24728 19864 24734 19916
rect 10137 19839 10195 19845
rect 10137 19805 10149 19839
rect 10183 19805 10195 19839
rect 10137 19799 10195 19805
rect 10781 19839 10839 19845
rect 10781 19805 10793 19839
rect 10827 19836 10839 19839
rect 11698 19836 11704 19848
rect 10827 19808 11704 19836
rect 10827 19805 10839 19808
rect 10781 19799 10839 19805
rect 9953 19703 10011 19709
rect 9953 19669 9965 19703
rect 9999 19700 10011 19703
rect 10042 19700 10048 19712
rect 9999 19672 10048 19700
rect 9999 19669 10011 19672
rect 9953 19663 10011 19669
rect 10042 19660 10048 19672
rect 10100 19700 10106 19712
rect 10152 19700 10180 19799
rect 11698 19796 11704 19808
rect 11756 19796 11762 19848
rect 14369 19839 14427 19845
rect 14369 19805 14381 19839
rect 14415 19836 14427 19839
rect 14458 19836 14464 19848
rect 14415 19808 14464 19836
rect 14415 19805 14427 19808
rect 14369 19799 14427 19805
rect 14458 19796 14464 19808
rect 14516 19796 14522 19848
rect 15286 19836 15292 19848
rect 15247 19808 15292 19836
rect 15286 19796 15292 19808
rect 15344 19796 15350 19848
rect 12250 19768 12256 19780
rect 12211 19740 12256 19768
rect 12250 19728 12256 19740
rect 12308 19728 12314 19780
rect 10100 19672 10180 19700
rect 10100 19660 10106 19672
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 10134 19456 10140 19508
rect 10192 19496 10198 19508
rect 10229 19499 10287 19505
rect 10229 19496 10241 19499
rect 10192 19468 10241 19496
rect 10192 19456 10198 19468
rect 10229 19465 10241 19468
rect 10275 19496 10287 19499
rect 10275 19468 10916 19496
rect 10275 19465 10287 19468
rect 10229 19459 10287 19465
rect 9953 19363 10011 19369
rect 9953 19329 9965 19363
rect 9999 19360 10011 19363
rect 10597 19363 10655 19369
rect 10597 19360 10609 19363
rect 9999 19332 10609 19360
rect 9999 19329 10011 19332
rect 9953 19323 10011 19329
rect 10597 19329 10609 19332
rect 10643 19360 10655 19363
rect 10686 19360 10692 19372
rect 10643 19332 10692 19360
rect 10643 19329 10655 19332
rect 10597 19323 10655 19329
rect 9125 19295 9183 19301
rect 9125 19261 9137 19295
rect 9171 19292 9183 19295
rect 9309 19295 9367 19301
rect 9309 19292 9321 19295
rect 9171 19264 9321 19292
rect 9171 19261 9183 19264
rect 9125 19255 9183 19261
rect 9309 19261 9321 19264
rect 9355 19292 9367 19295
rect 10226 19292 10232 19304
rect 9355 19264 10232 19292
rect 9355 19261 9367 19264
rect 9309 19255 9367 19261
rect 10226 19252 10232 19264
rect 10284 19252 10290 19304
rect 10612 19224 10640 19323
rect 10686 19320 10692 19332
rect 10744 19320 10750 19372
rect 10888 19369 10916 19468
rect 11698 19456 11704 19508
rect 11756 19496 11762 19508
rect 12621 19499 12679 19505
rect 12621 19496 12633 19499
rect 11756 19468 12633 19496
rect 11756 19456 11762 19468
rect 12621 19465 12633 19468
rect 12667 19465 12679 19499
rect 12621 19459 12679 19465
rect 13265 19499 13323 19505
rect 13265 19465 13277 19499
rect 13311 19496 13323 19499
rect 13538 19496 13544 19508
rect 13311 19468 13544 19496
rect 13311 19465 13323 19468
rect 13265 19459 13323 19465
rect 13538 19456 13544 19468
rect 13596 19496 13602 19508
rect 13814 19496 13820 19508
rect 13596 19468 13820 19496
rect 13596 19456 13602 19468
rect 13814 19456 13820 19468
rect 13872 19496 13878 19508
rect 14369 19499 14427 19505
rect 14369 19496 14381 19499
rect 13872 19468 14381 19496
rect 13872 19456 13878 19468
rect 14369 19465 14381 19468
rect 14415 19465 14427 19499
rect 15930 19496 15936 19508
rect 15891 19468 15936 19496
rect 14369 19459 14427 19465
rect 15930 19456 15936 19468
rect 15988 19456 15994 19508
rect 10873 19363 10931 19369
rect 10873 19329 10885 19363
rect 10919 19329 10931 19363
rect 10873 19323 10931 19329
rect 13449 19363 13507 19369
rect 13449 19329 13461 19363
rect 13495 19360 13507 19363
rect 13630 19360 13636 19372
rect 13495 19332 13636 19360
rect 13495 19329 13507 19332
rect 13449 19323 13507 19329
rect 13630 19320 13636 19332
rect 13688 19320 13694 19372
rect 16623 19363 16681 19369
rect 16623 19329 16635 19363
rect 16669 19360 16681 19363
rect 24581 19363 24639 19369
rect 24581 19360 24593 19363
rect 16669 19332 24593 19360
rect 16669 19329 16681 19332
rect 16623 19323 16681 19329
rect 24581 19329 24593 19332
rect 24627 19360 24639 19363
rect 24670 19360 24676 19372
rect 24627 19332 24676 19360
rect 24627 19329 24639 19332
rect 24581 19323 24639 19329
rect 24670 19320 24676 19332
rect 24728 19320 24734 19372
rect 16520 19295 16578 19301
rect 16520 19292 16532 19295
rect 15672 19264 16532 19292
rect 15672 19236 15700 19264
rect 16520 19261 16532 19264
rect 16566 19292 16578 19295
rect 16945 19295 17003 19301
rect 16945 19292 16957 19295
rect 16566 19264 16957 19292
rect 16566 19261 16578 19264
rect 16520 19255 16578 19261
rect 16945 19261 16957 19264
rect 16991 19261 17003 19295
rect 16945 19255 17003 19261
rect 10965 19227 11023 19233
rect 10965 19224 10977 19227
rect 10612 19196 10977 19224
rect 10965 19193 10977 19196
rect 11011 19193 11023 19227
rect 10965 19187 11023 19193
rect 11517 19227 11575 19233
rect 11517 19193 11529 19227
rect 11563 19224 11575 19227
rect 11606 19224 11612 19236
rect 11563 19196 11612 19224
rect 11563 19193 11575 19196
rect 11517 19187 11575 19193
rect 11606 19184 11612 19196
rect 11664 19184 11670 19236
rect 13538 19184 13544 19236
rect 13596 19224 13602 19236
rect 14093 19227 14151 19233
rect 13596 19196 13641 19224
rect 13596 19184 13602 19196
rect 14093 19193 14105 19227
rect 14139 19224 14151 19227
rect 15010 19224 15016 19236
rect 14139 19196 15016 19224
rect 14139 19193 14151 19196
rect 14093 19187 14151 19193
rect 15010 19184 15016 19196
rect 15068 19184 15074 19236
rect 15105 19227 15163 19233
rect 15105 19193 15117 19227
rect 15151 19224 15163 19227
rect 15286 19224 15292 19236
rect 15151 19196 15292 19224
rect 15151 19193 15163 19196
rect 15105 19187 15163 19193
rect 11330 19116 11336 19168
rect 11388 19156 11394 19168
rect 11793 19159 11851 19165
rect 11793 19156 11805 19159
rect 11388 19128 11805 19156
rect 11388 19116 11394 19128
rect 11793 19125 11805 19128
rect 11839 19125 11851 19159
rect 11793 19119 11851 19125
rect 11882 19116 11888 19168
rect 11940 19156 11946 19168
rect 12253 19159 12311 19165
rect 12253 19156 12265 19159
rect 11940 19128 12265 19156
rect 11940 19116 11946 19128
rect 12253 19125 12265 19128
rect 12299 19156 12311 19159
rect 13078 19156 13084 19168
rect 12299 19128 13084 19156
rect 12299 19125 12311 19128
rect 12253 19119 12311 19125
rect 13078 19116 13084 19128
rect 13136 19116 13142 19168
rect 14829 19159 14887 19165
rect 14829 19125 14841 19159
rect 14875 19156 14887 19159
rect 15120 19156 15148 19187
rect 15286 19184 15292 19196
rect 15344 19184 15350 19236
rect 15654 19224 15660 19236
rect 15615 19196 15660 19224
rect 15654 19184 15660 19196
rect 15712 19184 15718 19236
rect 14875 19128 15148 19156
rect 14875 19125 14887 19128
rect 14829 19119 14887 19125
rect 15378 19116 15384 19168
rect 15436 19156 15442 19168
rect 16666 19156 16672 19168
rect 15436 19128 16672 19156
rect 15436 19116 15442 19128
rect 16666 19116 16672 19128
rect 16724 19116 16730 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 13449 18955 13507 18961
rect 10790 18924 11744 18952
rect 10689 18887 10747 18893
rect 10689 18853 10701 18887
rect 10735 18884 10747 18887
rect 10790 18884 10818 18924
rect 11606 18884 11612 18896
rect 10735 18856 10818 18884
rect 11567 18856 11612 18884
rect 10735 18853 10747 18856
rect 10689 18847 10747 18853
rect 11606 18844 11612 18856
rect 11664 18844 11670 18896
rect 11716 18893 11744 18924
rect 13449 18921 13461 18955
rect 13495 18952 13507 18955
rect 13630 18952 13636 18964
rect 13495 18924 13636 18952
rect 13495 18921 13507 18924
rect 13449 18915 13507 18921
rect 13630 18912 13636 18924
rect 13688 18912 13694 18964
rect 15010 18952 15016 18964
rect 14971 18924 15016 18952
rect 15010 18912 15016 18924
rect 15068 18912 15074 18964
rect 15930 18952 15936 18964
rect 15488 18924 15936 18952
rect 15488 18896 15516 18924
rect 15930 18912 15936 18924
rect 15988 18912 15994 18964
rect 11701 18887 11759 18893
rect 11701 18853 11713 18887
rect 11747 18884 11759 18887
rect 11790 18884 11796 18896
rect 11747 18856 11796 18884
rect 11747 18853 11759 18856
rect 11701 18847 11759 18853
rect 11790 18844 11796 18856
rect 11848 18844 11854 18896
rect 12250 18884 12256 18896
rect 12211 18856 12256 18884
rect 12250 18844 12256 18856
rect 12308 18844 12314 18896
rect 13722 18844 13728 18896
rect 13780 18884 13786 18896
rect 13814 18884 13820 18896
rect 13780 18856 13820 18884
rect 13780 18844 13786 18856
rect 13814 18844 13820 18856
rect 13872 18884 13878 18896
rect 15470 18884 15476 18896
rect 13872 18856 13965 18884
rect 15383 18856 15476 18884
rect 13872 18844 13878 18856
rect 15470 18844 15476 18856
rect 15528 18844 15534 18896
rect 9674 18776 9680 18828
rect 9732 18816 9738 18828
rect 10597 18819 10655 18825
rect 10597 18816 10609 18819
rect 9732 18788 10609 18816
rect 9732 18776 9738 18788
rect 10597 18785 10609 18788
rect 10643 18816 10655 18819
rect 14369 18819 14427 18825
rect 10643 18788 11100 18816
rect 10643 18785 10655 18788
rect 10597 18779 10655 18785
rect 3418 18708 3424 18760
rect 3476 18748 3482 18760
rect 4246 18748 4252 18760
rect 3476 18720 4252 18748
rect 3476 18708 3482 18720
rect 4246 18708 4252 18720
rect 4304 18708 4310 18760
rect 9950 18708 9956 18760
rect 10008 18748 10014 18760
rect 10870 18748 10876 18760
rect 10008 18720 10876 18748
rect 10008 18708 10014 18720
rect 10870 18708 10876 18720
rect 10928 18748 10934 18760
rect 10965 18751 11023 18757
rect 10965 18748 10977 18751
rect 10928 18720 10977 18748
rect 10928 18708 10934 18720
rect 10965 18717 10977 18720
rect 11011 18717 11023 18751
rect 11072 18748 11100 18788
rect 14369 18785 14381 18819
rect 14415 18816 14427 18819
rect 14458 18816 14464 18828
rect 14415 18788 14464 18816
rect 14415 18785 14427 18788
rect 14369 18779 14427 18785
rect 14458 18776 14464 18788
rect 14516 18816 14522 18828
rect 14516 18788 15240 18816
rect 14516 18776 14522 18788
rect 11882 18748 11888 18760
rect 11072 18720 11888 18748
rect 10965 18711 11023 18717
rect 11882 18708 11888 18720
rect 11940 18708 11946 18760
rect 13722 18748 13728 18760
rect 13683 18720 13728 18748
rect 13722 18708 13728 18720
rect 13780 18748 13786 18760
rect 14642 18748 14648 18760
rect 13780 18720 14648 18748
rect 13780 18708 13786 18720
rect 14642 18708 14648 18720
rect 14700 18708 14706 18760
rect 15212 18748 15240 18788
rect 15378 18748 15384 18760
rect 15212 18720 15384 18748
rect 15378 18708 15384 18720
rect 15436 18708 15442 18760
rect 15654 18748 15660 18760
rect 15615 18720 15660 18748
rect 15654 18708 15660 18720
rect 15712 18708 15718 18760
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 9674 18408 9680 18420
rect 9635 18380 9680 18408
rect 9674 18368 9680 18380
rect 9732 18368 9738 18420
rect 9907 18411 9965 18417
rect 9907 18377 9919 18411
rect 9953 18408 9965 18411
rect 10042 18408 10048 18420
rect 9953 18380 10048 18408
rect 9953 18377 9965 18380
rect 9907 18371 9965 18377
rect 10042 18368 10048 18380
rect 10100 18368 10106 18420
rect 10134 18368 10140 18420
rect 10192 18408 10198 18420
rect 10597 18411 10655 18417
rect 10597 18408 10609 18411
rect 10192 18380 10609 18408
rect 10192 18368 10198 18380
rect 10597 18377 10609 18380
rect 10643 18377 10655 18411
rect 11790 18408 11796 18420
rect 11751 18380 11796 18408
rect 10597 18371 10655 18377
rect 4246 18300 4252 18352
rect 4304 18340 4310 18352
rect 4304 18312 9076 18340
rect 4304 18300 4310 18312
rect 7466 18272 7472 18284
rect 7427 18244 7472 18272
rect 7466 18232 7472 18244
rect 7524 18232 7530 18284
rect 8938 18272 8944 18284
rect 8899 18244 8944 18272
rect 8938 18232 8944 18244
rect 8996 18232 9002 18284
rect 2038 18164 2044 18216
rect 2096 18204 2102 18216
rect 6984 18207 7042 18213
rect 6984 18204 6996 18207
rect 2096 18176 6996 18204
rect 2096 18164 2102 18176
rect 6984 18173 6996 18176
rect 7030 18204 7042 18207
rect 7484 18204 7512 18232
rect 7030 18176 7512 18204
rect 9048 18204 9076 18312
rect 9804 18207 9862 18213
rect 9804 18204 9816 18207
rect 9048 18176 9816 18204
rect 7030 18173 7042 18176
rect 6984 18167 7042 18173
rect 9804 18173 9816 18176
rect 9850 18204 9862 18207
rect 10229 18207 10287 18213
rect 10229 18204 10241 18207
rect 9850 18176 10241 18204
rect 9850 18173 9862 18176
rect 9804 18167 9862 18173
rect 10229 18173 10241 18176
rect 10275 18173 10287 18207
rect 10229 18167 10287 18173
rect 8294 18136 8300 18148
rect 8255 18108 8300 18136
rect 8294 18096 8300 18108
rect 8352 18096 8358 18148
rect 8389 18139 8447 18145
rect 8389 18105 8401 18139
rect 8435 18105 8447 18139
rect 10612 18136 10640 18371
rect 11790 18368 11796 18380
rect 11848 18368 11854 18420
rect 13081 18411 13139 18417
rect 13081 18377 13093 18411
rect 13127 18408 13139 18411
rect 13722 18408 13728 18420
rect 13127 18380 13728 18408
rect 13127 18377 13139 18380
rect 13081 18371 13139 18377
rect 13722 18368 13728 18380
rect 13780 18368 13786 18420
rect 15289 18411 15347 18417
rect 15289 18377 15301 18411
rect 15335 18408 15347 18411
rect 15470 18408 15476 18420
rect 15335 18380 15476 18408
rect 15335 18377 15347 18380
rect 15289 18371 15347 18377
rect 15470 18368 15476 18380
rect 15528 18368 15534 18420
rect 14826 18340 14832 18352
rect 14787 18312 14832 18340
rect 14826 18300 14832 18312
rect 14884 18300 14890 18352
rect 15378 18300 15384 18352
rect 15436 18340 15442 18352
rect 16761 18343 16819 18349
rect 16761 18340 16773 18343
rect 15436 18312 16773 18340
rect 15436 18300 15442 18312
rect 16761 18309 16773 18312
rect 16807 18309 16819 18343
rect 16761 18303 16819 18309
rect 10870 18272 10876 18284
rect 10831 18244 10876 18272
rect 10870 18232 10876 18244
rect 10928 18232 10934 18284
rect 11517 18275 11575 18281
rect 11517 18241 11529 18275
rect 11563 18272 11575 18275
rect 11606 18272 11612 18284
rect 11563 18244 11612 18272
rect 11563 18241 11575 18244
rect 11517 18235 11575 18241
rect 11606 18232 11612 18244
rect 11664 18272 11670 18284
rect 12161 18275 12219 18281
rect 12161 18272 12173 18275
rect 11664 18244 12173 18272
rect 11664 18232 11670 18244
rect 12161 18241 12173 18244
rect 12207 18241 12219 18275
rect 12161 18235 12219 18241
rect 14090 18232 14096 18284
rect 14148 18272 14154 18284
rect 14277 18275 14335 18281
rect 14277 18272 14289 18275
rect 14148 18244 14289 18272
rect 14148 18232 14154 18244
rect 14277 18241 14289 18244
rect 14323 18272 14335 18275
rect 14458 18272 14464 18284
rect 14323 18244 14464 18272
rect 14323 18241 14335 18244
rect 14277 18235 14335 18241
rect 14458 18232 14464 18244
rect 14516 18232 14522 18284
rect 13224 18207 13282 18213
rect 13224 18173 13236 18207
rect 13270 18204 13282 18207
rect 13630 18204 13636 18216
rect 13270 18176 13636 18204
rect 13270 18173 13282 18176
rect 13224 18167 13282 18173
rect 13630 18164 13636 18176
rect 13688 18164 13694 18216
rect 15657 18207 15715 18213
rect 15657 18173 15669 18207
rect 15703 18204 15715 18207
rect 15841 18207 15899 18213
rect 15841 18204 15853 18207
rect 15703 18176 15853 18204
rect 15703 18173 15715 18176
rect 15657 18167 15715 18173
rect 15841 18173 15853 18176
rect 15887 18204 15899 18207
rect 16206 18204 16212 18216
rect 15887 18176 16212 18204
rect 15887 18173 15899 18176
rect 15841 18167 15899 18173
rect 16206 18164 16212 18176
rect 16264 18164 16270 18216
rect 10965 18139 11023 18145
rect 10965 18136 10977 18139
rect 10612 18108 10977 18136
rect 8389 18099 8447 18105
rect 10965 18105 10977 18108
rect 11011 18136 11023 18139
rect 11330 18136 11336 18148
rect 11011 18108 11336 18136
rect 11011 18105 11023 18108
rect 10965 18099 11023 18105
rect 7055 18071 7113 18077
rect 7055 18037 7067 18071
rect 7101 18068 7113 18071
rect 7190 18068 7196 18080
rect 7101 18040 7196 18068
rect 7101 18037 7113 18040
rect 7055 18031 7113 18037
rect 7190 18028 7196 18040
rect 7248 18028 7254 18080
rect 7466 18028 7472 18080
rect 7524 18068 7530 18080
rect 8021 18071 8079 18077
rect 8021 18068 8033 18071
rect 7524 18040 8033 18068
rect 7524 18028 7530 18040
rect 8021 18037 8033 18040
rect 8067 18068 8079 18071
rect 8404 18068 8432 18099
rect 11330 18096 11336 18108
rect 11388 18096 11394 18148
rect 13311 18139 13369 18145
rect 13311 18105 13323 18139
rect 13357 18136 13369 18139
rect 14274 18136 14280 18148
rect 13357 18108 14280 18136
rect 13357 18105 13369 18108
rect 13311 18099 13369 18105
rect 14274 18096 14280 18108
rect 14332 18096 14338 18148
rect 14369 18139 14427 18145
rect 14369 18105 14381 18139
rect 14415 18105 14427 18139
rect 14369 18099 14427 18105
rect 8067 18040 8432 18068
rect 8067 18037 8079 18040
rect 8021 18031 8079 18037
rect 13814 18028 13820 18080
rect 13872 18068 13878 18080
rect 14001 18071 14059 18077
rect 14001 18068 14013 18071
rect 13872 18040 14013 18068
rect 13872 18028 13878 18040
rect 14001 18037 14013 18040
rect 14047 18068 14059 18071
rect 14384 18068 14412 18099
rect 16022 18068 16028 18080
rect 14047 18040 14412 18068
rect 15983 18040 16028 18068
rect 14047 18037 14059 18040
rect 14001 18031 14059 18037
rect 16022 18028 16028 18040
rect 16080 18028 16086 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 7101 17867 7159 17873
rect 7101 17833 7113 17867
rect 7147 17864 7159 17867
rect 7190 17864 7196 17876
rect 7147 17836 7196 17864
rect 7147 17833 7159 17836
rect 7101 17827 7159 17833
rect 7190 17824 7196 17836
rect 7248 17824 7254 17876
rect 11330 17864 11336 17876
rect 11291 17836 11336 17864
rect 11330 17824 11336 17836
rect 11388 17824 11394 17876
rect 12526 17864 12532 17876
rect 12487 17836 12532 17864
rect 12526 17824 12532 17836
rect 12584 17824 12590 17876
rect 13078 17864 13084 17876
rect 13039 17836 13084 17864
rect 13078 17824 13084 17836
rect 13136 17824 13142 17876
rect 14090 17864 14096 17876
rect 14051 17836 14096 17864
rect 14090 17824 14096 17836
rect 14148 17824 14154 17876
rect 14458 17864 14464 17876
rect 14419 17836 14464 17864
rect 14458 17824 14464 17836
rect 14516 17824 14522 17876
rect 7374 17796 7380 17808
rect 7335 17768 7380 17796
rect 7374 17756 7380 17768
rect 7432 17756 7438 17808
rect 9766 17756 9772 17808
rect 9824 17796 9830 17808
rect 10734 17799 10792 17805
rect 10734 17796 10746 17799
rect 9824 17768 10746 17796
rect 9824 17756 9830 17768
rect 10734 17765 10746 17768
rect 10780 17765 10792 17799
rect 10734 17759 10792 17765
rect 13725 17799 13783 17805
rect 13725 17765 13737 17799
rect 13771 17796 13783 17799
rect 13814 17796 13820 17808
rect 13771 17768 13820 17796
rect 13771 17765 13783 17768
rect 13725 17759 13783 17765
rect 13814 17756 13820 17768
rect 13872 17756 13878 17808
rect 15378 17796 15384 17808
rect 15339 17768 15384 17796
rect 15378 17756 15384 17768
rect 15436 17756 15442 17808
rect 15473 17799 15531 17805
rect 15473 17765 15485 17799
rect 15519 17796 15531 17799
rect 16022 17796 16028 17808
rect 15519 17768 16028 17796
rect 15519 17765 15531 17768
rect 15473 17759 15531 17765
rect 16022 17756 16028 17768
rect 16080 17756 16086 17808
rect 17034 17796 17040 17808
rect 16995 17768 17040 17796
rect 17034 17756 17040 17768
rect 17092 17756 17098 17808
rect 4893 17731 4951 17737
rect 4893 17697 4905 17731
rect 4939 17728 4951 17731
rect 5074 17728 5080 17740
rect 4939 17700 5080 17728
rect 4939 17697 4951 17700
rect 4893 17691 4951 17697
rect 5074 17688 5080 17700
rect 5132 17688 5138 17740
rect 13354 17688 13360 17740
rect 13412 17728 13418 17740
rect 13906 17728 13912 17740
rect 13412 17700 13912 17728
rect 13412 17688 13418 17700
rect 13906 17688 13912 17700
rect 13964 17688 13970 17740
rect 7282 17660 7288 17672
rect 7243 17632 7288 17660
rect 7282 17620 7288 17632
rect 7340 17620 7346 17672
rect 7650 17660 7656 17672
rect 7611 17632 7656 17660
rect 7650 17620 7656 17632
rect 7708 17660 7714 17672
rect 8205 17663 8263 17669
rect 8205 17660 8217 17663
rect 7708 17632 8217 17660
rect 7708 17620 7714 17632
rect 8205 17629 8217 17632
rect 8251 17660 8263 17663
rect 8294 17660 8300 17672
rect 8251 17632 8300 17660
rect 8251 17629 8263 17632
rect 8205 17623 8263 17629
rect 8294 17620 8300 17632
rect 8352 17620 8358 17672
rect 10413 17663 10471 17669
rect 10413 17629 10425 17663
rect 10459 17660 10471 17663
rect 11422 17660 11428 17672
rect 10459 17632 11428 17660
rect 10459 17629 10471 17632
rect 10413 17623 10471 17629
rect 11422 17620 11428 17632
rect 11480 17620 11486 17672
rect 12161 17663 12219 17669
rect 12161 17629 12173 17663
rect 12207 17629 12219 17663
rect 12161 17623 12219 17629
rect 16025 17663 16083 17669
rect 16025 17629 16037 17663
rect 16071 17660 16083 17663
rect 16758 17660 16764 17672
rect 16071 17632 16764 17660
rect 16071 17629 16083 17632
rect 16025 17623 16083 17629
rect 5123 17527 5181 17533
rect 5123 17493 5135 17527
rect 5169 17524 5181 17527
rect 8110 17524 8116 17536
rect 5169 17496 8116 17524
rect 5169 17493 5181 17496
rect 5123 17487 5181 17493
rect 8110 17484 8116 17496
rect 8168 17484 8174 17536
rect 8938 17524 8944 17536
rect 8899 17496 8944 17524
rect 8938 17484 8944 17496
rect 8996 17484 9002 17536
rect 11790 17484 11796 17536
rect 11848 17524 11854 17536
rect 11977 17527 12035 17533
rect 11977 17524 11989 17527
rect 11848 17496 11989 17524
rect 11848 17484 11854 17496
rect 11977 17493 11989 17496
rect 12023 17524 12035 17527
rect 12176 17524 12204 17623
rect 16758 17620 16764 17632
rect 16816 17660 16822 17672
rect 16945 17663 17003 17669
rect 16945 17660 16957 17663
rect 16816 17632 16957 17660
rect 16816 17620 16822 17632
rect 16945 17629 16957 17632
rect 16991 17629 17003 17663
rect 17586 17660 17592 17672
rect 17547 17632 17592 17660
rect 16945 17623 17003 17629
rect 17586 17620 17592 17632
rect 17644 17620 17650 17672
rect 14274 17552 14280 17604
rect 14332 17592 14338 17604
rect 16393 17595 16451 17601
rect 16393 17592 16405 17595
rect 14332 17564 16405 17592
rect 14332 17552 14338 17564
rect 16393 17561 16405 17564
rect 16439 17592 16451 17595
rect 16482 17592 16488 17604
rect 16439 17564 16488 17592
rect 16439 17561 16451 17564
rect 16393 17555 16451 17561
rect 16482 17552 16488 17564
rect 16540 17552 16546 17604
rect 12023 17496 12204 17524
rect 12023 17493 12035 17496
rect 11977 17487 12035 17493
rect 22738 17484 22744 17536
rect 22796 17524 22802 17536
rect 23934 17524 23940 17536
rect 22796 17496 23940 17524
rect 22796 17484 22802 17496
rect 23934 17484 23940 17496
rect 23992 17484 23998 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 5074 17320 5080 17332
rect 5035 17292 5080 17320
rect 5074 17280 5080 17292
rect 5132 17280 5138 17332
rect 6641 17323 6699 17329
rect 6641 17289 6653 17323
rect 6687 17320 6699 17323
rect 6822 17320 6828 17332
rect 6687 17292 6828 17320
rect 6687 17289 6699 17292
rect 6641 17283 6699 17289
rect 6822 17280 6828 17292
rect 6880 17320 6886 17332
rect 7282 17320 7288 17332
rect 6880 17292 7288 17320
rect 6880 17280 6886 17292
rect 7282 17280 7288 17292
rect 7340 17280 7346 17332
rect 13814 17280 13820 17332
rect 13872 17320 13878 17332
rect 13872 17292 13917 17320
rect 13872 17280 13878 17292
rect 15470 17280 15476 17332
rect 15528 17320 15534 17332
rect 15565 17323 15623 17329
rect 15565 17320 15577 17323
rect 15528 17292 15577 17320
rect 15528 17280 15534 17292
rect 15565 17289 15577 17292
rect 15611 17289 15623 17323
rect 16206 17320 16212 17332
rect 16167 17292 16212 17320
rect 15565 17283 15623 17289
rect 16206 17280 16212 17292
rect 16264 17280 16270 17332
rect 17034 17280 17040 17332
rect 17092 17320 17098 17332
rect 17405 17323 17463 17329
rect 17405 17320 17417 17323
rect 17092 17292 17417 17320
rect 17092 17280 17098 17292
rect 17405 17289 17417 17292
rect 17451 17289 17463 17323
rect 17405 17283 17463 17289
rect 24765 17323 24823 17329
rect 24765 17289 24777 17323
rect 24811 17320 24823 17323
rect 25406 17320 25412 17332
rect 24811 17292 25412 17320
rect 24811 17289 24823 17292
rect 24765 17283 24823 17289
rect 25406 17280 25412 17292
rect 25464 17280 25470 17332
rect 6730 17212 6736 17264
rect 6788 17252 6794 17264
rect 8573 17255 8631 17261
rect 8573 17252 8585 17255
rect 6788 17224 8585 17252
rect 6788 17212 6794 17224
rect 8573 17221 8585 17224
rect 8619 17252 8631 17255
rect 8665 17255 8723 17261
rect 8665 17252 8677 17255
rect 8619 17224 8677 17252
rect 8619 17221 8631 17224
rect 8573 17215 8631 17221
rect 8665 17221 8677 17224
rect 8711 17221 8723 17255
rect 8665 17215 8723 17221
rect 15933 17255 15991 17261
rect 15933 17221 15945 17255
rect 15979 17252 15991 17255
rect 16022 17252 16028 17264
rect 15979 17224 16028 17252
rect 15979 17221 15991 17224
rect 15933 17215 15991 17221
rect 16022 17212 16028 17224
rect 16080 17252 16086 17264
rect 17770 17252 17776 17264
rect 16080 17224 17776 17252
rect 16080 17212 16086 17224
rect 17770 17212 17776 17224
rect 17828 17212 17834 17264
rect 7190 17144 7196 17196
rect 7248 17184 7254 17196
rect 7377 17187 7435 17193
rect 7377 17184 7389 17187
rect 7248 17156 7389 17184
rect 7248 17144 7254 17156
rect 7377 17153 7389 17156
rect 7423 17153 7435 17187
rect 7377 17147 7435 17153
rect 8021 17187 8079 17193
rect 8021 17153 8033 17187
rect 8067 17184 8079 17187
rect 8294 17184 8300 17196
rect 8067 17156 8300 17184
rect 8067 17153 8079 17156
rect 8021 17147 8079 17153
rect 8294 17144 8300 17156
rect 8352 17184 8358 17196
rect 8938 17184 8944 17196
rect 8352 17156 8944 17184
rect 8352 17144 8358 17156
rect 8938 17144 8944 17156
rect 8996 17144 9002 17196
rect 9030 17144 9036 17196
rect 9088 17184 9094 17196
rect 9217 17187 9275 17193
rect 9217 17184 9229 17187
rect 9088 17156 9229 17184
rect 9088 17144 9094 17156
rect 9217 17153 9229 17156
rect 9263 17153 9275 17187
rect 16482 17184 16488 17196
rect 9217 17147 9275 17153
rect 12728 17156 14228 17184
rect 16443 17156 16488 17184
rect 10597 17119 10655 17125
rect 10597 17085 10609 17119
rect 10643 17116 10655 17119
rect 12161 17119 12219 17125
rect 12161 17116 12173 17119
rect 10643 17088 12173 17116
rect 10643 17085 10655 17088
rect 10597 17079 10655 17085
rect 12161 17085 12173 17088
rect 12207 17116 12219 17119
rect 12526 17116 12532 17128
rect 12207 17088 12532 17116
rect 12207 17085 12219 17088
rect 12161 17079 12219 17085
rect 12526 17076 12532 17088
rect 12584 17116 12590 17128
rect 12728 17125 12756 17156
rect 12713 17119 12771 17125
rect 12713 17116 12725 17119
rect 12584 17088 12725 17116
rect 12584 17076 12590 17088
rect 12713 17085 12725 17088
rect 12759 17085 12771 17119
rect 12713 17079 12771 17085
rect 12897 17119 12955 17125
rect 12897 17085 12909 17119
rect 12943 17116 12955 17119
rect 13814 17116 13820 17128
rect 12943 17088 13820 17116
rect 12943 17085 12955 17088
rect 12897 17079 12955 17085
rect 7469 17051 7527 17057
rect 7469 17017 7481 17051
rect 7515 17017 7527 17051
rect 7469 17011 7527 17017
rect 8573 17051 8631 17057
rect 8573 17017 8585 17051
rect 8619 17048 8631 17051
rect 9033 17051 9091 17057
rect 9033 17048 9045 17051
rect 8619 17020 9045 17048
rect 8619 17017 8631 17020
rect 8573 17011 8631 17017
rect 9033 17017 9045 17020
rect 9079 17048 9091 17051
rect 9214 17048 9220 17060
rect 9079 17020 9220 17048
rect 9079 17017 9091 17020
rect 9033 17011 9091 17017
rect 7193 16983 7251 16989
rect 7193 16949 7205 16983
rect 7239 16980 7251 16983
rect 7282 16980 7288 16992
rect 7239 16952 7288 16980
rect 7239 16949 7251 16952
rect 7193 16943 7251 16949
rect 7282 16940 7288 16952
rect 7340 16980 7346 16992
rect 7484 16980 7512 17011
rect 9214 17008 9220 17020
rect 9272 17008 9278 17060
rect 10137 17051 10195 17057
rect 10137 17017 10149 17051
rect 10183 17048 10195 17051
rect 11146 17048 11152 17060
rect 10183 17020 11152 17048
rect 10183 17017 10195 17020
rect 10137 17011 10195 17017
rect 11146 17008 11152 17020
rect 11204 17008 11210 17060
rect 12728 17048 12756 17079
rect 13814 17076 13820 17088
rect 13872 17116 13878 17128
rect 14093 17119 14151 17125
rect 14093 17116 14105 17119
rect 13872 17088 14105 17116
rect 13872 17076 13878 17088
rect 14093 17085 14105 17088
rect 14139 17085 14151 17119
rect 14093 17079 14151 17085
rect 13218 17051 13276 17057
rect 13218 17048 13230 17051
rect 12728 17020 13230 17048
rect 13218 17017 13230 17020
rect 13264 17017 13276 17051
rect 14200 17048 14228 17156
rect 16482 17144 16488 17156
rect 16540 17144 16546 17196
rect 16758 17184 16764 17196
rect 16719 17156 16764 17184
rect 16758 17144 16764 17156
rect 16816 17144 16822 17196
rect 14642 17116 14648 17128
rect 14603 17088 14648 17116
rect 14642 17076 14648 17088
rect 14700 17076 14706 17128
rect 24210 17076 24216 17128
rect 24268 17116 24274 17128
rect 24581 17119 24639 17125
rect 24581 17116 24593 17119
rect 24268 17088 24593 17116
rect 24268 17076 24274 17088
rect 24581 17085 24593 17088
rect 24627 17116 24639 17119
rect 25133 17119 25191 17125
rect 25133 17116 25145 17119
rect 24627 17088 25145 17116
rect 24627 17085 24639 17088
rect 24581 17079 24639 17085
rect 25133 17085 25145 17088
rect 25179 17085 25191 17119
rect 25133 17079 25191 17085
rect 14550 17048 14556 17060
rect 14200 17020 14556 17048
rect 13218 17011 13276 17017
rect 14550 17008 14556 17020
rect 14608 17048 14614 17060
rect 14966 17051 15024 17057
rect 14966 17048 14978 17051
rect 14608 17020 14978 17048
rect 14608 17008 14614 17020
rect 14966 17017 14978 17020
rect 15012 17017 15024 17051
rect 14966 17011 15024 17017
rect 16577 17051 16635 17057
rect 16577 17017 16589 17051
rect 16623 17017 16635 17051
rect 16577 17011 16635 17017
rect 8386 16980 8392 16992
rect 7340 16952 7512 16980
rect 8347 16952 8392 16980
rect 7340 16940 7346 16952
rect 8386 16940 8392 16952
rect 8444 16940 8450 16992
rect 9766 16940 9772 16992
rect 9824 16980 9830 16992
rect 10413 16983 10471 16989
rect 10413 16980 10425 16983
rect 9824 16952 10425 16980
rect 9824 16940 9830 16952
rect 10413 16949 10425 16952
rect 10459 16980 10471 16983
rect 10597 16983 10655 16989
rect 10597 16980 10609 16983
rect 10459 16952 10609 16980
rect 10459 16949 10471 16952
rect 10413 16943 10471 16949
rect 10597 16949 10609 16952
rect 10643 16949 10655 16983
rect 10778 16980 10784 16992
rect 10739 16952 10784 16980
rect 10597 16943 10655 16949
rect 10778 16940 10784 16952
rect 10836 16940 10842 16992
rect 11241 16983 11299 16989
rect 11241 16949 11253 16983
rect 11287 16980 11299 16983
rect 11422 16980 11428 16992
rect 11287 16952 11428 16980
rect 11287 16949 11299 16952
rect 11241 16943 11299 16949
rect 11422 16940 11428 16952
rect 11480 16940 11486 16992
rect 11882 16980 11888 16992
rect 11843 16952 11888 16980
rect 11882 16940 11888 16952
rect 11940 16940 11946 16992
rect 16206 16940 16212 16992
rect 16264 16980 16270 16992
rect 16592 16980 16620 17011
rect 18046 16980 18052 16992
rect 16264 16952 16620 16980
rect 18007 16952 18052 16980
rect 16264 16940 16270 16952
rect 18046 16940 18052 16952
rect 18104 16940 18110 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 11517 16779 11575 16785
rect 11517 16776 11529 16779
rect 11072 16748 11529 16776
rect 6733 16711 6791 16717
rect 6733 16677 6745 16711
rect 6779 16708 6791 16711
rect 7466 16708 7472 16720
rect 6779 16680 7472 16708
rect 6779 16677 6791 16680
rect 6733 16671 6791 16677
rect 7466 16668 7472 16680
rect 7524 16668 7530 16720
rect 7742 16708 7748 16720
rect 7703 16680 7748 16708
rect 7742 16668 7748 16680
rect 7800 16668 7806 16720
rect 8294 16708 8300 16720
rect 8255 16680 8300 16708
rect 8294 16668 8300 16680
rect 8352 16668 8358 16720
rect 6638 16640 6644 16652
rect 6599 16612 6644 16640
rect 6638 16600 6644 16612
rect 6696 16600 6702 16652
rect 9125 16643 9183 16649
rect 9125 16609 9137 16643
rect 9171 16640 9183 16643
rect 9493 16643 9551 16649
rect 9493 16640 9505 16643
rect 9171 16612 9505 16640
rect 9171 16609 9183 16612
rect 9125 16603 9183 16609
rect 9493 16609 9505 16612
rect 9539 16640 9551 16643
rect 9953 16643 10011 16649
rect 9953 16640 9965 16643
rect 9539 16612 9965 16640
rect 9539 16609 9551 16612
rect 9493 16603 9551 16609
rect 9953 16609 9965 16612
rect 9999 16640 10011 16643
rect 10134 16640 10140 16652
rect 9999 16612 10140 16640
rect 9999 16609 10011 16612
rect 9953 16603 10011 16609
rect 10134 16600 10140 16612
rect 10192 16600 10198 16652
rect 10410 16640 10416 16652
rect 10371 16612 10416 16640
rect 10410 16600 10416 16612
rect 10468 16600 10474 16652
rect 11072 16649 11100 16748
rect 11517 16745 11529 16748
rect 11563 16776 11575 16779
rect 14642 16776 14648 16788
rect 11563 16748 13400 16776
rect 11563 16745 11575 16748
rect 11517 16739 11575 16745
rect 11149 16711 11207 16717
rect 11149 16677 11161 16711
rect 11195 16708 11207 16711
rect 11790 16708 11796 16720
rect 11195 16680 11796 16708
rect 11195 16677 11207 16680
rect 11149 16671 11207 16677
rect 11790 16668 11796 16680
rect 11848 16668 11854 16720
rect 11882 16668 11888 16720
rect 11940 16708 11946 16720
rect 12618 16708 12624 16720
rect 11940 16680 12624 16708
rect 11940 16668 11946 16680
rect 12268 16649 12296 16680
rect 12618 16668 12624 16680
rect 12676 16668 12682 16720
rect 10505 16643 10563 16649
rect 10505 16609 10517 16643
rect 10551 16609 10563 16643
rect 10505 16603 10563 16609
rect 11057 16643 11115 16649
rect 11057 16609 11069 16643
rect 11103 16609 11115 16643
rect 11057 16603 11115 16609
rect 12253 16643 12311 16649
rect 12253 16609 12265 16643
rect 12299 16609 12311 16643
rect 12253 16603 12311 16609
rect 12437 16643 12495 16649
rect 12437 16609 12449 16643
rect 12483 16609 12495 16643
rect 12802 16640 12808 16652
rect 12763 16612 12808 16640
rect 12437 16603 12495 16609
rect 7466 16532 7472 16584
rect 7524 16572 7530 16584
rect 7653 16575 7711 16581
rect 7653 16572 7665 16575
rect 7524 16544 7665 16572
rect 7524 16532 7530 16544
rect 7653 16541 7665 16544
rect 7699 16541 7711 16575
rect 10520 16572 10548 16603
rect 10778 16572 10784 16584
rect 7653 16535 7711 16541
rect 8680 16544 10784 16572
rect 8680 16448 8708 16544
rect 10778 16532 10784 16544
rect 10836 16532 10842 16584
rect 12452 16572 12480 16603
rect 12802 16600 12808 16612
rect 12860 16600 12866 16652
rect 13372 16649 13400 16748
rect 13786 16748 14648 16776
rect 13449 16711 13507 16717
rect 13449 16677 13461 16711
rect 13495 16708 13507 16711
rect 13786 16708 13814 16748
rect 14642 16736 14648 16748
rect 14700 16736 14706 16788
rect 15378 16736 15384 16788
rect 15436 16776 15442 16788
rect 15473 16779 15531 16785
rect 15473 16776 15485 16779
rect 15436 16748 15485 16776
rect 15436 16736 15442 16748
rect 15473 16745 15485 16748
rect 15519 16745 15531 16779
rect 15473 16739 15531 16745
rect 16758 16736 16764 16788
rect 16816 16776 16822 16788
rect 17129 16779 17187 16785
rect 17129 16776 17141 16779
rect 16816 16748 17141 16776
rect 16816 16736 16822 16748
rect 17129 16745 17141 16748
rect 17175 16745 17187 16779
rect 17129 16739 17187 16745
rect 13495 16680 13814 16708
rect 13495 16677 13507 16680
rect 13449 16671 13507 16677
rect 13906 16668 13912 16720
rect 13964 16708 13970 16720
rect 14093 16711 14151 16717
rect 14093 16708 14105 16711
rect 13964 16680 14105 16708
rect 13964 16668 13970 16680
rect 14093 16677 14105 16680
rect 14139 16677 14151 16711
rect 14093 16671 14151 16677
rect 16206 16668 16212 16720
rect 16264 16708 16270 16720
rect 16301 16711 16359 16717
rect 16301 16708 16313 16711
rect 16264 16680 16313 16708
rect 16264 16668 16270 16680
rect 16301 16677 16313 16680
rect 16347 16677 16359 16711
rect 16301 16671 16359 16677
rect 17770 16668 17776 16720
rect 17828 16708 17834 16720
rect 17865 16711 17923 16717
rect 17865 16708 17877 16711
rect 17828 16680 17877 16708
rect 17828 16668 17834 16680
rect 17865 16677 17877 16680
rect 17911 16677 17923 16711
rect 17865 16671 17923 16677
rect 13357 16643 13415 16649
rect 13357 16609 13369 16643
rect 13403 16640 13415 16643
rect 13630 16640 13636 16652
rect 13403 16612 13636 16640
rect 13403 16609 13415 16612
rect 13357 16603 13415 16609
rect 13630 16600 13636 16612
rect 13688 16600 13694 16652
rect 11808 16544 12480 16572
rect 16209 16575 16267 16581
rect 7282 16436 7288 16448
rect 7243 16408 7288 16436
rect 7282 16396 7288 16408
rect 7340 16396 7346 16448
rect 8662 16436 8668 16448
rect 8623 16408 8668 16436
rect 8662 16396 8668 16408
rect 8720 16396 8726 16448
rect 11698 16396 11704 16448
rect 11756 16436 11762 16448
rect 11808 16445 11836 16544
rect 16209 16541 16221 16575
rect 16255 16572 16267 16575
rect 17034 16572 17040 16584
rect 16255 16544 17040 16572
rect 16255 16541 16267 16544
rect 16209 16535 16267 16541
rect 17034 16532 17040 16544
rect 17092 16532 17098 16584
rect 17773 16575 17831 16581
rect 17773 16541 17785 16575
rect 17819 16572 17831 16575
rect 18046 16572 18052 16584
rect 17819 16544 18052 16572
rect 17819 16541 17831 16544
rect 17773 16535 17831 16541
rect 18046 16532 18052 16544
rect 18104 16572 18110 16584
rect 18506 16572 18512 16584
rect 18104 16544 18512 16572
rect 18104 16532 18110 16544
rect 18506 16532 18512 16544
rect 18564 16532 18570 16584
rect 16761 16507 16819 16513
rect 16761 16473 16773 16507
rect 16807 16504 16819 16507
rect 17126 16504 17132 16516
rect 16807 16476 17132 16504
rect 16807 16473 16819 16476
rect 16761 16467 16819 16473
rect 17126 16464 17132 16476
rect 17184 16504 17190 16516
rect 18325 16507 18383 16513
rect 18325 16504 18337 16507
rect 17184 16476 18337 16504
rect 17184 16464 17190 16476
rect 18325 16473 18337 16476
rect 18371 16473 18383 16507
rect 18325 16467 18383 16473
rect 11793 16439 11851 16445
rect 11793 16436 11805 16439
rect 11756 16408 11805 16436
rect 11756 16396 11762 16408
rect 11793 16405 11805 16408
rect 11839 16405 11851 16439
rect 11793 16399 11851 16405
rect 13446 16396 13452 16448
rect 13504 16436 13510 16448
rect 13725 16439 13783 16445
rect 13725 16436 13737 16439
rect 13504 16408 13737 16436
rect 13504 16396 13510 16408
rect 13725 16405 13737 16408
rect 13771 16405 13783 16439
rect 13725 16399 13783 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 6638 16232 6644 16244
rect 6599 16204 6644 16232
rect 6638 16192 6644 16204
rect 6696 16192 6702 16244
rect 7653 16235 7711 16241
rect 7653 16201 7665 16235
rect 7699 16232 7711 16235
rect 7742 16232 7748 16244
rect 7699 16204 7748 16232
rect 7699 16201 7711 16204
rect 7653 16195 7711 16201
rect 7742 16192 7748 16204
rect 7800 16192 7806 16244
rect 9214 16232 9220 16244
rect 9175 16204 9220 16232
rect 9214 16192 9220 16204
rect 9272 16192 9278 16244
rect 16206 16232 16212 16244
rect 16167 16204 16212 16232
rect 16206 16192 16212 16204
rect 16264 16192 16270 16244
rect 17770 16232 17776 16244
rect 17731 16204 17776 16232
rect 17770 16192 17776 16204
rect 17828 16192 17834 16244
rect 18506 16232 18512 16244
rect 18467 16204 18512 16232
rect 18506 16192 18512 16204
rect 18564 16192 18570 16244
rect 24762 16232 24768 16244
rect 24723 16204 24768 16232
rect 24762 16192 24768 16204
rect 24820 16192 24826 16244
rect 6273 16167 6331 16173
rect 6273 16133 6285 16167
rect 6319 16164 6331 16167
rect 8478 16164 8484 16176
rect 6319 16136 8484 16164
rect 6319 16133 6331 16136
rect 6273 16127 6331 16133
rect 5772 16031 5830 16037
rect 5772 15997 5784 16031
rect 5818 16028 5830 16031
rect 6086 16028 6092 16040
rect 5818 16000 6092 16028
rect 5818 15997 5830 16000
rect 5772 15991 5830 15997
rect 6086 15988 6092 16000
rect 6144 16028 6150 16040
rect 6288 16028 6316 16127
rect 8478 16124 8484 16136
rect 8536 16124 8542 16176
rect 11422 16164 11428 16176
rect 11383 16136 11428 16164
rect 11422 16124 11428 16136
rect 11480 16124 11486 16176
rect 13814 16124 13820 16176
rect 13872 16164 13878 16176
rect 15657 16167 15715 16173
rect 13872 16136 13917 16164
rect 13872 16124 13878 16136
rect 15657 16133 15669 16167
rect 15703 16164 15715 16167
rect 16942 16164 16948 16176
rect 15703 16136 16948 16164
rect 15703 16133 15715 16136
rect 15657 16127 15715 16133
rect 16942 16124 16948 16136
rect 17000 16124 17006 16176
rect 6822 16096 6828 16108
rect 6783 16068 6828 16096
rect 6822 16056 6828 16068
rect 6880 16056 6886 16108
rect 10336 16068 12664 16096
rect 6144 16000 6316 16028
rect 8297 16031 8355 16037
rect 6144 15988 6150 16000
rect 8297 15997 8309 16031
rect 8343 16028 8355 16031
rect 8386 16028 8392 16040
rect 8343 16000 8392 16028
rect 8343 15997 8355 16000
rect 8297 15991 8355 15997
rect 8386 15988 8392 16000
rect 8444 16028 8450 16040
rect 8754 16028 8760 16040
rect 8444 16000 8760 16028
rect 8444 15988 8450 16000
rect 8754 15988 8760 16000
rect 8812 15988 8818 16040
rect 10134 15988 10140 16040
rect 10192 16028 10198 16040
rect 10336 16037 10364 16068
rect 12636 16040 12664 16068
rect 15378 16056 15384 16108
rect 15436 16096 15442 16108
rect 19334 16096 19340 16108
rect 15436 16068 19340 16096
rect 15436 16056 15442 16068
rect 19334 16056 19340 16068
rect 19392 16056 19398 16108
rect 10321 16031 10379 16037
rect 10321 16028 10333 16031
rect 10192 16000 10333 16028
rect 10192 15988 10198 16000
rect 10321 15997 10333 16000
rect 10367 15997 10379 16031
rect 10321 15991 10379 15997
rect 10505 16031 10563 16037
rect 10505 15997 10517 16031
rect 10551 15997 10563 16031
rect 10505 15991 10563 15997
rect 5859 15963 5917 15969
rect 5859 15929 5871 15963
rect 5905 15960 5917 15963
rect 7466 15960 7472 15972
rect 5905 15932 7472 15960
rect 5905 15929 5917 15932
rect 5859 15923 5917 15929
rect 7466 15920 7472 15932
rect 7524 15920 7530 15972
rect 8202 15960 8208 15972
rect 8115 15932 8208 15960
rect 8202 15920 8208 15932
rect 8260 15960 8266 15972
rect 8659 15963 8717 15969
rect 8659 15960 8671 15963
rect 8260 15932 8671 15960
rect 8260 15920 8266 15932
rect 8659 15929 8671 15932
rect 8705 15960 8717 15963
rect 9766 15960 9772 15972
rect 8705 15932 9772 15960
rect 8705 15929 8717 15932
rect 8659 15923 8717 15929
rect 9766 15920 9772 15932
rect 9824 15920 9830 15972
rect 10410 15960 10416 15972
rect 9876 15932 10416 15960
rect 9122 15852 9128 15904
rect 9180 15892 9186 15904
rect 9876 15901 9904 15932
rect 10410 15920 10416 15932
rect 10468 15960 10474 15972
rect 10520 15960 10548 15991
rect 10778 15988 10784 16040
rect 10836 16028 10842 16040
rect 10873 16031 10931 16037
rect 10873 16028 10885 16031
rect 10836 16000 10885 16028
rect 10836 15988 10842 16000
rect 10873 15997 10885 16000
rect 10919 15997 10931 16031
rect 10873 15991 10931 15997
rect 11146 15988 11152 16040
rect 11204 16028 11210 16040
rect 11241 16031 11299 16037
rect 11241 16028 11253 16031
rect 11204 16000 11253 16028
rect 11204 15988 11210 16000
rect 11241 15997 11253 16000
rect 11287 15997 11299 16031
rect 12618 16028 12624 16040
rect 12579 16000 12624 16028
rect 11241 15991 11299 15997
rect 12618 15988 12624 16000
rect 12676 15988 12682 16040
rect 12894 16028 12900 16040
rect 12855 16000 12900 16028
rect 12894 15988 12900 16000
rect 12952 15988 12958 16040
rect 13265 16031 13323 16037
rect 13265 15997 13277 16031
rect 13311 15997 13323 16031
rect 13265 15991 13323 15997
rect 11698 15960 11704 15972
rect 10468 15932 11704 15960
rect 10468 15920 10474 15932
rect 11698 15920 11704 15932
rect 11756 15920 11762 15972
rect 12802 15960 12808 15972
rect 12176 15932 12808 15960
rect 9493 15895 9551 15901
rect 9493 15892 9505 15895
rect 9180 15864 9505 15892
rect 9180 15852 9186 15864
rect 9493 15861 9505 15864
rect 9539 15892 9551 15895
rect 9861 15895 9919 15901
rect 9861 15892 9873 15895
rect 9539 15864 9873 15892
rect 9539 15861 9551 15864
rect 9493 15855 9551 15861
rect 9861 15861 9873 15864
rect 9907 15861 9919 15895
rect 11882 15892 11888 15904
rect 11843 15864 11888 15892
rect 9861 15855 9919 15861
rect 11882 15852 11888 15864
rect 11940 15892 11946 15904
rect 12176 15901 12204 15932
rect 12802 15920 12808 15932
rect 12860 15960 12866 15972
rect 13280 15960 13308 15991
rect 13446 15988 13452 16040
rect 13504 16028 13510 16040
rect 13633 16031 13691 16037
rect 13633 16028 13645 16031
rect 13504 16000 13645 16028
rect 13504 15988 13510 16000
rect 13633 15997 13645 16000
rect 13679 15997 13691 16031
rect 14734 16028 14740 16040
rect 14695 16000 14740 16028
rect 13633 15991 13691 15997
rect 14734 15988 14740 16000
rect 14792 15988 14798 16040
rect 17586 15988 17592 16040
rect 17644 16028 17650 16040
rect 18084 16031 18142 16037
rect 18084 16028 18096 16031
rect 17644 16000 18096 16028
rect 17644 15988 17650 16000
rect 18084 15997 18096 16000
rect 18130 16028 18142 16031
rect 18877 16031 18935 16037
rect 18877 16028 18889 16031
rect 18130 16000 18889 16028
rect 18130 15997 18142 16000
rect 18084 15991 18142 15997
rect 18877 15997 18889 16000
rect 18923 15997 18935 16031
rect 18877 15991 18935 15997
rect 24026 15988 24032 16040
rect 24084 16028 24090 16040
rect 24581 16031 24639 16037
rect 24581 16028 24593 16031
rect 24084 16000 24593 16028
rect 24084 15988 24090 16000
rect 24581 15997 24593 16000
rect 24627 16028 24639 16031
rect 25133 16031 25191 16037
rect 25133 16028 25145 16031
rect 24627 16000 25145 16028
rect 24627 15997 24639 16000
rect 24581 15991 24639 15997
rect 25133 15997 25145 16000
rect 25179 15997 25191 16031
rect 25133 15991 25191 15997
rect 14185 15963 14243 15969
rect 14185 15960 14197 15963
rect 12860 15932 13308 15960
rect 13786 15932 14197 15960
rect 12860 15920 12866 15932
rect 12161 15895 12219 15901
rect 12161 15892 12173 15895
rect 11940 15864 12173 15892
rect 11940 15852 11946 15864
rect 12161 15861 12173 15864
rect 12207 15861 12219 15895
rect 12161 15855 12219 15861
rect 12894 15852 12900 15904
rect 12952 15892 12958 15904
rect 13786 15892 13814 15932
rect 14185 15929 14197 15932
rect 14231 15929 14243 15963
rect 14185 15923 14243 15929
rect 14550 15920 14556 15972
rect 14608 15960 14614 15972
rect 14645 15963 14703 15969
rect 14645 15960 14657 15963
rect 14608 15932 14657 15960
rect 14608 15920 14614 15932
rect 14645 15929 14657 15932
rect 14691 15960 14703 15963
rect 15099 15963 15157 15969
rect 15099 15960 15111 15963
rect 14691 15932 15111 15960
rect 14691 15929 14703 15932
rect 14645 15923 14703 15929
rect 15099 15929 15111 15932
rect 15145 15960 15157 15963
rect 15746 15960 15752 15972
rect 15145 15932 15752 15960
rect 15145 15929 15157 15932
rect 15099 15923 15157 15929
rect 15746 15920 15752 15932
rect 15804 15920 15810 15972
rect 18187 15963 18245 15969
rect 18187 15929 18199 15963
rect 18233 15960 18245 15963
rect 19702 15960 19708 15972
rect 18233 15932 19708 15960
rect 18233 15929 18245 15932
rect 18187 15923 18245 15929
rect 19702 15920 19708 15932
rect 19760 15920 19766 15972
rect 16482 15892 16488 15904
rect 12952 15864 13814 15892
rect 16443 15864 16488 15892
rect 12952 15852 12958 15864
rect 16482 15852 16488 15864
rect 16540 15852 16546 15904
rect 17034 15892 17040 15904
rect 16995 15864 17040 15892
rect 17034 15852 17040 15864
rect 17092 15852 17098 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 7466 15688 7472 15700
rect 7427 15660 7472 15688
rect 7466 15648 7472 15660
rect 7524 15648 7530 15700
rect 7742 15648 7748 15700
rect 7800 15688 7806 15700
rect 8573 15691 8631 15697
rect 8573 15688 8585 15691
rect 7800 15660 8585 15688
rect 7800 15648 7806 15660
rect 8573 15657 8585 15660
rect 8619 15657 8631 15691
rect 8573 15651 8631 15657
rect 8754 15648 8760 15700
rect 8812 15688 8818 15700
rect 10045 15691 10103 15697
rect 10045 15688 10057 15691
rect 8812 15660 10057 15688
rect 8812 15648 8818 15660
rect 10045 15657 10057 15660
rect 10091 15657 10103 15691
rect 11698 15688 11704 15700
rect 11659 15660 11704 15688
rect 10045 15651 10103 15657
rect 11698 15648 11704 15660
rect 11756 15648 11762 15700
rect 12618 15648 12624 15700
rect 12676 15688 12682 15700
rect 14001 15691 14059 15697
rect 14001 15688 14013 15691
rect 12676 15660 14013 15688
rect 12676 15648 12682 15660
rect 14001 15657 14013 15660
rect 14047 15657 14059 15691
rect 16206 15688 16212 15700
rect 16167 15660 16212 15688
rect 14001 15651 14059 15657
rect 16206 15648 16212 15660
rect 16264 15648 16270 15700
rect 17034 15648 17040 15700
rect 17092 15688 17098 15700
rect 18739 15691 18797 15697
rect 18739 15688 18751 15691
rect 17092 15660 18751 15688
rect 17092 15648 17098 15660
rect 18739 15657 18751 15660
rect 18785 15657 18797 15691
rect 18739 15651 18797 15657
rect 6825 15623 6883 15629
rect 6825 15589 6837 15623
rect 6871 15620 6883 15623
rect 7282 15620 7288 15632
rect 6871 15592 7288 15620
rect 6871 15589 6883 15592
rect 6825 15583 6883 15589
rect 7282 15580 7288 15592
rect 7340 15580 7346 15632
rect 6638 15512 6644 15564
rect 6696 15552 6702 15564
rect 6733 15555 6791 15561
rect 6733 15552 6745 15555
rect 6696 15524 6745 15552
rect 6696 15512 6702 15524
rect 6733 15521 6745 15524
rect 6779 15552 6791 15555
rect 7190 15552 7196 15564
rect 6779 15524 7196 15552
rect 6779 15521 6791 15524
rect 6733 15515 6791 15521
rect 7190 15512 7196 15524
rect 7248 15552 7254 15564
rect 7760 15552 7788 15648
rect 8015 15623 8073 15629
rect 8015 15589 8027 15623
rect 8061 15620 8073 15623
rect 8202 15620 8208 15632
rect 8061 15592 8208 15620
rect 8061 15589 8073 15592
rect 8015 15583 8073 15589
rect 8202 15580 8208 15592
rect 8260 15580 8266 15632
rect 11716 15620 11744 15648
rect 15651 15623 15709 15629
rect 11716 15592 12756 15620
rect 7248 15524 7788 15552
rect 9125 15555 9183 15561
rect 7248 15512 7254 15524
rect 9125 15521 9137 15555
rect 9171 15552 9183 15555
rect 10134 15552 10140 15564
rect 9171 15524 10140 15552
rect 9171 15521 9183 15524
rect 9125 15515 9183 15521
rect 10134 15512 10140 15524
rect 10192 15512 10198 15564
rect 10686 15552 10692 15564
rect 10647 15524 10692 15552
rect 10686 15512 10692 15524
rect 10744 15512 10750 15564
rect 10778 15512 10784 15564
rect 10836 15552 10842 15564
rect 11330 15552 11336 15564
rect 10836 15524 10881 15552
rect 11291 15524 11336 15552
rect 10836 15512 10842 15524
rect 11330 15512 11336 15524
rect 11388 15512 11394 15564
rect 12161 15555 12219 15561
rect 12161 15521 12173 15555
rect 12207 15552 12219 15555
rect 12434 15552 12440 15564
rect 12207 15524 12440 15552
rect 12207 15521 12219 15524
rect 12161 15515 12219 15521
rect 12434 15512 12440 15524
rect 12492 15512 12498 15564
rect 12728 15561 12756 15592
rect 15651 15589 15663 15623
rect 15697 15620 15709 15623
rect 15746 15620 15752 15632
rect 15697 15592 15752 15620
rect 15697 15589 15709 15592
rect 15651 15583 15709 15589
rect 15746 15580 15752 15592
rect 15804 15580 15810 15632
rect 17218 15620 17224 15632
rect 17179 15592 17224 15620
rect 17218 15580 17224 15592
rect 17276 15580 17282 15632
rect 12713 15555 12771 15561
rect 12713 15521 12725 15555
rect 12759 15552 12771 15555
rect 12894 15552 12900 15564
rect 12759 15524 12900 15552
rect 12759 15521 12771 15524
rect 12713 15515 12771 15521
rect 12894 15512 12900 15524
rect 12952 15512 12958 15564
rect 13078 15552 13084 15564
rect 13039 15524 13084 15552
rect 13078 15512 13084 15524
rect 13136 15512 13142 15564
rect 13446 15552 13452 15564
rect 13407 15524 13452 15552
rect 13446 15512 13452 15524
rect 13504 15512 13510 15564
rect 18601 15555 18659 15561
rect 18601 15521 18613 15555
rect 18647 15552 18659 15555
rect 18690 15552 18696 15564
rect 18647 15524 18696 15552
rect 18647 15521 18659 15524
rect 18601 15515 18659 15521
rect 18690 15512 18696 15524
rect 18748 15512 18754 15564
rect 7653 15487 7711 15493
rect 7653 15453 7665 15487
rect 7699 15484 7711 15487
rect 8478 15484 8484 15496
rect 7699 15456 8484 15484
rect 7699 15453 7711 15456
rect 7653 15447 7711 15453
rect 8478 15444 8484 15456
rect 8536 15444 8542 15496
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15484 13783 15487
rect 15289 15487 15347 15493
rect 15289 15484 15301 15487
rect 13771 15456 15301 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 15289 15453 15301 15456
rect 15335 15484 15347 15487
rect 16114 15484 16120 15496
rect 15335 15456 16120 15484
rect 15335 15453 15347 15456
rect 15289 15447 15347 15453
rect 16114 15444 16120 15456
rect 16172 15444 16178 15496
rect 17126 15484 17132 15496
rect 17087 15456 17132 15484
rect 17126 15444 17132 15456
rect 17184 15444 17190 15496
rect 17586 15484 17592 15496
rect 17547 15456 17592 15484
rect 17586 15444 17592 15456
rect 17644 15444 17650 15496
rect 9490 15348 9496 15360
rect 9451 15320 9496 15348
rect 9490 15308 9496 15320
rect 9548 15308 9554 15360
rect 13906 15308 13912 15360
rect 13964 15348 13970 15360
rect 14734 15348 14740 15360
rect 13964 15320 14740 15348
rect 13964 15308 13970 15320
rect 14734 15308 14740 15320
rect 14792 15308 14798 15360
rect 18046 15348 18052 15360
rect 18007 15320 18052 15348
rect 18046 15308 18052 15320
rect 18104 15308 18110 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 6181 15147 6239 15153
rect 6181 15113 6193 15147
rect 6227 15144 6239 15147
rect 6638 15144 6644 15156
rect 6227 15116 6644 15144
rect 6227 15113 6239 15116
rect 6181 15107 6239 15113
rect 6638 15104 6644 15116
rect 6696 15104 6702 15156
rect 8018 15104 8024 15156
rect 8076 15144 8082 15156
rect 8113 15147 8171 15153
rect 8113 15144 8125 15147
rect 8076 15116 8125 15144
rect 8076 15104 8082 15116
rect 8113 15113 8125 15116
rect 8159 15144 8171 15147
rect 8202 15144 8208 15156
rect 8159 15116 8208 15144
rect 8159 15113 8171 15116
rect 8113 15107 8171 15113
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 9122 15144 9128 15156
rect 9083 15116 9128 15144
rect 9122 15104 9128 15116
rect 9180 15104 9186 15156
rect 16114 15144 16120 15156
rect 16075 15116 16120 15144
rect 16114 15104 16120 15116
rect 16172 15104 16178 15156
rect 17126 15104 17132 15156
rect 17184 15144 17190 15156
rect 17681 15147 17739 15153
rect 17681 15144 17693 15147
rect 17184 15116 17693 15144
rect 17184 15104 17190 15116
rect 17681 15113 17693 15116
rect 17727 15113 17739 15147
rect 17681 15107 17739 15113
rect 7650 15076 7656 15088
rect 7611 15048 7656 15076
rect 7650 15036 7656 15048
rect 7708 15036 7714 15088
rect 12434 15036 12440 15088
rect 12492 15076 12498 15088
rect 14185 15079 14243 15085
rect 14185 15076 14197 15079
rect 12492 15048 14197 15076
rect 12492 15036 12498 15048
rect 14185 15045 14197 15048
rect 14231 15045 14243 15079
rect 14185 15039 14243 15045
rect 13906 15008 13912 15020
rect 13867 14980 13912 15008
rect 13906 14968 13912 14980
rect 13964 14968 13970 15020
rect 15286 15008 15292 15020
rect 15247 14980 15292 15008
rect 15286 14968 15292 14980
rect 15344 14968 15350 15020
rect 17037 15011 17095 15017
rect 17037 14977 17049 15011
rect 17083 15008 17095 15011
rect 17218 15008 17224 15020
rect 17083 14980 17224 15008
rect 17083 14977 17095 14980
rect 17037 14971 17095 14977
rect 17218 14968 17224 14980
rect 17276 15008 17282 15020
rect 17313 15011 17371 15017
rect 17313 15008 17325 15011
rect 17276 14980 17325 15008
rect 17276 14968 17282 14980
rect 17313 14977 17325 14980
rect 17359 14977 17371 15011
rect 17313 14971 17371 14977
rect 17954 14968 17960 15020
rect 18012 15008 18018 15020
rect 19061 15011 19119 15017
rect 19061 15008 19073 15011
rect 18012 14980 19073 15008
rect 18012 14968 18018 14980
rect 19061 14977 19073 14980
rect 19107 14977 19119 15011
rect 19061 14971 19119 14977
rect 8849 14943 8907 14949
rect 8849 14909 8861 14943
rect 8895 14940 8907 14943
rect 8941 14943 8999 14949
rect 8941 14940 8953 14943
rect 8895 14912 8953 14940
rect 8895 14909 8907 14912
rect 8849 14903 8907 14909
rect 8941 14909 8953 14912
rect 8987 14940 8999 14943
rect 9398 14940 9404 14952
rect 8987 14912 9404 14940
rect 8987 14909 8999 14912
rect 8941 14903 8999 14909
rect 9398 14900 9404 14912
rect 9456 14900 9462 14952
rect 10134 14940 10140 14952
rect 10095 14912 10140 14940
rect 10134 14900 10140 14912
rect 10192 14900 10198 14952
rect 10686 14940 10692 14952
rect 10647 14912 10692 14940
rect 10686 14900 10692 14912
rect 10744 14900 10750 14952
rect 10778 14900 10784 14952
rect 10836 14940 10842 14952
rect 11146 14940 11152 14952
rect 10836 14912 10881 14940
rect 11107 14912 11152 14940
rect 10836 14900 10842 14912
rect 11146 14900 11152 14912
rect 11204 14900 11210 14952
rect 12434 14940 12440 14952
rect 12395 14912 12440 14940
rect 12434 14900 12440 14912
rect 12492 14900 12498 14952
rect 12894 14940 12900 14952
rect 12855 14912 12900 14940
rect 12894 14900 12900 14912
rect 12952 14900 12958 14952
rect 13265 14943 13323 14949
rect 13265 14909 13277 14943
rect 13311 14909 13323 14943
rect 13630 14940 13636 14952
rect 13591 14912 13636 14940
rect 13265 14903 13323 14909
rect 7098 14872 7104 14884
rect 7059 14844 7104 14872
rect 7098 14832 7104 14844
rect 7156 14832 7162 14884
rect 7190 14832 7196 14884
rect 7248 14872 7254 14884
rect 8478 14872 8484 14884
rect 7248 14844 7293 14872
rect 8391 14844 8484 14872
rect 7248 14832 7254 14844
rect 8478 14832 8484 14844
rect 8536 14872 8542 14884
rect 10796 14872 10824 14900
rect 11701 14875 11759 14881
rect 11701 14872 11713 14875
rect 8536 14844 10088 14872
rect 10796 14844 11713 14872
rect 8536 14832 8542 14844
rect 9398 14804 9404 14816
rect 9359 14776 9404 14804
rect 9398 14764 9404 14776
rect 9456 14804 9462 14816
rect 10060 14813 10088 14844
rect 11701 14841 11713 14844
rect 11747 14872 11759 14875
rect 12161 14875 12219 14881
rect 12161 14872 12173 14875
rect 11747 14844 12173 14872
rect 11747 14841 11759 14844
rect 11701 14835 11759 14841
rect 12161 14841 12173 14844
rect 12207 14872 12219 14875
rect 13078 14872 13084 14884
rect 12207 14844 13084 14872
rect 12207 14841 12219 14844
rect 12161 14835 12219 14841
rect 13078 14832 13084 14844
rect 13136 14872 13142 14884
rect 13280 14872 13308 14903
rect 13630 14900 13636 14912
rect 13688 14900 13694 14952
rect 16850 14940 16856 14952
rect 16811 14912 16856 14940
rect 16850 14900 16856 14912
rect 16908 14900 16914 14952
rect 16942 14900 16948 14952
rect 17000 14940 17006 14952
rect 18046 14940 18052 14952
rect 18104 14949 18110 14952
rect 18104 14943 18142 14949
rect 17000 14912 18052 14940
rect 17000 14900 17006 14912
rect 18046 14900 18052 14912
rect 18130 14909 18142 14943
rect 18104 14903 18142 14909
rect 18104 14900 18110 14903
rect 14826 14872 14832 14884
rect 13136 14844 13308 14872
rect 14787 14844 14832 14872
rect 13136 14832 13142 14844
rect 14826 14832 14832 14844
rect 14884 14832 14890 14884
rect 14921 14875 14979 14881
rect 14921 14841 14933 14875
rect 14967 14841 14979 14875
rect 14921 14835 14979 14841
rect 18187 14875 18245 14881
rect 18187 14841 18199 14875
rect 18233 14872 18245 14875
rect 19702 14872 19708 14884
rect 18233 14844 19708 14872
rect 18233 14841 18245 14844
rect 18187 14835 18245 14841
rect 9769 14807 9827 14813
rect 9769 14804 9781 14807
rect 9456 14776 9781 14804
rect 9456 14764 9462 14776
rect 9769 14773 9781 14776
rect 9815 14773 9827 14807
rect 9769 14767 9827 14773
rect 10045 14807 10103 14813
rect 10045 14773 10057 14807
rect 10091 14773 10103 14807
rect 10045 14767 10103 14773
rect 14274 14764 14280 14816
rect 14332 14804 14338 14816
rect 14645 14807 14703 14813
rect 14645 14804 14657 14807
rect 14332 14776 14657 14804
rect 14332 14764 14338 14776
rect 14645 14773 14657 14776
rect 14691 14804 14703 14807
rect 14936 14804 14964 14835
rect 19702 14832 19708 14844
rect 19760 14832 19766 14884
rect 15746 14804 15752 14816
rect 14691 14776 14964 14804
rect 15707 14776 15752 14804
rect 14691 14773 14703 14776
rect 14645 14767 14703 14773
rect 15746 14764 15752 14776
rect 15804 14764 15810 14816
rect 18690 14804 18696 14816
rect 18651 14776 18696 14804
rect 18690 14764 18696 14776
rect 18748 14764 18754 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 9125 14603 9183 14609
rect 9125 14569 9137 14603
rect 9171 14600 9183 14603
rect 10134 14600 10140 14612
rect 9171 14572 10140 14600
rect 9171 14569 9183 14572
rect 9125 14563 9183 14569
rect 10134 14560 10140 14572
rect 10192 14600 10198 14612
rect 11241 14603 11299 14609
rect 11241 14600 11253 14603
rect 10192 14572 11253 14600
rect 10192 14560 10198 14572
rect 11241 14569 11253 14572
rect 11287 14569 11299 14603
rect 11241 14563 11299 14569
rect 11698 14560 11704 14612
rect 11756 14600 11762 14612
rect 11885 14603 11943 14609
rect 11885 14600 11897 14603
rect 11756 14572 11897 14600
rect 11756 14560 11762 14572
rect 11885 14569 11897 14572
rect 11931 14569 11943 14603
rect 13078 14600 13084 14612
rect 13039 14572 13084 14600
rect 11885 14563 11943 14569
rect 13078 14560 13084 14572
rect 13136 14560 13142 14612
rect 14826 14600 14832 14612
rect 14787 14572 14832 14600
rect 14826 14560 14832 14572
rect 14884 14600 14890 14612
rect 15427 14603 15485 14609
rect 15427 14600 15439 14603
rect 14884 14572 15439 14600
rect 14884 14560 14890 14572
rect 15427 14569 15439 14572
rect 15473 14569 15485 14603
rect 15427 14563 15485 14569
rect 16393 14603 16451 14609
rect 16393 14569 16405 14603
rect 16439 14600 16451 14603
rect 16850 14600 16856 14612
rect 16439 14572 16856 14600
rect 16439 14569 16451 14572
rect 16393 14563 16451 14569
rect 16850 14560 16856 14572
rect 16908 14560 16914 14612
rect 24762 14600 24768 14612
rect 24723 14572 24768 14600
rect 24762 14560 24768 14572
rect 24820 14560 24826 14612
rect 9214 14492 9220 14544
rect 9272 14532 9278 14544
rect 9490 14532 9496 14544
rect 9272 14504 9496 14532
rect 9272 14492 9278 14504
rect 9490 14492 9496 14504
rect 9548 14532 9554 14544
rect 9953 14535 10011 14541
rect 9953 14532 9965 14535
rect 9548 14504 9965 14532
rect 9548 14492 9554 14504
rect 9953 14501 9965 14504
rect 9999 14532 10011 14535
rect 11330 14532 11336 14544
rect 9999 14504 11336 14532
rect 9999 14501 10011 14504
rect 9953 14495 10011 14501
rect 11330 14492 11336 14504
rect 11388 14532 11394 14544
rect 11609 14535 11667 14541
rect 11609 14532 11621 14535
rect 11388 14504 11621 14532
rect 11388 14492 11394 14504
rect 11609 14501 11621 14504
rect 11655 14532 11667 14535
rect 13630 14532 13636 14544
rect 11655 14504 13636 14532
rect 11655 14501 11667 14504
rect 11609 14495 11667 14501
rect 13630 14492 13636 14504
rect 13688 14492 13694 14544
rect 16482 14492 16488 14544
rect 16540 14532 16546 14544
rect 16669 14535 16727 14541
rect 16669 14532 16681 14535
rect 16540 14504 16681 14532
rect 16540 14492 16546 14504
rect 16669 14501 16681 14504
rect 16715 14501 16727 14535
rect 16669 14495 16727 14501
rect 16761 14535 16819 14541
rect 16761 14501 16773 14535
rect 16807 14532 16819 14535
rect 17034 14532 17040 14544
rect 16807 14504 17040 14532
rect 16807 14501 16819 14504
rect 16761 14495 16819 14501
rect 17034 14492 17040 14504
rect 17092 14492 17098 14544
rect 6546 14424 6552 14476
rect 6604 14464 6610 14476
rect 6676 14467 6734 14473
rect 6676 14464 6688 14467
rect 6604 14436 6688 14464
rect 6604 14424 6610 14436
rect 6676 14433 6688 14436
rect 6722 14433 6734 14467
rect 6676 14427 6734 14433
rect 8180 14467 8238 14473
rect 8180 14433 8192 14467
rect 8226 14464 8238 14467
rect 8846 14464 8852 14476
rect 8226 14436 8852 14464
rect 8226 14433 8238 14436
rect 8180 14427 8238 14433
rect 8846 14424 8852 14436
rect 8904 14424 8910 14476
rect 10045 14467 10103 14473
rect 10045 14433 10057 14467
rect 10091 14464 10103 14467
rect 10134 14464 10140 14476
rect 10091 14436 10140 14464
rect 10091 14433 10103 14436
rect 10045 14427 10103 14433
rect 10134 14424 10140 14436
rect 10192 14424 10198 14476
rect 11054 14464 11060 14476
rect 11015 14436 11060 14464
rect 11054 14424 11060 14436
rect 11112 14424 11118 14476
rect 11698 14424 11704 14476
rect 11756 14464 11762 14476
rect 12069 14467 12127 14473
rect 12069 14464 12081 14467
rect 11756 14436 12081 14464
rect 11756 14424 11762 14436
rect 12069 14433 12081 14436
rect 12115 14433 12127 14467
rect 12069 14427 12127 14433
rect 12621 14467 12679 14473
rect 12621 14433 12633 14467
rect 12667 14464 12679 14467
rect 12894 14464 12900 14476
rect 12667 14436 12900 14464
rect 12667 14433 12679 14436
rect 12621 14427 12679 14433
rect 12894 14424 12900 14436
rect 12952 14424 12958 14476
rect 14274 14464 14280 14476
rect 14235 14436 14280 14464
rect 14274 14424 14280 14436
rect 14332 14424 14338 14476
rect 15356 14467 15414 14473
rect 15356 14433 15368 14467
rect 15402 14464 15414 14467
rect 15470 14464 15476 14476
rect 15402 14436 15476 14464
rect 15402 14433 15414 14436
rect 15356 14427 15414 14433
rect 15470 14424 15476 14436
rect 15528 14424 15534 14476
rect 17310 14424 17316 14476
rect 17368 14464 17374 14476
rect 18138 14464 18144 14476
rect 17368 14436 18144 14464
rect 17368 14424 17374 14436
rect 18138 14424 18144 14436
rect 18196 14424 18202 14476
rect 18506 14424 18512 14476
rect 18564 14464 18570 14476
rect 18601 14467 18659 14473
rect 18601 14464 18613 14467
rect 18564 14436 18613 14464
rect 18564 14424 18570 14436
rect 18601 14433 18613 14436
rect 18647 14433 18659 14467
rect 19702 14464 19708 14476
rect 19663 14436 19708 14464
rect 18601 14427 18659 14433
rect 19702 14424 19708 14436
rect 19760 14424 19766 14476
rect 24581 14467 24639 14473
rect 24581 14433 24593 14467
rect 24627 14464 24639 14467
rect 24670 14464 24676 14476
rect 24627 14436 24676 14464
rect 24627 14433 24639 14436
rect 24581 14427 24639 14433
rect 24670 14424 24676 14436
rect 24728 14424 24734 14476
rect 6362 14356 6368 14408
rect 6420 14396 6426 14408
rect 10505 14399 10563 14405
rect 10505 14396 10517 14399
rect 6420 14368 10517 14396
rect 6420 14356 6426 14368
rect 10505 14365 10517 14368
rect 10551 14396 10563 14399
rect 10778 14396 10784 14408
rect 10551 14368 10784 14396
rect 10551 14365 10563 14368
rect 10505 14359 10563 14365
rect 10778 14356 10784 14368
rect 10836 14356 10842 14408
rect 12805 14399 12863 14405
rect 12805 14365 12817 14399
rect 12851 14396 12863 14399
rect 14182 14396 14188 14408
rect 12851 14368 14188 14396
rect 12851 14365 12863 14368
rect 12805 14359 12863 14365
rect 14182 14356 14188 14368
rect 14240 14356 14246 14408
rect 14369 14399 14427 14405
rect 14369 14365 14381 14399
rect 14415 14396 14427 14399
rect 14642 14396 14648 14408
rect 14415 14368 14648 14396
rect 14415 14365 14427 14368
rect 14369 14359 14427 14365
rect 14642 14356 14648 14368
rect 14700 14356 14706 14408
rect 16942 14396 16948 14408
rect 16903 14368 16948 14396
rect 16942 14356 16948 14368
rect 17000 14356 17006 14408
rect 18782 14396 18788 14408
rect 18743 14368 18788 14396
rect 18782 14356 18788 14368
rect 18840 14356 18846 14408
rect 3878 14288 3884 14340
rect 3936 14328 3942 14340
rect 7098 14328 7104 14340
rect 3936 14300 7104 14328
rect 3936 14288 3942 14300
rect 7098 14288 7104 14300
rect 7156 14288 7162 14340
rect 9493 14331 9551 14337
rect 9493 14297 9505 14331
rect 9539 14328 9551 14331
rect 9582 14328 9588 14340
rect 9539 14300 9588 14328
rect 9539 14297 9551 14300
rect 9493 14291 9551 14297
rect 9582 14288 9588 14300
rect 9640 14328 9646 14340
rect 10229 14331 10287 14337
rect 10229 14328 10241 14331
rect 9640 14300 10241 14328
rect 9640 14288 9646 14300
rect 10229 14297 10241 14300
rect 10275 14328 10287 14331
rect 10962 14328 10968 14340
rect 10275 14300 10968 14328
rect 10275 14297 10287 14300
rect 10229 14291 10287 14297
rect 10962 14288 10968 14300
rect 11020 14328 11026 14340
rect 11146 14328 11152 14340
rect 11020 14300 11152 14328
rect 11020 14288 11026 14300
rect 11146 14288 11152 14300
rect 11204 14328 11210 14340
rect 13446 14328 13452 14340
rect 11204 14300 13452 14328
rect 11204 14288 11210 14300
rect 13446 14288 13452 14300
rect 13504 14288 13510 14340
rect 6546 14220 6552 14272
rect 6604 14260 6610 14272
rect 6779 14263 6837 14269
rect 6779 14260 6791 14263
rect 6604 14232 6791 14260
rect 6604 14220 6610 14232
rect 6779 14229 6791 14232
rect 6825 14229 6837 14263
rect 7834 14260 7840 14272
rect 7747 14232 7840 14260
rect 6779 14223 6837 14229
rect 7834 14220 7840 14232
rect 7892 14260 7898 14272
rect 8251 14263 8309 14269
rect 8251 14260 8263 14263
rect 7892 14232 8263 14260
rect 7892 14220 7898 14232
rect 8251 14229 8263 14232
rect 8297 14229 8309 14263
rect 8251 14223 8309 14229
rect 16025 14263 16083 14269
rect 16025 14229 16037 14263
rect 16071 14260 16083 14263
rect 16206 14260 16212 14272
rect 16071 14232 16212 14260
rect 16071 14229 16083 14232
rect 16025 14223 16083 14229
rect 16206 14220 16212 14232
rect 16264 14220 16270 14272
rect 19889 14263 19947 14269
rect 19889 14229 19901 14263
rect 19935 14260 19947 14263
rect 20070 14260 20076 14272
rect 19935 14232 20076 14260
rect 19935 14229 19947 14232
rect 19889 14223 19947 14229
rect 20070 14220 20076 14232
rect 20128 14220 20134 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 14093 14059 14151 14065
rect 14093 14025 14105 14059
rect 14139 14056 14151 14059
rect 14274 14056 14280 14068
rect 14139 14028 14280 14056
rect 14139 14025 14151 14028
rect 14093 14019 14151 14025
rect 14274 14016 14280 14028
rect 14332 14056 14338 14068
rect 14369 14059 14427 14065
rect 14369 14056 14381 14059
rect 14332 14028 14381 14056
rect 14332 14016 14338 14028
rect 14369 14025 14381 14028
rect 14415 14025 14427 14059
rect 14369 14019 14427 14025
rect 14829 14059 14887 14065
rect 14829 14025 14841 14059
rect 14875 14056 14887 14059
rect 15286 14056 15292 14068
rect 14875 14028 15292 14056
rect 14875 14025 14887 14028
rect 14829 14019 14887 14025
rect 15286 14016 15292 14028
rect 15344 14016 15350 14068
rect 15378 14016 15384 14068
rect 15436 14056 15442 14068
rect 15436 14028 15481 14056
rect 15436 14016 15442 14028
rect 18138 14016 18144 14068
rect 18196 14056 18202 14068
rect 18969 14059 19027 14065
rect 18969 14056 18981 14059
rect 18196 14028 18981 14056
rect 18196 14016 18202 14028
rect 18969 14025 18981 14028
rect 19015 14056 19027 14059
rect 19061 14059 19119 14065
rect 19061 14056 19073 14059
rect 19015 14028 19073 14056
rect 19015 14025 19027 14028
rect 18969 14019 19027 14025
rect 19061 14025 19073 14028
rect 19107 14025 19119 14059
rect 19061 14019 19119 14025
rect 24581 14059 24639 14065
rect 24581 14025 24593 14059
rect 24627 14056 24639 14059
rect 24670 14056 24676 14068
rect 24627 14028 24676 14056
rect 24627 14025 24639 14028
rect 24581 14019 24639 14025
rect 24670 14016 24676 14028
rect 24728 14056 24734 14068
rect 27614 14056 27620 14068
rect 24728 14028 27620 14056
rect 24728 14016 24734 14028
rect 27614 14016 27620 14028
rect 27672 14016 27678 14068
rect 9398 13948 9404 14000
rect 9456 13988 9462 14000
rect 10686 13988 10692 14000
rect 9456 13960 10692 13988
rect 9456 13948 9462 13960
rect 10686 13948 10692 13960
rect 10744 13988 10750 14000
rect 11238 13988 11244 14000
rect 10744 13960 11244 13988
rect 10744 13948 10750 13960
rect 11238 13948 11244 13960
rect 11296 13948 11302 14000
rect 20070 13988 20076 14000
rect 18616 13960 20076 13988
rect 7834 13920 7840 13932
rect 7795 13892 7840 13920
rect 7834 13880 7840 13892
rect 7892 13880 7898 13932
rect 8202 13920 8208 13932
rect 8163 13892 8208 13920
rect 8202 13880 8208 13892
rect 8260 13880 8266 13932
rect 9950 13880 9956 13932
rect 10008 13920 10014 13932
rect 10008 13892 13952 13920
rect 10008 13880 10014 13892
rect 1464 13855 1522 13861
rect 1464 13821 1476 13855
rect 1510 13852 1522 13855
rect 1854 13852 1860 13864
rect 1510 13824 1860 13852
rect 1510 13821 1522 13824
rect 1464 13815 1522 13821
rect 1854 13812 1860 13824
rect 1912 13812 1918 13864
rect 9306 13852 9312 13864
rect 9267 13824 9312 13852
rect 9306 13812 9312 13824
rect 9364 13812 9370 13864
rect 9674 13852 9680 13864
rect 9635 13824 9680 13852
rect 9674 13812 9680 13824
rect 9732 13812 9738 13864
rect 11054 13812 11060 13864
rect 11112 13852 11118 13864
rect 11149 13855 11207 13861
rect 11149 13852 11161 13855
rect 11112 13824 11161 13852
rect 11112 13812 11118 13824
rect 11149 13821 11161 13824
rect 11195 13852 11207 13855
rect 12066 13852 12072 13864
rect 11195 13824 12072 13852
rect 11195 13821 11207 13824
rect 11149 13815 11207 13821
rect 12066 13812 12072 13824
rect 12124 13812 12130 13864
rect 13173 13855 13231 13861
rect 13173 13821 13185 13855
rect 13219 13852 13231 13855
rect 13814 13852 13820 13864
rect 13219 13824 13820 13852
rect 13219 13821 13231 13824
rect 13173 13815 13231 13821
rect 13814 13812 13820 13824
rect 13872 13812 13878 13864
rect 13924 13796 13952 13892
rect 15286 13880 15292 13932
rect 15344 13920 15350 13932
rect 16117 13923 16175 13929
rect 16117 13920 16129 13923
rect 15344 13892 16129 13920
rect 15344 13880 15350 13892
rect 16117 13889 16129 13892
rect 16163 13889 16175 13923
rect 16117 13883 16175 13889
rect 16761 13923 16819 13929
rect 16761 13889 16773 13923
rect 16807 13920 16819 13923
rect 16942 13920 16948 13932
rect 16807 13892 16948 13920
rect 16807 13889 16819 13892
rect 16761 13883 16819 13889
rect 16942 13880 16948 13892
rect 17000 13880 17006 13932
rect 17681 13923 17739 13929
rect 17681 13889 17693 13923
rect 17727 13920 17739 13923
rect 18616 13920 18644 13960
rect 20070 13948 20076 13960
rect 20128 13948 20134 14000
rect 22738 13948 22744 14000
rect 22796 13988 22802 14000
rect 24811 13991 24869 13997
rect 24811 13988 24823 13991
rect 22796 13960 24823 13988
rect 22796 13948 22802 13960
rect 24811 13957 24823 13960
rect 24857 13957 24869 13991
rect 24811 13951 24869 13957
rect 17727 13892 18644 13920
rect 17727 13889 17739 13892
rect 17681 13883 17739 13889
rect 14988 13855 15046 13861
rect 14988 13821 15000 13855
rect 15034 13852 15046 13855
rect 15378 13852 15384 13864
rect 15034 13824 15384 13852
rect 15034 13821 15046 13824
rect 14988 13815 15046 13821
rect 15378 13812 15384 13824
rect 15436 13812 15442 13864
rect 18616 13861 18644 13892
rect 18690 13880 18696 13932
rect 18748 13920 18754 13932
rect 19702 13920 19708 13932
rect 18748 13892 19708 13920
rect 18748 13880 18754 13892
rect 19702 13880 19708 13892
rect 19760 13880 19766 13932
rect 24596 13892 25268 13920
rect 20254 13861 20260 13864
rect 18325 13855 18383 13861
rect 18325 13821 18337 13855
rect 18371 13821 18383 13855
rect 18325 13815 18383 13821
rect 18601 13855 18659 13861
rect 18601 13821 18613 13855
rect 18647 13821 18659 13855
rect 20232 13855 20260 13861
rect 20232 13852 20244 13855
rect 20167 13824 20244 13852
rect 18601 13815 18659 13821
rect 20232 13821 20244 13824
rect 20312 13852 20318 13864
rect 20625 13855 20683 13861
rect 20625 13852 20637 13855
rect 20312 13824 20637 13852
rect 20232 13815 20260 13821
rect 4154 13744 4160 13796
rect 4212 13784 4218 13796
rect 6638 13784 6644 13796
rect 4212 13756 6644 13784
rect 4212 13744 4218 13756
rect 6638 13744 6644 13756
rect 6696 13784 6702 13796
rect 7009 13787 7067 13793
rect 7009 13784 7021 13787
rect 6696 13756 7021 13784
rect 6696 13744 6702 13756
rect 7009 13753 7021 13756
rect 7055 13753 7067 13787
rect 7009 13747 7067 13753
rect 7653 13787 7711 13793
rect 7653 13753 7665 13787
rect 7699 13784 7711 13787
rect 7929 13787 7987 13793
rect 7929 13784 7941 13787
rect 7699 13756 7941 13784
rect 7699 13753 7711 13756
rect 7653 13747 7711 13753
rect 7929 13753 7941 13756
rect 7975 13784 7987 13787
rect 8570 13784 8576 13796
rect 7975 13756 8576 13784
rect 7975 13753 7987 13756
rect 7929 13747 7987 13753
rect 1535 13719 1593 13725
rect 1535 13685 1547 13719
rect 1581 13716 1593 13719
rect 6178 13716 6184 13728
rect 1581 13688 6184 13716
rect 1581 13685 1593 13688
rect 1535 13679 1593 13685
rect 6178 13676 6184 13688
rect 6236 13676 6242 13728
rect 7024 13716 7052 13747
rect 8570 13744 8576 13756
rect 8628 13744 8634 13796
rect 9766 13784 9772 13796
rect 8680 13756 9772 13784
rect 8680 13716 8708 13756
rect 9766 13744 9772 13756
rect 9824 13744 9830 13796
rect 10134 13744 10140 13796
rect 10192 13784 10198 13796
rect 10321 13787 10379 13793
rect 10321 13784 10333 13787
rect 10192 13756 10333 13784
rect 10192 13744 10198 13756
rect 10321 13753 10333 13756
rect 10367 13753 10379 13787
rect 10321 13747 10379 13753
rect 11698 13744 11704 13796
rect 11756 13784 11762 13796
rect 12161 13787 12219 13793
rect 12161 13784 12173 13787
rect 11756 13756 12173 13784
rect 11756 13744 11762 13756
rect 12161 13753 12173 13756
rect 12207 13784 12219 13787
rect 13354 13784 13360 13796
rect 12207 13756 13360 13784
rect 12207 13753 12219 13756
rect 12161 13747 12219 13753
rect 13354 13744 13360 13756
rect 13412 13744 13418 13796
rect 13906 13744 13912 13796
rect 13964 13784 13970 13796
rect 15470 13784 15476 13796
rect 13964 13756 15476 13784
rect 13964 13744 13970 13756
rect 15470 13744 15476 13756
rect 15528 13784 15534 13796
rect 15749 13787 15807 13793
rect 15749 13784 15761 13787
rect 15528 13756 15761 13784
rect 15528 13744 15534 13756
rect 15749 13753 15761 13756
rect 15795 13753 15807 13787
rect 16206 13784 16212 13796
rect 16167 13756 16212 13784
rect 15749 13747 15807 13753
rect 16206 13744 16212 13756
rect 16264 13744 16270 13796
rect 17126 13744 17132 13796
rect 17184 13784 17190 13796
rect 17773 13787 17831 13793
rect 17773 13784 17785 13787
rect 17184 13756 17785 13784
rect 17184 13744 17190 13756
rect 17773 13753 17785 13756
rect 17819 13753 17831 13787
rect 18340 13784 18368 13815
rect 20254 13812 20260 13815
rect 20312 13812 20318 13824
rect 20625 13821 20637 13824
rect 20671 13821 20683 13855
rect 20625 13815 20683 13821
rect 21244 13855 21302 13861
rect 21244 13821 21256 13855
rect 21290 13852 21302 13855
rect 22624 13855 22682 13861
rect 21290 13824 21496 13852
rect 21290 13821 21302 13824
rect 21244 13815 21302 13821
rect 17773 13747 17831 13753
rect 18202 13756 18368 13784
rect 18969 13787 19027 13793
rect 8846 13716 8852 13728
rect 7024 13688 8708 13716
rect 8807 13688 8852 13716
rect 8846 13676 8852 13688
rect 8904 13676 8910 13728
rect 9030 13676 9036 13728
rect 9088 13716 9094 13728
rect 9125 13719 9183 13725
rect 9125 13716 9137 13719
rect 9088 13688 9137 13716
rect 9088 13676 9094 13688
rect 9125 13685 9137 13688
rect 9171 13716 9183 13719
rect 9674 13716 9680 13728
rect 9171 13688 9680 13716
rect 9171 13685 9183 13688
rect 9125 13679 9183 13685
rect 9674 13676 9680 13688
rect 9732 13676 9738 13728
rect 11330 13716 11336 13728
rect 11291 13688 11336 13716
rect 11330 13676 11336 13688
rect 11388 13676 11394 13728
rect 12713 13719 12771 13725
rect 12713 13685 12725 13719
rect 12759 13716 12771 13719
rect 12894 13716 12900 13728
rect 12759 13688 12900 13716
rect 12759 13685 12771 13688
rect 12713 13679 12771 13685
rect 12894 13676 12900 13688
rect 12952 13676 12958 13728
rect 13081 13719 13139 13725
rect 13081 13685 13093 13719
rect 13127 13716 13139 13719
rect 13538 13716 13544 13728
rect 13127 13688 13544 13716
rect 13127 13685 13139 13688
rect 13081 13679 13139 13685
rect 13538 13676 13544 13688
rect 13596 13676 13602 13728
rect 14826 13676 14832 13728
rect 14884 13716 14890 13728
rect 15059 13719 15117 13725
rect 15059 13716 15071 13719
rect 14884 13688 15071 13716
rect 14884 13676 14890 13688
rect 15059 13685 15071 13688
rect 15105 13685 15117 13719
rect 17034 13716 17040 13728
rect 16995 13688 17040 13716
rect 15059 13679 15117 13685
rect 17034 13676 17040 13688
rect 17092 13676 17098 13728
rect 17494 13716 17500 13728
rect 17455 13688 17500 13716
rect 17494 13676 17500 13688
rect 17552 13716 17558 13728
rect 17681 13719 17739 13725
rect 17681 13716 17693 13719
rect 17552 13688 17693 13716
rect 17552 13676 17558 13688
rect 17681 13685 17693 13688
rect 17727 13685 17739 13719
rect 17788 13716 17816 13747
rect 18202 13716 18230 13756
rect 18969 13753 18981 13787
rect 19015 13784 19027 13787
rect 21082 13784 21088 13796
rect 19015 13756 21088 13784
rect 19015 13753 19027 13756
rect 18969 13747 19027 13753
rect 21082 13744 21088 13756
rect 21140 13744 21146 13796
rect 21468 13784 21496 13824
rect 22624 13821 22636 13855
rect 22670 13852 22682 13855
rect 24596 13852 24624 13892
rect 24708 13855 24766 13861
rect 24708 13852 24720 13855
rect 22670 13824 23152 13852
rect 24596 13824 24720 13852
rect 22670 13821 22682 13824
rect 22624 13815 22682 13821
rect 21542 13784 21548 13796
rect 21468 13756 21548 13784
rect 21542 13744 21548 13756
rect 21600 13784 21606 13796
rect 23124 13793 23152 13824
rect 24708 13821 24720 13824
rect 24754 13821 24766 13855
rect 24708 13815 24766 13821
rect 21637 13787 21695 13793
rect 21637 13784 21649 13787
rect 21600 13756 21649 13784
rect 21600 13744 21606 13756
rect 21637 13753 21649 13756
rect 21683 13753 21695 13787
rect 23109 13787 23167 13793
rect 23109 13784 23121 13787
rect 23019 13756 23121 13784
rect 21637 13747 21695 13753
rect 23109 13753 23121 13756
rect 23155 13784 23167 13787
rect 23382 13784 23388 13796
rect 23155 13756 23388 13784
rect 23155 13753 23167 13756
rect 23109 13747 23167 13753
rect 23382 13744 23388 13756
rect 23440 13744 23446 13796
rect 25240 13793 25268 13892
rect 25225 13787 25283 13793
rect 25225 13784 25237 13787
rect 25135 13756 25237 13784
rect 25225 13753 25237 13756
rect 25271 13784 25283 13787
rect 25682 13784 25688 13796
rect 25271 13756 25688 13784
rect 25271 13753 25283 13756
rect 25225 13747 25283 13753
rect 25682 13744 25688 13756
rect 25740 13744 25746 13796
rect 18322 13716 18328 13728
rect 17788 13688 18230 13716
rect 18283 13688 18328 13716
rect 17681 13679 17739 13685
rect 18322 13676 18328 13688
rect 18380 13676 18386 13728
rect 18414 13676 18420 13728
rect 18472 13716 18478 13728
rect 20303 13719 20361 13725
rect 20303 13716 20315 13719
rect 18472 13688 20315 13716
rect 18472 13676 18478 13688
rect 20303 13685 20315 13688
rect 20349 13685 20361 13719
rect 20303 13679 20361 13685
rect 21315 13719 21373 13725
rect 21315 13685 21327 13719
rect 21361 13716 21373 13719
rect 22278 13716 22284 13728
rect 21361 13688 22284 13716
rect 21361 13685 21373 13688
rect 21315 13679 21373 13685
rect 22278 13676 22284 13688
rect 22336 13676 22342 13728
rect 22462 13676 22468 13728
rect 22520 13716 22526 13728
rect 22695 13719 22753 13725
rect 22695 13716 22707 13719
rect 22520 13688 22707 13716
rect 22520 13676 22526 13688
rect 22695 13685 22707 13688
rect 22741 13685 22753 13719
rect 22695 13679 22753 13685
rect 23661 13719 23719 13725
rect 23661 13685 23673 13719
rect 23707 13716 23719 13719
rect 23750 13716 23756 13728
rect 23707 13688 23756 13716
rect 23707 13685 23719 13688
rect 23661 13679 23719 13685
rect 23750 13676 23756 13688
rect 23808 13676 23814 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 9674 13472 9680 13524
rect 9732 13512 9738 13524
rect 9732 13484 9904 13512
rect 9732 13472 9738 13484
rect 6365 13447 6423 13453
rect 6365 13413 6377 13447
rect 6411 13444 6423 13447
rect 6546 13444 6552 13456
rect 6411 13416 6552 13444
rect 6411 13413 6423 13416
rect 6365 13407 6423 13413
rect 6546 13404 6552 13416
rect 6604 13404 6610 13456
rect 6638 13404 6644 13456
rect 6696 13444 6702 13456
rect 6696 13416 6741 13444
rect 6696 13404 6702 13416
rect 7650 13404 7656 13456
rect 7708 13444 7714 13456
rect 8205 13447 8263 13453
rect 8205 13444 8217 13447
rect 7708 13416 8217 13444
rect 7708 13404 7714 13416
rect 8205 13413 8217 13416
rect 8251 13444 8263 13447
rect 9306 13444 9312 13456
rect 8251 13416 9312 13444
rect 8251 13413 8263 13416
rect 8205 13407 8263 13413
rect 9306 13404 9312 13416
rect 9364 13404 9370 13456
rect 9876 13453 9904 13484
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 13872 13484 13917 13512
rect 13872 13472 13878 13484
rect 16482 13472 16488 13524
rect 16540 13512 16546 13524
rect 16577 13515 16635 13521
rect 16577 13512 16589 13515
rect 16540 13484 16589 13512
rect 16540 13472 16546 13484
rect 16577 13481 16589 13484
rect 16623 13481 16635 13515
rect 16577 13475 16635 13481
rect 17586 13472 17592 13524
rect 17644 13512 17650 13524
rect 18693 13515 18751 13521
rect 18693 13512 18705 13515
rect 17644 13484 18705 13512
rect 17644 13472 17650 13484
rect 18693 13481 18705 13484
rect 18739 13481 18751 13515
rect 18693 13475 18751 13481
rect 20806 13472 20812 13524
rect 20864 13512 20870 13524
rect 20993 13515 21051 13521
rect 20993 13512 21005 13515
rect 20864 13484 21005 13512
rect 20864 13472 20870 13484
rect 20993 13481 21005 13484
rect 21039 13481 21051 13515
rect 20993 13475 21051 13481
rect 22646 13472 22652 13524
rect 22704 13521 22710 13524
rect 22704 13515 22753 13521
rect 22704 13481 22707 13515
rect 22741 13481 22753 13515
rect 22704 13475 22753 13481
rect 22704 13472 22710 13475
rect 9861 13447 9919 13453
rect 9861 13413 9873 13447
rect 9907 13413 9919 13447
rect 9861 13407 9919 13413
rect 9950 13404 9956 13456
rect 10008 13444 10014 13456
rect 11057 13447 11115 13453
rect 11057 13444 11069 13447
rect 10008 13416 11069 13444
rect 10008 13404 10014 13416
rect 11057 13413 11069 13416
rect 11103 13413 11115 13447
rect 11057 13407 11115 13413
rect 13538 13404 13544 13456
rect 13596 13444 13602 13456
rect 15610 13447 15668 13453
rect 15610 13444 15622 13447
rect 13596 13416 15622 13444
rect 13596 13404 13602 13416
rect 15610 13413 15622 13416
rect 15656 13444 15668 13447
rect 15746 13444 15752 13456
rect 15656 13416 15752 13444
rect 15656 13413 15668 13416
rect 15610 13407 15668 13413
rect 15746 13404 15752 13416
rect 15804 13404 15810 13456
rect 17034 13444 17040 13456
rect 16995 13416 17040 13444
rect 17034 13404 17040 13416
rect 17092 13404 17098 13456
rect 17218 13404 17224 13456
rect 17276 13444 17282 13456
rect 18233 13447 18291 13453
rect 18233 13444 18245 13447
rect 17276 13416 18245 13444
rect 17276 13404 17282 13416
rect 18233 13413 18245 13416
rect 18279 13444 18291 13447
rect 18506 13444 18512 13456
rect 18279 13416 18512 13444
rect 18279 13413 18291 13416
rect 18233 13407 18291 13413
rect 18506 13404 18512 13416
rect 18564 13444 18570 13456
rect 18564 13416 19104 13444
rect 18564 13404 18570 13416
rect 19076 13388 19104 13416
rect 8754 13336 8760 13388
rect 8812 13376 8818 13388
rect 9490 13376 9496 13388
rect 8812 13348 9496 13376
rect 8812 13336 8818 13348
rect 9490 13336 9496 13348
rect 9548 13336 9554 13388
rect 11698 13336 11704 13388
rect 11756 13376 11762 13388
rect 12066 13376 12072 13388
rect 11756 13348 12072 13376
rect 11756 13336 11762 13348
rect 12066 13336 12072 13348
rect 12124 13336 12130 13388
rect 12526 13376 12532 13388
rect 12487 13348 12532 13376
rect 12526 13336 12532 13348
rect 12584 13336 12590 13388
rect 13081 13379 13139 13385
rect 13081 13345 13093 13379
rect 13127 13376 13139 13379
rect 13262 13376 13268 13388
rect 13127 13348 13268 13376
rect 13127 13345 13139 13348
rect 13081 13339 13139 13345
rect 13262 13336 13268 13348
rect 13320 13336 13326 13388
rect 13449 13379 13507 13385
rect 13449 13345 13461 13379
rect 13495 13376 13507 13379
rect 13630 13376 13636 13388
rect 13495 13348 13636 13376
rect 13495 13345 13507 13348
rect 13449 13339 13507 13345
rect 13630 13336 13636 13348
rect 13688 13336 13694 13388
rect 16206 13376 16212 13388
rect 16119 13348 16212 13376
rect 16206 13336 16212 13348
rect 16264 13376 16270 13388
rect 17402 13376 17408 13388
rect 16264 13348 17408 13376
rect 16264 13336 16270 13348
rect 17402 13336 17408 13348
rect 17460 13336 17466 13388
rect 18874 13376 18880 13388
rect 18835 13348 18880 13376
rect 18874 13336 18880 13348
rect 18932 13336 18938 13388
rect 19058 13376 19064 13388
rect 18971 13348 19064 13376
rect 19058 13336 19064 13348
rect 19116 13336 19122 13388
rect 20901 13379 20959 13385
rect 20901 13345 20913 13379
rect 20947 13345 20959 13379
rect 20901 13339 20959 13345
rect 8110 13308 8116 13320
rect 8071 13280 8116 13308
rect 8110 13268 8116 13280
rect 8168 13268 8174 13320
rect 8202 13268 8208 13320
rect 8260 13308 8266 13320
rect 9769 13311 9827 13317
rect 9769 13308 9781 13311
rect 8260 13280 9781 13308
rect 8260 13268 8266 13280
rect 9769 13277 9781 13280
rect 9815 13308 9827 13311
rect 9950 13308 9956 13320
rect 9815 13280 9956 13308
rect 9815 13277 9827 13280
rect 9769 13271 9827 13277
rect 9950 13268 9956 13280
rect 10008 13268 10014 13320
rect 10045 13311 10103 13317
rect 10045 13277 10057 13311
rect 10091 13277 10103 13311
rect 10045 13271 10103 13277
rect 13541 13311 13599 13317
rect 13541 13277 13553 13311
rect 13587 13308 13599 13311
rect 15289 13311 15347 13317
rect 15289 13308 15301 13311
rect 13587 13280 15301 13308
rect 13587 13277 13599 13280
rect 13541 13271 13599 13277
rect 15289 13277 15301 13280
rect 15335 13308 15347 13311
rect 15378 13308 15384 13320
rect 15335 13280 15384 13308
rect 15335 13277 15347 13280
rect 15289 13271 15347 13277
rect 7101 13243 7159 13249
rect 7101 13209 7113 13243
rect 7147 13240 7159 13243
rect 8220 13240 8248 13268
rect 8662 13240 8668 13252
rect 7147 13212 8248 13240
rect 8575 13212 8668 13240
rect 7147 13209 7159 13212
rect 7101 13203 7159 13209
rect 8662 13200 8668 13212
rect 8720 13240 8726 13252
rect 10060 13240 10088 13271
rect 15378 13268 15384 13280
rect 15436 13268 15442 13320
rect 18892 13308 18920 13336
rect 20916 13308 20944 13339
rect 21266 13336 21272 13388
rect 21324 13376 21330 13388
rect 21361 13379 21419 13385
rect 21361 13376 21373 13379
rect 21324 13348 21373 13376
rect 21324 13336 21330 13348
rect 21361 13345 21373 13348
rect 21407 13345 21419 13379
rect 21361 13339 21419 13345
rect 22624 13379 22682 13385
rect 22624 13345 22636 13379
rect 22670 13376 22682 13379
rect 22830 13376 22836 13388
rect 22670 13348 22836 13376
rect 22670 13345 22682 13348
rect 22624 13339 22682 13345
rect 22830 13336 22836 13348
rect 22888 13336 22894 13388
rect 23636 13379 23694 13385
rect 23636 13345 23648 13379
rect 23682 13376 23694 13379
rect 24210 13376 24216 13388
rect 23682 13348 24216 13376
rect 23682 13345 23694 13348
rect 23636 13339 23694 13345
rect 24210 13336 24216 13348
rect 24268 13336 24274 13388
rect 24648 13379 24706 13385
rect 24648 13345 24660 13379
rect 24694 13376 24706 13379
rect 25222 13376 25228 13388
rect 24694 13348 25228 13376
rect 24694 13345 24706 13348
rect 24648 13339 24706 13345
rect 25222 13336 25228 13348
rect 25280 13336 25286 13388
rect 22186 13308 22192 13320
rect 18892 13280 22192 13308
rect 22186 13268 22192 13280
rect 22244 13268 22250 13320
rect 8720 13212 10088 13240
rect 10781 13243 10839 13249
rect 8720 13200 8726 13212
rect 10781 13209 10793 13243
rect 10827 13240 10839 13243
rect 11054 13240 11060 13252
rect 10827 13212 11060 13240
rect 10827 13209 10839 13212
rect 10781 13203 10839 13209
rect 11054 13200 11060 13212
rect 11112 13200 11118 13252
rect 11606 13200 11612 13252
rect 11664 13240 11670 13252
rect 18690 13240 18696 13252
rect 11664 13212 18696 13240
rect 11664 13200 11670 13212
rect 18690 13200 18696 13212
rect 18748 13200 18754 13252
rect 7926 13172 7932 13184
rect 7887 13144 7932 13172
rect 7926 13132 7932 13144
rect 7984 13132 7990 13184
rect 9030 13172 9036 13184
rect 8991 13144 9036 13172
rect 9030 13132 9036 13144
rect 9088 13132 9094 13184
rect 9490 13172 9496 13184
rect 9451 13144 9496 13172
rect 9490 13132 9496 13144
rect 9548 13132 9554 13184
rect 10962 13132 10968 13184
rect 11020 13172 11026 13184
rect 11517 13175 11575 13181
rect 11517 13172 11529 13175
rect 11020 13144 11529 13172
rect 11020 13132 11026 13144
rect 11517 13141 11529 13144
rect 11563 13141 11575 13175
rect 11517 13135 11575 13141
rect 11698 13132 11704 13184
rect 11756 13172 11762 13184
rect 11885 13175 11943 13181
rect 11885 13172 11897 13175
rect 11756 13144 11897 13172
rect 11756 13132 11762 13144
rect 11885 13141 11897 13144
rect 11931 13141 11943 13175
rect 11885 13135 11943 13141
rect 14274 13132 14280 13184
rect 14332 13172 14338 13184
rect 17494 13172 17500 13184
rect 14332 13144 17500 13172
rect 14332 13132 14338 13144
rect 17494 13132 17500 13144
rect 17552 13132 17558 13184
rect 20162 13132 20168 13184
rect 20220 13172 20226 13184
rect 23707 13175 23765 13181
rect 23707 13172 23719 13175
rect 20220 13144 23719 13172
rect 20220 13132 20226 13144
rect 23707 13141 23719 13144
rect 23753 13141 23765 13175
rect 23707 13135 23765 13141
rect 24026 13132 24032 13184
rect 24084 13172 24090 13184
rect 24719 13175 24777 13181
rect 24719 13172 24731 13175
rect 24084 13144 24731 13172
rect 24084 13132 24090 13144
rect 24719 13141 24731 13144
rect 24765 13141 24777 13175
rect 24719 13135 24777 13141
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 7650 12968 7656 12980
rect 7611 12940 7656 12968
rect 7650 12928 7656 12940
rect 7708 12928 7714 12980
rect 8018 12968 8024 12980
rect 7979 12940 8024 12968
rect 8018 12928 8024 12940
rect 8076 12928 8082 12980
rect 9030 12968 9036 12980
rect 8991 12940 9036 12968
rect 9030 12928 9036 12940
rect 9088 12928 9094 12980
rect 11238 12928 11244 12980
rect 11296 12968 11302 12980
rect 11793 12971 11851 12977
rect 11793 12968 11805 12971
rect 11296 12940 11805 12968
rect 11296 12928 11302 12940
rect 11793 12937 11805 12940
rect 11839 12968 11851 12971
rect 12161 12971 12219 12977
rect 12161 12968 12173 12971
rect 11839 12940 12173 12968
rect 11839 12937 11851 12940
rect 11793 12931 11851 12937
rect 12161 12937 12173 12940
rect 12207 12968 12219 12971
rect 12526 12968 12532 12980
rect 12207 12940 12532 12968
rect 12207 12937 12219 12940
rect 12161 12931 12219 12937
rect 12526 12928 12532 12940
rect 12584 12928 12590 12980
rect 14642 12968 14648 12980
rect 14603 12940 14648 12968
rect 14642 12928 14648 12940
rect 14700 12928 14706 12980
rect 15378 12928 15384 12980
rect 15436 12968 15442 12980
rect 16209 12971 16267 12977
rect 16209 12968 16221 12971
rect 15436 12940 16221 12968
rect 15436 12928 15442 12940
rect 16209 12937 16221 12940
rect 16255 12937 16267 12971
rect 17402 12968 17408 12980
rect 17363 12940 17408 12968
rect 16209 12931 16267 12937
rect 17402 12928 17408 12940
rect 17460 12928 17466 12980
rect 19058 12968 19064 12980
rect 19019 12940 19064 12968
rect 19058 12928 19064 12940
rect 19116 12928 19122 12980
rect 12434 12900 12440 12912
rect 11532 12872 12440 12900
rect 11532 12832 11560 12872
rect 12434 12860 12440 12872
rect 12492 12860 12498 12912
rect 13814 12860 13820 12912
rect 13872 12900 13878 12912
rect 13872 12872 13917 12900
rect 13872 12860 13878 12872
rect 14826 12860 14832 12912
rect 14884 12900 14890 12912
rect 14884 12872 14964 12900
rect 14884 12860 14890 12872
rect 14936 12841 14964 12872
rect 15746 12860 15752 12912
rect 15804 12900 15810 12912
rect 15841 12903 15899 12909
rect 15841 12900 15853 12903
rect 15804 12872 15853 12900
rect 15804 12860 15810 12872
rect 15841 12869 15853 12872
rect 15887 12869 15899 12903
rect 15841 12863 15899 12869
rect 16942 12860 16948 12912
rect 17000 12900 17006 12912
rect 17000 12872 18736 12900
rect 17000 12860 17006 12872
rect 14185 12835 14243 12841
rect 14185 12832 14197 12835
rect 10152 12804 11560 12832
rect 12452 12804 14197 12832
rect 5077 12767 5135 12773
rect 5077 12733 5089 12767
rect 5123 12764 5135 12767
rect 5810 12764 5816 12776
rect 5123 12736 5816 12764
rect 5123 12733 5135 12736
rect 5077 12727 5135 12733
rect 5810 12724 5816 12736
rect 5868 12724 5874 12776
rect 7926 12724 7932 12776
rect 7984 12764 7990 12776
rect 8113 12767 8171 12773
rect 8113 12764 8125 12767
rect 7984 12736 8125 12764
rect 7984 12724 7990 12736
rect 8113 12733 8125 12736
rect 8159 12764 8171 12767
rect 9401 12767 9459 12773
rect 8159 12736 8708 12764
rect 8159 12733 8171 12736
rect 8113 12727 8171 12733
rect 5905 12699 5963 12705
rect 5905 12665 5917 12699
rect 5951 12696 5963 12699
rect 6457 12699 6515 12705
rect 6457 12696 6469 12699
rect 5951 12668 6469 12696
rect 5951 12665 5963 12668
rect 5905 12659 5963 12665
rect 6457 12665 6469 12668
rect 6503 12696 6515 12699
rect 6638 12696 6644 12708
rect 6503 12668 6644 12696
rect 6503 12665 6515 12668
rect 6457 12659 6515 12665
rect 6638 12656 6644 12668
rect 6696 12656 6702 12708
rect 8018 12656 8024 12708
rect 8076 12696 8082 12708
rect 8434 12699 8492 12705
rect 8434 12696 8446 12699
rect 8076 12668 8446 12696
rect 8076 12656 8082 12668
rect 8434 12665 8446 12668
rect 8480 12665 8492 12699
rect 8680 12696 8708 12736
rect 9401 12733 9413 12767
rect 9447 12764 9459 12767
rect 10042 12764 10048 12776
rect 9447 12736 10048 12764
rect 9447 12733 9459 12736
rect 9401 12727 9459 12733
rect 10042 12724 10048 12736
rect 10100 12764 10106 12776
rect 10152 12773 10180 12804
rect 10137 12767 10195 12773
rect 10137 12764 10149 12767
rect 10100 12736 10149 12764
rect 10100 12724 10106 12736
rect 10137 12733 10149 12736
rect 10183 12733 10195 12767
rect 10594 12764 10600 12776
rect 10555 12736 10600 12764
rect 10137 12727 10195 12733
rect 10594 12724 10600 12736
rect 10652 12724 10658 12776
rect 10778 12764 10784 12776
rect 10739 12736 10784 12764
rect 10778 12724 10784 12736
rect 10836 12724 10842 12776
rect 11054 12764 11060 12776
rect 11015 12736 11060 12764
rect 11054 12724 11060 12736
rect 11112 12724 11118 12776
rect 11698 12724 11704 12776
rect 11756 12764 11762 12776
rect 12452 12773 12480 12804
rect 14185 12801 14197 12804
rect 14231 12801 14243 12835
rect 14185 12795 14243 12801
rect 14921 12835 14979 12841
rect 14921 12801 14933 12835
rect 14967 12801 14979 12835
rect 15286 12832 15292 12844
rect 15247 12804 15292 12832
rect 14921 12795 14979 12801
rect 15286 12792 15292 12804
rect 15344 12792 15350 12844
rect 16482 12832 16488 12844
rect 16443 12804 16488 12832
rect 16482 12792 16488 12804
rect 16540 12792 16546 12844
rect 16758 12832 16764 12844
rect 16719 12804 16764 12832
rect 16758 12792 16764 12804
rect 16816 12792 16822 12844
rect 18598 12832 18604 12844
rect 18559 12804 18604 12832
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 18708 12832 18736 12872
rect 19426 12860 19432 12912
rect 19484 12900 19490 12912
rect 23799 12903 23857 12909
rect 23799 12900 23811 12903
rect 19484 12872 23811 12900
rect 19484 12860 19490 12872
rect 23799 12869 23811 12872
rect 23845 12869 23857 12903
rect 24581 12903 24639 12909
rect 24581 12900 24593 12903
rect 23799 12863 23857 12869
rect 24044 12872 24593 12900
rect 21269 12835 21327 12841
rect 21269 12832 21281 12835
rect 18708 12804 19840 12832
rect 12437 12767 12495 12773
rect 12437 12764 12449 12767
rect 11756 12736 12449 12764
rect 11756 12724 11762 12736
rect 12437 12733 12449 12736
rect 12483 12733 12495 12767
rect 12437 12727 12495 12733
rect 12526 12724 12532 12776
rect 12584 12764 12590 12776
rect 12897 12767 12955 12773
rect 12897 12764 12909 12767
rect 12584 12736 12909 12764
rect 12584 12724 12590 12736
rect 12897 12733 12909 12736
rect 12943 12733 12955 12767
rect 13262 12764 13268 12776
rect 13223 12736 13268 12764
rect 12897 12727 12955 12733
rect 13262 12724 13268 12736
rect 13320 12724 13326 12776
rect 13446 12724 13452 12776
rect 13504 12764 13510 12776
rect 19812 12773 19840 12804
rect 20364 12804 21281 12832
rect 13633 12767 13691 12773
rect 13633 12764 13645 12767
rect 13504 12736 13645 12764
rect 13504 12724 13510 12736
rect 13633 12733 13645 12736
rect 13679 12733 13691 12767
rect 13633 12727 13691 12733
rect 19797 12767 19855 12773
rect 19797 12733 19809 12767
rect 19843 12764 19855 12767
rect 19889 12767 19947 12773
rect 19889 12764 19901 12767
rect 19843 12736 19901 12764
rect 19843 12733 19855 12736
rect 19797 12727 19855 12733
rect 19889 12733 19901 12736
rect 19935 12733 19947 12767
rect 19889 12727 19947 12733
rect 20070 12724 20076 12776
rect 20128 12764 20134 12776
rect 20364 12773 20392 12804
rect 21269 12801 21281 12804
rect 21315 12832 21327 12835
rect 21358 12832 21364 12844
rect 21315 12804 21364 12832
rect 21315 12801 21327 12804
rect 21269 12795 21327 12801
rect 21358 12792 21364 12804
rect 21416 12832 21422 12844
rect 21416 12804 21956 12832
rect 21416 12792 21422 12804
rect 20349 12767 20407 12773
rect 20349 12764 20361 12767
rect 20128 12736 20361 12764
rect 20128 12724 20134 12736
rect 20349 12733 20361 12736
rect 20395 12733 20407 12767
rect 20349 12727 20407 12733
rect 21082 12724 21088 12776
rect 21140 12764 21146 12776
rect 21928 12773 21956 12804
rect 21453 12767 21511 12773
rect 21453 12764 21465 12767
rect 21140 12736 21465 12764
rect 21140 12724 21146 12736
rect 21453 12733 21465 12736
rect 21499 12733 21511 12767
rect 21453 12727 21511 12733
rect 21913 12767 21971 12773
rect 21913 12733 21925 12767
rect 21959 12733 21971 12767
rect 21913 12727 21971 12733
rect 23728 12767 23786 12773
rect 23728 12733 23740 12767
rect 23774 12764 23786 12767
rect 24044 12764 24072 12872
rect 24581 12869 24593 12872
rect 24627 12900 24639 12903
rect 25958 12900 25964 12912
rect 24627 12872 25964 12900
rect 24627 12869 24639 12872
rect 24581 12863 24639 12869
rect 25958 12860 25964 12872
rect 26016 12860 26022 12912
rect 25222 12832 25228 12844
rect 25135 12804 25228 12832
rect 25222 12792 25228 12804
rect 25280 12832 25286 12844
rect 26326 12832 26332 12844
rect 25280 12804 26332 12832
rect 25280 12792 25286 12804
rect 26326 12792 26332 12804
rect 26384 12792 26390 12844
rect 23774 12736 24072 12764
rect 24740 12767 24798 12773
rect 23774 12733 23786 12736
rect 23728 12727 23786 12733
rect 24740 12733 24752 12767
rect 24786 12764 24798 12767
rect 24786 12736 25544 12764
rect 24786 12733 24798 12736
rect 24740 12727 24798 12733
rect 8680 12668 9904 12696
rect 8434 12659 8492 12665
rect 6822 12628 6828 12640
rect 6783 12600 6828 12628
rect 6822 12588 6828 12600
rect 6880 12588 6886 12640
rect 9766 12628 9772 12640
rect 9727 12600 9772 12628
rect 9766 12588 9772 12600
rect 9824 12588 9830 12640
rect 9876 12628 9904 12668
rect 14642 12656 14648 12708
rect 14700 12696 14706 12708
rect 15013 12699 15071 12705
rect 15013 12696 15025 12699
rect 14700 12668 15025 12696
rect 14700 12656 14706 12668
rect 15013 12665 15025 12668
rect 15059 12665 15071 12699
rect 15013 12659 15071 12665
rect 16577 12699 16635 12705
rect 16577 12665 16589 12699
rect 16623 12665 16635 12699
rect 18138 12696 18144 12708
rect 18099 12668 18144 12696
rect 16577 12659 16635 12665
rect 9953 12631 10011 12637
rect 9953 12628 9965 12631
rect 9876 12600 9965 12628
rect 9953 12597 9965 12600
rect 9999 12597 10011 12631
rect 9953 12591 10011 12597
rect 16206 12588 16212 12640
rect 16264 12628 16270 12640
rect 16592 12628 16620 12659
rect 18138 12656 18144 12668
rect 18196 12656 18202 12708
rect 18233 12699 18291 12705
rect 18233 12665 18245 12699
rect 18279 12665 18291 12699
rect 18233 12659 18291 12665
rect 20625 12699 20683 12705
rect 20625 12665 20637 12699
rect 20671 12696 20683 12699
rect 21174 12696 21180 12708
rect 20671 12668 21180 12696
rect 20671 12665 20683 12668
rect 20625 12659 20683 12665
rect 17773 12631 17831 12637
rect 17773 12628 17785 12631
rect 16264 12600 17785 12628
rect 16264 12588 16270 12600
rect 17773 12597 17785 12600
rect 17819 12628 17831 12631
rect 18248 12628 18276 12659
rect 21174 12656 21180 12668
rect 21232 12656 21238 12708
rect 24949 12699 25007 12705
rect 24949 12665 24961 12699
rect 24995 12696 25007 12699
rect 25314 12696 25320 12708
rect 24995 12668 25320 12696
rect 24995 12665 25007 12668
rect 24949 12659 25007 12665
rect 25314 12656 25320 12668
rect 25372 12656 25378 12708
rect 25516 12640 25544 12736
rect 17819 12600 18276 12628
rect 17819 12597 17831 12600
rect 17773 12591 17831 12597
rect 20530 12588 20536 12640
rect 20588 12628 20594 12640
rect 20901 12631 20959 12637
rect 20901 12628 20913 12631
rect 20588 12600 20913 12628
rect 20588 12588 20594 12600
rect 20901 12597 20913 12600
rect 20947 12628 20959 12631
rect 21266 12628 21272 12640
rect 20947 12600 21272 12628
rect 20947 12597 20959 12600
rect 20901 12591 20959 12597
rect 21266 12588 21272 12600
rect 21324 12588 21330 12640
rect 21726 12628 21732 12640
rect 21687 12600 21732 12628
rect 21726 12588 21732 12600
rect 21784 12588 21790 12640
rect 22186 12588 22192 12640
rect 22244 12628 22250 12640
rect 22465 12631 22523 12637
rect 22465 12628 22477 12631
rect 22244 12600 22477 12628
rect 22244 12588 22250 12600
rect 22465 12597 22477 12600
rect 22511 12597 22523 12631
rect 22830 12628 22836 12640
rect 22791 12600 22836 12628
rect 22465 12591 22523 12597
rect 22830 12588 22836 12600
rect 22888 12588 22894 12640
rect 24210 12628 24216 12640
rect 24123 12600 24216 12628
rect 24210 12588 24216 12600
rect 24268 12628 24274 12640
rect 25130 12628 25136 12640
rect 24268 12600 25136 12628
rect 24268 12588 24274 12600
rect 25130 12588 25136 12600
rect 25188 12588 25194 12640
rect 25498 12628 25504 12640
rect 25459 12600 25504 12628
rect 25498 12588 25504 12600
rect 25556 12588 25562 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 6822 12384 6828 12436
rect 6880 12424 6886 12436
rect 7101 12427 7159 12433
rect 7101 12424 7113 12427
rect 6880 12396 7113 12424
rect 6880 12384 6886 12396
rect 7101 12393 7113 12396
rect 7147 12393 7159 12427
rect 7558 12424 7564 12436
rect 7471 12396 7564 12424
rect 7101 12387 7159 12393
rect 7558 12384 7564 12396
rect 7616 12424 7622 12436
rect 8110 12424 8116 12436
rect 7616 12396 8116 12424
rect 7616 12384 7622 12396
rect 8110 12384 8116 12396
rect 8168 12384 8174 12436
rect 9861 12427 9919 12433
rect 9861 12424 9873 12427
rect 8449 12396 9873 12424
rect 5810 12316 5816 12368
rect 5868 12356 5874 12368
rect 6178 12356 6184 12368
rect 5868 12328 6184 12356
rect 5868 12316 5874 12328
rect 6178 12316 6184 12328
rect 6236 12356 6242 12368
rect 6273 12359 6331 12365
rect 6273 12356 6285 12359
rect 6236 12328 6285 12356
rect 6236 12316 6242 12328
rect 6273 12325 6285 12328
rect 6319 12356 6331 12359
rect 6917 12359 6975 12365
rect 6917 12356 6929 12359
rect 6319 12328 6929 12356
rect 6319 12325 6331 12328
rect 6273 12319 6331 12325
rect 6917 12325 6929 12328
rect 6963 12325 6975 12359
rect 6917 12319 6975 12325
rect 7906 12359 7964 12365
rect 7906 12325 7918 12359
rect 7952 12356 7964 12359
rect 8018 12356 8024 12368
rect 7952 12328 8024 12356
rect 7952 12325 7964 12328
rect 7906 12319 7964 12325
rect 8018 12316 8024 12328
rect 8076 12316 8082 12368
rect 6825 12291 6883 12297
rect 6825 12257 6837 12291
rect 6871 12288 6883 12291
rect 7558 12288 7564 12300
rect 6871 12260 7564 12288
rect 6871 12257 6883 12260
rect 6825 12251 6883 12257
rect 7558 12248 7564 12260
rect 7616 12248 7622 12300
rect 7653 12291 7711 12297
rect 7653 12257 7665 12291
rect 7699 12288 7711 12291
rect 7742 12288 7748 12300
rect 7699 12260 7748 12288
rect 7699 12257 7711 12260
rect 7653 12251 7711 12257
rect 7742 12248 7748 12260
rect 7800 12288 7806 12300
rect 8449 12288 8477 12396
rect 9861 12393 9873 12396
rect 9907 12393 9919 12427
rect 14826 12424 14832 12436
rect 14787 12396 14832 12424
rect 9861 12387 9919 12393
rect 14826 12384 14832 12396
rect 14884 12384 14890 12436
rect 15427 12427 15485 12433
rect 15427 12393 15439 12427
rect 15473 12424 15485 12427
rect 17681 12427 17739 12433
rect 17681 12424 17693 12427
rect 15473 12396 17693 12424
rect 15473 12393 15485 12396
rect 15427 12387 15485 12393
rect 17681 12393 17693 12396
rect 17727 12424 17739 12427
rect 18138 12424 18144 12436
rect 17727 12396 18144 12424
rect 17727 12393 17739 12396
rect 17681 12387 17739 12393
rect 18138 12384 18144 12396
rect 18196 12384 18202 12436
rect 19518 12384 19524 12436
rect 19576 12424 19582 12436
rect 19705 12427 19763 12433
rect 19705 12424 19717 12427
rect 19576 12396 19717 12424
rect 19576 12384 19582 12396
rect 19705 12393 19717 12396
rect 19751 12393 19763 12427
rect 19705 12387 19763 12393
rect 21082 12384 21088 12436
rect 21140 12424 21146 12436
rect 21913 12427 21971 12433
rect 21913 12424 21925 12427
rect 21140 12396 21925 12424
rect 21140 12384 21146 12396
rect 21913 12393 21925 12396
rect 21959 12393 21971 12427
rect 22554 12424 22560 12436
rect 22515 12396 22560 12424
rect 21913 12387 21971 12393
rect 22554 12384 22560 12396
rect 22612 12384 22618 12436
rect 9125 12359 9183 12365
rect 9125 12325 9137 12359
rect 9171 12356 9183 12359
rect 9582 12356 9588 12368
rect 9171 12328 9588 12356
rect 9171 12325 9183 12328
rect 9125 12319 9183 12325
rect 9582 12316 9588 12328
rect 9640 12356 9646 12368
rect 9640 12328 11008 12356
rect 9640 12316 9646 12328
rect 8570 12288 8576 12300
rect 7800 12260 8477 12288
rect 8531 12260 8576 12288
rect 7800 12248 7806 12260
rect 8570 12248 8576 12260
rect 8628 12248 8634 12300
rect 10042 12288 10048 12300
rect 10003 12260 10048 12288
rect 10042 12248 10048 12260
rect 10100 12248 10106 12300
rect 10229 12291 10287 12297
rect 10229 12257 10241 12291
rect 10275 12257 10287 12291
rect 10594 12288 10600 12300
rect 10555 12260 10600 12288
rect 10229 12251 10287 12257
rect 5534 12180 5540 12232
rect 5592 12220 5598 12232
rect 6181 12223 6239 12229
rect 6181 12220 6193 12223
rect 5592 12192 6193 12220
rect 5592 12180 5598 12192
rect 6181 12189 6193 12192
rect 6227 12189 6239 12223
rect 6181 12183 6239 12189
rect 6917 12223 6975 12229
rect 6917 12189 6929 12223
rect 6963 12220 6975 12223
rect 8588 12220 8616 12248
rect 6963 12192 8616 12220
rect 6963 12189 6975 12192
rect 6917 12183 6975 12189
rect 9766 12180 9772 12232
rect 9824 12220 9830 12232
rect 10244 12220 10272 12251
rect 10594 12248 10600 12260
rect 10652 12288 10658 12300
rect 10778 12288 10784 12300
rect 10652 12260 10784 12288
rect 10652 12248 10658 12260
rect 10778 12248 10784 12260
rect 10836 12248 10842 12300
rect 10980 12297 11008 12328
rect 13722 12316 13728 12368
rect 13780 12356 13786 12368
rect 13817 12359 13875 12365
rect 13817 12356 13829 12359
rect 13780 12328 13829 12356
rect 13780 12316 13786 12328
rect 13817 12325 13829 12328
rect 13863 12356 13875 12359
rect 16114 12356 16120 12368
rect 13863 12328 16120 12356
rect 13863 12325 13875 12328
rect 13817 12319 13875 12325
rect 16114 12316 16120 12328
rect 16172 12316 16178 12368
rect 16482 12356 16488 12368
rect 16443 12328 16488 12356
rect 16482 12316 16488 12328
rect 16540 12316 16546 12368
rect 16574 12316 16580 12368
rect 16632 12356 16638 12368
rect 17313 12359 17371 12365
rect 17313 12356 17325 12359
rect 16632 12328 17325 12356
rect 16632 12316 16638 12328
rect 17313 12325 17325 12328
rect 17359 12325 17371 12359
rect 17954 12356 17960 12368
rect 17915 12328 17960 12356
rect 17313 12319 17371 12325
rect 17954 12316 17960 12328
rect 18012 12316 18018 12368
rect 18046 12316 18052 12368
rect 18104 12356 18110 12368
rect 24670 12356 24676 12368
rect 18104 12328 18149 12356
rect 24111 12328 24676 12356
rect 18104 12316 18110 12328
rect 10965 12291 11023 12297
rect 10965 12257 10977 12291
rect 11011 12257 11023 12291
rect 10965 12251 11023 12257
rect 12713 12291 12771 12297
rect 12713 12257 12725 12291
rect 12759 12288 12771 12291
rect 13078 12288 13084 12300
rect 12759 12260 13084 12288
rect 12759 12257 12771 12260
rect 12713 12251 12771 12257
rect 13078 12248 13084 12260
rect 13136 12248 13142 12300
rect 14642 12248 14648 12300
rect 14700 12288 14706 12300
rect 15197 12291 15255 12297
rect 15197 12288 15209 12291
rect 14700 12260 15209 12288
rect 14700 12248 14706 12260
rect 15197 12257 15209 12260
rect 15243 12257 15255 12291
rect 15746 12288 15752 12300
rect 15707 12260 15752 12288
rect 15197 12251 15255 12257
rect 15746 12248 15752 12260
rect 15804 12248 15810 12300
rect 19242 12248 19248 12300
rect 19300 12288 19306 12300
rect 19464 12291 19522 12297
rect 19464 12288 19476 12291
rect 19300 12260 19476 12288
rect 19300 12248 19306 12260
rect 19464 12257 19476 12260
rect 19510 12257 19522 12291
rect 20898 12288 20904 12300
rect 20859 12260 20904 12288
rect 19464 12251 19522 12257
rect 20898 12248 20904 12260
rect 20956 12248 20962 12300
rect 21358 12288 21364 12300
rect 21319 12260 21364 12288
rect 21358 12248 21364 12260
rect 21416 12248 21422 12300
rect 22186 12248 22192 12300
rect 22244 12288 22250 12300
rect 22465 12291 22523 12297
rect 22465 12288 22477 12291
rect 22244 12260 22477 12288
rect 22244 12248 22250 12260
rect 22465 12257 22477 12260
rect 22511 12257 22523 12291
rect 22922 12288 22928 12300
rect 22883 12260 22928 12288
rect 22465 12251 22523 12257
rect 22922 12248 22928 12260
rect 22980 12248 22986 12300
rect 23014 12248 23020 12300
rect 23072 12288 23078 12300
rect 24111 12297 24139 12328
rect 24670 12316 24676 12328
rect 24728 12356 24734 12368
rect 27614 12356 27620 12368
rect 24728 12328 27620 12356
rect 24728 12316 24734 12328
rect 27614 12316 27620 12328
rect 27672 12316 27678 12368
rect 24096 12291 24154 12297
rect 24096 12288 24108 12291
rect 23072 12260 24108 12288
rect 23072 12248 23078 12260
rect 24096 12257 24108 12260
rect 24142 12257 24154 12291
rect 24096 12251 24154 12257
rect 25108 12291 25166 12297
rect 25108 12257 25120 12291
rect 25154 12288 25166 12291
rect 25866 12288 25872 12300
rect 25154 12260 25872 12288
rect 25154 12257 25166 12260
rect 25108 12251 25166 12257
rect 25866 12248 25872 12260
rect 25924 12248 25930 12300
rect 10686 12220 10692 12232
rect 9824 12192 10692 12220
rect 9824 12180 9830 12192
rect 10686 12180 10692 12192
rect 10744 12180 10750 12232
rect 11974 12180 11980 12232
rect 12032 12220 12038 12232
rect 13725 12223 13783 12229
rect 13725 12220 13737 12223
rect 12032 12192 13737 12220
rect 12032 12180 12038 12192
rect 13725 12189 13737 12192
rect 13771 12220 13783 12223
rect 13998 12220 14004 12232
rect 13771 12192 14004 12220
rect 13771 12189 13783 12192
rect 13725 12183 13783 12189
rect 13998 12180 14004 12192
rect 14056 12180 14062 12232
rect 14369 12223 14427 12229
rect 14369 12189 14381 12223
rect 14415 12220 14427 12223
rect 16393 12223 16451 12229
rect 16393 12220 16405 12223
rect 14415 12192 16405 12220
rect 14415 12189 14427 12192
rect 14369 12183 14427 12189
rect 16393 12189 16405 12192
rect 16439 12220 16451 12223
rect 16758 12220 16764 12232
rect 16439 12192 16764 12220
rect 16439 12189 16451 12192
rect 16393 12183 16451 12189
rect 16758 12180 16764 12192
rect 16816 12180 16822 12232
rect 17034 12220 17040 12232
rect 16995 12192 17040 12220
rect 17034 12180 17040 12192
rect 17092 12180 17098 12232
rect 19889 12223 19947 12229
rect 19889 12189 19901 12223
rect 19935 12220 19947 12223
rect 20070 12220 20076 12232
rect 19935 12192 20076 12220
rect 19935 12189 19947 12192
rect 19889 12183 19947 12189
rect 20070 12180 20076 12192
rect 20128 12180 20134 12232
rect 21634 12220 21640 12232
rect 21595 12192 21640 12220
rect 21634 12180 21640 12192
rect 21692 12180 21698 12232
rect 6454 12112 6460 12164
rect 6512 12152 6518 12164
rect 9214 12152 9220 12164
rect 6512 12124 9220 12152
rect 6512 12112 6518 12124
rect 9214 12112 9220 12124
rect 9272 12152 9278 12164
rect 11054 12152 11060 12164
rect 9272 12124 11060 12152
rect 9272 12112 9278 12124
rect 11054 12112 11060 12124
rect 11112 12152 11118 12164
rect 11517 12155 11575 12161
rect 11517 12152 11529 12155
rect 11112 12124 11529 12152
rect 11112 12112 11118 12124
rect 11517 12121 11529 12124
rect 11563 12121 11575 12155
rect 13081 12155 13139 12161
rect 13081 12152 13093 12155
rect 11517 12115 11575 12121
rect 11900 12124 13093 12152
rect 9493 12087 9551 12093
rect 9493 12053 9505 12087
rect 9539 12084 9551 12087
rect 9766 12084 9772 12096
rect 9539 12056 9772 12084
rect 9539 12053 9551 12056
rect 9493 12047 9551 12053
rect 9766 12044 9772 12056
rect 9824 12044 9830 12096
rect 10778 12044 10784 12096
rect 10836 12084 10842 12096
rect 11900 12093 11928 12124
rect 13081 12121 13093 12124
rect 13127 12152 13139 12155
rect 13262 12152 13268 12164
rect 13127 12124 13268 12152
rect 13127 12121 13139 12124
rect 13081 12115 13139 12121
rect 13262 12112 13268 12124
rect 13320 12112 13326 12164
rect 18509 12155 18567 12161
rect 18509 12121 18521 12155
rect 18555 12152 18567 12155
rect 18598 12152 18604 12164
rect 18555 12124 18604 12152
rect 18555 12121 18567 12124
rect 18509 12115 18567 12121
rect 18598 12112 18604 12124
rect 18656 12152 18662 12164
rect 18656 12124 19380 12152
rect 18656 12112 18662 12124
rect 19352 12096 19380 12124
rect 11885 12087 11943 12093
rect 11885 12084 11897 12087
rect 10836 12056 11897 12084
rect 10836 12044 10842 12056
rect 11885 12053 11897 12056
rect 11931 12053 11943 12087
rect 12342 12084 12348 12096
rect 12303 12056 12348 12084
rect 11885 12047 11943 12053
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 16206 12084 16212 12096
rect 16167 12056 16212 12084
rect 16206 12044 16212 12056
rect 16264 12044 16270 12096
rect 16574 12044 16580 12096
rect 16632 12084 16638 12096
rect 18874 12084 18880 12096
rect 16632 12056 18880 12084
rect 16632 12044 16638 12056
rect 18874 12044 18880 12056
rect 18932 12044 18938 12096
rect 19334 12084 19340 12096
rect 19295 12056 19340 12084
rect 19334 12044 19340 12056
rect 19392 12044 19398 12096
rect 20622 12084 20628 12096
rect 20583 12056 20628 12084
rect 20622 12044 20628 12056
rect 20680 12044 20686 12096
rect 23566 12044 23572 12096
rect 23624 12084 23630 12096
rect 24167 12087 24225 12093
rect 24167 12084 24179 12087
rect 23624 12056 24179 12084
rect 23624 12044 23630 12056
rect 24167 12053 24179 12056
rect 24213 12053 24225 12087
rect 24167 12047 24225 12053
rect 24762 12044 24768 12096
rect 24820 12084 24826 12096
rect 25179 12087 25237 12093
rect 25179 12084 25191 12087
rect 24820 12056 25191 12084
rect 24820 12044 24826 12056
rect 25179 12053 25191 12056
rect 25225 12053 25237 12087
rect 25179 12047 25237 12053
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 5905 11883 5963 11889
rect 5905 11849 5917 11883
rect 5951 11880 5963 11883
rect 6454 11880 6460 11892
rect 5951 11852 6460 11880
rect 5951 11849 5963 11852
rect 5905 11843 5963 11849
rect 6454 11840 6460 11852
rect 6512 11840 6518 11892
rect 6638 11880 6644 11892
rect 6599 11852 6644 11880
rect 6638 11840 6644 11852
rect 6696 11840 6702 11892
rect 7929 11883 7987 11889
rect 7929 11849 7941 11883
rect 7975 11880 7987 11883
rect 8018 11880 8024 11892
rect 7975 11852 8024 11880
rect 7975 11849 7987 11852
rect 7929 11843 7987 11849
rect 8018 11840 8024 11852
rect 8076 11840 8082 11892
rect 8757 11883 8815 11889
rect 8757 11849 8769 11883
rect 8803 11880 8815 11883
rect 10042 11880 10048 11892
rect 8803 11852 10048 11880
rect 8803 11849 8815 11852
rect 8757 11843 8815 11849
rect 10042 11840 10048 11852
rect 10100 11840 10106 11892
rect 12253 11883 12311 11889
rect 12253 11849 12265 11883
rect 12299 11880 12311 11883
rect 12342 11880 12348 11892
rect 12299 11852 12348 11880
rect 12299 11849 12311 11852
rect 12253 11843 12311 11849
rect 12342 11840 12348 11852
rect 12400 11840 12406 11892
rect 14277 11883 14335 11889
rect 14277 11849 14289 11883
rect 14323 11880 14335 11883
rect 14366 11880 14372 11892
rect 14323 11852 14372 11880
rect 14323 11849 14335 11852
rect 14277 11843 14335 11849
rect 14366 11840 14372 11852
rect 14424 11840 14430 11892
rect 16209 11883 16267 11889
rect 16209 11849 16221 11883
rect 16255 11880 16267 11883
rect 16482 11880 16488 11892
rect 16255 11852 16488 11880
rect 16255 11849 16267 11852
rect 16209 11843 16267 11849
rect 16482 11840 16488 11852
rect 16540 11840 16546 11892
rect 17865 11883 17923 11889
rect 17865 11849 17877 11883
rect 17911 11880 17923 11883
rect 17954 11880 17960 11892
rect 17911 11852 17960 11880
rect 17911 11849 17923 11852
rect 17865 11843 17923 11849
rect 17954 11840 17960 11852
rect 18012 11840 18018 11892
rect 19150 11840 19156 11892
rect 19208 11880 19214 11892
rect 20898 11880 20904 11892
rect 19208 11852 20904 11880
rect 19208 11840 19214 11852
rect 20898 11840 20904 11852
rect 20956 11840 20962 11892
rect 21358 11840 21364 11892
rect 21416 11880 21422 11892
rect 22189 11883 22247 11889
rect 22189 11880 22201 11883
rect 21416 11852 22201 11880
rect 21416 11840 21422 11852
rect 22189 11849 22201 11852
rect 22235 11880 22247 11883
rect 22557 11883 22615 11889
rect 22557 11880 22569 11883
rect 22235 11852 22569 11880
rect 22235 11849 22247 11852
rect 22189 11843 22247 11849
rect 22557 11849 22569 11852
rect 22603 11880 22615 11883
rect 22922 11880 22928 11892
rect 22603 11852 22928 11880
rect 22603 11849 22615 11852
rect 22557 11843 22615 11849
rect 22922 11840 22928 11852
rect 22980 11840 22986 11892
rect 24118 11840 24124 11892
rect 24176 11880 24182 11892
rect 24213 11883 24271 11889
rect 24213 11880 24225 11883
rect 24176 11852 24225 11880
rect 24176 11840 24182 11852
rect 24213 11849 24225 11852
rect 24259 11849 24271 11883
rect 24213 11843 24271 11849
rect 24489 11883 24547 11889
rect 24489 11849 24501 11883
rect 24535 11880 24547 11883
rect 24670 11880 24676 11892
rect 24535 11852 24676 11880
rect 24535 11849 24547 11852
rect 24489 11843 24547 11849
rect 24670 11840 24676 11852
rect 24728 11840 24734 11892
rect 6822 11772 6828 11824
rect 6880 11812 6886 11824
rect 9125 11815 9183 11821
rect 6880 11784 6960 11812
rect 6880 11772 6886 11784
rect 6932 11753 6960 11784
rect 9125 11781 9137 11815
rect 9171 11812 9183 11815
rect 9309 11815 9367 11821
rect 9309 11812 9321 11815
rect 9171 11784 9321 11812
rect 9171 11781 9183 11784
rect 9125 11775 9183 11781
rect 9309 11781 9321 11784
rect 9355 11812 9367 11815
rect 9398 11812 9404 11824
rect 9355 11784 9404 11812
rect 9355 11781 9367 11784
rect 9309 11775 9367 11781
rect 9398 11772 9404 11784
rect 9456 11772 9462 11824
rect 9490 11772 9496 11824
rect 9548 11772 9554 11824
rect 10137 11815 10195 11821
rect 10137 11781 10149 11815
rect 10183 11812 10195 11815
rect 13449 11815 13507 11821
rect 13449 11812 13461 11815
rect 10183 11784 11100 11812
rect 10183 11781 10195 11784
rect 10137 11775 10195 11781
rect 6917 11747 6975 11753
rect 6917 11713 6929 11747
rect 6963 11713 6975 11747
rect 7558 11744 7564 11756
rect 7519 11716 7564 11744
rect 6917 11707 6975 11713
rect 7558 11704 7564 11716
rect 7616 11704 7622 11756
rect 8846 11704 8852 11756
rect 8904 11744 8910 11756
rect 9508 11744 9536 11772
rect 10594 11744 10600 11756
rect 8904 11716 10600 11744
rect 8904 11704 8910 11716
rect 10594 11704 10600 11716
rect 10652 11704 10658 11756
rect 5721 11679 5779 11685
rect 5721 11645 5733 11679
rect 5767 11676 5779 11679
rect 6181 11679 6239 11685
rect 6181 11676 6193 11679
rect 5767 11648 6193 11676
rect 5767 11645 5779 11648
rect 5721 11639 5779 11645
rect 6181 11645 6193 11648
rect 6227 11676 6239 11679
rect 6730 11676 6736 11688
rect 6227 11648 6736 11676
rect 6227 11645 6239 11648
rect 6181 11639 6239 11645
rect 6730 11636 6736 11648
rect 6788 11636 6794 11688
rect 9214 11676 9220 11688
rect 9175 11648 9220 11676
rect 9214 11636 9220 11648
rect 9272 11636 9278 11688
rect 9493 11679 9551 11685
rect 9493 11645 9505 11679
rect 9539 11676 9551 11679
rect 10137 11679 10195 11685
rect 10137 11676 10149 11679
rect 9539 11648 10149 11676
rect 9539 11645 9551 11648
rect 9493 11639 9551 11645
rect 10137 11645 10149 11648
rect 10183 11645 10195 11679
rect 10778 11676 10784 11688
rect 10137 11639 10195 11645
rect 10244 11648 10784 11676
rect 6638 11568 6644 11620
rect 6696 11608 6702 11620
rect 7009 11611 7067 11617
rect 7009 11608 7021 11611
rect 6696 11580 7021 11608
rect 6696 11568 6702 11580
rect 7009 11577 7021 11580
rect 7055 11577 7067 11611
rect 7009 11571 7067 11577
rect 7190 11568 7196 11620
rect 7248 11608 7254 11620
rect 8389 11611 8447 11617
rect 8389 11608 8401 11611
rect 7248 11580 8401 11608
rect 7248 11568 7254 11580
rect 8389 11577 8401 11580
rect 8435 11608 8447 11611
rect 9508 11608 9536 11639
rect 9950 11608 9956 11620
rect 8435 11580 9536 11608
rect 9911 11580 9956 11608
rect 8435 11577 8447 11580
rect 8389 11571 8447 11577
rect 9950 11568 9956 11580
rect 10008 11568 10014 11620
rect 4338 11500 4344 11552
rect 4396 11540 4402 11552
rect 5534 11540 5540 11552
rect 4396 11512 5540 11540
rect 4396 11500 4402 11512
rect 5534 11500 5540 11512
rect 5592 11500 5598 11552
rect 9858 11500 9864 11552
rect 9916 11540 9922 11552
rect 10244 11549 10272 11648
rect 10778 11636 10784 11648
rect 10836 11636 10842 11688
rect 11072 11685 11100 11784
rect 12544 11784 13461 11812
rect 11330 11704 11336 11756
rect 11388 11744 11394 11756
rect 12544 11753 12572 11784
rect 13449 11781 13461 11784
rect 13495 11781 13507 11815
rect 13449 11775 13507 11781
rect 17034 11772 17040 11824
rect 17092 11812 17098 11824
rect 18693 11815 18751 11821
rect 18693 11812 18705 11815
rect 17092 11784 18705 11812
rect 17092 11772 17098 11784
rect 18693 11781 18705 11784
rect 18739 11812 18751 11815
rect 19242 11812 19248 11824
rect 18739 11784 19248 11812
rect 18739 11781 18751 11784
rect 18693 11775 18751 11781
rect 19242 11772 19248 11784
rect 19300 11772 19306 11824
rect 20070 11772 20076 11824
rect 20128 11812 20134 11824
rect 21821 11815 21879 11821
rect 21821 11812 21833 11815
rect 20128 11784 21833 11812
rect 20128 11772 20134 11784
rect 21821 11781 21833 11784
rect 21867 11781 21879 11815
rect 21821 11775 21879 11781
rect 12529 11747 12587 11753
rect 12529 11744 12541 11747
rect 11388 11716 12541 11744
rect 11388 11704 11394 11716
rect 12529 11713 12541 11716
rect 12575 11713 12587 11747
rect 13170 11744 13176 11756
rect 13131 11716 13176 11744
rect 12529 11707 12587 11713
rect 13170 11704 13176 11716
rect 13228 11704 13234 11756
rect 14182 11704 14188 11756
rect 14240 11744 14246 11756
rect 15289 11747 15347 11753
rect 15289 11744 15301 11747
rect 14240 11716 15301 11744
rect 14240 11704 14246 11716
rect 15289 11713 15301 11716
rect 15335 11744 15347 11747
rect 16853 11747 16911 11753
rect 16853 11744 16865 11747
rect 15335 11716 16865 11744
rect 15335 11713 15347 11716
rect 15289 11707 15347 11713
rect 16853 11713 16865 11716
rect 16899 11713 16911 11747
rect 16853 11707 16911 11713
rect 18141 11747 18199 11753
rect 18141 11713 18153 11747
rect 18187 11744 18199 11747
rect 19334 11744 19340 11756
rect 18187 11716 19340 11744
rect 18187 11713 18199 11716
rect 18141 11707 18199 11713
rect 19334 11704 19340 11716
rect 19392 11744 19398 11756
rect 19981 11747 20039 11753
rect 19981 11744 19993 11747
rect 19392 11716 19993 11744
rect 19392 11704 19398 11716
rect 19981 11713 19993 11716
rect 20027 11713 20039 11747
rect 19981 11707 20039 11713
rect 10873 11679 10931 11685
rect 10873 11645 10885 11679
rect 10919 11645 10931 11679
rect 10873 11639 10931 11645
rect 11057 11679 11115 11685
rect 11057 11645 11069 11679
rect 11103 11645 11115 11679
rect 11057 11639 11115 11645
rect 11517 11679 11575 11685
rect 11517 11645 11529 11679
rect 11563 11676 11575 11679
rect 11606 11676 11612 11688
rect 11563 11648 11612 11676
rect 11563 11645 11575 11648
rect 11517 11639 11575 11645
rect 10229 11543 10287 11549
rect 10229 11540 10241 11543
rect 9916 11512 10241 11540
rect 9916 11500 9922 11512
rect 10229 11509 10241 11512
rect 10275 11509 10287 11543
rect 10686 11540 10692 11552
rect 10647 11512 10692 11540
rect 10229 11503 10287 11509
rect 10686 11500 10692 11512
rect 10744 11540 10750 11552
rect 10888 11540 10916 11639
rect 11072 11608 11100 11639
rect 11606 11636 11612 11648
rect 11664 11636 11670 11688
rect 14090 11676 14096 11688
rect 14051 11648 14096 11676
rect 14090 11636 14096 11648
rect 14148 11676 14154 11688
rect 14645 11679 14703 11685
rect 14645 11676 14657 11679
rect 14148 11648 14657 11676
rect 14148 11636 14154 11648
rect 14645 11645 14657 11648
rect 14691 11645 14703 11679
rect 14645 11639 14703 11645
rect 16114 11636 16120 11688
rect 16172 11676 16178 11688
rect 17405 11679 17463 11685
rect 17405 11676 17417 11679
rect 16172 11648 17417 11676
rect 16172 11636 16178 11648
rect 17405 11645 17417 11648
rect 17451 11676 17463 11679
rect 17954 11676 17960 11688
rect 17451 11648 17960 11676
rect 17451 11645 17463 11648
rect 17405 11639 17463 11645
rect 17954 11636 17960 11648
rect 18012 11636 18018 11688
rect 22186 11636 22192 11688
rect 22244 11676 22250 11688
rect 22925 11679 22983 11685
rect 22925 11676 22937 11679
rect 22244 11648 22937 11676
rect 22244 11636 22250 11648
rect 22925 11645 22937 11648
rect 22971 11645 22983 11679
rect 22925 11639 22983 11645
rect 23290 11636 23296 11688
rect 23348 11676 23354 11688
rect 24004 11679 24062 11685
rect 24004 11676 24016 11679
rect 23348 11648 24016 11676
rect 23348 11636 23354 11648
rect 24004 11645 24016 11648
rect 24050 11676 24062 11679
rect 24118 11676 24124 11688
rect 24050 11648 24124 11676
rect 24050 11645 24062 11648
rect 24004 11639 24062 11645
rect 24118 11636 24124 11648
rect 24176 11676 24182 11688
rect 24765 11679 24823 11685
rect 24765 11676 24777 11679
rect 24176 11648 24777 11676
rect 24176 11636 24182 11648
rect 24765 11645 24777 11648
rect 24811 11645 24823 11679
rect 24765 11639 24823 11645
rect 25016 11679 25074 11685
rect 25016 11645 25028 11679
rect 25062 11676 25074 11679
rect 25062 11648 25544 11676
rect 25062 11645 25074 11648
rect 25016 11639 25074 11645
rect 12621 11611 12679 11617
rect 11072 11580 11928 11608
rect 11900 11549 11928 11580
rect 12621 11577 12633 11611
rect 12667 11577 12679 11611
rect 12621 11571 12679 11577
rect 15651 11611 15709 11617
rect 15651 11577 15663 11611
rect 15697 11608 15709 11611
rect 15746 11608 15752 11620
rect 15697 11580 15752 11608
rect 15697 11577 15709 11580
rect 15651 11571 15709 11577
rect 10744 11512 10916 11540
rect 11885 11543 11943 11549
rect 10744 11500 10750 11512
rect 11885 11509 11897 11543
rect 11931 11540 11943 11543
rect 12066 11540 12072 11552
rect 11931 11512 12072 11540
rect 11931 11509 11943 11512
rect 11885 11503 11943 11509
rect 12066 11500 12072 11512
rect 12124 11500 12130 11552
rect 12342 11500 12348 11552
rect 12400 11540 12406 11552
rect 12636 11540 12664 11571
rect 15746 11568 15752 11580
rect 15804 11568 15810 11620
rect 18233 11611 18291 11617
rect 18233 11577 18245 11611
rect 18279 11577 18291 11611
rect 18233 11571 18291 11577
rect 12400 11512 12664 11540
rect 12400 11500 12406 11512
rect 13814 11500 13820 11552
rect 13872 11540 13878 11552
rect 13872 11512 13917 11540
rect 13872 11500 13878 11512
rect 14642 11500 14648 11552
rect 14700 11540 14706 11552
rect 15105 11543 15163 11549
rect 15105 11540 15117 11543
rect 14700 11512 15117 11540
rect 14700 11500 14706 11512
rect 15105 11509 15117 11512
rect 15151 11509 15163 11543
rect 15105 11503 15163 11509
rect 17954 11500 17960 11552
rect 18012 11540 18018 11552
rect 18248 11540 18276 11571
rect 19518 11568 19524 11620
rect 19576 11608 19582 11620
rect 19705 11611 19763 11617
rect 19705 11608 19717 11611
rect 19576 11580 19717 11608
rect 19576 11568 19582 11580
rect 19705 11577 19717 11580
rect 19751 11577 19763 11611
rect 19705 11571 19763 11577
rect 19797 11611 19855 11617
rect 19797 11577 19809 11611
rect 19843 11577 19855 11611
rect 19797 11571 19855 11577
rect 19061 11543 19119 11549
rect 19061 11540 19073 11543
rect 18012 11512 19073 11540
rect 18012 11500 18018 11512
rect 19061 11509 19073 11512
rect 19107 11509 19119 11543
rect 19426 11540 19432 11552
rect 19339 11512 19432 11540
rect 19061 11503 19119 11509
rect 19426 11500 19432 11512
rect 19484 11540 19490 11552
rect 19812 11540 19840 11571
rect 20622 11568 20628 11620
rect 20680 11608 20686 11620
rect 21269 11611 21327 11617
rect 21269 11608 21281 11611
rect 20680 11580 21281 11608
rect 20680 11568 20686 11580
rect 21269 11577 21281 11580
rect 21315 11577 21327 11611
rect 21269 11571 21327 11577
rect 21358 11568 21364 11620
rect 21416 11608 21422 11620
rect 25516 11617 25544 11648
rect 25501 11611 25559 11617
rect 21416 11580 21461 11608
rect 21416 11568 21422 11580
rect 25501 11577 25513 11611
rect 25547 11608 25559 11611
rect 26142 11608 26148 11620
rect 25547 11580 26148 11608
rect 25547 11577 25559 11580
rect 25501 11571 25559 11577
rect 26142 11568 26148 11580
rect 26200 11568 26206 11620
rect 19484 11512 19840 11540
rect 19484 11500 19490 11512
rect 24946 11500 24952 11552
rect 25004 11540 25010 11552
rect 25087 11543 25145 11549
rect 25087 11540 25099 11543
rect 25004 11512 25099 11540
rect 25004 11500 25010 11512
rect 25087 11509 25099 11512
rect 25133 11509 25145 11543
rect 25866 11540 25872 11552
rect 25827 11512 25872 11540
rect 25087 11503 25145 11509
rect 25866 11500 25872 11512
rect 25924 11500 25930 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 6178 11336 6184 11348
rect 6139 11308 6184 11336
rect 6178 11296 6184 11308
rect 6236 11296 6242 11348
rect 7742 11336 7748 11348
rect 7703 11308 7748 11336
rect 7742 11296 7748 11308
rect 7800 11296 7806 11348
rect 12526 11336 12532 11348
rect 12487 11308 12532 11336
rect 12526 11296 12532 11308
rect 12584 11296 12590 11348
rect 13078 11336 13084 11348
rect 13039 11308 13084 11336
rect 13078 11296 13084 11308
rect 13136 11336 13142 11348
rect 13814 11336 13820 11348
rect 13136 11308 13820 11336
rect 13136 11296 13142 11308
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 13998 11336 14004 11348
rect 13959 11308 14004 11336
rect 13998 11296 14004 11308
rect 14056 11296 14062 11348
rect 16114 11296 16120 11348
rect 16172 11336 16178 11348
rect 16209 11339 16267 11345
rect 16209 11336 16221 11339
rect 16172 11308 16221 11336
rect 16172 11296 16178 11308
rect 16209 11305 16221 11308
rect 16255 11305 16267 11339
rect 16209 11299 16267 11305
rect 16577 11339 16635 11345
rect 16577 11305 16589 11339
rect 16623 11336 16635 11339
rect 16758 11336 16764 11348
rect 16623 11308 16764 11336
rect 16623 11305 16635 11308
rect 16577 11299 16635 11305
rect 16758 11296 16764 11308
rect 16816 11296 16822 11348
rect 17954 11336 17960 11348
rect 17915 11308 17960 11336
rect 17954 11296 17960 11308
rect 18012 11296 18018 11348
rect 18693 11339 18751 11345
rect 18693 11305 18705 11339
rect 18739 11336 18751 11339
rect 18782 11336 18788 11348
rect 18739 11308 18788 11336
rect 18739 11305 18751 11308
rect 18693 11299 18751 11305
rect 18782 11296 18788 11308
rect 18840 11296 18846 11348
rect 21174 11296 21180 11348
rect 21232 11336 21238 11348
rect 21913 11339 21971 11345
rect 21913 11336 21925 11339
rect 21232 11308 21925 11336
rect 21232 11296 21238 11308
rect 21913 11305 21925 11308
rect 21959 11305 21971 11339
rect 21913 11299 21971 11305
rect 22002 11296 22008 11348
rect 22060 11336 22066 11348
rect 24213 11339 24271 11345
rect 24213 11336 24225 11339
rect 22060 11308 24225 11336
rect 22060 11296 22066 11308
rect 24213 11305 24225 11308
rect 24259 11305 24271 11339
rect 24213 11299 24271 11305
rect 8021 11271 8079 11277
rect 8021 11237 8033 11271
rect 8067 11268 8079 11271
rect 8386 11268 8392 11280
rect 8067 11240 8392 11268
rect 8067 11237 8079 11240
rect 8021 11231 8079 11237
rect 8386 11228 8392 11240
rect 8444 11228 8450 11280
rect 9766 11228 9772 11280
rect 9824 11268 9830 11280
rect 11882 11268 11888 11280
rect 9824 11240 10364 11268
rect 9824 11228 9830 11240
rect 1464 11203 1522 11209
rect 1464 11169 1476 11203
rect 1510 11200 1522 11203
rect 1578 11200 1584 11212
rect 1510 11172 1584 11200
rect 1510 11169 1522 11172
rect 1464 11163 1522 11169
rect 1578 11160 1584 11172
rect 1636 11160 1642 11212
rect 6876 11203 6934 11209
rect 6876 11169 6888 11203
rect 6922 11200 6934 11203
rect 7098 11200 7104 11212
rect 6922 11172 7104 11200
rect 6922 11169 6934 11172
rect 6876 11163 6934 11169
rect 7098 11160 7104 11172
rect 7156 11160 7162 11212
rect 10042 11200 10048 11212
rect 10003 11172 10048 11200
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 10336 11209 10364 11240
rect 10888 11240 11888 11268
rect 10321 11203 10379 11209
rect 10321 11169 10333 11203
rect 10367 11169 10379 11203
rect 10321 11163 10379 11169
rect 10410 11160 10416 11212
rect 10468 11200 10474 11212
rect 10888 11209 10916 11240
rect 11882 11228 11888 11240
rect 11940 11228 11946 11280
rect 13722 11268 13728 11280
rect 13683 11240 13728 11268
rect 13722 11228 13728 11240
rect 13780 11228 13786 11280
rect 15651 11271 15709 11277
rect 15651 11237 15663 11271
rect 15697 11268 15709 11271
rect 15746 11268 15752 11280
rect 15697 11240 15752 11268
rect 15697 11237 15709 11240
rect 15651 11231 15709 11237
rect 15746 11228 15752 11240
rect 15804 11268 15810 11280
rect 17358 11271 17416 11277
rect 17358 11268 17370 11271
rect 15804 11240 17370 11268
rect 15804 11228 15810 11240
rect 17358 11237 17370 11240
rect 17404 11268 17416 11271
rect 17678 11268 17684 11280
rect 17404 11240 17684 11268
rect 17404 11237 17416 11240
rect 17358 11231 17416 11237
rect 17678 11228 17684 11240
rect 17736 11268 17742 11280
rect 18233 11271 18291 11277
rect 18233 11268 18245 11271
rect 17736 11240 18245 11268
rect 17736 11228 17742 11240
rect 18233 11237 18245 11240
rect 18279 11237 18291 11271
rect 18966 11268 18972 11280
rect 18927 11240 18972 11268
rect 18233 11231 18291 11237
rect 18966 11228 18972 11240
rect 19024 11228 19030 11280
rect 19242 11228 19248 11280
rect 19300 11268 19306 11280
rect 19521 11271 19579 11277
rect 19521 11268 19533 11271
rect 19300 11240 19533 11268
rect 19300 11228 19306 11240
rect 19521 11237 19533 11240
rect 19567 11268 19579 11271
rect 20165 11271 20223 11277
rect 20165 11268 20177 11271
rect 19567 11240 20177 11268
rect 19567 11237 19579 11240
rect 19521 11231 19579 11237
rect 20165 11237 20177 11240
rect 20211 11237 20223 11271
rect 22738 11268 22744 11280
rect 22699 11240 22744 11268
rect 20165 11231 20223 11237
rect 22738 11228 22744 11240
rect 22796 11228 22802 11280
rect 23290 11268 23296 11280
rect 23251 11240 23296 11268
rect 23290 11228 23296 11240
rect 23348 11228 23354 11280
rect 10873 11203 10931 11209
rect 10873 11200 10885 11203
rect 10468 11172 10885 11200
rect 10468 11160 10474 11172
rect 10873 11169 10885 11172
rect 10919 11169 10931 11203
rect 10873 11163 10931 11169
rect 11149 11203 11207 11209
rect 11149 11169 11161 11203
rect 11195 11169 11207 11203
rect 11149 11163 11207 11169
rect 14252 11203 14310 11209
rect 14252 11169 14264 11203
rect 14298 11200 14310 11203
rect 14550 11200 14556 11212
rect 14298 11172 14556 11200
rect 14298 11169 14310 11172
rect 14252 11163 14310 11169
rect 6963 11135 7021 11141
rect 6963 11101 6975 11135
rect 7009 11132 7021 11135
rect 7282 11132 7288 11144
rect 7009 11104 7288 11132
rect 7009 11101 7021 11104
rect 6963 11095 7021 11101
rect 7282 11092 7288 11104
rect 7340 11132 7346 11144
rect 7929 11135 7987 11141
rect 7929 11132 7941 11135
rect 7340 11104 7941 11132
rect 7340 11092 7346 11104
rect 7929 11101 7941 11104
rect 7975 11101 7987 11135
rect 8202 11132 8208 11144
rect 8163 11104 8208 11132
rect 7929 11095 7987 11101
rect 8202 11092 8208 11104
rect 8260 11092 8266 11144
rect 9214 11092 9220 11144
rect 9272 11132 9278 11144
rect 9309 11135 9367 11141
rect 9309 11132 9321 11135
rect 9272 11104 9321 11132
rect 9272 11092 9278 11104
rect 9309 11101 9321 11104
rect 9355 11132 9367 11135
rect 10428 11132 10456 11160
rect 9355 11104 10456 11132
rect 9355 11101 9367 11104
rect 9309 11095 9367 11101
rect 11164 11076 11192 11163
rect 14550 11160 14556 11172
rect 14608 11160 14614 11212
rect 17037 11203 17095 11209
rect 17037 11169 17049 11203
rect 17083 11200 17095 11203
rect 17586 11200 17592 11212
rect 17083 11172 17592 11200
rect 17083 11169 17095 11172
rect 17037 11163 17095 11169
rect 17586 11160 17592 11172
rect 17644 11160 17650 11212
rect 21082 11200 21088 11212
rect 21043 11172 21088 11200
rect 21082 11160 21088 11172
rect 21140 11160 21146 11212
rect 21266 11160 21272 11212
rect 21324 11200 21330 11212
rect 21361 11203 21419 11209
rect 21361 11200 21373 11203
rect 21324 11172 21373 11200
rect 21324 11160 21330 11172
rect 21361 11169 21373 11172
rect 21407 11169 21419 11203
rect 24210 11200 24216 11212
rect 21361 11163 21419 11169
rect 23446 11172 24216 11200
rect 11333 11135 11391 11141
rect 11333 11101 11345 11135
rect 11379 11132 11391 11135
rect 11790 11132 11796 11144
rect 11379 11104 11796 11132
rect 11379 11101 11391 11104
rect 11333 11095 11391 11101
rect 11790 11092 11796 11104
rect 11848 11132 11854 11144
rect 12161 11135 12219 11141
rect 12161 11132 12173 11135
rect 11848 11104 12173 11132
rect 11848 11092 11854 11104
rect 12161 11101 12173 11104
rect 12207 11101 12219 11135
rect 15286 11132 15292 11144
rect 15247 11104 15292 11132
rect 12161 11095 12219 11101
rect 15286 11092 15292 11104
rect 15344 11092 15350 11144
rect 18874 11132 18880 11144
rect 18787 11104 18880 11132
rect 18874 11092 18880 11104
rect 18932 11132 18938 11144
rect 20070 11132 20076 11144
rect 18932 11104 20076 11132
rect 18932 11092 18938 11104
rect 20070 11092 20076 11104
rect 20128 11092 20134 11144
rect 21100 11132 21128 11160
rect 21637 11135 21695 11141
rect 21100 11104 21588 11132
rect 6730 11024 6736 11076
rect 6788 11064 6794 11076
rect 11146 11064 11152 11076
rect 6788 11036 11152 11064
rect 6788 11024 6794 11036
rect 11146 11024 11152 11036
rect 11204 11064 11210 11076
rect 11422 11064 11428 11076
rect 11204 11036 11428 11064
rect 11204 11024 11210 11036
rect 11422 11024 11428 11036
rect 11480 11024 11486 11076
rect 18046 11024 18052 11076
rect 18104 11064 18110 11076
rect 20625 11067 20683 11073
rect 20625 11064 20637 11067
rect 18104 11036 20637 11064
rect 18104 11024 18110 11036
rect 20625 11033 20637 11036
rect 20671 11064 20683 11067
rect 21358 11064 21364 11076
rect 20671 11036 21364 11064
rect 20671 11033 20683 11036
rect 20625 11027 20683 11033
rect 21358 11024 21364 11036
rect 21416 11024 21422 11076
rect 21560 11064 21588 11104
rect 21637 11101 21649 11135
rect 21683 11132 21695 11135
rect 21818 11132 21824 11144
rect 21683 11104 21824 11132
rect 21683 11101 21695 11104
rect 21637 11095 21695 11101
rect 21818 11092 21824 11104
rect 21876 11092 21882 11144
rect 22649 11135 22707 11141
rect 22649 11101 22661 11135
rect 22695 11132 22707 11135
rect 22922 11132 22928 11144
rect 22695 11104 22928 11132
rect 22695 11101 22707 11104
rect 22649 11095 22707 11101
rect 22922 11092 22928 11104
rect 22980 11092 22986 11144
rect 23446 11064 23474 11172
rect 24210 11160 24216 11172
rect 24268 11160 24274 11212
rect 24581 11203 24639 11209
rect 24581 11169 24593 11203
rect 24627 11169 24639 11203
rect 24581 11163 24639 11169
rect 24596 11132 24624 11163
rect 24670 11132 24676 11144
rect 21560 11036 23474 11064
rect 23584 11104 24676 11132
rect 1535 10999 1593 11005
rect 1535 10965 1547 10999
rect 1581 10996 1593 10999
rect 5994 10996 6000 11008
rect 1581 10968 6000 10996
rect 1581 10965 1593 10968
rect 1535 10959 1593 10965
rect 5994 10956 6000 10968
rect 6052 10956 6058 11008
rect 7374 10996 7380 11008
rect 7335 10968 7380 10996
rect 7374 10956 7380 10968
rect 7432 10956 7438 11008
rect 8846 10996 8852 11008
rect 8807 10968 8852 10996
rect 8846 10956 8852 10968
rect 8904 10956 8910 11008
rect 9122 10956 9128 11008
rect 9180 10996 9186 11008
rect 9766 10996 9772 11008
rect 9180 10968 9772 10996
rect 9180 10956 9186 10968
rect 9766 10956 9772 10968
rect 9824 10956 9830 11008
rect 14323 10999 14381 11005
rect 14323 10965 14335 10999
rect 14369 10996 14381 10999
rect 14734 10996 14740 11008
rect 14369 10968 14740 10996
rect 14369 10965 14381 10968
rect 14323 10959 14381 10965
rect 14734 10956 14740 10968
rect 14792 10956 14798 11008
rect 14826 10956 14832 11008
rect 14884 10996 14890 11008
rect 15013 10999 15071 11005
rect 15013 10996 15025 10999
rect 14884 10968 15025 10996
rect 14884 10956 14890 10968
rect 15013 10965 15025 10968
rect 15059 10965 15071 10999
rect 15013 10959 15071 10965
rect 18690 10956 18696 11008
rect 18748 10996 18754 11008
rect 19518 10996 19524 11008
rect 18748 10968 19524 10996
rect 18748 10956 18754 10968
rect 19518 10956 19524 10968
rect 19576 10996 19582 11008
rect 19797 10999 19855 11005
rect 19797 10996 19809 10999
rect 19576 10968 19809 10996
rect 19576 10956 19582 10968
rect 19797 10965 19809 10968
rect 19843 10965 19855 10999
rect 19797 10959 19855 10965
rect 20530 10956 20536 11008
rect 20588 10996 20594 11008
rect 23584 10996 23612 11104
rect 24670 11092 24676 11104
rect 24728 11092 24734 11144
rect 20588 10968 23612 10996
rect 23753 10999 23811 11005
rect 20588 10956 20594 10968
rect 23753 10965 23765 10999
rect 23799 10996 23811 10999
rect 23842 10996 23848 11008
rect 23799 10968 23848 10996
rect 23799 10965 23811 10968
rect 23753 10959 23811 10965
rect 23842 10956 23848 10968
rect 23900 10956 23906 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1578 10792 1584 10804
rect 1539 10764 1584 10792
rect 1578 10752 1584 10764
rect 1636 10752 1642 10804
rect 6086 10752 6092 10804
rect 6144 10792 6150 10804
rect 8757 10795 8815 10801
rect 8757 10792 8769 10795
rect 6144 10764 8769 10792
rect 6144 10752 6150 10764
rect 8757 10761 8769 10764
rect 8803 10792 8815 10795
rect 9122 10792 9128 10804
rect 8803 10764 9128 10792
rect 8803 10761 8815 10764
rect 8757 10755 8815 10761
rect 9122 10752 9128 10764
rect 9180 10752 9186 10804
rect 9217 10795 9275 10801
rect 9217 10761 9229 10795
rect 9263 10792 9275 10795
rect 9674 10792 9680 10804
rect 9263 10764 9680 10792
rect 9263 10761 9275 10764
rect 9217 10755 9275 10761
rect 9674 10752 9680 10764
rect 9732 10792 9738 10804
rect 10134 10792 10140 10804
rect 9732 10764 10140 10792
rect 9732 10752 9738 10764
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 11422 10792 11428 10804
rect 11383 10764 11428 10792
rect 11422 10752 11428 10764
rect 11480 10752 11486 10804
rect 11790 10792 11796 10804
rect 11751 10764 11796 10792
rect 11790 10752 11796 10764
rect 11848 10752 11854 10804
rect 12253 10795 12311 10801
rect 12253 10761 12265 10795
rect 12299 10792 12311 10795
rect 12526 10792 12532 10804
rect 12299 10764 12532 10792
rect 12299 10761 12311 10764
rect 12253 10755 12311 10761
rect 12526 10752 12532 10764
rect 12584 10792 12590 10804
rect 15197 10795 15255 10801
rect 15197 10792 15209 10795
rect 12584 10764 15209 10792
rect 12584 10752 12590 10764
rect 15197 10761 15209 10764
rect 15243 10792 15255 10795
rect 15746 10792 15752 10804
rect 15243 10764 15752 10792
rect 15243 10761 15255 10764
rect 15197 10755 15255 10761
rect 15746 10752 15752 10764
rect 15804 10752 15810 10804
rect 16991 10795 17049 10801
rect 16991 10761 17003 10795
rect 17037 10792 17049 10795
rect 18690 10792 18696 10804
rect 17037 10764 18696 10792
rect 17037 10761 17049 10764
rect 16991 10755 17049 10761
rect 18690 10752 18696 10764
rect 18748 10752 18754 10804
rect 18966 10792 18972 10804
rect 18927 10764 18972 10792
rect 18966 10752 18972 10764
rect 19024 10792 19030 10804
rect 19245 10795 19303 10801
rect 19245 10792 19257 10795
rect 19024 10764 19257 10792
rect 19024 10752 19030 10764
rect 19245 10761 19257 10764
rect 19291 10761 19303 10795
rect 19245 10755 19303 10761
rect 19935 10795 19993 10801
rect 19935 10761 19947 10795
rect 19981 10792 19993 10795
rect 20622 10792 20628 10804
rect 19981 10764 20628 10792
rect 19981 10761 19993 10764
rect 19935 10755 19993 10761
rect 20622 10752 20628 10764
rect 20680 10752 20686 10804
rect 20717 10795 20775 10801
rect 20717 10761 20729 10795
rect 20763 10792 20775 10795
rect 21266 10792 21272 10804
rect 20763 10764 21272 10792
rect 20763 10761 20775 10764
rect 20717 10755 20775 10761
rect 21266 10752 21272 10764
rect 21324 10752 21330 10804
rect 22097 10795 22155 10801
rect 22097 10761 22109 10795
rect 22143 10792 22155 10795
rect 22649 10795 22707 10801
rect 22649 10792 22661 10795
rect 22143 10764 22661 10792
rect 22143 10761 22155 10764
rect 22097 10755 22155 10761
rect 22649 10761 22661 10764
rect 22695 10792 22707 10795
rect 22738 10792 22744 10804
rect 22695 10764 22744 10792
rect 22695 10761 22707 10764
rect 22649 10755 22707 10761
rect 22738 10752 22744 10764
rect 22796 10752 22802 10804
rect 24670 10792 24676 10804
rect 24631 10764 24676 10792
rect 24670 10752 24676 10764
rect 24728 10752 24734 10804
rect 5905 10727 5963 10733
rect 5905 10693 5917 10727
rect 5951 10724 5963 10727
rect 9306 10724 9312 10736
rect 5951 10696 9312 10724
rect 5951 10693 5963 10696
rect 5905 10687 5963 10693
rect 9306 10684 9312 10696
rect 9364 10684 9370 10736
rect 9950 10684 9956 10736
rect 10008 10724 10014 10736
rect 13817 10727 13875 10733
rect 13817 10724 13829 10727
rect 10008 10696 13829 10724
rect 10008 10684 10014 10696
rect 13817 10693 13829 10696
rect 13863 10693 13875 10727
rect 13817 10687 13875 10693
rect 6273 10659 6331 10665
rect 6273 10625 6285 10659
rect 6319 10656 6331 10659
rect 7190 10656 7196 10668
rect 6319 10628 7196 10656
rect 6319 10625 6331 10628
rect 6273 10619 6331 10625
rect 5721 10591 5779 10597
rect 5721 10557 5733 10591
rect 5767 10588 5779 10591
rect 6288 10588 6316 10619
rect 7190 10616 7196 10628
rect 7248 10616 7254 10668
rect 8202 10616 8208 10668
rect 8260 10656 8266 10668
rect 12529 10659 12587 10665
rect 12529 10656 12541 10659
rect 8260 10628 12541 10656
rect 8260 10616 8266 10628
rect 12529 10625 12541 10628
rect 12575 10656 12587 10659
rect 12802 10656 12808 10668
rect 12575 10628 12808 10656
rect 12575 10625 12587 10628
rect 12529 10619 12587 10625
rect 12802 10616 12808 10628
rect 12860 10616 12866 10668
rect 13170 10656 13176 10668
rect 13131 10628 13176 10656
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 5767 10560 6316 10588
rect 5767 10557 5779 10560
rect 5721 10551 5779 10557
rect 7374 10548 7380 10600
rect 7432 10588 7438 10600
rect 7561 10591 7619 10597
rect 7561 10588 7573 10591
rect 7432 10560 7573 10588
rect 7432 10548 7438 10560
rect 7561 10557 7573 10560
rect 7607 10588 7619 10591
rect 9585 10591 9643 10597
rect 7607 10560 9260 10588
rect 7607 10557 7619 10560
rect 7561 10551 7619 10557
rect 7469 10523 7527 10529
rect 7469 10489 7481 10523
rect 7515 10520 7527 10523
rect 7923 10523 7981 10529
rect 7923 10520 7935 10523
rect 7515 10492 7935 10520
rect 7515 10489 7527 10492
rect 7469 10483 7527 10489
rect 7923 10489 7935 10492
rect 7969 10520 7981 10523
rect 8018 10520 8024 10532
rect 7969 10492 8024 10520
rect 7969 10489 7981 10492
rect 7923 10483 7981 10489
rect 8018 10480 8024 10492
rect 8076 10480 8082 10532
rect 7098 10452 7104 10464
rect 7059 10424 7104 10452
rect 7098 10412 7104 10424
rect 7156 10412 7162 10464
rect 8478 10452 8484 10464
rect 8439 10424 8484 10452
rect 8478 10412 8484 10424
rect 8536 10412 8542 10464
rect 9232 10452 9260 10560
rect 9585 10557 9597 10591
rect 9631 10557 9643 10591
rect 9766 10588 9772 10600
rect 9727 10560 9772 10588
rect 9585 10551 9643 10557
rect 9306 10480 9312 10532
rect 9364 10520 9370 10532
rect 9600 10520 9628 10551
rect 9766 10548 9772 10560
rect 9824 10548 9830 10600
rect 9950 10548 9956 10600
rect 10008 10588 10014 10600
rect 10321 10591 10379 10597
rect 10321 10588 10333 10591
rect 10008 10560 10333 10588
rect 10008 10548 10014 10560
rect 10321 10557 10333 10560
rect 10367 10588 10379 10591
rect 10410 10588 10416 10600
rect 10367 10560 10416 10588
rect 10367 10557 10379 10560
rect 10321 10551 10379 10557
rect 10410 10548 10416 10560
rect 10468 10548 10474 10600
rect 10505 10591 10563 10597
rect 10505 10557 10517 10591
rect 10551 10557 10563 10591
rect 13832 10588 13860 10687
rect 15286 10684 15292 10736
rect 15344 10724 15350 10736
rect 16669 10727 16727 10733
rect 16669 10724 16681 10727
rect 15344 10696 16681 10724
rect 15344 10684 15350 10696
rect 16669 10693 16681 10696
rect 16715 10693 16727 10727
rect 17678 10724 17684 10736
rect 17639 10696 17684 10724
rect 16669 10687 16727 10693
rect 17678 10684 17684 10696
rect 17736 10684 17742 10736
rect 19705 10727 19763 10733
rect 19705 10693 19717 10727
rect 19751 10724 19763 10727
rect 20070 10724 20076 10736
rect 19751 10696 20076 10724
rect 19751 10693 19763 10696
rect 19705 10687 19763 10693
rect 20070 10684 20076 10696
rect 20128 10684 20134 10736
rect 20349 10727 20407 10733
rect 20349 10693 20361 10727
rect 20395 10724 20407 10727
rect 23014 10724 23020 10736
rect 20395 10696 23020 10724
rect 20395 10693 20407 10696
rect 20349 10687 20407 10693
rect 16025 10659 16083 10665
rect 16025 10625 16037 10659
rect 16071 10656 16083 10659
rect 16758 10656 16764 10668
rect 16071 10628 16764 10656
rect 16071 10625 16083 10628
rect 16025 10619 16083 10625
rect 16758 10616 16764 10628
rect 16816 10616 16822 10668
rect 18049 10659 18107 10665
rect 18049 10625 18061 10659
rect 18095 10656 18107 10659
rect 18782 10656 18788 10668
rect 18095 10628 18788 10656
rect 18095 10625 18107 10628
rect 18049 10619 18107 10625
rect 18782 10616 18788 10628
rect 18840 10616 18846 10668
rect 14001 10591 14059 10597
rect 14001 10588 14013 10591
rect 13832 10560 14013 10588
rect 10505 10551 10563 10557
rect 14001 10557 14013 10560
rect 14047 10557 14059 10591
rect 14001 10551 14059 10557
rect 10042 10520 10048 10532
rect 9364 10492 10048 10520
rect 9364 10480 9370 10492
rect 10042 10480 10048 10492
rect 10100 10480 10106 10532
rect 10134 10480 10140 10532
rect 10192 10520 10198 10532
rect 10520 10520 10548 10551
rect 16666 10548 16672 10600
rect 16724 10588 16730 10600
rect 16888 10591 16946 10597
rect 16888 10588 16900 10591
rect 16724 10560 16900 10588
rect 16724 10548 16730 10560
rect 16888 10557 16900 10560
rect 16934 10588 16946 10591
rect 17313 10591 17371 10597
rect 17313 10588 17325 10591
rect 16934 10560 17325 10588
rect 16934 10557 16946 10560
rect 16888 10551 16946 10557
rect 17313 10557 17325 10560
rect 17359 10557 17371 10591
rect 17313 10551 17371 10557
rect 19864 10591 19922 10597
rect 19864 10557 19876 10591
rect 19910 10588 19922 10591
rect 20364 10588 20392 10687
rect 23014 10684 23020 10696
rect 23072 10684 23078 10736
rect 21174 10656 21180 10668
rect 21135 10628 21180 10656
rect 21174 10616 21180 10628
rect 21232 10616 21238 10668
rect 23753 10659 23811 10665
rect 23753 10625 23765 10659
rect 23799 10656 23811 10659
rect 23842 10656 23848 10668
rect 23799 10628 23848 10656
rect 23799 10625 23811 10628
rect 23753 10619 23811 10625
rect 23842 10616 23848 10628
rect 23900 10616 23906 10668
rect 24026 10656 24032 10668
rect 23987 10628 24032 10656
rect 24026 10616 24032 10628
rect 24084 10616 24090 10668
rect 19910 10560 20392 10588
rect 19910 10557 19922 10560
rect 19864 10551 19922 10557
rect 20622 10548 20628 10600
rect 20680 10588 20686 10600
rect 22922 10588 22928 10600
rect 20680 10560 22928 10588
rect 20680 10548 20686 10560
rect 22922 10548 22928 10560
rect 22980 10548 22986 10600
rect 24854 10548 24860 10600
rect 24912 10588 24918 10600
rect 25260 10591 25318 10597
rect 25260 10588 25272 10591
rect 24912 10560 25272 10588
rect 24912 10548 24918 10560
rect 25260 10557 25272 10560
rect 25306 10588 25318 10591
rect 25685 10591 25743 10597
rect 25685 10588 25697 10591
rect 25306 10560 25697 10588
rect 25306 10557 25318 10560
rect 25260 10551 25318 10557
rect 25685 10557 25697 10560
rect 25731 10557 25743 10591
rect 25685 10551 25743 10557
rect 10192 10492 10548 10520
rect 10192 10480 10198 10492
rect 12618 10480 12624 10532
rect 12676 10520 12682 10532
rect 12986 10520 12992 10532
rect 12676 10492 12992 10520
rect 12676 10480 12682 10492
rect 12986 10480 12992 10492
rect 13044 10480 13050 10532
rect 13170 10480 13176 10532
rect 13228 10520 13234 10532
rect 14826 10520 14832 10532
rect 13228 10492 14832 10520
rect 13228 10480 13234 10492
rect 14826 10480 14832 10492
rect 14884 10520 14890 10532
rect 15381 10523 15439 10529
rect 15381 10520 15393 10523
rect 14884 10492 15393 10520
rect 14884 10480 14890 10492
rect 15381 10489 15393 10492
rect 15427 10489 15439 10523
rect 15381 10483 15439 10489
rect 15473 10523 15531 10529
rect 15473 10489 15485 10523
rect 15519 10520 15531 10523
rect 15519 10492 16436 10520
rect 15519 10489 15531 10492
rect 15473 10483 15531 10489
rect 16408 10464 16436 10492
rect 17678 10480 17684 10532
rect 17736 10520 17742 10532
rect 18370 10523 18428 10529
rect 18370 10520 18382 10523
rect 17736 10492 18382 10520
rect 17736 10480 17742 10492
rect 18370 10489 18382 10492
rect 18416 10520 18428 10523
rect 20993 10523 21051 10529
rect 20993 10520 21005 10523
rect 18416 10492 21005 10520
rect 18416 10489 18428 10492
rect 18370 10483 18428 10489
rect 20993 10489 21005 10492
rect 21039 10520 21051 10523
rect 21450 10520 21456 10532
rect 21039 10492 21456 10520
rect 21039 10489 21051 10492
rect 20993 10483 21051 10489
rect 21450 10480 21456 10492
rect 21508 10529 21514 10532
rect 21508 10523 21556 10529
rect 21508 10489 21510 10523
rect 21544 10489 21556 10523
rect 21508 10483 21556 10489
rect 21508 10480 21514 10483
rect 23106 10480 23112 10532
rect 23164 10520 23170 10532
rect 23385 10523 23443 10529
rect 23385 10520 23397 10523
rect 23164 10492 23397 10520
rect 23164 10480 23170 10492
rect 23385 10489 23397 10492
rect 23431 10520 23443 10523
rect 23845 10523 23903 10529
rect 23431 10492 23679 10520
rect 23431 10489 23443 10492
rect 23385 10483 23443 10489
rect 9401 10455 9459 10461
rect 9401 10452 9413 10455
rect 9232 10424 9413 10452
rect 9401 10421 9413 10424
rect 9447 10421 9459 10455
rect 9401 10415 9459 10421
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 11057 10455 11115 10461
rect 11057 10452 11069 10455
rect 9824 10424 11069 10452
rect 9824 10412 9830 10424
rect 11057 10421 11069 10424
rect 11103 10421 11115 10455
rect 14182 10452 14188 10464
rect 14143 10424 14188 10452
rect 11057 10415 11115 10421
rect 14182 10412 14188 10424
rect 14240 10412 14246 10464
rect 14550 10452 14556 10464
rect 14511 10424 14556 10452
rect 14550 10412 14556 10424
rect 14608 10412 14614 10464
rect 16390 10452 16396 10464
rect 16351 10424 16396 10452
rect 16390 10412 16396 10424
rect 16448 10412 16454 10464
rect 23651 10452 23679 10492
rect 23845 10489 23857 10523
rect 23891 10489 23903 10523
rect 23845 10483 23903 10489
rect 23860 10452 23888 10483
rect 23934 10480 23940 10532
rect 23992 10520 23998 10532
rect 24670 10520 24676 10532
rect 23992 10492 24676 10520
rect 23992 10480 23998 10492
rect 24670 10480 24676 10492
rect 24728 10480 24734 10532
rect 23651 10424 23888 10452
rect 25363 10455 25421 10461
rect 25363 10421 25375 10455
rect 25409 10452 25421 10455
rect 25590 10452 25596 10464
rect 25409 10424 25596 10452
rect 25409 10421 25421 10424
rect 25363 10415 25421 10421
rect 25590 10412 25596 10424
rect 25648 10412 25654 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 7282 10248 7288 10260
rect 7243 10220 7288 10248
rect 7282 10208 7288 10220
rect 7340 10208 7346 10260
rect 9033 10251 9091 10257
rect 9033 10217 9045 10251
rect 9079 10248 9091 10251
rect 9306 10248 9312 10260
rect 9079 10220 9312 10248
rect 9079 10217 9091 10220
rect 9033 10211 9091 10217
rect 9306 10208 9312 10220
rect 9364 10208 9370 10260
rect 9401 10251 9459 10257
rect 9401 10217 9413 10251
rect 9447 10248 9459 10251
rect 9950 10248 9956 10260
rect 9447 10220 9956 10248
rect 9447 10217 9459 10220
rect 9401 10211 9459 10217
rect 9950 10208 9956 10220
rect 10008 10208 10014 10260
rect 10042 10208 10048 10260
rect 10100 10248 10106 10260
rect 10597 10251 10655 10257
rect 10597 10248 10609 10251
rect 10100 10220 10609 10248
rect 10100 10208 10106 10220
rect 10597 10217 10609 10220
rect 10643 10217 10655 10251
rect 10597 10211 10655 10217
rect 12529 10251 12587 10257
rect 12529 10217 12541 10251
rect 12575 10248 12587 10251
rect 12618 10248 12624 10260
rect 12575 10220 12624 10248
rect 12575 10217 12587 10220
rect 12529 10211 12587 10217
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 12802 10248 12808 10260
rect 12763 10220 12808 10248
rect 12802 10208 12808 10220
rect 12860 10208 12866 10260
rect 15562 10248 15568 10260
rect 15523 10220 15568 10248
rect 15562 10208 15568 10220
rect 15620 10208 15626 10260
rect 17405 10251 17463 10257
rect 17405 10217 17417 10251
rect 17451 10248 17463 10251
rect 17586 10248 17592 10260
rect 17451 10220 17592 10248
rect 17451 10217 17463 10220
rect 17405 10211 17463 10217
rect 17586 10208 17592 10220
rect 17644 10208 17650 10260
rect 19426 10248 19432 10260
rect 18248 10220 19432 10248
rect 7558 10180 7564 10192
rect 7519 10152 7564 10180
rect 7558 10140 7564 10152
rect 7616 10140 7622 10192
rect 8113 10183 8171 10189
rect 8113 10149 8125 10183
rect 8159 10180 8171 10183
rect 8202 10180 8208 10192
rect 8159 10152 8208 10180
rect 8159 10149 8171 10152
rect 8113 10143 8171 10149
rect 8202 10140 8208 10152
rect 8260 10140 8266 10192
rect 14182 10140 14188 10192
rect 14240 10180 14246 10192
rect 14826 10180 14832 10192
rect 14240 10152 14832 10180
rect 14240 10140 14246 10152
rect 14826 10140 14832 10152
rect 14884 10180 14890 10192
rect 17218 10180 17224 10192
rect 14884 10152 17224 10180
rect 14884 10140 14890 10152
rect 106 10072 112 10124
rect 164 10112 170 10124
rect 4798 10112 4804 10124
rect 4856 10121 4862 10124
rect 4856 10115 4894 10121
rect 164 10084 4804 10112
rect 164 10072 170 10084
rect 4798 10072 4804 10084
rect 4882 10081 4894 10115
rect 4856 10075 4894 10081
rect 4856 10072 4862 10075
rect 5534 10072 5540 10124
rect 5592 10112 5598 10124
rect 5813 10115 5871 10121
rect 5813 10112 5825 10115
rect 5592 10084 5825 10112
rect 5592 10072 5598 10084
rect 5813 10081 5825 10084
rect 5859 10081 5871 10115
rect 5813 10075 5871 10081
rect 6365 10115 6423 10121
rect 6365 10081 6377 10115
rect 6411 10112 6423 10115
rect 6546 10112 6552 10124
rect 6411 10084 6552 10112
rect 6411 10081 6423 10084
rect 6365 10075 6423 10081
rect 6546 10072 6552 10084
rect 6604 10072 6610 10124
rect 10134 10112 10140 10124
rect 10095 10084 10140 10112
rect 10134 10072 10140 10084
rect 10192 10112 10198 10124
rect 10686 10112 10692 10124
rect 10192 10084 10692 10112
rect 10192 10072 10198 10084
rect 10686 10072 10692 10084
rect 10744 10072 10750 10124
rect 11790 10112 11796 10124
rect 11751 10084 11796 10112
rect 11790 10072 11796 10084
rect 11848 10072 11854 10124
rect 13906 10112 13912 10124
rect 13867 10084 13912 10112
rect 13906 10072 13912 10084
rect 13964 10072 13970 10124
rect 14093 10115 14151 10121
rect 14093 10081 14105 10115
rect 14139 10112 14151 10115
rect 14274 10112 14280 10124
rect 14139 10084 14280 10112
rect 14139 10081 14151 10084
rect 14093 10075 14151 10081
rect 14274 10072 14280 10084
rect 14332 10072 14338 10124
rect 15470 10112 15476 10124
rect 15431 10084 15476 10112
rect 15470 10072 15476 10084
rect 15528 10072 15534 10124
rect 15856 10121 15884 10152
rect 17218 10140 17224 10152
rect 17276 10140 17282 10192
rect 18138 10140 18144 10192
rect 18196 10180 18202 10192
rect 18248 10189 18276 10220
rect 19426 10208 19432 10220
rect 19484 10208 19490 10260
rect 21082 10248 21088 10260
rect 21043 10220 21088 10248
rect 21082 10208 21088 10220
rect 21140 10208 21146 10260
rect 22465 10251 22523 10257
rect 22465 10217 22477 10251
rect 22511 10248 22523 10251
rect 23290 10248 23296 10260
rect 22511 10220 23296 10248
rect 22511 10217 22523 10220
rect 22465 10211 22523 10217
rect 23290 10208 23296 10220
rect 23348 10248 23354 10260
rect 23348 10220 23520 10248
rect 23348 10208 23354 10220
rect 18233 10183 18291 10189
rect 18233 10180 18245 10183
rect 18196 10152 18245 10180
rect 18196 10140 18202 10152
rect 18233 10149 18245 10152
rect 18279 10149 18291 10183
rect 18233 10143 18291 10149
rect 18785 10183 18843 10189
rect 18785 10149 18797 10183
rect 18831 10180 18843 10183
rect 18874 10180 18880 10192
rect 18831 10152 18880 10180
rect 18831 10149 18843 10152
rect 18785 10143 18843 10149
rect 18874 10140 18880 10152
rect 18932 10140 18938 10192
rect 21450 10140 21456 10192
rect 21508 10180 21514 10192
rect 23492 10189 23520 10220
rect 24210 10208 24216 10260
rect 24268 10248 24274 10260
rect 24305 10251 24363 10257
rect 24305 10248 24317 10251
rect 24268 10220 24317 10248
rect 24268 10208 24274 10220
rect 24305 10217 24317 10220
rect 24351 10217 24363 10251
rect 24305 10211 24363 10217
rect 21866 10183 21924 10189
rect 21866 10180 21878 10183
rect 21508 10152 21878 10180
rect 21508 10140 21514 10152
rect 21866 10149 21878 10152
rect 21912 10149 21924 10183
rect 21866 10143 21924 10149
rect 23477 10183 23535 10189
rect 23477 10149 23489 10183
rect 23523 10149 23535 10183
rect 23477 10143 23535 10149
rect 24029 10183 24087 10189
rect 24029 10149 24041 10183
rect 24075 10180 24087 10183
rect 24118 10180 24124 10192
rect 24075 10152 24124 10180
rect 24075 10149 24087 10152
rect 24029 10143 24087 10149
rect 24118 10140 24124 10152
rect 24176 10140 24182 10192
rect 24946 10180 24952 10192
rect 24228 10152 24952 10180
rect 24228 10124 24256 10152
rect 24946 10140 24952 10152
rect 25004 10140 25010 10192
rect 25041 10183 25099 10189
rect 25041 10149 25053 10183
rect 25087 10180 25099 10183
rect 25222 10180 25228 10192
rect 25087 10152 25228 10180
rect 25087 10149 25099 10152
rect 25041 10143 25099 10149
rect 25222 10140 25228 10152
rect 25280 10140 25286 10192
rect 15841 10115 15899 10121
rect 15841 10081 15853 10115
rect 15887 10081 15899 10115
rect 16850 10112 16856 10124
rect 16811 10084 16856 10112
rect 15841 10075 15899 10081
rect 16850 10072 16856 10084
rect 16908 10072 16914 10124
rect 19058 10072 19064 10124
rect 19116 10112 19122 10124
rect 19702 10121 19708 10124
rect 19648 10115 19708 10121
rect 19648 10112 19660 10115
rect 19116 10084 19660 10112
rect 19116 10072 19122 10084
rect 19648 10081 19660 10084
rect 19694 10081 19708 10115
rect 19648 10075 19708 10081
rect 19702 10072 19708 10075
rect 19760 10072 19766 10124
rect 20714 10072 20720 10124
rect 20772 10112 20778 10124
rect 21545 10115 21603 10121
rect 21545 10112 21557 10115
rect 20772 10084 21557 10112
rect 20772 10072 20778 10084
rect 21545 10081 21557 10084
rect 21591 10112 21603 10115
rect 22554 10112 22560 10124
rect 21591 10084 22560 10112
rect 21591 10081 21603 10084
rect 21545 10075 21603 10081
rect 22554 10072 22560 10084
rect 22612 10072 22618 10124
rect 24210 10072 24216 10124
rect 24268 10072 24274 10124
rect 6454 10044 6460 10056
rect 6415 10016 6460 10044
rect 6454 10004 6460 10016
rect 6512 10004 6518 10056
rect 7466 10044 7472 10056
rect 7427 10016 7472 10044
rect 7466 10004 7472 10016
rect 7524 10004 7530 10056
rect 11149 10047 11207 10053
rect 11149 10044 11161 10047
rect 8449 10016 11161 10044
rect 7006 9936 7012 9988
rect 7064 9976 7070 9988
rect 8449 9976 8477 10016
rect 11149 10013 11161 10016
rect 11195 10044 11207 10047
rect 11606 10044 11612 10056
rect 11195 10016 11612 10044
rect 11195 10013 11207 10016
rect 11149 10007 11207 10013
rect 11606 10004 11612 10016
rect 11664 10004 11670 10056
rect 14366 10044 14372 10056
rect 14327 10016 14372 10044
rect 14366 10004 14372 10016
rect 14424 10004 14430 10056
rect 17494 10004 17500 10056
rect 17552 10044 17558 10056
rect 18141 10047 18199 10053
rect 18141 10044 18153 10047
rect 17552 10016 18153 10044
rect 17552 10004 17558 10016
rect 18141 10013 18153 10016
rect 18187 10013 18199 10047
rect 18141 10007 18199 10013
rect 22833 10047 22891 10053
rect 22833 10013 22845 10047
rect 22879 10044 22891 10047
rect 23385 10047 23443 10053
rect 23385 10044 23397 10047
rect 22879 10016 23397 10044
rect 22879 10013 22891 10016
rect 22833 10007 22891 10013
rect 23385 10013 23397 10016
rect 23431 10044 23443 10047
rect 24026 10044 24032 10056
rect 23431 10016 24032 10044
rect 23431 10013 23443 10016
rect 23385 10007 23443 10013
rect 24026 10004 24032 10016
rect 24084 10004 24090 10056
rect 24946 10044 24952 10056
rect 24907 10016 24952 10044
rect 24946 10004 24952 10016
rect 25004 10004 25010 10056
rect 25225 10047 25283 10053
rect 25225 10044 25237 10047
rect 25056 10016 25237 10044
rect 7064 9948 8477 9976
rect 7064 9936 7070 9948
rect 9398 9936 9404 9988
rect 9456 9976 9462 9988
rect 10321 9979 10379 9985
rect 10321 9976 10333 9979
rect 9456 9948 10333 9976
rect 9456 9936 9462 9948
rect 10321 9945 10333 9948
rect 10367 9945 10379 9979
rect 10321 9939 10379 9945
rect 14458 9936 14464 9988
rect 14516 9976 14522 9988
rect 20530 9976 20536 9988
rect 14516 9948 20536 9976
rect 14516 9936 14522 9948
rect 20530 9936 20536 9948
rect 20588 9936 20594 9988
rect 22922 9936 22928 9988
rect 22980 9976 22986 9988
rect 25056 9976 25084 10016
rect 25225 10013 25237 10016
rect 25271 10013 25283 10047
rect 25225 10007 25283 10013
rect 22980 9948 23888 9976
rect 22980 9936 22986 9948
rect 4062 9868 4068 9920
rect 4120 9908 4126 9920
rect 4939 9911 4997 9917
rect 4939 9908 4951 9911
rect 4120 9880 4951 9908
rect 4120 9868 4126 9880
rect 4939 9877 4951 9880
rect 4985 9877 4997 9911
rect 4939 9871 4997 9877
rect 7190 9868 7196 9920
rect 7248 9908 7254 9920
rect 8389 9911 8447 9917
rect 8389 9908 8401 9911
rect 7248 9880 8401 9908
rect 7248 9868 7254 9880
rect 8389 9877 8401 9880
rect 8435 9908 8447 9911
rect 8478 9908 8484 9920
rect 8435 9880 8484 9908
rect 8435 9877 8447 9880
rect 8389 9871 8447 9877
rect 8478 9868 8484 9880
rect 8536 9868 8542 9920
rect 13538 9908 13544 9920
rect 13499 9880 13544 9908
rect 13538 9868 13544 9880
rect 13596 9868 13602 9920
rect 15105 9911 15163 9917
rect 15105 9877 15117 9911
rect 15151 9908 15163 9911
rect 15378 9908 15384 9920
rect 15151 9880 15384 9908
rect 15151 9877 15163 9880
rect 15105 9871 15163 9877
rect 15378 9868 15384 9880
rect 15436 9868 15442 9920
rect 16991 9911 17049 9917
rect 16991 9877 17003 9911
rect 17037 9908 17049 9911
rect 17218 9908 17224 9920
rect 17037 9880 17224 9908
rect 17037 9877 17049 9880
rect 16991 9871 17049 9877
rect 17218 9868 17224 9880
rect 17276 9868 17282 9920
rect 19150 9868 19156 9920
rect 19208 9908 19214 9920
rect 19751 9911 19809 9917
rect 19751 9908 19763 9911
rect 19208 9880 19763 9908
rect 19208 9868 19214 9880
rect 19751 9877 19763 9880
rect 19797 9877 19809 9911
rect 23198 9908 23204 9920
rect 23159 9880 23204 9908
rect 19751 9871 19809 9877
rect 23198 9868 23204 9880
rect 23256 9868 23262 9920
rect 23382 9868 23388 9920
rect 23440 9908 23446 9920
rect 23658 9908 23664 9920
rect 23440 9880 23664 9908
rect 23440 9868 23446 9880
rect 23658 9868 23664 9880
rect 23716 9868 23722 9920
rect 23860 9908 23888 9948
rect 24044 9948 25084 9976
rect 24044 9908 24072 9948
rect 23860 9880 24072 9908
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 4798 9704 4804 9716
rect 4759 9676 4804 9704
rect 4798 9664 4804 9676
rect 4856 9664 4862 9716
rect 6546 9704 6552 9716
rect 6507 9676 6552 9704
rect 6546 9664 6552 9676
rect 6604 9664 6610 9716
rect 12575 9707 12633 9713
rect 12575 9673 12587 9707
rect 12621 9704 12633 9707
rect 12710 9704 12716 9716
rect 12621 9676 12716 9704
rect 12621 9673 12633 9676
rect 12575 9667 12633 9673
rect 12710 9664 12716 9676
rect 12768 9664 12774 9716
rect 13354 9664 13360 9716
rect 13412 9704 13418 9716
rect 13630 9704 13636 9716
rect 13412 9676 13636 9704
rect 13412 9664 13418 9676
rect 13630 9664 13636 9676
rect 13688 9664 13694 9716
rect 15289 9707 15347 9713
rect 15289 9673 15301 9707
rect 15335 9704 15347 9707
rect 15746 9704 15752 9716
rect 15335 9676 15752 9704
rect 15335 9673 15347 9676
rect 15289 9667 15347 9673
rect 15746 9664 15752 9676
rect 15804 9664 15810 9716
rect 17678 9664 17684 9716
rect 17736 9704 17742 9716
rect 18325 9707 18383 9713
rect 18325 9704 18337 9707
rect 17736 9676 18337 9704
rect 17736 9664 17742 9676
rect 18325 9673 18337 9676
rect 18371 9673 18383 9707
rect 19702 9704 19708 9716
rect 19663 9676 19708 9704
rect 18325 9667 18383 9673
rect 10597 9639 10655 9645
rect 10597 9636 10609 9639
rect 8404 9608 10609 9636
rect 7558 9528 7564 9580
rect 7616 9568 7622 9580
rect 7837 9571 7895 9577
rect 7837 9568 7849 9571
rect 7616 9540 7849 9568
rect 7616 9528 7622 9540
rect 7837 9537 7849 9540
rect 7883 9568 7895 9571
rect 8113 9571 8171 9577
rect 8113 9568 8125 9571
rect 7883 9540 8125 9568
rect 7883 9537 7895 9540
rect 7837 9531 7895 9537
rect 8113 9537 8125 9540
rect 8159 9537 8171 9571
rect 8113 9531 8171 9537
rect 5629 9503 5687 9509
rect 5629 9469 5641 9503
rect 5675 9500 5687 9503
rect 5721 9503 5779 9509
rect 5721 9500 5733 9503
rect 5675 9472 5733 9500
rect 5675 9469 5687 9472
rect 5629 9463 5687 9469
rect 5721 9469 5733 9472
rect 5767 9500 5779 9503
rect 7006 9500 7012 9512
rect 5767 9472 7012 9500
rect 5767 9469 5779 9472
rect 5721 9463 5779 9469
rect 7006 9460 7012 9472
rect 7064 9460 7070 9512
rect 7190 9500 7196 9512
rect 7151 9472 7196 9500
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 5534 9392 5540 9444
rect 5592 9432 5598 9444
rect 6181 9435 6239 9441
rect 6181 9432 6193 9435
rect 5592 9404 6193 9432
rect 5592 9392 5598 9404
rect 6181 9401 6193 9404
rect 6227 9432 6239 9435
rect 8404 9432 8432 9608
rect 10597 9605 10609 9608
rect 10643 9636 10655 9639
rect 11238 9636 11244 9648
rect 10643 9608 11244 9636
rect 10643 9605 10655 9608
rect 10597 9599 10655 9605
rect 11238 9596 11244 9608
rect 11296 9596 11302 9648
rect 13722 9596 13728 9648
rect 13780 9636 13786 9648
rect 16942 9636 16948 9648
rect 13780 9608 16948 9636
rect 13780 9596 13786 9608
rect 16942 9596 16948 9608
rect 17000 9596 17006 9648
rect 18340 9636 18368 9667
rect 19702 9664 19708 9676
rect 19760 9664 19766 9716
rect 21450 9664 21456 9716
rect 21508 9704 21514 9716
rect 21545 9707 21603 9713
rect 21545 9704 21557 9707
rect 21508 9676 21557 9704
rect 21508 9664 21514 9676
rect 21545 9673 21557 9676
rect 21591 9673 21603 9707
rect 21545 9667 21603 9673
rect 23842 9664 23848 9716
rect 23900 9704 23906 9716
rect 25363 9707 25421 9713
rect 25363 9704 25375 9707
rect 23900 9676 25375 9704
rect 23900 9664 23906 9676
rect 25363 9673 25375 9676
rect 25409 9673 25421 9707
rect 25363 9667 25421 9673
rect 19429 9639 19487 9645
rect 18340 9608 18644 9636
rect 8754 9528 8760 9580
rect 8812 9568 8818 9580
rect 8812 9540 12547 9568
rect 8812 9528 8818 9540
rect 8665 9503 8723 9509
rect 8665 9500 8677 9503
rect 6227 9404 8432 9432
rect 8496 9472 8677 9500
rect 6227 9401 6239 9404
rect 6181 9395 6239 9401
rect 5905 9367 5963 9373
rect 5905 9333 5917 9367
rect 5951 9364 5963 9367
rect 5994 9364 6000 9376
rect 5951 9336 6000 9364
rect 5951 9333 5963 9336
rect 5905 9327 5963 9333
rect 5994 9324 6000 9336
rect 6052 9324 6058 9376
rect 7834 9324 7840 9376
rect 7892 9364 7898 9376
rect 8496 9373 8524 9472
rect 8665 9469 8677 9472
rect 8711 9469 8723 9503
rect 8665 9463 8723 9469
rect 9217 9503 9275 9509
rect 9217 9469 9229 9503
rect 9263 9500 9275 9503
rect 9306 9500 9312 9512
rect 9263 9472 9312 9500
rect 9263 9469 9275 9472
rect 9217 9463 9275 9469
rect 9306 9460 9312 9472
rect 9364 9460 9370 9512
rect 11054 9500 11060 9512
rect 11015 9472 11060 9500
rect 11054 9460 11060 9472
rect 11112 9460 11118 9512
rect 11238 9500 11244 9512
rect 11199 9472 11244 9500
rect 11238 9460 11244 9472
rect 11296 9460 11302 9512
rect 12519 9509 12547 9540
rect 13538 9528 13544 9580
rect 13596 9568 13602 9580
rect 17865 9571 17923 9577
rect 13596 9540 13952 9568
rect 13596 9528 13602 9540
rect 12504 9503 12562 9509
rect 12504 9469 12516 9503
rect 12550 9500 12562 9503
rect 12894 9500 12900 9512
rect 12550 9472 12900 9500
rect 12550 9469 12562 9472
rect 12504 9463 12562 9469
rect 12894 9460 12900 9472
rect 12952 9460 12958 9512
rect 13924 9509 13952 9540
rect 17865 9537 17877 9571
rect 17911 9568 17923 9571
rect 18322 9568 18328 9580
rect 17911 9540 18328 9568
rect 17911 9537 17923 9540
rect 17865 9531 17923 9537
rect 18322 9528 18328 9540
rect 18380 9568 18386 9580
rect 18509 9571 18567 9577
rect 18509 9568 18521 9571
rect 18380 9540 18521 9568
rect 18380 9528 18386 9540
rect 18509 9537 18521 9540
rect 18555 9537 18567 9571
rect 18509 9531 18567 9537
rect 13449 9503 13507 9509
rect 13449 9500 13461 9503
rect 13280 9472 13461 9500
rect 10134 9392 10140 9444
rect 10192 9432 10198 9444
rect 10229 9435 10287 9441
rect 10229 9432 10241 9435
rect 10192 9404 10241 9432
rect 10192 9392 10198 9404
rect 10229 9401 10241 9404
rect 10275 9432 10287 9435
rect 11514 9432 11520 9444
rect 10275 9404 10732 9432
rect 11475 9404 11520 9432
rect 10275 9401 10287 9404
rect 10229 9395 10287 9401
rect 8481 9367 8539 9373
rect 8481 9364 8493 9367
rect 7892 9336 8493 9364
rect 7892 9324 7898 9336
rect 8481 9333 8493 9336
rect 8527 9333 8539 9367
rect 8754 9364 8760 9376
rect 8715 9336 8760 9364
rect 8481 9327 8539 9333
rect 8754 9324 8760 9336
rect 8812 9324 8818 9376
rect 10704 9364 10732 9404
rect 11514 9392 11520 9404
rect 11572 9392 11578 9444
rect 11790 9364 11796 9376
rect 10704 9336 11796 9364
rect 11790 9324 11796 9336
rect 11848 9364 11854 9376
rect 11885 9367 11943 9373
rect 11885 9364 11897 9367
rect 11848 9336 11897 9364
rect 11848 9324 11854 9336
rect 11885 9333 11897 9336
rect 11931 9364 11943 9367
rect 12342 9364 12348 9376
rect 11931 9336 12348 9364
rect 11931 9333 11943 9336
rect 11885 9327 11943 9333
rect 12342 9324 12348 9336
rect 12400 9324 12406 9376
rect 13078 9324 13084 9376
rect 13136 9364 13142 9376
rect 13280 9373 13308 9472
rect 13449 9469 13461 9472
rect 13495 9469 13507 9503
rect 13449 9463 13507 9469
rect 13909 9503 13967 9509
rect 13909 9469 13921 9503
rect 13955 9500 13967 9503
rect 14090 9500 14096 9512
rect 13955 9472 14096 9500
rect 13955 9469 13967 9472
rect 13909 9463 13967 9469
rect 14090 9460 14096 9472
rect 14148 9460 14154 9512
rect 15378 9500 15384 9512
rect 15339 9472 15384 9500
rect 15378 9460 15384 9472
rect 15436 9460 15442 9512
rect 16206 9460 16212 9512
rect 16264 9500 16270 9512
rect 16301 9503 16359 9509
rect 16301 9500 16313 9503
rect 16264 9472 16313 9500
rect 16264 9460 16270 9472
rect 16301 9469 16313 9472
rect 16347 9500 16359 9503
rect 18046 9500 18052 9512
rect 16347 9472 18052 9500
rect 16347 9469 16359 9472
rect 16301 9463 16359 9469
rect 18046 9460 18052 9472
rect 18104 9460 18110 9512
rect 14182 9432 14188 9444
rect 14143 9404 14188 9432
rect 14182 9392 14188 9404
rect 14240 9392 14246 9444
rect 14553 9435 14611 9441
rect 14553 9401 14565 9435
rect 14599 9432 14611 9435
rect 14921 9435 14979 9441
rect 14921 9432 14933 9435
rect 14599 9404 14933 9432
rect 14599 9401 14611 9404
rect 14553 9395 14611 9401
rect 14921 9401 14933 9404
rect 14967 9432 14979 9435
rect 15630 9435 15688 9441
rect 14967 9404 15332 9432
rect 14967 9401 14979 9404
rect 14921 9395 14979 9401
rect 13265 9367 13323 9373
rect 13265 9364 13277 9367
rect 13136 9336 13277 9364
rect 13136 9324 13142 9336
rect 13265 9333 13277 9336
rect 13311 9364 13323 9367
rect 13906 9364 13912 9376
rect 13311 9336 13912 9364
rect 13311 9333 13323 9336
rect 13265 9327 13323 9333
rect 13906 9324 13912 9336
rect 13964 9364 13970 9376
rect 14568 9364 14596 9395
rect 13964 9336 14596 9364
rect 15304 9364 15332 9404
rect 15630 9401 15642 9435
rect 15676 9432 15688 9435
rect 15746 9432 15752 9444
rect 15676 9404 15752 9432
rect 15676 9401 15688 9404
rect 15630 9395 15688 9401
rect 15746 9392 15752 9404
rect 15804 9392 15810 9444
rect 15838 9392 15844 9444
rect 15896 9432 15902 9444
rect 16114 9432 16120 9444
rect 15896 9404 16120 9432
rect 15896 9392 15902 9404
rect 16114 9392 16120 9404
rect 16172 9432 16178 9444
rect 16850 9432 16856 9444
rect 16172 9404 16856 9432
rect 16172 9392 16178 9404
rect 16850 9392 16856 9404
rect 16908 9392 16914 9444
rect 18616 9432 18644 9608
rect 19429 9605 19441 9639
rect 19475 9636 19487 9639
rect 20165 9639 20223 9645
rect 20165 9636 20177 9639
rect 19475 9608 20177 9636
rect 19475 9605 19487 9608
rect 19429 9599 19487 9605
rect 20165 9605 20177 9608
rect 20211 9636 20223 9639
rect 20530 9636 20536 9648
rect 20211 9608 20536 9636
rect 20211 9605 20223 9608
rect 20165 9599 20223 9605
rect 20530 9596 20536 9608
rect 20588 9636 20594 9648
rect 23106 9636 23112 9648
rect 20588 9608 23112 9636
rect 20588 9596 20594 9608
rect 23106 9596 23112 9608
rect 23164 9596 23170 9648
rect 24949 9639 25007 9645
rect 24949 9605 24961 9639
rect 24995 9636 25007 9639
rect 25222 9636 25228 9648
rect 24995 9608 25228 9636
rect 24995 9605 25007 9608
rect 24949 9599 25007 9605
rect 25222 9596 25228 9608
rect 25280 9596 25286 9648
rect 19978 9528 19984 9580
rect 20036 9568 20042 9580
rect 20349 9571 20407 9577
rect 20349 9568 20361 9571
rect 20036 9540 20361 9568
rect 20036 9528 20042 9540
rect 20349 9537 20361 9540
rect 20395 9537 20407 9571
rect 20622 9568 20628 9580
rect 20583 9540 20628 9568
rect 20349 9531 20407 9537
rect 20622 9528 20628 9540
rect 20680 9528 20686 9580
rect 21726 9528 21732 9580
rect 21784 9568 21790 9580
rect 21821 9571 21879 9577
rect 21821 9568 21833 9571
rect 21784 9540 21833 9568
rect 21784 9528 21790 9540
rect 21821 9537 21833 9540
rect 21867 9537 21879 9571
rect 21821 9531 21879 9537
rect 23198 9528 23204 9580
rect 23256 9568 23262 9580
rect 23753 9571 23811 9577
rect 23753 9568 23765 9571
rect 23256 9540 23765 9568
rect 23256 9528 23262 9540
rect 23753 9537 23765 9540
rect 23799 9568 23811 9571
rect 23934 9568 23940 9580
rect 23799 9540 23940 9568
rect 23799 9537 23811 9540
rect 23753 9531 23811 9537
rect 23934 9528 23940 9540
rect 23992 9528 23998 9580
rect 24118 9568 24124 9580
rect 24079 9540 24124 9568
rect 24118 9528 24124 9540
rect 24176 9528 24182 9580
rect 24670 9460 24676 9512
rect 24728 9500 24734 9512
rect 25260 9503 25318 9509
rect 25260 9500 25272 9503
rect 24728 9472 25272 9500
rect 24728 9460 24734 9472
rect 25260 9469 25272 9472
rect 25306 9500 25318 9503
rect 25685 9503 25743 9509
rect 25685 9500 25697 9503
rect 25306 9472 25697 9500
rect 25306 9469 25318 9472
rect 25260 9463 25318 9469
rect 25685 9469 25697 9472
rect 25731 9469 25743 9503
rect 25685 9463 25743 9469
rect 18871 9435 18929 9441
rect 18871 9432 18883 9435
rect 18616 9404 18883 9432
rect 18871 9401 18883 9404
rect 18917 9432 18929 9435
rect 18966 9432 18972 9444
rect 18917 9404 18972 9432
rect 18917 9401 18929 9404
rect 18871 9395 18929 9401
rect 18966 9392 18972 9404
rect 19024 9392 19030 9444
rect 20441 9435 20499 9441
rect 20441 9401 20453 9435
rect 20487 9432 20499 9435
rect 20530 9432 20536 9444
rect 20487 9404 20536 9432
rect 20487 9401 20499 9404
rect 20441 9395 20499 9401
rect 20530 9392 20536 9404
rect 20588 9392 20594 9444
rect 21450 9392 21456 9444
rect 21508 9432 21514 9444
rect 22186 9441 22192 9444
rect 22142 9435 22192 9441
rect 22142 9432 22154 9435
rect 21508 9404 22154 9432
rect 21508 9392 21514 9404
rect 22142 9401 22154 9404
rect 22188 9401 22192 9435
rect 22142 9395 22192 9401
rect 22186 9392 22192 9395
rect 22244 9432 22250 9444
rect 23017 9435 23075 9441
rect 23017 9432 23029 9435
rect 22244 9404 23029 9432
rect 22244 9392 22250 9404
rect 23017 9401 23029 9404
rect 23063 9401 23075 9435
rect 23017 9395 23075 9401
rect 23845 9435 23903 9441
rect 23845 9401 23857 9435
rect 23891 9401 23903 9435
rect 23845 9395 23903 9401
rect 15470 9364 15476 9376
rect 15304 9336 15476 9364
rect 13964 9324 13970 9336
rect 15470 9324 15476 9336
rect 15528 9364 15534 9376
rect 16298 9364 16304 9376
rect 15528 9336 16304 9364
rect 15528 9324 15534 9336
rect 16298 9324 16304 9336
rect 16356 9324 16362 9376
rect 17494 9364 17500 9376
rect 17455 9336 17500 9364
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 22741 9367 22799 9373
rect 22741 9333 22753 9367
rect 22787 9364 22799 9367
rect 23385 9367 23443 9373
rect 23385 9364 23397 9367
rect 22787 9336 23397 9364
rect 22787 9333 22799 9336
rect 22741 9327 22799 9333
rect 23385 9333 23397 9336
rect 23431 9364 23443 9367
rect 23860 9364 23888 9395
rect 23431 9336 23888 9364
rect 23431 9333 23443 9336
rect 23385 9327 23443 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 5169 9163 5227 9169
rect 5169 9160 5181 9163
rect 4120 9132 5181 9160
rect 4120 9120 4126 9132
rect 5169 9129 5181 9132
rect 5215 9160 5227 9163
rect 5258 9160 5264 9172
rect 5215 9132 5264 9160
rect 5215 9129 5227 9132
rect 5169 9123 5227 9129
rect 5258 9120 5264 9132
rect 5316 9120 5322 9172
rect 7190 9160 7196 9172
rect 7151 9132 7196 9160
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 9861 9163 9919 9169
rect 9861 9129 9873 9163
rect 9907 9160 9919 9163
rect 9950 9160 9956 9172
rect 9907 9132 9956 9160
rect 9907 9129 9919 9132
rect 9861 9123 9919 9129
rect 9950 9120 9956 9132
rect 10008 9120 10014 9172
rect 13909 9163 13967 9169
rect 13909 9129 13921 9163
rect 13955 9160 13967 9163
rect 14274 9160 14280 9172
rect 13955 9132 14280 9160
rect 13955 9129 13967 9132
rect 13909 9123 13967 9129
rect 14274 9120 14280 9132
rect 14332 9120 14338 9172
rect 14826 9120 14832 9172
rect 14884 9160 14890 9172
rect 15013 9163 15071 9169
rect 15013 9160 15025 9163
rect 14884 9132 15025 9160
rect 14884 9120 14890 9132
rect 15013 9129 15025 9132
rect 15059 9160 15071 9163
rect 15746 9160 15752 9172
rect 15059 9132 15752 9160
rect 15059 9129 15071 9132
rect 15013 9123 15071 9129
rect 15746 9120 15752 9132
rect 15804 9120 15810 9172
rect 15838 9120 15844 9172
rect 15896 9160 15902 9172
rect 15933 9163 15991 9169
rect 15933 9160 15945 9163
rect 15896 9132 15945 9160
rect 15896 9120 15902 9132
rect 15933 9129 15945 9132
rect 15979 9129 15991 9163
rect 15933 9123 15991 9129
rect 16390 9120 16396 9172
rect 16448 9160 16454 9172
rect 16485 9163 16543 9169
rect 16485 9160 16497 9163
rect 16448 9132 16497 9160
rect 16448 9120 16454 9132
rect 16485 9129 16497 9132
rect 16531 9160 16543 9163
rect 18138 9160 18144 9172
rect 16531 9132 18144 9160
rect 16531 9129 16543 9132
rect 16485 9123 16543 9129
rect 18138 9120 18144 9132
rect 18196 9120 18202 9172
rect 19978 9120 19984 9172
rect 20036 9160 20042 9172
rect 20257 9163 20315 9169
rect 20257 9160 20269 9163
rect 20036 9132 20269 9160
rect 20036 9120 20042 9132
rect 20257 9129 20269 9132
rect 20303 9129 20315 9163
rect 20714 9160 20720 9172
rect 20675 9132 20720 9160
rect 20257 9123 20315 9129
rect 20714 9120 20720 9132
rect 20772 9120 20778 9172
rect 21726 9160 21732 9172
rect 21687 9132 21732 9160
rect 21726 9120 21732 9132
rect 21784 9120 21790 9172
rect 22186 9120 22192 9172
rect 22244 9160 22250 9172
rect 22281 9163 22339 9169
rect 22281 9160 22293 9163
rect 22244 9132 22293 9160
rect 22244 9120 22250 9132
rect 22281 9129 22293 9132
rect 22327 9129 22339 9163
rect 22281 9123 22339 9129
rect 22833 9163 22891 9169
rect 22833 9129 22845 9163
rect 22879 9160 22891 9163
rect 23474 9160 23480 9172
rect 22879 9132 23480 9160
rect 22879 9129 22891 9132
rect 22833 9123 22891 9129
rect 23474 9120 23480 9132
rect 23532 9160 23538 9172
rect 24670 9160 24676 9172
rect 23532 9132 24676 9160
rect 23532 9120 23538 9132
rect 4706 9052 4712 9104
rect 4764 9092 4770 9104
rect 6178 9092 6184 9104
rect 4764 9064 6184 9092
rect 4764 9052 4770 9064
rect 6178 9052 6184 9064
rect 6236 9052 6242 9104
rect 6270 9052 6276 9104
rect 6328 9092 6334 9104
rect 7929 9095 7987 9101
rect 6328 9064 6373 9092
rect 6328 9052 6334 9064
rect 7929 9061 7941 9095
rect 7975 9092 7987 9095
rect 8202 9092 8208 9104
rect 7975 9064 8208 9092
rect 7975 9061 7987 9064
rect 7929 9055 7987 9061
rect 8202 9052 8208 9064
rect 8260 9052 8266 9104
rect 12526 9052 12532 9104
rect 12584 9092 12590 9104
rect 12942 9095 13000 9101
rect 12942 9092 12954 9095
rect 12584 9064 12954 9092
rect 12584 9052 12590 9064
rect 12942 9061 12954 9064
rect 12988 9061 13000 9095
rect 18871 9095 18929 9101
rect 12942 9055 13000 9061
rect 13786 9064 15700 9092
rect 9398 8984 9404 9036
rect 9456 9024 9462 9036
rect 9677 9027 9735 9033
rect 9677 9024 9689 9027
rect 9456 8996 9689 9024
rect 9456 8984 9462 8996
rect 9677 8993 9689 8996
rect 9723 8993 9735 9027
rect 11054 9024 11060 9036
rect 11015 8996 11060 9024
rect 9677 8987 9735 8993
rect 11054 8984 11060 8996
rect 11112 8984 11118 9036
rect 11422 8984 11428 9036
rect 11480 9024 11486 9036
rect 11517 9027 11575 9033
rect 11517 9024 11529 9027
rect 11480 8996 11529 9024
rect 11480 8984 11486 8996
rect 11517 8993 11529 8996
rect 11563 9024 11575 9027
rect 13786 9024 13814 9064
rect 15562 9024 15568 9036
rect 11563 8996 13814 9024
rect 15523 8996 15568 9024
rect 11563 8993 11575 8996
rect 11517 8987 11575 8993
rect 15562 8984 15568 8996
rect 15620 8984 15626 9036
rect 15672 9024 15700 9064
rect 18871 9061 18883 9095
rect 18917 9092 18929 9095
rect 18966 9092 18972 9104
rect 18917 9064 18972 9092
rect 18917 9061 18929 9064
rect 18871 9055 18929 9061
rect 18966 9052 18972 9064
rect 19024 9052 19030 9104
rect 23290 9092 23296 9104
rect 23251 9064 23296 9092
rect 23290 9052 23296 9064
rect 23348 9052 23354 9104
rect 23750 9092 23756 9104
rect 23711 9064 23756 9092
rect 23750 9052 23756 9064
rect 23808 9052 23814 9104
rect 23860 9101 23888 9132
rect 24670 9120 24676 9132
rect 24728 9160 24734 9172
rect 24765 9163 24823 9169
rect 24765 9160 24777 9163
rect 24728 9132 24777 9160
rect 24728 9120 24734 9132
rect 24765 9129 24777 9132
rect 24811 9160 24823 9163
rect 25222 9160 25228 9172
rect 24811 9132 25228 9160
rect 24811 9129 24823 9132
rect 24765 9123 24823 9129
rect 25222 9120 25228 9132
rect 25280 9120 25286 9172
rect 23845 9095 23903 9101
rect 23845 9061 23857 9095
rect 23891 9061 23903 9095
rect 23845 9055 23903 9061
rect 17310 9024 17316 9036
rect 15672 8996 17316 9024
rect 17310 8984 17316 8996
rect 17368 8984 17374 9036
rect 17564 9027 17622 9033
rect 17564 8993 17576 9027
rect 17610 9024 17622 9027
rect 17678 9024 17684 9036
rect 17610 8996 17684 9024
rect 17610 8993 17622 8996
rect 17564 8987 17622 8993
rect 17678 8984 17684 8996
rect 17736 8984 17742 9036
rect 20438 8984 20444 9036
rect 20496 9024 20502 9036
rect 20898 9024 20904 9036
rect 20956 9033 20962 9036
rect 20956 9027 20994 9033
rect 20496 8996 20904 9024
rect 20496 8984 20502 8996
rect 20898 8984 20904 8996
rect 20982 8993 20994 9027
rect 20956 8987 20994 8993
rect 20956 8984 20962 8987
rect 21634 8984 21640 9036
rect 21692 9024 21698 9036
rect 21913 9027 21971 9033
rect 21913 9024 21925 9027
rect 21692 8996 21925 9024
rect 21692 8984 21698 8996
rect 21913 8993 21925 8996
rect 21959 8993 21971 9027
rect 21913 8987 21971 8993
rect 25292 9027 25350 9033
rect 25292 8993 25304 9027
rect 25338 9024 25350 9027
rect 25498 9024 25504 9036
rect 25338 8996 25504 9024
rect 25338 8993 25350 8996
rect 25292 8987 25350 8993
rect 25498 8984 25504 8996
rect 25556 8984 25562 9036
rect 6454 8956 6460 8968
rect 6415 8928 6460 8956
rect 6454 8916 6460 8928
rect 6512 8956 6518 8968
rect 8113 8959 8171 8965
rect 8113 8956 8125 8959
rect 6512 8928 8125 8956
rect 6512 8916 6518 8928
rect 8113 8925 8125 8928
rect 8159 8956 8171 8959
rect 9030 8956 9036 8968
rect 8159 8928 9036 8956
rect 8159 8925 8171 8928
rect 8113 8919 8171 8925
rect 9030 8916 9036 8928
rect 9088 8916 9094 8968
rect 11793 8959 11851 8965
rect 11793 8925 11805 8959
rect 11839 8956 11851 8959
rect 12621 8959 12679 8965
rect 12621 8956 12633 8959
rect 11839 8928 12633 8956
rect 11839 8925 11851 8928
rect 11793 8919 11851 8925
rect 12621 8925 12633 8928
rect 12667 8956 12679 8959
rect 12710 8956 12716 8968
rect 12667 8928 12716 8956
rect 12667 8925 12679 8928
rect 12621 8919 12679 8925
rect 12710 8916 12716 8928
rect 12768 8916 12774 8968
rect 14366 8916 14372 8968
rect 14424 8956 14430 8968
rect 18509 8959 18567 8965
rect 18509 8956 18521 8959
rect 14424 8928 18521 8956
rect 14424 8916 14430 8928
rect 18509 8925 18521 8928
rect 18555 8956 18567 8959
rect 18690 8956 18696 8968
rect 18555 8928 18696 8956
rect 18555 8925 18567 8928
rect 18509 8919 18567 8925
rect 18690 8916 18696 8928
rect 18748 8916 18754 8968
rect 24026 8956 24032 8968
rect 23987 8928 24032 8956
rect 24026 8916 24032 8928
rect 24084 8916 24090 8968
rect 7466 8888 7472 8900
rect 6840 8860 7472 8888
rect 3694 8780 3700 8832
rect 3752 8820 3758 8832
rect 6840 8820 6868 8860
rect 7466 8848 7472 8860
rect 7524 8848 7530 8900
rect 8662 8888 8668 8900
rect 8623 8860 8668 8888
rect 8662 8848 8668 8860
rect 8720 8848 8726 8900
rect 8938 8848 8944 8900
rect 8996 8888 9002 8900
rect 19705 8891 19763 8897
rect 19705 8888 19717 8891
rect 8996 8860 19717 8888
rect 8996 8848 9002 8860
rect 19705 8857 19717 8860
rect 19751 8888 19763 8891
rect 19794 8888 19800 8900
rect 19751 8860 19800 8888
rect 19751 8857 19763 8860
rect 19705 8851 19763 8857
rect 19794 8848 19800 8860
rect 19852 8848 19858 8900
rect 21174 8888 21180 8900
rect 21135 8860 21180 8888
rect 21174 8848 21180 8860
rect 21232 8848 21238 8900
rect 24946 8848 24952 8900
rect 25004 8888 25010 8900
rect 25133 8891 25191 8897
rect 25133 8888 25145 8891
rect 25004 8860 25145 8888
rect 25004 8848 25010 8860
rect 25133 8857 25145 8860
rect 25179 8888 25191 8891
rect 25314 8888 25320 8900
rect 25179 8860 25320 8888
rect 25179 8857 25191 8860
rect 25133 8851 25191 8857
rect 25314 8848 25320 8860
rect 25372 8848 25378 8900
rect 3752 8792 6868 8820
rect 9125 8823 9183 8829
rect 3752 8780 3758 8792
rect 9125 8789 9137 8823
rect 9171 8820 9183 8823
rect 9306 8820 9312 8832
rect 9171 8792 9312 8820
rect 9171 8789 9183 8792
rect 9125 8783 9183 8789
rect 9306 8780 9312 8792
rect 9364 8780 9370 8832
rect 9950 8780 9956 8832
rect 10008 8820 10014 8832
rect 10137 8823 10195 8829
rect 10137 8820 10149 8823
rect 10008 8792 10149 8820
rect 10008 8780 10014 8792
rect 10137 8789 10149 8792
rect 10183 8820 10195 8823
rect 10781 8823 10839 8829
rect 10781 8820 10793 8823
rect 10183 8792 10793 8820
rect 10183 8789 10195 8792
rect 10137 8783 10195 8789
rect 10781 8789 10793 8792
rect 10827 8820 10839 8823
rect 11054 8820 11060 8832
rect 10827 8792 11060 8820
rect 10827 8789 10839 8792
rect 10781 8783 10839 8789
rect 11054 8780 11060 8792
rect 11112 8780 11118 8832
rect 12158 8780 12164 8832
rect 12216 8820 12222 8832
rect 12526 8820 12532 8832
rect 12216 8792 12532 8820
rect 12216 8780 12222 8792
rect 12526 8780 12532 8792
rect 12584 8780 12590 8832
rect 13541 8823 13599 8829
rect 13541 8789 13553 8823
rect 13587 8820 13599 8823
rect 13998 8820 14004 8832
rect 13587 8792 14004 8820
rect 13587 8789 13599 8792
rect 13541 8783 13599 8789
rect 13998 8780 14004 8792
rect 14056 8780 14062 8832
rect 14274 8820 14280 8832
rect 14235 8792 14280 8820
rect 14274 8780 14280 8792
rect 14332 8780 14338 8832
rect 17405 8823 17463 8829
rect 17405 8789 17417 8823
rect 17451 8820 17463 8823
rect 17635 8823 17693 8829
rect 17635 8820 17647 8823
rect 17451 8792 17647 8820
rect 17451 8789 17463 8792
rect 17405 8783 17463 8789
rect 17635 8789 17647 8792
rect 17681 8820 17693 8823
rect 17954 8820 17960 8832
rect 17681 8792 17960 8820
rect 17681 8789 17693 8792
rect 17635 8783 17693 8789
rect 17954 8780 17960 8792
rect 18012 8780 18018 8832
rect 19426 8820 19432 8832
rect 19387 8792 19432 8820
rect 19426 8780 19432 8792
rect 19484 8780 19490 8832
rect 21450 8820 21456 8832
rect 21411 8792 21456 8820
rect 21450 8780 21456 8792
rect 21508 8780 21514 8832
rect 25406 8820 25412 8832
rect 25367 8792 25412 8820
rect 25406 8780 25412 8792
rect 25464 8780 25470 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 6178 8576 6184 8628
rect 6236 8616 6242 8628
rect 6549 8619 6607 8625
rect 6549 8616 6561 8619
rect 6236 8588 6561 8616
rect 6236 8576 6242 8588
rect 6549 8585 6561 8588
rect 6595 8585 6607 8619
rect 8018 8616 8024 8628
rect 7979 8588 8024 8616
rect 6549 8579 6607 8585
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 8202 8576 8208 8628
rect 8260 8616 8266 8628
rect 9033 8619 9091 8625
rect 9033 8616 9045 8619
rect 8260 8588 9045 8616
rect 8260 8576 8266 8588
rect 9033 8585 9045 8588
rect 9079 8585 9091 8619
rect 11054 8616 11060 8628
rect 11015 8588 11060 8616
rect 9033 8579 9091 8585
rect 11054 8576 11060 8588
rect 11112 8576 11118 8628
rect 11514 8576 11520 8628
rect 11572 8616 11578 8628
rect 11793 8619 11851 8625
rect 11793 8616 11805 8619
rect 11572 8588 11805 8616
rect 11572 8576 11578 8588
rect 11793 8585 11805 8588
rect 11839 8585 11851 8619
rect 13998 8616 14004 8628
rect 13959 8588 14004 8616
rect 11793 8579 11851 8585
rect 8938 8548 8944 8560
rect 4126 8520 8944 8548
rect 106 8372 112 8424
rect 164 8412 170 8424
rect 1432 8415 1490 8421
rect 1432 8412 1444 8415
rect 164 8384 1444 8412
rect 164 8372 170 8384
rect 1432 8381 1444 8384
rect 1478 8412 1490 8415
rect 1857 8415 1915 8421
rect 1857 8412 1869 8415
rect 1478 8384 1869 8412
rect 1478 8381 1490 8384
rect 1432 8375 1490 8381
rect 1857 8381 1869 8384
rect 1903 8381 1915 8415
rect 1857 8375 1915 8381
rect 1535 8347 1593 8353
rect 1535 8313 1547 8347
rect 1581 8344 1593 8347
rect 4126 8344 4154 8520
rect 8938 8508 8944 8520
rect 8996 8508 9002 8560
rect 9766 8548 9772 8560
rect 9679 8520 9772 8548
rect 9766 8508 9772 8520
rect 9824 8548 9830 8560
rect 9824 8520 10548 8548
rect 9824 8508 9830 8520
rect 5258 8480 5264 8492
rect 5219 8452 5264 8480
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8480 5963 8483
rect 6454 8480 6460 8492
rect 5951 8452 6460 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 6454 8440 6460 8452
rect 6512 8440 6518 8492
rect 7742 8440 7748 8492
rect 7800 8480 7806 8492
rect 8113 8483 8171 8489
rect 8113 8480 8125 8483
rect 7800 8452 8125 8480
rect 7800 8440 7806 8452
rect 8113 8449 8125 8452
rect 8159 8480 8171 8483
rect 10413 8483 10471 8489
rect 10413 8480 10425 8483
rect 8159 8452 10425 8480
rect 8159 8449 8171 8452
rect 8113 8443 8171 8449
rect 10413 8449 10425 8452
rect 10459 8449 10471 8483
rect 10413 8443 10471 8449
rect 7101 8415 7159 8421
rect 7101 8381 7113 8415
rect 7147 8412 7159 8415
rect 7190 8412 7196 8424
rect 7147 8384 7196 8412
rect 7147 8381 7159 8384
rect 7101 8375 7159 8381
rect 7190 8372 7196 8384
rect 7248 8412 7254 8424
rect 7561 8415 7619 8421
rect 7561 8412 7573 8415
rect 7248 8384 7573 8412
rect 7248 8372 7254 8384
rect 7561 8381 7573 8384
rect 7607 8381 7619 8415
rect 9950 8412 9956 8424
rect 9911 8384 9956 8412
rect 7561 8375 7619 8381
rect 9950 8372 9956 8384
rect 10008 8372 10014 8424
rect 10321 8415 10379 8421
rect 10321 8381 10333 8415
rect 10367 8412 10379 8415
rect 10520 8412 10548 8520
rect 11808 8480 11836 8579
rect 13998 8576 14004 8588
rect 14056 8576 14062 8628
rect 15289 8619 15347 8625
rect 15289 8585 15301 8619
rect 15335 8616 15347 8619
rect 15562 8616 15568 8628
rect 15335 8588 15568 8616
rect 15335 8585 15347 8588
rect 15289 8579 15347 8585
rect 15562 8576 15568 8588
rect 15620 8576 15626 8628
rect 15657 8619 15715 8625
rect 15657 8585 15669 8619
rect 15703 8616 15715 8619
rect 15838 8616 15844 8628
rect 15703 8588 15844 8616
rect 15703 8585 15715 8588
rect 15657 8579 15715 8585
rect 15838 8576 15844 8588
rect 15896 8576 15902 8628
rect 20898 8616 20904 8628
rect 20859 8588 20904 8616
rect 20898 8576 20904 8588
rect 20956 8576 20962 8628
rect 21634 8576 21640 8628
rect 21692 8616 21698 8628
rect 22649 8619 22707 8625
rect 22649 8616 22661 8619
rect 21692 8588 22661 8616
rect 21692 8576 21698 8588
rect 22649 8585 22661 8588
rect 22695 8585 22707 8619
rect 22649 8579 22707 8585
rect 23474 8576 23480 8628
rect 23532 8616 23538 8628
rect 23532 8588 23577 8616
rect 23532 8576 23538 8588
rect 23750 8576 23756 8628
rect 23808 8616 23814 8628
rect 23845 8619 23903 8625
rect 23845 8616 23857 8619
rect 23808 8588 23857 8616
rect 23808 8576 23814 8588
rect 23845 8585 23857 8588
rect 23891 8585 23903 8619
rect 23845 8579 23903 8585
rect 23934 8576 23940 8628
rect 23992 8616 23998 8628
rect 25409 8619 25467 8625
rect 23992 8588 24992 8616
rect 23992 8576 23998 8588
rect 24964 8560 24992 8588
rect 25409 8585 25421 8619
rect 25455 8616 25467 8619
rect 25498 8616 25504 8628
rect 25455 8588 25504 8616
rect 25455 8585 25467 8588
rect 25409 8579 25467 8585
rect 25498 8576 25504 8588
rect 25556 8576 25562 8628
rect 12894 8508 12900 8560
rect 12952 8548 12958 8560
rect 21913 8551 21971 8557
rect 12952 8520 14596 8548
rect 12952 8508 12958 8520
rect 12437 8483 12495 8489
rect 12437 8480 12449 8483
rect 11808 8452 12449 8480
rect 12437 8449 12449 8452
rect 12483 8449 12495 8483
rect 14274 8480 14280 8492
rect 14235 8452 14280 8480
rect 12437 8443 12495 8449
rect 14274 8440 14280 8452
rect 14332 8440 14338 8492
rect 14568 8489 14596 8520
rect 21913 8517 21925 8551
rect 21959 8548 21971 8551
rect 24026 8548 24032 8560
rect 21959 8520 24032 8548
rect 21959 8517 21971 8520
rect 21913 8511 21971 8517
rect 24026 8508 24032 8520
rect 24084 8508 24090 8560
rect 24946 8548 24952 8560
rect 24859 8520 24952 8548
rect 24946 8508 24952 8520
rect 25004 8508 25010 8560
rect 14553 8483 14611 8489
rect 14553 8449 14565 8483
rect 14599 8449 14611 8483
rect 14553 8443 14611 8449
rect 17954 8440 17960 8492
rect 18012 8480 18018 8492
rect 18233 8483 18291 8489
rect 18233 8480 18245 8483
rect 18012 8452 18245 8480
rect 18012 8440 18018 8452
rect 18233 8449 18245 8452
rect 18279 8449 18291 8483
rect 18874 8480 18880 8492
rect 18835 8452 18880 8480
rect 18233 8443 18291 8449
rect 18874 8440 18880 8452
rect 18932 8440 18938 8492
rect 19794 8480 19800 8492
rect 19755 8452 19800 8480
rect 19794 8440 19800 8452
rect 19852 8440 19858 8492
rect 20441 8483 20499 8489
rect 20441 8449 20453 8483
rect 20487 8480 20499 8483
rect 20622 8480 20628 8492
rect 20487 8452 20628 8480
rect 20487 8449 20499 8452
rect 20441 8443 20499 8449
rect 20622 8440 20628 8452
rect 20680 8440 20686 8492
rect 21174 8440 21180 8492
rect 21232 8480 21238 8492
rect 21361 8483 21419 8489
rect 21361 8480 21373 8483
rect 21232 8452 21373 8480
rect 21232 8440 21238 8452
rect 21361 8449 21373 8452
rect 21407 8480 21419 8483
rect 23017 8483 23075 8489
rect 23017 8480 23029 8483
rect 21407 8452 23029 8480
rect 21407 8449 21419 8452
rect 21361 8443 21419 8449
rect 23017 8449 23029 8452
rect 23063 8449 23075 8483
rect 23017 8443 23075 8449
rect 24397 8483 24455 8489
rect 24397 8449 24409 8483
rect 24443 8480 24455 8483
rect 25406 8480 25412 8492
rect 24443 8452 25412 8480
rect 24443 8449 24455 8452
rect 24397 8443 24455 8449
rect 25406 8440 25412 8452
rect 25464 8480 25470 8492
rect 25685 8483 25743 8489
rect 25685 8480 25697 8483
rect 25464 8452 25697 8480
rect 25464 8440 25470 8452
rect 25685 8449 25697 8452
rect 25731 8449 25743 8483
rect 25685 8443 25743 8449
rect 13722 8412 13728 8424
rect 10367 8384 13728 8412
rect 10367 8381 10379 8384
rect 10321 8375 10379 8381
rect 13722 8372 13728 8384
rect 13780 8372 13786 8424
rect 16666 8412 16672 8424
rect 16627 8384 16672 8412
rect 16666 8372 16672 8384
rect 16724 8372 16730 8424
rect 16945 8415 17003 8421
rect 16945 8381 16957 8415
rect 16991 8412 17003 8415
rect 17862 8412 17868 8424
rect 16991 8384 17868 8412
rect 16991 8381 17003 8384
rect 16945 8375 17003 8381
rect 1581 8316 4154 8344
rect 5077 8347 5135 8353
rect 1581 8313 1593 8316
rect 1535 8307 1593 8313
rect 5077 8313 5089 8347
rect 5123 8344 5135 8347
rect 5350 8344 5356 8356
rect 5123 8316 5356 8344
rect 5123 8313 5135 8316
rect 5077 8307 5135 8313
rect 5350 8304 5356 8316
rect 5408 8304 5414 8356
rect 6270 8344 6276 8356
rect 6183 8316 6276 8344
rect 6270 8304 6276 8316
rect 6328 8344 6334 8356
rect 6328 8316 7420 8344
rect 6328 8304 6334 8316
rect 5442 8236 5448 8288
rect 5500 8276 5506 8288
rect 7282 8276 7288 8288
rect 5500 8248 7288 8276
rect 5500 8236 5506 8248
rect 7282 8236 7288 8248
rect 7340 8236 7346 8288
rect 7392 8276 7420 8316
rect 8018 8304 8024 8356
rect 8076 8344 8082 8356
rect 8434 8347 8492 8353
rect 8434 8344 8446 8347
rect 8076 8316 8446 8344
rect 8076 8304 8082 8316
rect 8434 8313 8446 8316
rect 8480 8313 8492 8347
rect 8434 8307 8492 8313
rect 8588 8316 12296 8344
rect 8588 8276 8616 8316
rect 9398 8276 9404 8288
rect 7392 8248 8616 8276
rect 9359 8248 9404 8276
rect 9398 8236 9404 8248
rect 9456 8236 9462 8288
rect 9490 8236 9496 8288
rect 9548 8276 9554 8288
rect 9766 8276 9772 8288
rect 9548 8248 9772 8276
rect 9548 8236 9554 8248
rect 9766 8236 9772 8248
rect 9824 8236 9830 8288
rect 10778 8236 10784 8288
rect 10836 8276 10842 8288
rect 11422 8276 11428 8288
rect 10836 8248 11428 8276
rect 10836 8236 10842 8248
rect 11422 8236 11428 8248
rect 11480 8236 11486 8288
rect 12158 8276 12164 8288
rect 12119 8248 12164 8276
rect 12158 8236 12164 8248
rect 12216 8236 12222 8288
rect 12268 8276 12296 8316
rect 12526 8304 12532 8356
rect 12584 8344 12590 8356
rect 12758 8347 12816 8353
rect 12758 8344 12770 8347
rect 12584 8316 12770 8344
rect 12584 8304 12590 8316
rect 12758 8313 12770 8316
rect 12804 8313 12816 8347
rect 12758 8307 12816 8313
rect 13998 8304 14004 8356
rect 14056 8344 14062 8356
rect 14369 8347 14427 8353
rect 14369 8344 14381 8347
rect 14056 8316 14381 8344
rect 14056 8304 14062 8316
rect 14369 8313 14381 8316
rect 14415 8313 14427 8347
rect 14369 8307 14427 8313
rect 16301 8347 16359 8353
rect 16301 8313 16313 8347
rect 16347 8344 16359 8347
rect 16482 8344 16488 8356
rect 16347 8316 16488 8344
rect 16347 8313 16359 8316
rect 16301 8307 16359 8313
rect 16482 8304 16488 8316
rect 16540 8344 16546 8356
rect 16960 8344 16988 8375
rect 17862 8372 17868 8384
rect 17920 8372 17926 8424
rect 22186 8372 22192 8424
rect 22244 8412 22250 8424
rect 22281 8415 22339 8421
rect 22281 8412 22293 8415
rect 22244 8384 22293 8412
rect 22244 8372 22250 8384
rect 22281 8381 22293 8384
rect 22327 8381 22339 8415
rect 22281 8375 22339 8381
rect 16540 8316 16988 8344
rect 17129 8347 17187 8353
rect 16540 8304 16546 8316
rect 17129 8313 17141 8347
rect 17175 8344 17187 8347
rect 17954 8344 17960 8356
rect 17175 8316 17960 8344
rect 17175 8313 17187 8316
rect 17129 8307 17187 8313
rect 17954 8304 17960 8316
rect 18012 8304 18018 8356
rect 18046 8304 18052 8356
rect 18104 8344 18110 8356
rect 18325 8347 18383 8353
rect 18325 8344 18337 8347
rect 18104 8316 18337 8344
rect 18104 8304 18110 8316
rect 18325 8313 18337 8316
rect 18371 8313 18383 8347
rect 18325 8307 18383 8313
rect 19426 8304 19432 8356
rect 19484 8344 19490 8356
rect 19613 8347 19671 8353
rect 19613 8344 19625 8347
rect 19484 8316 19625 8344
rect 19484 8304 19490 8316
rect 19613 8313 19625 8316
rect 19659 8344 19671 8347
rect 19889 8347 19947 8353
rect 19889 8344 19901 8347
rect 19659 8316 19901 8344
rect 19659 8313 19671 8316
rect 19613 8307 19671 8313
rect 19889 8313 19901 8316
rect 19935 8313 19947 8347
rect 21450 8344 21456 8356
rect 21363 8316 21456 8344
rect 19889 8307 19947 8313
rect 13354 8276 13360 8288
rect 12268 8248 13360 8276
rect 13354 8236 13360 8248
rect 13412 8236 13418 8288
rect 17589 8279 17647 8285
rect 17589 8245 17601 8279
rect 17635 8276 17647 8279
rect 17678 8276 17684 8288
rect 17635 8248 17684 8276
rect 17635 8245 17647 8248
rect 17589 8239 17647 8245
rect 17678 8236 17684 8248
rect 17736 8236 17742 8288
rect 18966 8236 18972 8288
rect 19024 8276 19030 8288
rect 19153 8279 19211 8285
rect 19153 8276 19165 8279
rect 19024 8248 19165 8276
rect 19024 8236 19030 8248
rect 19153 8245 19165 8248
rect 19199 8245 19211 8279
rect 19904 8276 19932 8307
rect 21450 8304 21456 8316
rect 21508 8344 21514 8356
rect 23658 8344 23664 8356
rect 21508 8316 22416 8344
rect 21508 8304 21514 8316
rect 21468 8276 21496 8304
rect 19904 8248 21496 8276
rect 22388 8276 22416 8316
rect 23446 8316 23664 8344
rect 23446 8276 23474 8316
rect 23658 8304 23664 8316
rect 23716 8304 23722 8356
rect 24489 8347 24547 8353
rect 24489 8313 24501 8347
rect 24535 8344 24547 8347
rect 24670 8344 24676 8356
rect 24535 8316 24676 8344
rect 24535 8313 24547 8316
rect 24489 8307 24547 8313
rect 24670 8304 24676 8316
rect 24728 8304 24734 8356
rect 22388 8248 23474 8276
rect 19153 8239 19211 8245
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 5350 8032 5356 8084
rect 5408 8072 5414 8084
rect 7006 8072 7012 8084
rect 5408 8044 7012 8072
rect 5408 8032 5414 8044
rect 7006 8032 7012 8044
rect 7064 8072 7070 8084
rect 7285 8075 7343 8081
rect 7285 8072 7297 8075
rect 7064 8044 7297 8072
rect 7064 8032 7070 8044
rect 7285 8041 7297 8044
rect 7331 8041 7343 8075
rect 7742 8072 7748 8084
rect 7703 8044 7748 8072
rect 7285 8035 7343 8041
rect 6178 7964 6184 8016
rect 6236 8004 6242 8016
rect 6457 8007 6515 8013
rect 6457 8004 6469 8007
rect 6236 7976 6469 8004
rect 6236 7964 6242 7976
rect 6457 7973 6469 7976
rect 6503 7973 6515 8007
rect 7300 8004 7328 8035
rect 7742 8032 7748 8044
rect 7800 8032 7806 8084
rect 9030 8072 9036 8084
rect 7944 8044 8892 8072
rect 8991 8044 9036 8072
rect 7944 8004 7972 8044
rect 7300 7976 7972 8004
rect 6457 7967 6515 7973
rect 8018 7964 8024 8016
rect 8076 8004 8082 8016
rect 8158 8007 8216 8013
rect 8158 8004 8170 8007
rect 8076 7976 8170 8004
rect 8076 7964 8082 7976
rect 8158 7973 8170 7976
rect 8204 7973 8216 8007
rect 8864 8004 8892 8044
rect 9030 8032 9036 8044
rect 9088 8032 9094 8084
rect 12434 8072 12440 8084
rect 9646 8044 12440 8072
rect 9646 8004 9674 8044
rect 12434 8032 12440 8044
rect 12492 8032 12498 8084
rect 12710 8072 12716 8084
rect 12671 8044 12716 8072
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 15378 8072 15384 8084
rect 15339 8044 15384 8072
rect 15378 8032 15384 8044
rect 15436 8032 15442 8084
rect 16482 8072 16488 8084
rect 16443 8044 16488 8072
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 18046 8072 18052 8084
rect 18007 8044 18052 8072
rect 18046 8032 18052 8044
rect 18104 8032 18110 8084
rect 18690 8072 18696 8084
rect 18651 8044 18696 8072
rect 18690 8032 18696 8044
rect 18748 8032 18754 8084
rect 19150 8072 19156 8084
rect 19111 8044 19156 8072
rect 19150 8032 19156 8044
rect 19208 8032 19214 8084
rect 21082 8032 21088 8084
rect 21140 8072 21146 8084
rect 23658 8072 23664 8084
rect 21140 8044 22876 8072
rect 23619 8044 23664 8072
rect 21140 8032 21146 8044
rect 8864 7976 9674 8004
rect 11879 8007 11937 8013
rect 8158 7967 8216 7973
rect 11879 7973 11891 8007
rect 11925 8004 11937 8007
rect 12158 8004 12164 8016
rect 11925 7976 12164 8004
rect 11925 7973 11937 7976
rect 11879 7967 11937 7973
rect 12158 7964 12164 7976
rect 12216 7964 12222 8016
rect 13354 7964 13360 8016
rect 13412 8004 13418 8016
rect 13817 8007 13875 8013
rect 13817 8004 13829 8007
rect 13412 7976 13829 8004
rect 13412 7964 13418 7976
rect 13817 7973 13829 7976
rect 13863 7973 13875 8007
rect 21174 8004 21180 8016
rect 13817 7967 13875 7973
rect 15304 7976 16988 8004
rect 15304 7948 15332 7976
rect 5166 7896 5172 7948
rect 5224 7936 5230 7948
rect 5296 7939 5354 7945
rect 5296 7936 5308 7939
rect 5224 7908 5308 7936
rect 5224 7896 5230 7908
rect 5296 7905 5308 7908
rect 5342 7905 5354 7939
rect 5296 7899 5354 7905
rect 7837 7939 7895 7945
rect 7837 7905 7849 7939
rect 7883 7936 7895 7939
rect 7926 7936 7932 7948
rect 7883 7908 7932 7936
rect 7883 7905 7895 7908
rect 7837 7899 7895 7905
rect 7926 7896 7932 7908
rect 7984 7936 7990 7948
rect 8754 7936 8760 7948
rect 7984 7908 8760 7936
rect 7984 7896 7990 7908
rect 8754 7896 8760 7908
rect 8812 7896 8818 7948
rect 9950 7936 9956 7948
rect 9416 7908 9956 7936
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7868 4307 7871
rect 6365 7871 6423 7877
rect 6365 7868 6377 7871
rect 4295 7840 6377 7868
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 6365 7837 6377 7840
rect 6411 7868 6423 7871
rect 6546 7868 6552 7880
rect 6411 7840 6552 7868
rect 6411 7837 6423 7840
rect 6365 7831 6423 7837
rect 6546 7828 6552 7840
rect 6604 7828 6610 7880
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7868 7067 7871
rect 7374 7868 7380 7880
rect 7055 7840 7380 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 7374 7828 7380 7840
rect 7432 7828 7438 7880
rect 5399 7735 5457 7741
rect 5399 7701 5411 7735
rect 5445 7732 5457 7735
rect 6089 7735 6147 7741
rect 6089 7732 6101 7735
rect 5445 7704 6101 7732
rect 5445 7701 5457 7704
rect 5399 7695 5457 7701
rect 6089 7701 6101 7704
rect 6135 7732 6147 7735
rect 6638 7732 6644 7744
rect 6135 7704 6644 7732
rect 6135 7701 6147 7704
rect 6089 7695 6147 7701
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 8754 7732 8760 7744
rect 8715 7704 8760 7732
rect 8754 7692 8760 7704
rect 8812 7692 8818 7744
rect 9306 7692 9312 7744
rect 9364 7732 9370 7744
rect 9416 7741 9444 7908
rect 9950 7896 9956 7908
rect 10008 7896 10014 7948
rect 10134 7896 10140 7948
rect 10192 7936 10198 7948
rect 10413 7939 10471 7945
rect 10413 7936 10425 7939
rect 10192 7908 10425 7936
rect 10192 7896 10198 7908
rect 10413 7905 10425 7908
rect 10459 7905 10471 7939
rect 15286 7936 15292 7948
rect 15247 7908 15292 7936
rect 10413 7899 10471 7905
rect 15286 7896 15292 7908
rect 15344 7896 15350 7948
rect 15746 7936 15752 7948
rect 15707 7908 15752 7936
rect 15746 7896 15752 7908
rect 15804 7896 15810 7948
rect 16960 7945 16988 7976
rect 19812 7976 21180 8004
rect 19812 7948 19840 7976
rect 21174 7964 21180 7976
rect 21232 7964 21238 8016
rect 21269 8007 21327 8013
rect 21269 7973 21281 8007
rect 21315 8004 21327 8007
rect 21450 8004 21456 8016
rect 21315 7976 21456 8004
rect 21315 7973 21327 7976
rect 21269 7967 21327 7973
rect 21450 7964 21456 7976
rect 21508 7964 21514 8016
rect 22848 8013 22876 8044
rect 23658 8032 23664 8044
rect 23716 8032 23722 8084
rect 22833 8007 22891 8013
rect 22833 7973 22845 8007
rect 22879 8004 22891 8007
rect 23382 8004 23388 8016
rect 22879 7976 23388 8004
rect 22879 7973 22891 7976
rect 22833 7967 22891 7973
rect 23382 7964 23388 7976
rect 23440 7964 23446 8016
rect 23474 7964 23480 8016
rect 23532 8004 23538 8016
rect 24397 8007 24455 8013
rect 24397 8004 24409 8007
rect 23532 7976 24409 8004
rect 23532 7964 23538 7976
rect 24397 7973 24409 7976
rect 24443 8004 24455 8007
rect 24670 8004 24676 8016
rect 24443 7976 24676 8004
rect 24443 7973 24455 7976
rect 24397 7967 24455 7973
rect 24670 7964 24676 7976
rect 24728 7964 24734 8016
rect 24946 8004 24952 8016
rect 24907 7976 24952 8004
rect 24946 7964 24952 7976
rect 25004 7964 25010 8016
rect 16945 7939 17003 7945
rect 16945 7905 16957 7939
rect 16991 7936 17003 7939
rect 17126 7936 17132 7948
rect 16991 7908 17132 7936
rect 16991 7905 17003 7908
rect 16945 7899 17003 7905
rect 17126 7896 17132 7908
rect 17184 7936 17190 7948
rect 17402 7936 17408 7948
rect 17184 7908 17408 7936
rect 17184 7896 17190 7908
rect 17402 7896 17408 7908
rect 17460 7896 17466 7948
rect 17497 7939 17555 7945
rect 17497 7905 17509 7939
rect 17543 7936 17555 7939
rect 17862 7936 17868 7948
rect 17543 7908 17868 7936
rect 17543 7905 17555 7908
rect 17497 7899 17555 7905
rect 17862 7896 17868 7908
rect 17920 7896 17926 7948
rect 19242 7936 19248 7948
rect 19203 7908 19248 7936
rect 19242 7896 19248 7908
rect 19300 7896 19306 7948
rect 19794 7936 19800 7948
rect 19707 7908 19800 7936
rect 19794 7896 19800 7908
rect 19852 7896 19858 7948
rect 10689 7871 10747 7877
rect 10689 7837 10701 7871
rect 10735 7868 10747 7871
rect 11517 7871 11575 7877
rect 11517 7868 11529 7871
rect 10735 7840 11529 7868
rect 10735 7837 10747 7840
rect 10689 7831 10747 7837
rect 11517 7837 11529 7840
rect 11563 7868 11575 7871
rect 11882 7868 11888 7880
rect 11563 7840 11888 7868
rect 11563 7837 11575 7840
rect 11517 7831 11575 7837
rect 11882 7828 11888 7840
rect 11940 7828 11946 7880
rect 13541 7871 13599 7877
rect 13541 7837 13553 7871
rect 13587 7868 13599 7871
rect 13722 7868 13728 7880
rect 13587 7840 13728 7868
rect 13587 7837 13599 7840
rect 13541 7831 13599 7837
rect 13722 7828 13728 7840
rect 13780 7828 13786 7880
rect 17586 7868 17592 7880
rect 17547 7840 17592 7868
rect 17586 7828 17592 7840
rect 17644 7828 17650 7880
rect 19978 7868 19984 7880
rect 19939 7840 19984 7868
rect 19978 7828 19984 7840
rect 20036 7828 20042 7880
rect 21174 7868 21180 7880
rect 21135 7840 21180 7868
rect 21174 7828 21180 7840
rect 21232 7828 21238 7880
rect 21453 7871 21511 7877
rect 21453 7837 21465 7871
rect 21499 7837 21511 7871
rect 21453 7831 21511 7837
rect 22741 7871 22799 7877
rect 22741 7837 22753 7871
rect 22787 7868 22799 7871
rect 23106 7868 23112 7880
rect 22787 7840 23112 7868
rect 22787 7837 22799 7840
rect 22741 7831 22799 7837
rect 14274 7800 14280 7812
rect 14235 7772 14280 7800
rect 14274 7760 14280 7772
rect 14332 7760 14338 7812
rect 14642 7760 14648 7812
rect 14700 7800 14706 7812
rect 16666 7800 16672 7812
rect 14700 7772 16672 7800
rect 14700 7760 14706 7772
rect 16666 7760 16672 7772
rect 16724 7800 16730 7812
rect 16761 7803 16819 7809
rect 16761 7800 16773 7803
rect 16724 7772 16773 7800
rect 16724 7760 16730 7772
rect 16761 7769 16773 7772
rect 16807 7769 16819 7803
rect 16761 7763 16819 7769
rect 20254 7760 20260 7812
rect 20312 7800 20318 7812
rect 20898 7800 20904 7812
rect 20312 7772 20904 7800
rect 20312 7760 20318 7772
rect 20898 7760 20904 7772
rect 20956 7800 20962 7812
rect 21468 7800 21496 7831
rect 23106 7828 23112 7840
rect 23164 7828 23170 7880
rect 24305 7871 24363 7877
rect 24305 7837 24317 7871
rect 24351 7868 24363 7871
rect 25038 7868 25044 7880
rect 24351 7840 25044 7868
rect 24351 7837 24363 7840
rect 24305 7831 24363 7837
rect 25038 7828 25044 7840
rect 25096 7828 25102 7880
rect 20956 7772 21496 7800
rect 23293 7803 23351 7809
rect 20956 7760 20962 7772
rect 23293 7769 23305 7803
rect 23339 7769 23351 7803
rect 23293 7763 23351 7769
rect 9401 7735 9459 7741
rect 9401 7732 9413 7735
rect 9364 7704 9413 7732
rect 9364 7692 9370 7704
rect 9401 7701 9413 7704
rect 9447 7701 9459 7735
rect 9401 7695 9459 7701
rect 18417 7735 18475 7741
rect 18417 7701 18429 7735
rect 18463 7732 18475 7735
rect 18506 7732 18512 7744
rect 18463 7704 18512 7732
rect 18463 7701 18475 7704
rect 18417 7695 18475 7701
rect 18506 7692 18512 7704
rect 18564 7692 18570 7744
rect 22094 7732 22100 7744
rect 22055 7704 22100 7732
rect 22094 7692 22100 7704
rect 22152 7692 22158 7744
rect 22738 7692 22744 7744
rect 22796 7732 22802 7744
rect 23308 7732 23336 7763
rect 24118 7732 24124 7744
rect 22796 7704 23336 7732
rect 24079 7704 24124 7732
rect 22796 7692 22802 7704
rect 24118 7692 24124 7704
rect 24176 7692 24182 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1394 7488 1400 7540
rect 1452 7528 1458 7540
rect 4154 7528 4160 7540
rect 1452 7500 4160 7528
rect 1452 7488 1458 7500
rect 4154 7488 4160 7500
rect 4212 7488 4218 7540
rect 5166 7528 5172 7540
rect 4540 7500 5172 7528
rect 3786 7420 3792 7472
rect 3844 7460 3850 7472
rect 4540 7460 4568 7500
rect 5166 7488 5172 7500
rect 5224 7528 5230 7540
rect 5261 7531 5319 7537
rect 5261 7528 5273 7531
rect 5224 7500 5273 7528
rect 5224 7488 5230 7500
rect 5261 7497 5273 7500
rect 5307 7497 5319 7531
rect 5261 7491 5319 7497
rect 5350 7488 5356 7540
rect 5408 7528 5414 7540
rect 5534 7528 5540 7540
rect 5408 7500 5540 7528
rect 5408 7488 5414 7500
rect 5534 7488 5540 7500
rect 5592 7488 5598 7540
rect 6546 7528 6552 7540
rect 6507 7500 6552 7528
rect 6546 7488 6552 7500
rect 6604 7488 6610 7540
rect 7929 7531 7987 7537
rect 7929 7497 7941 7531
rect 7975 7528 7987 7531
rect 8018 7528 8024 7540
rect 7975 7500 8024 7528
rect 7975 7497 7987 7500
rect 7929 7491 7987 7497
rect 8018 7488 8024 7500
rect 8076 7488 8082 7540
rect 11882 7528 11888 7540
rect 11843 7500 11888 7528
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 12434 7488 12440 7540
rect 12492 7528 12498 7540
rect 13541 7531 13599 7537
rect 13541 7528 13553 7531
rect 12492 7500 13553 7528
rect 12492 7488 12498 7500
rect 13541 7497 13553 7500
rect 13587 7528 13599 7531
rect 13633 7531 13691 7537
rect 13633 7528 13645 7531
rect 13587 7500 13645 7528
rect 13587 7497 13599 7500
rect 13541 7491 13599 7497
rect 13633 7497 13645 7500
rect 13679 7497 13691 7531
rect 13633 7491 13691 7497
rect 13722 7488 13728 7540
rect 13780 7528 13786 7540
rect 15519 7531 15577 7537
rect 15519 7528 15531 7531
rect 13780 7500 15531 7528
rect 13780 7488 13786 7500
rect 15519 7497 15531 7500
rect 15565 7497 15577 7531
rect 17402 7528 17408 7540
rect 17363 7500 17408 7528
rect 15519 7491 15577 7497
rect 17402 7488 17408 7500
rect 17460 7488 17466 7540
rect 17862 7528 17868 7540
rect 17775 7500 17868 7528
rect 17862 7488 17868 7500
rect 17920 7528 17926 7540
rect 19794 7528 19800 7540
rect 17920 7500 19800 7528
rect 17920 7488 17926 7500
rect 19794 7488 19800 7500
rect 19852 7488 19858 7540
rect 23382 7528 23388 7540
rect 23343 7500 23388 7528
rect 23382 7488 23388 7500
rect 23440 7488 23446 7540
rect 24118 7488 24124 7540
rect 24176 7528 24182 7540
rect 25363 7531 25421 7537
rect 25363 7528 25375 7531
rect 24176 7500 25375 7528
rect 24176 7488 24182 7500
rect 25363 7497 25375 7500
rect 25409 7497 25421 7531
rect 25363 7491 25421 7497
rect 3844 7432 4568 7460
rect 4617 7463 4675 7469
rect 3844 7420 3850 7432
rect 4617 7429 4629 7463
rect 4663 7460 4675 7463
rect 11974 7460 11980 7472
rect 4663 7432 11980 7460
rect 4663 7429 4675 7432
rect 4617 7423 4675 7429
rect 4724 7333 4752 7432
rect 11974 7420 11980 7432
rect 12032 7420 12038 7472
rect 14826 7460 14832 7472
rect 14787 7432 14832 7460
rect 14826 7420 14832 7432
rect 14884 7420 14890 7472
rect 15838 7420 15844 7472
rect 15896 7460 15902 7472
rect 20990 7460 20996 7472
rect 15896 7432 20996 7460
rect 15896 7420 15902 7432
rect 20990 7420 20996 7432
rect 21048 7420 21054 7472
rect 6638 7352 6644 7404
rect 6696 7392 6702 7404
rect 6917 7395 6975 7401
rect 6917 7392 6929 7395
rect 6696 7364 6929 7392
rect 6696 7352 6702 7364
rect 6917 7361 6929 7364
rect 6963 7361 6975 7395
rect 6917 7355 6975 7361
rect 8662 7352 8668 7404
rect 8720 7392 8726 7404
rect 8757 7395 8815 7401
rect 8757 7392 8769 7395
rect 8720 7364 8769 7392
rect 8720 7352 8726 7364
rect 8757 7361 8769 7364
rect 8803 7361 8815 7395
rect 10965 7395 11023 7401
rect 10965 7392 10977 7395
rect 8757 7355 8815 7361
rect 9968 7364 10977 7392
rect 4709 7327 4767 7333
rect 4709 7293 4721 7327
rect 4755 7293 4767 7327
rect 4709 7287 4767 7293
rect 5534 7284 5540 7336
rect 5592 7324 5598 7336
rect 5788 7327 5846 7333
rect 5788 7324 5800 7327
rect 5592 7296 5800 7324
rect 5592 7284 5598 7296
rect 5788 7293 5800 7296
rect 5834 7324 5846 7327
rect 6273 7327 6331 7333
rect 6273 7324 6285 7327
rect 5834 7296 6285 7324
rect 5834 7293 5846 7296
rect 5788 7287 5846 7293
rect 6273 7293 6285 7296
rect 6319 7324 6331 7327
rect 6730 7324 6736 7336
rect 6319 7296 6736 7324
rect 6319 7293 6331 7296
rect 6273 7287 6331 7293
rect 6730 7284 6736 7296
rect 6788 7284 6794 7336
rect 9306 7284 9312 7336
rect 9364 7324 9370 7336
rect 9968 7333 9996 7364
rect 10965 7361 10977 7364
rect 11011 7361 11023 7395
rect 14274 7392 14280 7404
rect 14235 7364 14280 7392
rect 10965 7355 11023 7361
rect 14274 7352 14280 7364
rect 14332 7352 14338 7404
rect 16301 7395 16359 7401
rect 16301 7361 16313 7395
rect 16347 7392 16359 7395
rect 16942 7392 16948 7404
rect 16347 7364 16948 7392
rect 16347 7361 16359 7364
rect 16301 7355 16359 7361
rect 9953 7327 10011 7333
rect 9953 7324 9965 7327
rect 9364 7296 9965 7324
rect 9364 7284 9370 7296
rect 9953 7293 9965 7296
rect 9999 7293 10011 7327
rect 9953 7287 10011 7293
rect 10413 7327 10471 7333
rect 10413 7293 10425 7327
rect 10459 7293 10471 7327
rect 10413 7287 10471 7293
rect 12856 7327 12914 7333
rect 12856 7293 12868 7327
rect 12902 7324 12914 7327
rect 13354 7324 13360 7336
rect 12902 7296 13360 7324
rect 12902 7293 12914 7296
rect 12856 7287 12914 7293
rect 4908 7228 6960 7256
rect 4908 7197 4936 7228
rect 4893 7191 4951 7197
rect 4893 7157 4905 7191
rect 4939 7157 4951 7191
rect 4893 7151 4951 7157
rect 5859 7191 5917 7197
rect 5859 7157 5871 7191
rect 5905 7188 5917 7191
rect 6086 7188 6092 7200
rect 5905 7160 6092 7188
rect 5905 7157 5917 7160
rect 5859 7151 5917 7157
rect 6086 7148 6092 7160
rect 6144 7148 6150 7200
rect 6932 7188 6960 7228
rect 7006 7216 7012 7268
rect 7064 7256 7070 7268
rect 7064 7228 7109 7256
rect 7064 7216 7070 7228
rect 7374 7216 7380 7268
rect 7432 7256 7438 7268
rect 7561 7259 7619 7265
rect 7561 7256 7573 7259
rect 7432 7228 7573 7256
rect 7432 7216 7438 7228
rect 7561 7225 7573 7228
rect 7607 7256 7619 7259
rect 8478 7256 8484 7268
rect 7607 7228 8484 7256
rect 7607 7225 7619 7228
rect 7561 7219 7619 7225
rect 8478 7216 8484 7228
rect 8536 7216 8542 7268
rect 8573 7259 8631 7265
rect 8573 7225 8585 7259
rect 8619 7256 8631 7259
rect 8754 7256 8760 7268
rect 8619 7228 8760 7256
rect 8619 7225 8631 7228
rect 8573 7219 8631 7225
rect 8110 7188 8116 7200
rect 6932 7160 8116 7188
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 8297 7191 8355 7197
rect 8297 7157 8309 7191
rect 8343 7188 8355 7191
rect 8588 7188 8616 7219
rect 8754 7216 8760 7228
rect 8812 7216 8818 7268
rect 10428 7256 10456 7287
rect 13354 7284 13360 7296
rect 13412 7284 13418 7336
rect 15448 7327 15506 7333
rect 15448 7293 15460 7327
rect 15494 7324 15506 7327
rect 15838 7324 15844 7336
rect 15494 7296 15844 7324
rect 15494 7293 15506 7296
rect 15448 7287 15506 7293
rect 15838 7284 15844 7296
rect 15896 7284 15902 7336
rect 16684 7333 16712 7364
rect 16942 7352 16948 7364
rect 17000 7352 17006 7404
rect 18417 7395 18475 7401
rect 18417 7361 18429 7395
rect 18463 7392 18475 7395
rect 19150 7392 19156 7404
rect 18463 7364 19156 7392
rect 18463 7361 18475 7364
rect 18417 7355 18475 7361
rect 19150 7352 19156 7364
rect 19208 7352 19214 7404
rect 20254 7392 20260 7404
rect 19812 7364 20260 7392
rect 16669 7327 16727 7333
rect 16669 7293 16681 7327
rect 16715 7293 16727 7327
rect 16850 7324 16856 7336
rect 16763 7296 16856 7324
rect 16669 7287 16727 7293
rect 16850 7284 16856 7296
rect 16908 7324 16914 7336
rect 17862 7324 17868 7336
rect 16908 7296 17868 7324
rect 16908 7284 16914 7296
rect 17862 7284 17868 7296
rect 17920 7284 17926 7336
rect 19061 7327 19119 7333
rect 19061 7293 19073 7327
rect 19107 7324 19119 7327
rect 19812 7324 19840 7364
rect 20254 7352 20260 7364
rect 20312 7392 20318 7404
rect 20717 7395 20775 7401
rect 20717 7392 20729 7395
rect 20312 7364 20729 7392
rect 20312 7352 20318 7364
rect 20717 7361 20729 7364
rect 20763 7361 20775 7395
rect 20717 7355 20775 7361
rect 23753 7395 23811 7401
rect 23753 7361 23765 7395
rect 23799 7392 23811 7395
rect 24136 7392 24164 7488
rect 24670 7460 24676 7472
rect 24631 7432 24676 7460
rect 24670 7420 24676 7432
rect 24728 7420 24734 7472
rect 25038 7460 25044 7472
rect 24999 7432 25044 7460
rect 25038 7420 25044 7432
rect 25096 7420 25102 7472
rect 23799 7364 24164 7392
rect 24397 7395 24455 7401
rect 23799 7361 23811 7364
rect 23753 7355 23811 7361
rect 24397 7361 24409 7395
rect 24443 7392 24455 7395
rect 24946 7392 24952 7404
rect 24443 7364 24952 7392
rect 24443 7361 24455 7364
rect 24397 7355 24455 7361
rect 24946 7352 24952 7364
rect 25004 7352 25010 7404
rect 19107 7296 19840 7324
rect 25292 7327 25350 7333
rect 19107 7293 19119 7296
rect 19061 7287 19119 7293
rect 25292 7293 25304 7327
rect 25338 7324 25350 7327
rect 25338 7296 25820 7324
rect 25338 7293 25350 7296
rect 25292 7287 25350 7293
rect 10686 7256 10692 7268
rect 9416 7228 10456 7256
rect 10647 7228 10692 7256
rect 8343 7160 8616 7188
rect 8343 7157 8355 7160
rect 8297 7151 8355 7157
rect 8846 7148 8852 7200
rect 8904 7188 8910 7200
rect 9416 7197 9444 7228
rect 10686 7216 10692 7228
rect 10744 7216 10750 7268
rect 12943 7259 13001 7265
rect 12943 7225 12955 7259
rect 12989 7256 13001 7259
rect 13906 7256 13912 7268
rect 12989 7228 13912 7256
rect 12989 7225 13001 7228
rect 12943 7219 13001 7225
rect 13906 7216 13912 7228
rect 13964 7216 13970 7268
rect 14001 7259 14059 7265
rect 14001 7225 14013 7259
rect 14047 7225 14059 7259
rect 14001 7219 14059 7225
rect 17129 7259 17187 7265
rect 17129 7225 17141 7259
rect 17175 7256 17187 7259
rect 18414 7256 18420 7268
rect 17175 7228 18420 7256
rect 17175 7225 17187 7228
rect 17129 7219 17187 7225
rect 9401 7191 9459 7197
rect 9401 7188 9413 7191
rect 8904 7160 9413 7188
rect 8904 7148 8910 7160
rect 9401 7157 9413 7160
rect 9447 7157 9459 7191
rect 9401 7151 9459 7157
rect 9861 7191 9919 7197
rect 9861 7157 9873 7191
rect 9907 7188 9919 7191
rect 10134 7188 10140 7200
rect 9907 7160 10140 7188
rect 9907 7157 9919 7160
rect 9861 7151 9919 7157
rect 10134 7148 10140 7160
rect 10192 7148 10198 7200
rect 11609 7191 11667 7197
rect 11609 7157 11621 7191
rect 11655 7188 11667 7191
rect 12158 7188 12164 7200
rect 11655 7160 12164 7188
rect 11655 7157 11667 7160
rect 11609 7151 11667 7157
rect 12158 7148 12164 7160
rect 12216 7188 12222 7200
rect 12710 7188 12716 7200
rect 12216 7160 12716 7188
rect 12216 7148 12222 7160
rect 12710 7148 12716 7160
rect 12768 7148 12774 7200
rect 13354 7188 13360 7200
rect 13315 7160 13360 7188
rect 13354 7148 13360 7160
rect 13412 7148 13418 7200
rect 13541 7191 13599 7197
rect 13541 7157 13553 7191
rect 13587 7188 13599 7191
rect 14016 7188 14044 7219
rect 18414 7216 18420 7228
rect 18472 7216 18478 7268
rect 18506 7216 18512 7268
rect 18564 7256 18570 7268
rect 18564 7228 18609 7256
rect 18564 7216 18570 7228
rect 19242 7216 19248 7268
rect 19300 7256 19306 7268
rect 19337 7259 19395 7265
rect 19337 7256 19349 7259
rect 19300 7228 19349 7256
rect 19300 7216 19306 7228
rect 19337 7225 19349 7228
rect 19383 7225 19395 7259
rect 20438 7256 20444 7268
rect 20399 7228 20444 7256
rect 19337 7219 19395 7225
rect 20438 7216 20444 7228
rect 20496 7216 20502 7268
rect 20533 7259 20591 7265
rect 20533 7225 20545 7259
rect 20579 7225 20591 7259
rect 20533 7219 20591 7225
rect 13587 7160 14044 7188
rect 13587 7157 13599 7160
rect 13541 7151 13599 7157
rect 14826 7148 14832 7200
rect 14884 7188 14890 7200
rect 15197 7191 15255 7197
rect 15197 7188 15209 7191
rect 14884 7160 15209 7188
rect 14884 7148 14890 7160
rect 15197 7157 15209 7160
rect 15243 7188 15255 7191
rect 15286 7188 15292 7200
rect 15243 7160 15292 7188
rect 15243 7157 15255 7160
rect 15197 7151 15255 7157
rect 15286 7148 15292 7160
rect 15344 7148 15350 7200
rect 20257 7191 20315 7197
rect 20257 7157 20269 7191
rect 20303 7188 20315 7191
rect 20548 7188 20576 7219
rect 21634 7216 21640 7268
rect 21692 7256 21698 7268
rect 22094 7256 22100 7268
rect 21692 7228 22100 7256
rect 21692 7216 21698 7228
rect 22094 7216 22100 7228
rect 22152 7216 22158 7268
rect 22189 7259 22247 7265
rect 22189 7225 22201 7259
rect 22235 7225 22247 7259
rect 22738 7256 22744 7268
rect 22699 7228 22744 7256
rect 22189 7219 22247 7225
rect 21082 7188 21088 7200
rect 20303 7160 21088 7188
rect 20303 7157 20315 7160
rect 20257 7151 20315 7157
rect 21082 7148 21088 7160
rect 21140 7148 21146 7200
rect 21450 7188 21456 7200
rect 21411 7160 21456 7188
rect 21450 7148 21456 7160
rect 21508 7148 21514 7200
rect 21726 7148 21732 7200
rect 21784 7188 21790 7200
rect 21821 7191 21879 7197
rect 21821 7188 21833 7191
rect 21784 7160 21833 7188
rect 21784 7148 21790 7160
rect 21821 7157 21833 7160
rect 21867 7188 21879 7191
rect 22204 7188 22232 7219
rect 22738 7216 22744 7228
rect 22796 7216 22802 7268
rect 23845 7259 23903 7265
rect 23845 7225 23857 7259
rect 23891 7225 23903 7259
rect 23845 7219 23903 7225
rect 23106 7188 23112 7200
rect 21867 7160 22232 7188
rect 23067 7160 23112 7188
rect 21867 7157 21879 7160
rect 21821 7151 21879 7157
rect 23106 7148 23112 7160
rect 23164 7148 23170 7200
rect 23658 7148 23664 7200
rect 23716 7188 23722 7200
rect 23860 7188 23888 7219
rect 25792 7197 25820 7296
rect 23716 7160 23888 7188
rect 25777 7191 25835 7197
rect 23716 7148 23722 7160
rect 25777 7157 25789 7191
rect 25823 7188 25835 7191
rect 25958 7188 25964 7200
rect 25823 7160 25964 7188
rect 25823 7157 25835 7160
rect 25777 7151 25835 7157
rect 25958 7148 25964 7160
rect 26016 7148 26022 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 658 6944 664 6996
rect 716 6984 722 6996
rect 5534 6984 5540 6996
rect 716 6956 5540 6984
rect 716 6944 722 6956
rect 5534 6944 5540 6956
rect 5592 6944 5598 6996
rect 6270 6984 6276 6996
rect 6231 6956 6276 6984
rect 6270 6944 6276 6956
rect 6328 6944 6334 6996
rect 8205 6987 8263 6993
rect 8205 6984 8217 6987
rect 6748 6956 8217 6984
rect 4617 6919 4675 6925
rect 4617 6885 4629 6919
rect 4663 6916 4675 6919
rect 5442 6916 5448 6928
rect 4663 6888 5448 6916
rect 4663 6885 4675 6888
rect 4617 6879 4675 6885
rect 4132 6851 4190 6857
rect 4132 6817 4144 6851
rect 4178 6848 4190 6851
rect 4706 6848 4712 6860
rect 4178 6820 4712 6848
rect 4178 6817 4190 6820
rect 4132 6811 4190 6817
rect 4706 6808 4712 6820
rect 4764 6808 4770 6860
rect 5092 6857 5120 6888
rect 5442 6876 5448 6888
rect 5500 6876 5506 6928
rect 6086 6876 6092 6928
rect 6144 6916 6150 6928
rect 6748 6925 6776 6956
rect 8205 6953 8217 6956
rect 8251 6953 8263 6987
rect 8205 6947 8263 6953
rect 8478 6944 8484 6996
rect 8536 6984 8542 6996
rect 10873 6987 10931 6993
rect 10873 6984 10885 6987
rect 8536 6956 10885 6984
rect 8536 6944 8542 6956
rect 10873 6953 10885 6956
rect 10919 6953 10931 6987
rect 11974 6984 11980 6996
rect 11935 6956 11980 6984
rect 10873 6947 10931 6953
rect 11974 6944 11980 6956
rect 12032 6944 12038 6996
rect 13446 6984 13452 6996
rect 13407 6956 13452 6984
rect 13446 6944 13452 6956
rect 13504 6944 13510 6996
rect 13906 6944 13912 6996
rect 13964 6984 13970 6996
rect 14645 6987 14703 6993
rect 14645 6984 14657 6987
rect 13964 6956 14657 6984
rect 13964 6944 13970 6956
rect 14645 6953 14657 6956
rect 14691 6953 14703 6987
rect 14645 6947 14703 6953
rect 14734 6944 14740 6996
rect 14792 6984 14798 6996
rect 15378 6984 15384 6996
rect 14792 6956 15384 6984
rect 14792 6944 14798 6956
rect 15378 6944 15384 6956
rect 15436 6984 15442 6996
rect 15473 6987 15531 6993
rect 15473 6984 15485 6987
rect 15436 6956 15485 6984
rect 15436 6944 15442 6956
rect 15473 6953 15485 6956
rect 15519 6953 15531 6987
rect 15473 6947 15531 6953
rect 17494 6944 17500 6996
rect 17552 6984 17558 6996
rect 19475 6987 19533 6993
rect 19475 6984 19487 6987
rect 17552 6956 19487 6984
rect 17552 6944 17558 6956
rect 19475 6953 19487 6956
rect 19521 6953 19533 6987
rect 21174 6984 21180 6996
rect 21135 6956 21180 6984
rect 19475 6947 19533 6953
rect 21174 6944 21180 6956
rect 21232 6944 21238 6996
rect 21450 6944 21456 6996
rect 21508 6984 21514 6996
rect 22741 6987 22799 6993
rect 22741 6984 22753 6987
rect 21508 6956 22753 6984
rect 21508 6944 21514 6956
rect 22741 6953 22753 6956
rect 22787 6953 22799 6987
rect 22741 6947 22799 6953
rect 23474 6944 23480 6996
rect 23532 6984 23538 6996
rect 23532 6956 25335 6984
rect 23532 6944 23538 6956
rect 6733 6919 6791 6925
rect 6733 6916 6745 6919
rect 6144 6888 6745 6916
rect 6144 6876 6150 6888
rect 6733 6885 6745 6888
rect 6779 6885 6791 6919
rect 6733 6879 6791 6885
rect 6825 6919 6883 6925
rect 6825 6885 6837 6919
rect 6871 6916 6883 6919
rect 7006 6916 7012 6928
rect 6871 6888 7012 6916
rect 6871 6885 6883 6888
rect 6825 6879 6883 6885
rect 7006 6876 7012 6888
rect 7064 6876 7070 6928
rect 7374 6916 7380 6928
rect 7335 6888 7380 6916
rect 7374 6876 7380 6888
rect 7432 6876 7438 6928
rect 7926 6916 7932 6928
rect 7887 6888 7932 6916
rect 7926 6876 7932 6888
rect 7984 6876 7990 6928
rect 8110 6876 8116 6928
rect 8168 6916 8174 6928
rect 9923 6919 9981 6925
rect 8168 6888 9720 6916
rect 8168 6876 8174 6888
rect 5077 6851 5135 6857
rect 5077 6817 5089 6851
rect 5123 6817 5135 6851
rect 5077 6811 5135 6817
rect 5353 6851 5411 6857
rect 5353 6817 5365 6851
rect 5399 6848 5411 6851
rect 5534 6848 5540 6860
rect 5399 6820 5540 6848
rect 5399 6817 5411 6820
rect 5353 6811 5411 6817
rect 4985 6783 5043 6789
rect 4985 6749 4997 6783
rect 5031 6780 5043 6783
rect 5368 6780 5396 6811
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 8573 6851 8631 6857
rect 8573 6817 8585 6851
rect 8619 6817 8631 6851
rect 9692 6848 9720 6888
rect 9923 6885 9935 6919
rect 9969 6916 9981 6919
rect 10042 6916 10048 6928
rect 9969 6888 10048 6916
rect 9969 6885 9981 6888
rect 9923 6879 9981 6885
rect 10042 6876 10048 6888
rect 10100 6876 10106 6928
rect 11422 6876 11428 6928
rect 11480 6916 11486 6928
rect 11480 6888 11560 6916
rect 11480 6876 11486 6888
rect 11532 6857 11560 6888
rect 13538 6876 13544 6928
rect 13596 6916 13602 6928
rect 13817 6919 13875 6925
rect 13817 6916 13829 6919
rect 13596 6888 13829 6916
rect 13596 6876 13602 6888
rect 13817 6885 13829 6888
rect 13863 6885 13875 6919
rect 13817 6879 13875 6885
rect 17678 6876 17684 6928
rect 17736 6916 17742 6928
rect 17910 6919 17968 6925
rect 17910 6916 17922 6919
rect 17736 6888 17922 6916
rect 17736 6876 17742 6888
rect 17910 6885 17922 6888
rect 17956 6916 17968 6919
rect 18785 6919 18843 6925
rect 18785 6916 18797 6919
rect 17956 6888 18797 6916
rect 17956 6885 17968 6888
rect 17910 6879 17968 6885
rect 18785 6885 18797 6888
rect 18831 6916 18843 6919
rect 18966 6916 18972 6928
rect 18831 6888 18972 6916
rect 18831 6885 18843 6888
rect 18785 6879 18843 6885
rect 18966 6876 18972 6888
rect 19024 6916 19030 6928
rect 19797 6919 19855 6925
rect 19797 6916 19809 6919
rect 19024 6888 19809 6916
rect 19024 6876 19030 6888
rect 19797 6885 19809 6888
rect 19843 6885 19855 6919
rect 22094 6916 22100 6928
rect 22055 6888 22100 6916
rect 19797 6879 19855 6885
rect 22094 6876 22100 6888
rect 22152 6876 22158 6928
rect 23842 6916 23848 6928
rect 23803 6888 23848 6916
rect 23842 6876 23848 6888
rect 23900 6876 23906 6928
rect 11517 6851 11575 6857
rect 8573 6811 8631 6817
rect 8680 6820 9628 6848
rect 9692 6820 11468 6848
rect 5031 6752 5396 6780
rect 5813 6783 5871 6789
rect 5031 6749 5043 6752
rect 4985 6743 5043 6749
rect 5813 6749 5825 6783
rect 5859 6780 5871 6783
rect 8294 6780 8300 6792
rect 5859 6752 8300 6780
rect 5859 6749 5871 6752
rect 5813 6743 5871 6749
rect 8294 6740 8300 6752
rect 8352 6780 8358 6792
rect 8588 6780 8616 6811
rect 8352 6752 8616 6780
rect 8352 6740 8358 6752
rect 4203 6715 4261 6721
rect 4203 6681 4215 6715
rect 4249 6712 4261 6715
rect 4798 6712 4804 6724
rect 4249 6684 4804 6712
rect 4249 6681 4261 6684
rect 4203 6675 4261 6681
rect 4798 6672 4804 6684
rect 4856 6672 4862 6724
rect 5074 6672 5080 6724
rect 5132 6712 5138 6724
rect 5169 6715 5227 6721
rect 5169 6712 5181 6715
rect 5132 6684 5181 6712
rect 5132 6672 5138 6684
rect 5169 6681 5181 6684
rect 5215 6712 5227 6715
rect 8680 6712 8708 6820
rect 5215 6684 8708 6712
rect 8757 6715 8815 6721
rect 5215 6681 5227 6684
rect 5169 6675 5227 6681
rect 8757 6681 8769 6715
rect 8803 6712 8815 6715
rect 9306 6712 9312 6724
rect 8803 6684 9312 6712
rect 8803 6681 8815 6684
rect 8757 6675 8815 6681
rect 9306 6672 9312 6684
rect 9364 6672 9370 6724
rect 9600 6712 9628 6820
rect 9677 6783 9735 6789
rect 9677 6749 9689 6783
rect 9723 6780 9735 6783
rect 10686 6780 10692 6792
rect 9723 6752 10692 6780
rect 9723 6749 9735 6752
rect 9677 6743 9735 6749
rect 10686 6740 10692 6752
rect 10744 6740 10750 6792
rect 11440 6780 11468 6820
rect 11517 6817 11529 6851
rect 11563 6817 11575 6851
rect 11517 6811 11575 6817
rect 11606 6808 11612 6860
rect 11664 6848 11670 6860
rect 11790 6848 11796 6860
rect 11664 6820 11709 6848
rect 11751 6820 11796 6848
rect 11664 6808 11670 6820
rect 11790 6808 11796 6820
rect 11848 6808 11854 6860
rect 16298 6848 16304 6860
rect 16259 6820 16304 6848
rect 16298 6808 16304 6820
rect 16356 6808 16362 6860
rect 16577 6851 16635 6857
rect 16577 6817 16589 6851
rect 16623 6848 16635 6851
rect 16850 6848 16856 6860
rect 16623 6820 16856 6848
rect 16623 6817 16635 6820
rect 16577 6811 16635 6817
rect 13170 6780 13176 6792
rect 11440 6752 13032 6780
rect 13083 6752 13176 6780
rect 12342 6712 12348 6724
rect 9600 6684 12348 6712
rect 12342 6672 12348 6684
rect 12400 6672 12406 6724
rect 13004 6712 13032 6752
rect 13170 6740 13176 6752
rect 13228 6780 13234 6792
rect 13725 6783 13783 6789
rect 13725 6780 13737 6783
rect 13228 6752 13737 6780
rect 13228 6740 13234 6752
rect 13725 6749 13737 6752
rect 13771 6749 13783 6783
rect 16592 6780 16620 6811
rect 16850 6808 16856 6820
rect 16908 6808 16914 6860
rect 17586 6848 17592 6860
rect 17547 6820 17592 6848
rect 17586 6808 17592 6820
rect 17644 6808 17650 6860
rect 19337 6851 19395 6857
rect 19337 6817 19349 6851
rect 19383 6848 19395 6851
rect 19426 6848 19432 6860
rect 19383 6820 19432 6848
rect 19383 6817 19395 6820
rect 19337 6811 19395 6817
rect 19426 6808 19432 6820
rect 19484 6808 19490 6860
rect 21818 6848 21824 6860
rect 21779 6820 21824 6848
rect 21818 6808 21824 6820
rect 21876 6808 21882 6860
rect 25307 6857 25335 6956
rect 25292 6851 25350 6857
rect 25292 6817 25304 6851
rect 25338 6848 25350 6851
rect 25774 6848 25780 6860
rect 25338 6820 25780 6848
rect 25338 6817 25350 6820
rect 25292 6811 25350 6817
rect 25774 6808 25780 6820
rect 25832 6808 25838 6860
rect 13725 6743 13783 6749
rect 14108 6752 16620 6780
rect 16761 6783 16819 6789
rect 14108 6712 14136 6752
rect 16761 6749 16773 6783
rect 16807 6780 16819 6783
rect 18046 6780 18052 6792
rect 16807 6752 18052 6780
rect 16807 6749 16819 6752
rect 16761 6743 16819 6749
rect 18046 6740 18052 6752
rect 18104 6740 18110 6792
rect 23198 6740 23204 6792
rect 23256 6780 23262 6792
rect 23753 6783 23811 6789
rect 23753 6780 23765 6783
rect 23256 6752 23765 6780
rect 23256 6740 23262 6752
rect 23753 6749 23765 6752
rect 23799 6749 23811 6783
rect 24026 6780 24032 6792
rect 23987 6752 24032 6780
rect 23753 6743 23811 6749
rect 24026 6740 24032 6752
rect 24084 6740 24090 6792
rect 14274 6712 14280 6724
rect 13004 6684 14136 6712
rect 14235 6684 14280 6712
rect 14274 6672 14280 6684
rect 14332 6672 14338 6724
rect 20438 6712 20444 6724
rect 20351 6684 20444 6712
rect 20438 6672 20444 6684
rect 20496 6712 20502 6724
rect 20496 6684 23474 6712
rect 20496 6672 20502 6684
rect 9214 6644 9220 6656
rect 9175 6616 9220 6644
rect 9214 6604 9220 6616
rect 9272 6604 9278 6656
rect 9582 6604 9588 6656
rect 9640 6644 9646 6656
rect 10597 6647 10655 6653
rect 10597 6644 10609 6647
rect 9640 6616 10609 6644
rect 9640 6604 9646 6616
rect 10597 6613 10609 6616
rect 10643 6644 10655 6647
rect 13354 6644 13360 6656
rect 10643 6616 13360 6644
rect 10643 6613 10655 6616
rect 10597 6607 10655 6613
rect 13354 6604 13360 6616
rect 13412 6604 13418 6656
rect 18506 6644 18512 6656
rect 18467 6616 18512 6644
rect 18506 6604 18512 6616
rect 18564 6604 18570 6656
rect 23446 6644 23474 6684
rect 25363 6647 25421 6653
rect 25363 6644 25375 6647
rect 23446 6616 25375 6644
rect 25363 6613 25375 6616
rect 25409 6613 25421 6647
rect 25363 6607 25421 6613
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 4706 6440 4712 6452
rect 4667 6412 4712 6440
rect 4706 6400 4712 6412
rect 4764 6400 4770 6452
rect 5074 6440 5080 6452
rect 5035 6412 5080 6440
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 6089 6443 6147 6449
rect 6089 6409 6101 6443
rect 6135 6440 6147 6443
rect 6641 6443 6699 6449
rect 6641 6440 6653 6443
rect 6135 6412 6653 6440
rect 6135 6409 6147 6412
rect 6089 6403 6147 6409
rect 6641 6409 6653 6412
rect 6687 6440 6699 6443
rect 7926 6440 7932 6452
rect 6687 6412 7932 6440
rect 6687 6409 6699 6412
rect 6641 6403 6699 6409
rect 7926 6400 7932 6412
rect 7984 6400 7990 6452
rect 8294 6440 8300 6452
rect 8255 6412 8300 6440
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 11606 6400 11612 6452
rect 11664 6440 11670 6452
rect 11793 6443 11851 6449
rect 11793 6440 11805 6443
rect 11664 6412 11805 6440
rect 11664 6400 11670 6412
rect 11793 6409 11805 6412
rect 11839 6409 11851 6443
rect 11793 6403 11851 6409
rect 12667 6443 12725 6449
rect 12667 6409 12679 6443
rect 12713 6440 12725 6443
rect 13170 6440 13176 6452
rect 12713 6412 13176 6440
rect 12713 6409 12725 6412
rect 12667 6403 12725 6409
rect 13170 6400 13176 6412
rect 13228 6400 13234 6452
rect 17034 6440 17040 6452
rect 13280 6412 16896 6440
rect 16995 6412 17040 6440
rect 5261 6375 5319 6381
rect 5261 6341 5273 6375
rect 5307 6372 5319 6375
rect 5994 6372 6000 6384
rect 5307 6344 6000 6372
rect 5307 6341 5319 6344
rect 5261 6335 5319 6341
rect 5994 6332 6000 6344
rect 6052 6372 6058 6384
rect 6181 6375 6239 6381
rect 6181 6372 6193 6375
rect 6052 6344 6193 6372
rect 6052 6332 6058 6344
rect 6181 6341 6193 6344
rect 6227 6372 6239 6375
rect 7374 6372 7380 6384
rect 6227 6344 7380 6372
rect 6227 6341 6239 6344
rect 6181 6335 6239 6341
rect 7374 6332 7380 6344
rect 7432 6332 7438 6384
rect 7466 6332 7472 6384
rect 7524 6372 7530 6384
rect 9214 6372 9220 6384
rect 7524 6344 9220 6372
rect 7524 6332 7530 6344
rect 9214 6332 9220 6344
rect 9272 6372 9278 6384
rect 9309 6375 9367 6381
rect 9309 6372 9321 6375
rect 9272 6344 9321 6372
rect 9272 6332 9278 6344
rect 9309 6341 9321 6344
rect 9355 6341 9367 6375
rect 9309 6335 9367 6341
rect 6362 6304 6368 6316
rect 5184 6276 6368 6304
rect 4203 6239 4261 6245
rect 4203 6205 4215 6239
rect 4249 6205 4261 6239
rect 4203 6199 4261 6205
rect 3970 6100 3976 6112
rect 3931 6072 3976 6100
rect 3970 6060 3976 6072
rect 4028 6100 4034 6112
rect 4218 6100 4246 6199
rect 4890 6196 4896 6248
rect 4948 6236 4954 6248
rect 5184 6245 5212 6276
rect 6362 6264 6368 6276
rect 6420 6264 6426 6316
rect 6454 6264 6460 6316
rect 6512 6304 6518 6316
rect 7193 6307 7251 6313
rect 7193 6304 7205 6307
rect 6512 6276 7205 6304
rect 6512 6264 6518 6276
rect 7193 6273 7205 6276
rect 7239 6273 7251 6307
rect 7193 6267 7251 6273
rect 7558 6264 7564 6316
rect 7616 6304 7622 6316
rect 7929 6307 7987 6313
rect 7929 6304 7941 6307
rect 7616 6276 7941 6304
rect 7616 6264 7622 6276
rect 7929 6273 7941 6276
rect 7975 6304 7987 6307
rect 9582 6304 9588 6316
rect 7975 6276 9588 6304
rect 7975 6273 7987 6276
rect 7929 6267 7987 6273
rect 9582 6264 9588 6276
rect 9640 6264 9646 6316
rect 11606 6304 11612 6316
rect 11440 6276 11612 6304
rect 5169 6239 5227 6245
rect 5169 6236 5181 6239
rect 4948 6208 5181 6236
rect 4948 6196 4954 6208
rect 5169 6205 5181 6208
rect 5215 6205 5227 6239
rect 5169 6199 5227 6205
rect 5445 6239 5503 6245
rect 5445 6205 5457 6239
rect 5491 6236 5503 6239
rect 5534 6236 5540 6248
rect 5491 6208 5540 6236
rect 5491 6205 5503 6208
rect 5445 6199 5503 6205
rect 5534 6196 5540 6208
rect 5592 6236 5598 6248
rect 11440 6245 11468 6276
rect 11606 6264 11612 6276
rect 11664 6304 11670 6316
rect 13280 6304 13308 6412
rect 13354 6332 13360 6384
rect 13412 6372 13418 6384
rect 16114 6372 16120 6384
rect 13412 6344 16120 6372
rect 13412 6332 13418 6344
rect 16114 6332 16120 6344
rect 16172 6332 16178 6384
rect 16298 6372 16304 6384
rect 16259 6344 16304 6372
rect 16298 6332 16304 6344
rect 16356 6332 16362 6384
rect 16758 6372 16764 6384
rect 16719 6344 16764 6372
rect 16758 6332 16764 6344
rect 16816 6332 16822 6384
rect 15378 6304 15384 6316
rect 11664 6276 13308 6304
rect 15339 6276 15384 6304
rect 11664 6264 11670 6276
rect 15378 6264 15384 6276
rect 15436 6264 15442 6316
rect 6089 6239 6147 6245
rect 6089 6236 6101 6239
rect 5592 6208 6101 6236
rect 5592 6196 5598 6208
rect 6089 6205 6101 6208
rect 6135 6205 6147 6239
rect 9217 6239 9275 6245
rect 9217 6236 9229 6239
rect 6089 6199 6147 6205
rect 8680 6208 9229 6236
rect 6454 6128 6460 6180
rect 6512 6168 6518 6180
rect 6914 6168 6920 6180
rect 6512 6140 6684 6168
rect 6875 6140 6920 6168
rect 6512 6128 6518 6140
rect 4028 6072 4246 6100
rect 4295 6103 4353 6109
rect 4028 6060 4034 6072
rect 4295 6069 4307 6103
rect 4341 6100 4353 6103
rect 4522 6100 4528 6112
rect 4341 6072 4528 6100
rect 4341 6069 4353 6072
rect 4295 6063 4353 6069
rect 4522 6060 4528 6072
rect 4580 6060 4586 6112
rect 5074 6060 5080 6112
rect 5132 6100 5138 6112
rect 5629 6103 5687 6109
rect 5629 6100 5641 6103
rect 5132 6072 5641 6100
rect 5132 6060 5138 6072
rect 5629 6069 5641 6072
rect 5675 6069 5687 6103
rect 6656 6100 6684 6140
rect 6914 6128 6920 6140
rect 6972 6128 6978 6180
rect 7006 6128 7012 6180
rect 7064 6168 7070 6180
rect 7558 6168 7564 6180
rect 7064 6140 7564 6168
rect 7064 6128 7070 6140
rect 7558 6128 7564 6140
rect 7616 6128 7622 6180
rect 8680 6112 8708 6208
rect 9217 6205 9229 6208
rect 9263 6205 9275 6239
rect 9217 6199 9275 6205
rect 9493 6239 9551 6245
rect 9493 6205 9505 6239
rect 9539 6205 9551 6239
rect 9493 6199 9551 6205
rect 10689 6239 10747 6245
rect 10689 6205 10701 6239
rect 10735 6236 10747 6239
rect 11425 6239 11483 6245
rect 11425 6236 11437 6239
rect 10735 6208 11437 6236
rect 10735 6205 10747 6208
rect 10689 6199 10747 6205
rect 11425 6205 11437 6208
rect 11471 6205 11483 6239
rect 11425 6199 11483 6205
rect 11517 6239 11575 6245
rect 11517 6205 11529 6239
rect 11563 6236 11575 6239
rect 11790 6236 11796 6248
rect 11563 6208 11796 6236
rect 11563 6205 11575 6208
rect 11517 6199 11575 6205
rect 8662 6100 8668 6112
rect 6656 6072 8668 6100
rect 5629 6063 5687 6069
rect 8662 6060 8668 6072
rect 8720 6060 8726 6112
rect 9030 6100 9036 6112
rect 8991 6072 9036 6100
rect 9030 6060 9036 6072
rect 9088 6100 9094 6112
rect 9508 6100 9536 6199
rect 11790 6196 11796 6208
rect 11848 6236 11854 6248
rect 12161 6239 12219 6245
rect 12161 6236 12173 6239
rect 11848 6208 12173 6236
rect 11848 6196 11854 6208
rect 12161 6205 12173 6208
rect 12207 6205 12219 6239
rect 12161 6199 12219 6205
rect 12596 6239 12654 6245
rect 12596 6205 12608 6239
rect 12642 6236 12654 6239
rect 13541 6239 13599 6245
rect 12642 6208 13124 6236
rect 12642 6205 12654 6208
rect 12596 6199 12654 6205
rect 9953 6171 10011 6177
rect 9953 6137 9965 6171
rect 9999 6168 10011 6171
rect 11238 6168 11244 6180
rect 9999 6140 11244 6168
rect 9999 6137 10011 6140
rect 9953 6131 10011 6137
rect 11238 6128 11244 6140
rect 11296 6128 11302 6180
rect 9088 6072 9536 6100
rect 9088 6060 9094 6072
rect 10042 6060 10048 6112
rect 10100 6100 10106 6112
rect 10321 6103 10379 6109
rect 10321 6100 10333 6103
rect 10100 6072 10333 6100
rect 10100 6060 10106 6072
rect 10321 6069 10333 6072
rect 10367 6100 10379 6103
rect 12710 6100 12716 6112
rect 10367 6072 12716 6100
rect 10367 6069 10379 6072
rect 10321 6063 10379 6069
rect 12710 6060 12716 6072
rect 12768 6060 12774 6112
rect 13096 6109 13124 6208
rect 13541 6205 13553 6239
rect 13587 6205 13599 6239
rect 13541 6199 13599 6205
rect 13081 6103 13139 6109
rect 13081 6069 13093 6103
rect 13127 6100 13139 6103
rect 13170 6100 13176 6112
rect 13127 6072 13176 6100
rect 13127 6069 13139 6072
rect 13081 6063 13139 6069
rect 13170 6060 13176 6072
rect 13228 6060 13234 6112
rect 13262 6060 13268 6112
rect 13320 6100 13326 6112
rect 13357 6103 13415 6109
rect 13357 6100 13369 6103
rect 13320 6072 13369 6100
rect 13320 6060 13326 6072
rect 13357 6069 13369 6072
rect 13403 6100 13415 6103
rect 13556 6100 13584 6199
rect 13814 6196 13820 6248
rect 13872 6236 13878 6248
rect 14090 6236 14096 6248
rect 13872 6208 14096 6236
rect 13872 6196 13878 6208
rect 14090 6196 14096 6208
rect 14148 6236 14154 6248
rect 16868 6245 16896 6412
rect 17034 6400 17040 6412
rect 17092 6400 17098 6452
rect 23293 6443 23351 6449
rect 23293 6409 23305 6443
rect 23339 6440 23351 6443
rect 23842 6440 23848 6452
rect 23339 6412 23848 6440
rect 23339 6409 23351 6412
rect 23293 6403 23351 6409
rect 23842 6400 23848 6412
rect 23900 6400 23906 6452
rect 25038 6400 25044 6452
rect 25096 6440 25102 6452
rect 25455 6443 25513 6449
rect 25455 6440 25467 6443
rect 25096 6412 25467 6440
rect 25096 6400 25102 6412
rect 25455 6409 25467 6412
rect 25501 6409 25513 6443
rect 25455 6403 25513 6409
rect 25866 6400 25872 6452
rect 25924 6440 25930 6452
rect 26145 6443 26203 6449
rect 26145 6440 26157 6443
rect 25924 6412 26157 6440
rect 25924 6400 25930 6412
rect 26145 6409 26157 6412
rect 26191 6409 26203 6443
rect 26145 6403 26203 6409
rect 19426 6372 19432 6384
rect 19339 6344 19432 6372
rect 19426 6332 19432 6344
rect 19484 6372 19490 6384
rect 23474 6372 23480 6384
rect 19484 6344 23480 6372
rect 19484 6332 19490 6344
rect 23474 6332 23480 6344
rect 23532 6332 23538 6384
rect 23566 6332 23572 6384
rect 23624 6372 23630 6384
rect 24765 6375 24823 6381
rect 24765 6372 24777 6375
rect 23624 6344 24777 6372
rect 23624 6332 23630 6344
rect 24765 6341 24777 6344
rect 24811 6341 24823 6375
rect 24765 6335 24823 6341
rect 18046 6304 18052 6316
rect 18007 6276 18052 6304
rect 18046 6264 18052 6276
rect 18104 6264 18110 6316
rect 18414 6264 18420 6316
rect 18472 6304 18478 6316
rect 19518 6304 19524 6316
rect 18472 6276 19524 6304
rect 18472 6264 18478 6276
rect 19518 6264 19524 6276
rect 19576 6304 19582 6316
rect 19797 6307 19855 6313
rect 19797 6304 19809 6307
rect 19576 6276 19809 6304
rect 19576 6264 19582 6276
rect 19797 6273 19809 6276
rect 19843 6273 19855 6307
rect 22186 6304 22192 6316
rect 19797 6267 19855 6273
rect 21836 6276 22192 6304
rect 14553 6239 14611 6245
rect 14553 6236 14565 6239
rect 14148 6208 14565 6236
rect 14148 6196 14154 6208
rect 14553 6205 14565 6208
rect 14599 6205 14611 6239
rect 14553 6199 14611 6205
rect 16853 6239 16911 6245
rect 16853 6205 16865 6239
rect 16899 6236 16911 6239
rect 17313 6239 17371 6245
rect 17313 6236 17325 6239
rect 16899 6208 17325 6236
rect 16899 6205 16911 6208
rect 16853 6199 16911 6205
rect 17313 6205 17325 6208
rect 17359 6205 17371 6239
rect 17313 6199 17371 6205
rect 17954 6196 17960 6248
rect 18012 6236 18018 6248
rect 21836 6245 21864 6276
rect 22186 6264 22192 6276
rect 22244 6264 22250 6316
rect 23842 6264 23848 6316
rect 23900 6304 23906 6316
rect 24026 6304 24032 6316
rect 23900 6276 24032 6304
rect 23900 6264 23906 6276
rect 24026 6264 24032 6276
rect 24084 6304 24090 6316
rect 24121 6307 24179 6313
rect 24121 6304 24133 6307
rect 24084 6276 24133 6304
rect 24084 6264 24090 6276
rect 24121 6273 24133 6276
rect 24167 6273 24179 6307
rect 24121 6267 24179 6273
rect 21821 6239 21879 6245
rect 21821 6236 21833 6239
rect 18012 6208 21833 6236
rect 18012 6196 18018 6208
rect 21821 6205 21833 6208
rect 21867 6205 21879 6239
rect 23293 6239 23351 6245
rect 23293 6236 23305 6239
rect 21821 6199 21879 6205
rect 21928 6208 23305 6236
rect 14277 6171 14335 6177
rect 14277 6137 14289 6171
rect 14323 6168 14335 6171
rect 15194 6168 15200 6180
rect 14323 6140 15200 6168
rect 14323 6137 14335 6140
rect 14277 6131 14335 6137
rect 15194 6128 15200 6140
rect 15252 6128 15258 6180
rect 15470 6128 15476 6180
rect 15528 6168 15534 6180
rect 16025 6171 16083 6177
rect 15528 6140 15573 6168
rect 15528 6128 15534 6140
rect 16025 6137 16037 6171
rect 16071 6168 16083 6171
rect 16758 6168 16764 6180
rect 16071 6140 16764 6168
rect 16071 6137 16083 6140
rect 16025 6131 16083 6137
rect 16758 6128 16764 6140
rect 16816 6128 16822 6180
rect 18370 6171 18428 6177
rect 18370 6168 18382 6171
rect 17696 6140 18382 6168
rect 17696 6112 17724 6140
rect 18370 6137 18382 6140
rect 18416 6168 18428 6171
rect 20118 6171 20176 6177
rect 20118 6168 20130 6171
rect 18416 6140 20130 6168
rect 18416 6137 18428 6140
rect 18370 6131 18428 6137
rect 20118 6137 20130 6140
rect 20164 6137 20176 6171
rect 21726 6168 21732 6180
rect 20118 6131 20176 6137
rect 20548 6140 21732 6168
rect 14826 6100 14832 6112
rect 13403 6072 14832 6100
rect 13403 6069 13415 6072
rect 13357 6063 13415 6069
rect 14826 6060 14832 6072
rect 14884 6060 14890 6112
rect 15105 6103 15163 6109
rect 15105 6069 15117 6103
rect 15151 6100 15163 6103
rect 15286 6100 15292 6112
rect 15151 6072 15292 6100
rect 15151 6069 15163 6072
rect 15105 6063 15163 6069
rect 15286 6060 15292 6072
rect 15344 6060 15350 6112
rect 15654 6060 15660 6112
rect 15712 6100 15718 6112
rect 17678 6100 17684 6112
rect 15712 6072 17684 6100
rect 15712 6060 15718 6072
rect 17678 6060 17684 6072
rect 17736 6060 17742 6112
rect 18230 6060 18236 6112
rect 18288 6100 18294 6112
rect 18969 6103 19027 6109
rect 18969 6100 18981 6103
rect 18288 6072 18981 6100
rect 18288 6060 18294 6072
rect 18969 6069 18981 6072
rect 19015 6100 19027 6103
rect 20548 6100 20576 6140
rect 21726 6128 21732 6140
rect 21784 6168 21790 6180
rect 21928 6168 21956 6208
rect 23293 6205 23305 6208
rect 23339 6236 23351 6239
rect 23385 6239 23443 6245
rect 23385 6236 23397 6239
rect 23339 6208 23397 6236
rect 23339 6205 23351 6208
rect 23293 6199 23351 6205
rect 23385 6205 23397 6208
rect 23431 6205 23443 6239
rect 23385 6199 23443 6205
rect 25384 6239 25442 6245
rect 25384 6205 25396 6239
rect 25430 6236 25442 6239
rect 25866 6236 25872 6248
rect 25430 6208 25872 6236
rect 25430 6205 25442 6208
rect 25384 6199 25442 6205
rect 25866 6196 25872 6208
rect 25924 6196 25930 6248
rect 21784 6140 21956 6168
rect 21784 6128 21790 6140
rect 23566 6128 23572 6180
rect 23624 6168 23630 6180
rect 23845 6171 23903 6177
rect 23845 6168 23857 6171
rect 23624 6140 23857 6168
rect 23624 6128 23630 6140
rect 23845 6137 23857 6140
rect 23891 6137 23903 6171
rect 23845 6131 23903 6137
rect 23937 6171 23995 6177
rect 23937 6137 23949 6171
rect 23983 6137 23995 6171
rect 23937 6131 23995 6137
rect 20714 6100 20720 6112
rect 19015 6072 20576 6100
rect 20675 6072 20720 6100
rect 19015 6069 19027 6072
rect 18969 6063 19027 6069
rect 20714 6060 20720 6072
rect 20772 6060 20778 6112
rect 21266 6100 21272 6112
rect 21227 6072 21272 6100
rect 21266 6060 21272 6072
rect 21324 6100 21330 6112
rect 21637 6103 21695 6109
rect 21637 6100 21649 6103
rect 21324 6072 21649 6100
rect 21324 6060 21330 6072
rect 21637 6069 21649 6072
rect 21683 6069 21695 6103
rect 21637 6063 21695 6069
rect 22094 6060 22100 6112
rect 22152 6100 22158 6112
rect 22189 6103 22247 6109
rect 22189 6100 22201 6103
rect 22152 6072 22201 6100
rect 22152 6060 22158 6072
rect 22189 6069 22201 6072
rect 22235 6069 22247 6103
rect 22189 6063 22247 6069
rect 22554 6060 22560 6112
rect 22612 6100 22618 6112
rect 22741 6103 22799 6109
rect 22741 6100 22753 6103
rect 22612 6072 22753 6100
rect 22612 6060 22618 6072
rect 22741 6069 22753 6072
rect 22787 6069 22799 6103
rect 22741 6063 22799 6069
rect 23109 6103 23167 6109
rect 23109 6069 23121 6103
rect 23155 6100 23167 6103
rect 23198 6100 23204 6112
rect 23155 6072 23204 6100
rect 23155 6069 23167 6072
rect 23109 6063 23167 6069
rect 23198 6060 23204 6072
rect 23256 6060 23262 6112
rect 23750 6060 23756 6112
rect 23808 6100 23814 6112
rect 23952 6100 23980 6131
rect 25774 6100 25780 6112
rect 23808 6072 23980 6100
rect 25735 6072 25780 6100
rect 23808 6060 23814 6072
rect 25774 6060 25780 6072
rect 25832 6060 25838 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 8481 5899 8539 5905
rect 8481 5896 8493 5899
rect 4126 5868 8493 5896
rect 3234 5828 3240 5840
rect 2976 5800 3240 5828
rect 2976 5769 3004 5800
rect 3234 5788 3240 5800
rect 3292 5828 3298 5840
rect 4126 5828 4154 5868
rect 8481 5865 8493 5868
rect 8527 5865 8539 5899
rect 8481 5859 8539 5865
rect 8662 5856 8668 5908
rect 8720 5896 8726 5908
rect 9033 5899 9091 5905
rect 9033 5896 9045 5899
rect 8720 5868 9045 5896
rect 8720 5856 8726 5868
rect 9033 5865 9045 5868
rect 9079 5865 9091 5899
rect 9033 5859 9091 5865
rect 3292 5800 4154 5828
rect 3292 5788 3298 5800
rect 4522 5788 4528 5840
rect 4580 5828 4586 5840
rect 6273 5831 6331 5837
rect 6273 5828 6285 5831
rect 4580 5800 6285 5828
rect 4580 5788 4586 5800
rect 6273 5797 6285 5800
rect 6319 5828 6331 5831
rect 6914 5828 6920 5840
rect 6319 5800 6920 5828
rect 6319 5797 6331 5800
rect 6273 5791 6331 5797
rect 6914 5788 6920 5800
rect 6972 5788 6978 5840
rect 7190 5828 7196 5840
rect 7151 5800 7196 5828
rect 7190 5788 7196 5800
rect 7248 5788 7254 5840
rect 7558 5828 7564 5840
rect 7519 5800 7564 5828
rect 7558 5788 7564 5800
rect 7616 5788 7622 5840
rect 7926 5828 7932 5840
rect 7839 5800 7932 5828
rect 7926 5788 7932 5800
rect 7984 5828 7990 5840
rect 7984 5800 8340 5828
rect 7984 5788 7990 5800
rect 2961 5763 3019 5769
rect 2961 5729 2973 5763
rect 3007 5729 3019 5763
rect 2961 5723 3019 5729
rect 4614 5720 4620 5772
rect 4672 5760 4678 5772
rect 4893 5763 4951 5769
rect 4893 5760 4905 5763
rect 4672 5732 4905 5760
rect 4672 5720 4678 5732
rect 4893 5729 4905 5732
rect 4939 5729 4951 5763
rect 5166 5760 5172 5772
rect 5127 5732 5172 5760
rect 4893 5723 4951 5729
rect 5166 5720 5172 5732
rect 5224 5720 5230 5772
rect 5997 5763 6055 5769
rect 5997 5729 6009 5763
rect 6043 5760 6055 5763
rect 6362 5760 6368 5772
rect 6043 5732 6368 5760
rect 6043 5729 6055 5732
rect 5997 5723 6055 5729
rect 6362 5720 6368 5732
rect 6420 5720 6426 5772
rect 6454 5720 6460 5772
rect 6512 5760 6518 5772
rect 6733 5763 6791 5769
rect 6512 5732 6557 5760
rect 6512 5720 6518 5732
rect 6733 5729 6745 5763
rect 6779 5729 6791 5763
rect 8018 5760 8024 5772
rect 7979 5732 8024 5760
rect 6733 5723 6791 5729
rect 4706 5652 4712 5704
rect 4764 5692 4770 5704
rect 4801 5695 4859 5701
rect 4801 5692 4813 5695
rect 4764 5664 4813 5692
rect 4764 5652 4770 5664
rect 4801 5661 4813 5664
rect 4847 5692 4859 5695
rect 5353 5695 5411 5701
rect 5353 5692 5365 5695
rect 4847 5664 5365 5692
rect 4847 5661 4859 5664
rect 4801 5655 4859 5661
rect 5353 5661 5365 5664
rect 5399 5661 5411 5695
rect 5353 5655 5411 5661
rect 6638 5652 6644 5704
rect 6696 5692 6702 5704
rect 6748 5692 6776 5723
rect 8018 5720 8024 5732
rect 8076 5720 8082 5772
rect 8312 5769 8340 5800
rect 8297 5763 8355 5769
rect 8297 5729 8309 5763
rect 8343 5760 8355 5763
rect 8386 5760 8392 5772
rect 8343 5732 8392 5760
rect 8343 5729 8355 5732
rect 8297 5723 8355 5729
rect 8386 5720 8392 5732
rect 8444 5720 8450 5772
rect 9048 5760 9076 5859
rect 9398 5856 9404 5908
rect 9456 5896 9462 5908
rect 10137 5899 10195 5905
rect 10137 5896 10149 5899
rect 9456 5868 10149 5896
rect 9456 5856 9462 5868
rect 10137 5865 10149 5868
rect 10183 5865 10195 5899
rect 10686 5896 10692 5908
rect 10647 5868 10692 5896
rect 10137 5859 10195 5865
rect 10686 5856 10692 5868
rect 10744 5856 10750 5908
rect 11422 5856 11428 5908
rect 11480 5896 11486 5908
rect 11517 5899 11575 5905
rect 11517 5896 11529 5899
rect 11480 5868 11529 5896
rect 11480 5856 11486 5868
rect 11517 5865 11529 5868
rect 11563 5865 11575 5899
rect 13538 5896 13544 5908
rect 13499 5868 13544 5896
rect 11517 5859 11575 5865
rect 13538 5856 13544 5868
rect 13596 5856 13602 5908
rect 15654 5896 15660 5908
rect 15615 5868 15660 5896
rect 15654 5856 15660 5868
rect 15712 5856 15718 5908
rect 17586 5896 17592 5908
rect 17547 5868 17592 5896
rect 17586 5856 17592 5868
rect 17644 5856 17650 5908
rect 18138 5856 18144 5908
rect 18196 5896 18202 5908
rect 18877 5899 18935 5905
rect 18877 5896 18889 5899
rect 18196 5868 18889 5896
rect 18196 5856 18202 5868
rect 18877 5865 18889 5868
rect 18923 5865 18935 5899
rect 19334 5896 19340 5908
rect 19295 5868 19340 5896
rect 18877 5859 18935 5865
rect 19334 5856 19340 5868
rect 19392 5856 19398 5908
rect 19518 5856 19524 5908
rect 19576 5896 19582 5908
rect 19889 5899 19947 5905
rect 19889 5896 19901 5899
rect 19576 5868 19901 5896
rect 19576 5856 19582 5868
rect 19889 5865 19901 5868
rect 19935 5865 19947 5899
rect 20254 5896 20260 5908
rect 20215 5868 20260 5896
rect 19889 5859 19947 5865
rect 20254 5856 20260 5868
rect 20312 5856 20318 5908
rect 21266 5896 21272 5908
rect 21227 5868 21272 5896
rect 21266 5856 21272 5868
rect 21324 5856 21330 5908
rect 21818 5856 21824 5908
rect 21876 5896 21882 5908
rect 22097 5899 22155 5905
rect 22097 5896 22109 5899
rect 21876 5868 22109 5896
rect 21876 5856 21882 5868
rect 22097 5865 22109 5868
rect 22143 5865 22155 5899
rect 22097 5859 22155 5865
rect 22186 5856 22192 5908
rect 22244 5896 22250 5908
rect 22465 5899 22523 5905
rect 22465 5896 22477 5899
rect 22244 5868 22477 5896
rect 22244 5856 22250 5868
rect 22465 5865 22477 5868
rect 22511 5865 22523 5899
rect 23106 5896 23112 5908
rect 23067 5868 23112 5896
rect 22465 5859 22523 5865
rect 23106 5856 23112 5868
rect 23164 5856 23170 5908
rect 23750 5896 23756 5908
rect 23711 5868 23756 5896
rect 23750 5856 23756 5868
rect 23808 5896 23814 5908
rect 23808 5868 24348 5896
rect 23808 5856 23814 5868
rect 13814 5788 13820 5840
rect 13872 5828 13878 5840
rect 13872 5800 13917 5828
rect 13872 5788 13878 5800
rect 17218 5788 17224 5840
rect 17276 5828 17282 5840
rect 17770 5828 17776 5840
rect 17276 5800 17776 5828
rect 17276 5788 17282 5800
rect 17770 5788 17776 5800
rect 17828 5828 17834 5840
rect 17957 5831 18015 5837
rect 17957 5828 17969 5831
rect 17828 5800 17969 5828
rect 17828 5788 17834 5800
rect 17957 5797 17969 5800
rect 18003 5797 18015 5831
rect 17957 5791 18015 5797
rect 18049 5831 18107 5837
rect 18049 5797 18061 5831
rect 18095 5828 18107 5831
rect 18230 5828 18236 5840
rect 18095 5800 18236 5828
rect 18095 5797 18107 5800
rect 18049 5791 18107 5797
rect 18230 5788 18236 5800
rect 18288 5788 18294 5840
rect 18601 5831 18659 5837
rect 18601 5797 18613 5831
rect 18647 5828 18659 5831
rect 20272 5828 20300 5856
rect 18647 5800 20300 5828
rect 21284 5828 21312 5856
rect 24210 5828 24216 5840
rect 21284 5800 22140 5828
rect 24171 5800 24216 5828
rect 18647 5797 18659 5800
rect 18601 5791 18659 5797
rect 22112 5772 22140 5800
rect 24210 5788 24216 5800
rect 24268 5788 24274 5840
rect 24320 5837 24348 5868
rect 24305 5831 24363 5837
rect 24305 5797 24317 5831
rect 24351 5828 24363 5831
rect 24670 5828 24676 5840
rect 24351 5800 24676 5828
rect 24351 5797 24363 5800
rect 24305 5791 24363 5797
rect 24670 5788 24676 5800
rect 24728 5788 24734 5840
rect 9677 5763 9735 5769
rect 9677 5760 9689 5763
rect 9048 5732 9689 5760
rect 9677 5729 9689 5732
rect 9723 5729 9735 5763
rect 9677 5723 9735 5729
rect 9953 5763 10011 5769
rect 9953 5729 9965 5763
rect 9999 5729 10011 5763
rect 9953 5723 10011 5729
rect 9030 5692 9036 5704
rect 6696 5664 9036 5692
rect 6696 5652 6702 5664
rect 9030 5652 9036 5664
rect 9088 5652 9094 5704
rect 9968 5692 9996 5723
rect 11330 5720 11336 5772
rect 11388 5760 11394 5772
rect 12069 5763 12127 5769
rect 12069 5760 12081 5763
rect 11388 5732 12081 5760
rect 11388 5720 11394 5732
rect 12069 5729 12081 5732
rect 12115 5729 12127 5763
rect 12069 5723 12127 5729
rect 12158 5720 12164 5772
rect 12216 5760 12222 5772
rect 12621 5763 12679 5769
rect 12621 5760 12633 5763
rect 12216 5732 12633 5760
rect 12216 5720 12222 5732
rect 12621 5729 12633 5732
rect 12667 5760 12679 5763
rect 13538 5760 13544 5772
rect 12667 5732 13544 5760
rect 12667 5729 12679 5732
rect 12621 5723 12679 5729
rect 13538 5720 13544 5732
rect 13596 5720 13602 5772
rect 15194 5720 15200 5772
rect 15252 5760 15258 5772
rect 15289 5763 15347 5769
rect 15289 5760 15301 5763
rect 15252 5732 15301 5760
rect 15252 5720 15258 5732
rect 15289 5729 15301 5732
rect 15335 5729 15347 5763
rect 19496 5763 19554 5769
rect 19496 5760 19508 5763
rect 15289 5723 15347 5729
rect 18616 5732 19508 5760
rect 12802 5692 12808 5704
rect 9416 5664 9996 5692
rect 12763 5664 12808 5692
rect 4982 5624 4988 5636
rect 4943 5596 4988 5624
rect 4982 5584 4988 5596
rect 5040 5584 5046 5636
rect 6546 5624 6552 5636
rect 6507 5596 6552 5624
rect 6546 5584 6552 5596
rect 6604 5584 6610 5636
rect 7374 5584 7380 5636
rect 7432 5624 7438 5636
rect 7926 5624 7932 5636
rect 7432 5596 7932 5624
rect 7432 5584 7438 5596
rect 7926 5584 7932 5596
rect 7984 5624 7990 5636
rect 8113 5627 8171 5633
rect 8113 5624 8125 5627
rect 7984 5596 8125 5624
rect 7984 5584 7990 5596
rect 8113 5593 8125 5596
rect 8159 5593 8171 5627
rect 8113 5587 8171 5593
rect 9416 5568 9444 5664
rect 12802 5652 12808 5664
rect 12860 5652 12866 5704
rect 13722 5692 13728 5704
rect 13683 5664 13728 5692
rect 13722 5652 13728 5664
rect 13780 5652 13786 5704
rect 14369 5695 14427 5701
rect 14369 5661 14381 5695
rect 14415 5692 14427 5695
rect 18616 5692 18644 5732
rect 19496 5729 19508 5732
rect 19542 5760 19554 5763
rect 19702 5760 19708 5772
rect 19542 5732 19708 5760
rect 19542 5729 19554 5732
rect 19496 5723 19554 5729
rect 19702 5720 19708 5732
rect 19760 5720 19766 5772
rect 19978 5720 19984 5772
rect 20036 5760 20042 5772
rect 20901 5763 20959 5769
rect 20901 5760 20913 5763
rect 20036 5732 20913 5760
rect 20036 5720 20042 5732
rect 20901 5729 20913 5732
rect 20947 5729 20959 5763
rect 20901 5723 20959 5729
rect 21082 5720 21088 5772
rect 21140 5760 21146 5772
rect 21818 5760 21824 5772
rect 21140 5732 21824 5760
rect 21140 5720 21146 5732
rect 21818 5720 21824 5732
rect 21876 5720 21882 5772
rect 22094 5720 22100 5772
rect 22152 5720 22158 5772
rect 14415 5664 18644 5692
rect 14415 5661 14427 5664
rect 14369 5655 14427 5661
rect 9766 5624 9772 5636
rect 9727 5596 9772 5624
rect 9766 5584 9772 5596
rect 9824 5584 9830 5636
rect 11698 5584 11704 5636
rect 11756 5624 11762 5636
rect 14384 5624 14412 5655
rect 21358 5652 21364 5704
rect 21416 5692 21422 5704
rect 22738 5692 22744 5704
rect 21416 5664 22744 5692
rect 21416 5652 21422 5664
rect 22738 5652 22744 5664
rect 22796 5692 22802 5704
rect 24489 5695 24547 5701
rect 22796 5664 23474 5692
rect 22796 5652 22802 5664
rect 11756 5596 14412 5624
rect 11756 5584 11762 5596
rect 16114 5584 16120 5636
rect 16172 5624 16178 5636
rect 16485 5627 16543 5633
rect 16485 5624 16497 5627
rect 16172 5596 16497 5624
rect 16172 5584 16178 5596
rect 16485 5593 16497 5596
rect 16531 5593 16543 5627
rect 23446 5624 23474 5664
rect 24489 5661 24501 5695
rect 24535 5661 24547 5695
rect 24489 5655 24547 5661
rect 24504 5624 24532 5655
rect 23446 5596 24532 5624
rect 16485 5587 16543 5593
rect 3145 5559 3203 5565
rect 3145 5525 3157 5559
rect 3191 5556 3203 5559
rect 5534 5556 5540 5568
rect 3191 5528 5540 5556
rect 3191 5525 3203 5528
rect 3145 5519 3203 5525
rect 5534 5516 5540 5528
rect 5592 5516 5598 5568
rect 9398 5556 9404 5568
rect 9359 5528 9404 5556
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 13078 5556 13084 5568
rect 13039 5528 13084 5556
rect 13078 5516 13084 5528
rect 13136 5516 13142 5568
rect 16206 5556 16212 5568
rect 16167 5528 16212 5556
rect 16206 5516 16212 5528
rect 16264 5516 16270 5568
rect 19334 5516 19340 5568
rect 19392 5556 19398 5568
rect 19567 5559 19625 5565
rect 19567 5556 19579 5559
rect 19392 5528 19579 5556
rect 19392 5516 19398 5528
rect 19567 5525 19579 5528
rect 19613 5525 19625 5559
rect 19567 5519 19625 5525
rect 23566 5516 23572 5568
rect 23624 5556 23630 5568
rect 25498 5556 25504 5568
rect 23624 5528 25504 5556
rect 23624 5516 23630 5528
rect 25498 5516 25504 5528
rect 25556 5516 25562 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1670 5352 1676 5364
rect 1631 5324 1676 5352
rect 1670 5312 1676 5324
rect 1728 5312 1734 5364
rect 3234 5352 3240 5364
rect 3195 5324 3240 5352
rect 3234 5312 3240 5324
rect 3292 5312 3298 5364
rect 3878 5312 3884 5364
rect 3936 5352 3942 5364
rect 3973 5355 4031 5361
rect 3973 5352 3985 5355
rect 3936 5324 3985 5352
rect 3936 5312 3942 5324
rect 3973 5321 3985 5324
rect 4019 5321 4031 5355
rect 3973 5315 4031 5321
rect 4617 5355 4675 5361
rect 4617 5321 4629 5355
rect 4663 5352 4675 5355
rect 5166 5352 5172 5364
rect 4663 5324 5172 5352
rect 4663 5321 4675 5324
rect 4617 5315 4675 5321
rect 5166 5312 5172 5324
rect 5224 5352 5230 5364
rect 9309 5355 9367 5361
rect 9309 5352 9321 5355
rect 5224 5324 9321 5352
rect 5224 5312 5230 5324
rect 9309 5321 9321 5324
rect 9355 5352 9367 5355
rect 9398 5352 9404 5364
rect 9355 5324 9404 5352
rect 9355 5321 9367 5324
rect 9309 5315 9367 5321
rect 9398 5312 9404 5324
rect 9456 5312 9462 5364
rect 11330 5312 11336 5364
rect 11388 5352 11394 5364
rect 12069 5355 12127 5361
rect 12069 5352 12081 5355
rect 11388 5324 12081 5352
rect 11388 5312 11394 5324
rect 12069 5321 12081 5324
rect 12115 5321 12127 5355
rect 12069 5315 12127 5321
rect 13541 5355 13599 5361
rect 13541 5321 13553 5355
rect 13587 5352 13599 5355
rect 13817 5355 13875 5361
rect 13817 5352 13829 5355
rect 13587 5324 13829 5352
rect 13587 5321 13599 5324
rect 13541 5315 13599 5321
rect 13817 5321 13829 5324
rect 13863 5352 13875 5355
rect 14458 5352 14464 5364
rect 13863 5324 14464 5352
rect 13863 5321 13875 5324
rect 13817 5315 13875 5321
rect 14458 5312 14464 5324
rect 14516 5312 14522 5364
rect 15197 5355 15255 5361
rect 15197 5321 15209 5355
rect 15243 5352 15255 5355
rect 15378 5352 15384 5364
rect 15243 5324 15384 5352
rect 15243 5321 15255 5324
rect 15197 5315 15255 5321
rect 15378 5312 15384 5324
rect 15436 5312 15442 5364
rect 17770 5352 17776 5364
rect 17731 5324 17776 5352
rect 17770 5312 17776 5324
rect 17828 5312 17834 5364
rect 18230 5352 18236 5364
rect 18191 5324 18236 5352
rect 18230 5312 18236 5324
rect 18288 5312 18294 5364
rect 19702 5352 19708 5364
rect 19663 5324 19708 5352
rect 19702 5312 19708 5324
rect 19760 5312 19766 5364
rect 19978 5312 19984 5364
rect 20036 5352 20042 5364
rect 20073 5355 20131 5361
rect 20073 5352 20085 5355
rect 20036 5324 20085 5352
rect 20036 5312 20042 5324
rect 20073 5321 20085 5324
rect 20119 5321 20131 5355
rect 21818 5352 21824 5364
rect 21779 5324 21824 5352
rect 20073 5315 20131 5321
rect 21818 5312 21824 5324
rect 21876 5312 21882 5364
rect 23198 5312 23204 5364
rect 23256 5352 23262 5364
rect 25363 5355 25421 5361
rect 25363 5352 25375 5355
rect 23256 5324 25375 5352
rect 23256 5312 23262 5324
rect 25363 5321 25375 5324
rect 25409 5321 25421 5355
rect 25363 5315 25421 5321
rect 25590 5312 25596 5364
rect 25648 5352 25654 5364
rect 25685 5355 25743 5361
rect 25685 5352 25697 5355
rect 25648 5324 25697 5352
rect 25648 5312 25654 5324
rect 25685 5321 25697 5324
rect 25731 5321 25743 5355
rect 25685 5315 25743 5321
rect 2869 5287 2927 5293
rect 2869 5253 2881 5287
rect 2915 5284 2927 5287
rect 3142 5284 3148 5296
rect 2915 5256 3148 5284
rect 2915 5253 2927 5256
rect 2869 5247 2927 5253
rect 3142 5244 3148 5256
rect 3200 5244 3206 5296
rect 3605 5287 3663 5293
rect 3605 5253 3617 5287
rect 3651 5284 3663 5287
rect 5074 5284 5080 5296
rect 3651 5256 5080 5284
rect 3651 5253 3663 5256
rect 3605 5247 3663 5253
rect 198 5108 204 5160
rect 256 5148 262 5160
rect 1432 5151 1490 5157
rect 1432 5148 1444 5151
rect 256 5120 1444 5148
rect 256 5108 262 5120
rect 1432 5117 1444 5120
rect 1478 5148 1490 5151
rect 1857 5151 1915 5157
rect 1857 5148 1869 5151
rect 1478 5120 1869 5148
rect 1478 5117 1490 5120
rect 1432 5111 1490 5117
rect 1857 5117 1869 5120
rect 1903 5117 1915 5151
rect 1857 5111 1915 5117
rect 2685 5151 2743 5157
rect 2685 5117 2697 5151
rect 2731 5148 2743 5151
rect 3620 5148 3648 5247
rect 5074 5244 5080 5256
rect 5132 5244 5138 5296
rect 6549 5287 6607 5293
rect 6549 5253 6561 5287
rect 6595 5284 6607 5287
rect 6638 5284 6644 5296
rect 6595 5256 6644 5284
rect 6595 5253 6607 5256
rect 6549 5247 6607 5253
rect 6638 5244 6644 5256
rect 6696 5244 6702 5296
rect 8018 5244 8024 5296
rect 8076 5284 8082 5296
rect 8481 5287 8539 5293
rect 8481 5284 8493 5287
rect 8076 5256 8493 5284
rect 8076 5244 8082 5256
rect 8481 5253 8493 5256
rect 8527 5284 8539 5287
rect 8757 5287 8815 5293
rect 8757 5284 8769 5287
rect 8527 5256 8769 5284
rect 8527 5253 8539 5256
rect 8481 5247 8539 5253
rect 8757 5253 8769 5256
rect 8803 5253 8815 5287
rect 8757 5247 8815 5253
rect 8846 5244 8852 5296
rect 8904 5284 8910 5296
rect 12253 5287 12311 5293
rect 12253 5284 12265 5287
rect 8904 5256 12265 5284
rect 8904 5244 8910 5256
rect 12253 5253 12265 5256
rect 12299 5253 12311 5287
rect 12253 5247 12311 5253
rect 12526 5244 12532 5296
rect 12584 5284 12590 5296
rect 19334 5284 19340 5296
rect 12584 5256 19340 5284
rect 12584 5244 12590 5256
rect 19334 5244 19340 5256
rect 19392 5244 19398 5296
rect 20254 5244 20260 5296
rect 20312 5284 20318 5296
rect 20898 5284 20904 5296
rect 20312 5256 20392 5284
rect 20859 5256 20904 5284
rect 20312 5244 20318 5256
rect 5629 5219 5687 5225
rect 5629 5185 5641 5219
rect 5675 5216 5687 5219
rect 5675 5188 6592 5216
rect 5675 5185 5687 5188
rect 5629 5179 5687 5185
rect 2731 5120 3648 5148
rect 3764 5151 3822 5157
rect 2731 5117 2743 5120
rect 2685 5111 2743 5117
rect 3764 5117 3776 5151
rect 3810 5148 3822 5151
rect 4706 5148 4712 5160
rect 3810 5120 4154 5148
rect 4667 5120 4712 5148
rect 3810 5117 3822 5120
rect 3764 5111 3822 5117
rect 4126 5080 4154 5120
rect 4706 5108 4712 5120
rect 4764 5108 4770 5160
rect 5258 5148 5264 5160
rect 5219 5120 5264 5148
rect 5258 5108 5264 5120
rect 5316 5148 5322 5160
rect 5756 5151 5814 5157
rect 5756 5148 5768 5151
rect 5316 5120 5768 5148
rect 5316 5108 5322 5120
rect 5756 5117 5768 5120
rect 5802 5117 5814 5151
rect 5756 5111 5814 5117
rect 6564 5092 6592 5188
rect 6914 5176 6920 5228
rect 6972 5216 6978 5228
rect 13541 5219 13599 5225
rect 13541 5216 13553 5219
rect 6972 5188 13553 5216
rect 6972 5176 6978 5188
rect 7466 5148 7472 5160
rect 7427 5120 7472 5148
rect 7466 5108 7472 5120
rect 7524 5108 7530 5160
rect 8113 5151 8171 5157
rect 8113 5117 8125 5151
rect 8159 5117 8171 5151
rect 8113 5111 8171 5117
rect 8941 5151 8999 5157
rect 8941 5117 8953 5151
rect 8987 5148 8999 5151
rect 9030 5148 9036 5160
rect 8987 5120 9036 5148
rect 8987 5117 8999 5120
rect 8941 5111 8999 5117
rect 4249 5083 4307 5089
rect 4249 5080 4261 5083
rect 4126 5052 4261 5080
rect 4249 5049 4261 5052
rect 4295 5080 4307 5083
rect 6178 5080 6184 5092
rect 4295 5052 6184 5080
rect 4295 5049 4307 5052
rect 4249 5043 4307 5049
rect 6178 5040 6184 5052
rect 6236 5040 6242 5092
rect 6546 5040 6552 5092
rect 6604 5080 6610 5092
rect 7377 5083 7435 5089
rect 7377 5080 7389 5083
rect 6604 5052 7389 5080
rect 6604 5040 6610 5052
rect 7377 5049 7389 5052
rect 7423 5080 7435 5083
rect 8128 5080 8156 5111
rect 9030 5108 9036 5120
rect 9088 5148 9094 5160
rect 9582 5148 9588 5160
rect 9088 5120 9588 5148
rect 9088 5108 9094 5120
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 10686 5108 10692 5160
rect 10744 5148 10750 5160
rect 10781 5151 10839 5157
rect 10781 5148 10793 5151
rect 10744 5120 10793 5148
rect 10744 5108 10750 5120
rect 10781 5117 10793 5120
rect 10827 5117 10839 5151
rect 10781 5111 10839 5117
rect 11333 5151 11391 5157
rect 11333 5117 11345 5151
rect 11379 5148 11391 5151
rect 12158 5148 12164 5160
rect 11379 5120 12164 5148
rect 11379 5117 11391 5120
rect 11333 5111 11391 5117
rect 12158 5108 12164 5120
rect 12216 5108 12222 5160
rect 12345 5151 12403 5157
rect 12345 5117 12357 5151
rect 12391 5148 12403 5151
rect 12713 5151 12771 5157
rect 12713 5148 12725 5151
rect 12391 5120 12725 5148
rect 12391 5117 12403 5120
rect 12345 5111 12403 5117
rect 12713 5117 12725 5120
rect 12759 5148 12771 5151
rect 13078 5148 13084 5160
rect 12759 5120 13084 5148
rect 12759 5117 12771 5120
rect 12713 5111 12771 5117
rect 13078 5108 13084 5120
rect 13136 5108 13142 5160
rect 13188 5157 13216 5188
rect 13541 5185 13553 5188
rect 13587 5185 13599 5219
rect 13541 5179 13599 5185
rect 14182 5176 14188 5228
rect 14240 5216 14246 5228
rect 14277 5219 14335 5225
rect 14277 5216 14289 5219
rect 14240 5188 14289 5216
rect 14240 5176 14246 5188
rect 14277 5185 14289 5188
rect 14323 5185 14335 5219
rect 16114 5216 16120 5228
rect 16075 5188 16120 5216
rect 14277 5179 14335 5185
rect 16114 5176 16120 5188
rect 16172 5176 16178 5228
rect 18785 5219 18843 5225
rect 18785 5185 18797 5219
rect 18831 5216 18843 5219
rect 19242 5216 19248 5228
rect 18831 5188 19248 5216
rect 18831 5185 18843 5188
rect 18785 5179 18843 5185
rect 19242 5176 19248 5188
rect 19300 5176 19306 5228
rect 20364 5225 20392 5256
rect 20898 5244 20904 5256
rect 20956 5244 20962 5296
rect 24670 5284 24676 5296
rect 24631 5256 24676 5284
rect 24670 5244 24676 5256
rect 24728 5244 24734 5296
rect 20349 5219 20407 5225
rect 20349 5185 20361 5219
rect 20395 5185 20407 5219
rect 20349 5179 20407 5185
rect 21174 5176 21180 5228
rect 21232 5216 21238 5228
rect 22373 5219 22431 5225
rect 22373 5216 22385 5219
rect 21232 5188 22385 5216
rect 21232 5176 21238 5188
rect 22373 5185 22385 5188
rect 22419 5216 22431 5219
rect 23842 5216 23848 5228
rect 22419 5188 23848 5216
rect 22419 5185 22431 5188
rect 22373 5179 22431 5185
rect 23842 5176 23848 5188
rect 23900 5176 23906 5228
rect 23934 5176 23940 5228
rect 23992 5216 23998 5228
rect 24029 5219 24087 5225
rect 24029 5216 24041 5219
rect 23992 5188 24041 5216
rect 23992 5176 23998 5188
rect 24029 5185 24041 5188
rect 24075 5185 24087 5219
rect 24029 5179 24087 5185
rect 13173 5151 13231 5157
rect 13173 5117 13185 5151
rect 13219 5117 13231 5151
rect 13173 5111 13231 5117
rect 13449 5151 13507 5157
rect 13449 5117 13461 5151
rect 13495 5148 13507 5151
rect 15746 5148 15752 5160
rect 13495 5120 15752 5148
rect 13495 5117 13507 5120
rect 13449 5111 13507 5117
rect 15746 5108 15752 5120
rect 15804 5108 15810 5160
rect 25292 5151 25350 5157
rect 25292 5117 25304 5151
rect 25338 5148 25350 5151
rect 25590 5148 25596 5160
rect 25338 5120 25596 5148
rect 25338 5117 25350 5120
rect 25292 5111 25350 5117
rect 25590 5108 25596 5120
rect 25648 5108 25654 5160
rect 9766 5080 9772 5092
rect 7423 5052 9772 5080
rect 7423 5049 7435 5052
rect 7377 5043 7435 5049
rect 9766 5040 9772 5052
rect 9824 5080 9830 5092
rect 10137 5083 10195 5089
rect 10137 5080 10149 5083
rect 9824 5052 10149 5080
rect 9824 5040 9830 5052
rect 10137 5049 10149 5052
rect 10183 5080 10195 5083
rect 11054 5080 11060 5092
rect 10183 5052 11060 5080
rect 10183 5049 10195 5052
rect 10137 5043 10195 5049
rect 11054 5040 11060 5052
rect 11112 5040 11118 5092
rect 11517 5083 11575 5089
rect 11517 5049 11529 5083
rect 11563 5080 11575 5083
rect 12250 5080 12256 5092
rect 11563 5052 12256 5080
rect 11563 5049 11575 5052
rect 11517 5043 11575 5049
rect 12250 5040 12256 5052
rect 12308 5040 12314 5092
rect 14598 5083 14656 5089
rect 14598 5080 14610 5083
rect 14108 5052 14610 5080
rect 4890 5012 4896 5024
rect 4851 4984 4896 5012
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 5859 5015 5917 5021
rect 5859 4981 5871 5015
rect 5905 5012 5917 5015
rect 6362 5012 6368 5024
rect 5905 4984 6368 5012
rect 5905 4981 5917 4984
rect 5859 4975 5917 4981
rect 6362 4972 6368 4984
rect 6420 4972 6426 5024
rect 8757 5015 8815 5021
rect 8757 4981 8769 5015
rect 8803 5012 8815 5015
rect 9858 5012 9864 5024
rect 8803 4984 9864 5012
rect 8803 4981 8815 4984
rect 8757 4975 8815 4981
rect 9858 4972 9864 4984
rect 9916 5012 9922 5024
rect 10042 5012 10048 5024
rect 9916 4984 10048 5012
rect 9916 4972 9922 4984
rect 10042 4972 10048 4984
rect 10100 4972 10106 5024
rect 10686 5012 10692 5024
rect 10647 4984 10692 5012
rect 10686 4972 10692 4984
rect 10744 4972 10750 5024
rect 12710 4972 12716 5024
rect 12768 5012 12774 5024
rect 14108 5021 14136 5052
rect 14598 5049 14610 5052
rect 14644 5080 14656 5083
rect 15473 5083 15531 5089
rect 15473 5080 15485 5083
rect 14644 5052 15485 5080
rect 14644 5049 14656 5052
rect 14598 5043 14656 5049
rect 15473 5049 15485 5052
rect 15519 5080 15531 5083
rect 15654 5080 15660 5092
rect 15519 5052 15660 5080
rect 15519 5049 15531 5052
rect 15473 5043 15531 5049
rect 15654 5040 15660 5052
rect 15712 5040 15718 5092
rect 16206 5040 16212 5092
rect 16264 5080 16270 5092
rect 16758 5080 16764 5092
rect 16264 5052 16357 5080
rect 16719 5052 16764 5080
rect 16264 5040 16270 5052
rect 16758 5040 16764 5052
rect 16816 5040 16822 5092
rect 18874 5040 18880 5092
rect 18932 5080 18938 5092
rect 19426 5080 19432 5092
rect 18932 5052 18977 5080
rect 19387 5052 19432 5080
rect 18932 5040 18938 5052
rect 19426 5040 19432 5052
rect 19484 5040 19490 5092
rect 20441 5083 20499 5089
rect 20441 5049 20453 5083
rect 20487 5080 20499 5083
rect 20714 5080 20720 5092
rect 20487 5052 20720 5080
rect 20487 5049 20499 5052
rect 20441 5043 20499 5049
rect 20714 5040 20720 5052
rect 20772 5040 20778 5092
rect 22094 5080 22100 5092
rect 22055 5052 22100 5080
rect 22094 5040 22100 5052
rect 22152 5040 22158 5092
rect 22189 5083 22247 5089
rect 22189 5049 22201 5083
rect 22235 5049 22247 5083
rect 23750 5080 23756 5092
rect 23711 5052 23756 5080
rect 22189 5043 22247 5049
rect 14093 5015 14151 5021
rect 14093 5012 14105 5015
rect 12768 4984 14105 5012
rect 12768 4972 12774 4984
rect 14093 4981 14105 4984
rect 14139 4981 14151 5015
rect 15838 5012 15844 5024
rect 15799 4984 15844 5012
rect 14093 4975 14151 4981
rect 15838 4972 15844 4984
rect 15896 5012 15902 5024
rect 16224 5012 16252 5040
rect 21266 5012 21272 5024
rect 15896 4984 16252 5012
rect 21227 4984 21272 5012
rect 15896 4972 15902 4984
rect 21266 4972 21272 4984
rect 21324 4972 21330 5024
rect 21818 4972 21824 5024
rect 21876 5012 21882 5024
rect 22204 5012 22232 5043
rect 23750 5040 23756 5052
rect 23808 5040 23814 5092
rect 23845 5083 23903 5089
rect 23845 5049 23857 5083
rect 23891 5049 23903 5083
rect 23845 5043 23903 5049
rect 23382 5012 23388 5024
rect 21876 4984 22232 5012
rect 23295 4984 23388 5012
rect 21876 4972 21882 4984
rect 23382 4972 23388 4984
rect 23440 5012 23446 5024
rect 23860 5012 23888 5043
rect 23440 4984 23888 5012
rect 23440 4972 23446 4984
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 3099 4811 3157 4817
rect 3099 4777 3111 4811
rect 3145 4808 3157 4811
rect 4338 4808 4344 4820
rect 3145 4780 4344 4808
rect 3145 4777 3157 4780
rect 3099 4771 3157 4777
rect 4338 4768 4344 4780
rect 4396 4768 4402 4820
rect 4433 4811 4491 4817
rect 4433 4777 4445 4811
rect 4479 4808 4491 4811
rect 4614 4808 4620 4820
rect 4479 4780 4620 4808
rect 4479 4777 4491 4780
rect 4433 4771 4491 4777
rect 4614 4768 4620 4780
rect 4672 4768 4678 4820
rect 4801 4811 4859 4817
rect 4801 4777 4813 4811
rect 4847 4808 4859 4811
rect 4982 4808 4988 4820
rect 4847 4780 4988 4808
rect 4847 4777 4859 4780
rect 4801 4771 4859 4777
rect 4982 4768 4988 4780
rect 5040 4808 5046 4820
rect 7466 4808 7472 4820
rect 5040 4780 7472 4808
rect 5040 4768 5046 4780
rect 7466 4768 7472 4780
rect 7524 4768 7530 4820
rect 7926 4808 7932 4820
rect 7887 4780 7932 4808
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 10778 4808 10784 4820
rect 8036 4780 10784 4808
rect 4632 4740 4660 4768
rect 6273 4743 6331 4749
rect 6273 4740 6285 4743
rect 4632 4712 6285 4740
rect 6273 4709 6285 4712
rect 6319 4740 6331 4743
rect 6454 4740 6460 4752
rect 6319 4712 6460 4740
rect 6319 4709 6331 4712
rect 6273 4703 6331 4709
rect 6454 4700 6460 4712
rect 6512 4700 6518 4752
rect 2866 4632 2872 4684
rect 2924 4672 2930 4684
rect 2996 4675 3054 4681
rect 2996 4672 3008 4675
rect 2924 4644 3008 4672
rect 2924 4632 2930 4644
rect 2996 4641 3008 4644
rect 3042 4641 3054 4675
rect 2996 4635 3054 4641
rect 4062 4632 4068 4684
rect 4120 4672 4126 4684
rect 4890 4672 4896 4684
rect 4120 4644 4896 4672
rect 4120 4632 4126 4644
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 5442 4672 5448 4684
rect 5403 4644 5448 4672
rect 5442 4632 5448 4644
rect 5500 4672 5506 4684
rect 6914 4672 6920 4684
rect 5500 4644 6920 4672
rect 5500 4632 5506 4644
rect 6914 4632 6920 4644
rect 6972 4632 6978 4684
rect 7098 4672 7104 4684
rect 7059 4644 7104 4672
rect 7098 4632 7104 4644
rect 7156 4632 7162 4684
rect 8036 4681 8064 4780
rect 10778 4768 10784 4780
rect 10836 4768 10842 4820
rect 10873 4811 10931 4817
rect 10873 4777 10885 4811
rect 10919 4808 10931 4811
rect 12158 4808 12164 4820
rect 10919 4780 12164 4808
rect 10919 4777 10931 4780
rect 10873 4771 10931 4777
rect 10888 4740 10916 4771
rect 12158 4768 12164 4780
rect 12216 4768 12222 4820
rect 12526 4808 12532 4820
rect 12487 4780 12532 4808
rect 12526 4768 12532 4780
rect 12584 4768 12590 4820
rect 13541 4811 13599 4817
rect 13541 4777 13553 4811
rect 13587 4808 13599 4811
rect 13814 4808 13820 4820
rect 13587 4780 13820 4808
rect 13587 4777 13599 4780
rect 13541 4771 13599 4777
rect 13814 4768 13820 4780
rect 13872 4808 13878 4820
rect 13872 4780 13917 4808
rect 13872 4768 13878 4780
rect 14182 4768 14188 4820
rect 14240 4808 14246 4820
rect 14277 4811 14335 4817
rect 14277 4808 14289 4811
rect 14240 4780 14289 4808
rect 14240 4768 14246 4780
rect 14277 4777 14289 4780
rect 14323 4777 14335 4811
rect 14277 4771 14335 4777
rect 15286 4768 15292 4820
rect 15344 4808 15350 4820
rect 15473 4811 15531 4817
rect 15473 4808 15485 4811
rect 15344 4780 15485 4808
rect 15344 4768 15350 4780
rect 15473 4777 15485 4780
rect 15519 4777 15531 4811
rect 15473 4771 15531 4777
rect 15654 4768 15660 4820
rect 15712 4808 15718 4820
rect 16758 4808 16764 4820
rect 15712 4780 16764 4808
rect 15712 4768 15718 4780
rect 16758 4768 16764 4780
rect 16816 4768 16822 4820
rect 17678 4768 17684 4820
rect 17736 4808 17742 4820
rect 18325 4811 18383 4817
rect 18325 4808 18337 4811
rect 17736 4780 18337 4808
rect 17736 4768 17742 4780
rect 18325 4777 18337 4780
rect 18371 4777 18383 4811
rect 18325 4771 18383 4777
rect 19518 4768 19524 4820
rect 19576 4808 19582 4820
rect 20162 4808 20168 4820
rect 19576 4780 20168 4808
rect 19576 4768 19582 4780
rect 20162 4768 20168 4780
rect 20220 4768 20226 4820
rect 20349 4811 20407 4817
rect 20349 4777 20361 4811
rect 20395 4808 20407 4811
rect 20714 4808 20720 4820
rect 20395 4780 20720 4808
rect 20395 4777 20407 4780
rect 20349 4771 20407 4777
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 22094 4768 22100 4820
rect 22152 4808 22158 4820
rect 22465 4811 22523 4817
rect 22465 4808 22477 4811
rect 22152 4780 22477 4808
rect 22152 4768 22158 4780
rect 22465 4777 22477 4780
rect 22511 4808 22523 4811
rect 23566 4808 23572 4820
rect 22511 4780 23572 4808
rect 22511 4777 22523 4780
rect 22465 4771 22523 4777
rect 23566 4768 23572 4780
rect 23624 4768 23630 4820
rect 24210 4808 24216 4820
rect 24171 4780 24216 4808
rect 24210 4768 24216 4780
rect 24268 4768 24274 4820
rect 8588 4712 10916 4740
rect 7561 4675 7619 4681
rect 7561 4641 7573 4675
rect 7607 4672 7619 4675
rect 8021 4675 8079 4681
rect 8021 4672 8033 4675
rect 7607 4644 8033 4672
rect 7607 4641 7619 4644
rect 7561 4635 7619 4641
rect 8021 4641 8033 4644
rect 8067 4641 8079 4675
rect 8021 4635 8079 4641
rect 8478 4632 8484 4684
rect 8536 4672 8542 4684
rect 8588 4681 8616 4712
rect 12710 4700 12716 4752
rect 12768 4740 12774 4752
rect 12942 4743 13000 4749
rect 12942 4740 12954 4743
rect 12768 4712 12954 4740
rect 12768 4700 12774 4712
rect 12942 4709 12954 4712
rect 12988 4709 13000 4743
rect 12942 4703 13000 4709
rect 15378 4700 15384 4752
rect 15436 4740 15442 4752
rect 16209 4743 16267 4749
rect 16209 4740 16221 4743
rect 15436 4712 16221 4740
rect 15436 4700 15442 4712
rect 16209 4709 16221 4712
rect 16255 4740 16267 4743
rect 16390 4740 16396 4752
rect 16255 4712 16396 4740
rect 16255 4709 16267 4712
rect 16209 4703 16267 4709
rect 16390 4700 16396 4712
rect 16448 4700 16454 4752
rect 19150 4740 19156 4752
rect 19111 4712 19156 4740
rect 19150 4700 19156 4712
rect 19208 4700 19214 4752
rect 21174 4700 21180 4752
rect 21232 4740 21238 4752
rect 21269 4743 21327 4749
rect 21269 4740 21281 4743
rect 21232 4712 21281 4740
rect 21232 4700 21238 4712
rect 21269 4709 21281 4712
rect 21315 4740 21327 4743
rect 22554 4740 22560 4752
rect 21315 4712 22560 4740
rect 21315 4709 21327 4712
rect 21269 4703 21327 4709
rect 22554 4700 22560 4712
rect 22612 4700 22618 4752
rect 22830 4740 22836 4752
rect 22791 4712 22836 4740
rect 22830 4700 22836 4712
rect 22888 4700 22894 4752
rect 24026 4700 24032 4752
rect 24084 4740 24090 4752
rect 24673 4743 24731 4749
rect 24673 4740 24685 4743
rect 24084 4712 24685 4740
rect 24084 4700 24090 4712
rect 24673 4709 24685 4712
rect 24719 4709 24731 4743
rect 24673 4703 24731 4709
rect 8573 4675 8631 4681
rect 8573 4672 8585 4675
rect 8536 4644 8585 4672
rect 8536 4632 8542 4644
rect 8573 4641 8585 4644
rect 8619 4641 8631 4675
rect 9674 4672 9680 4684
rect 9635 4644 9680 4672
rect 8573 4635 8631 4641
rect 9674 4632 9680 4644
rect 9732 4632 9738 4684
rect 9950 4672 9956 4684
rect 9911 4644 9956 4672
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 11238 4672 11244 4684
rect 11199 4644 11244 4672
rect 11238 4632 11244 4644
rect 11296 4632 11302 4684
rect 11790 4672 11796 4684
rect 11703 4644 11796 4672
rect 11790 4632 11796 4644
rect 11848 4672 11854 4684
rect 14550 4672 14556 4684
rect 11848 4644 14556 4672
rect 11848 4632 11854 4644
rect 14550 4632 14556 4644
rect 14608 4632 14614 4684
rect 14737 4675 14795 4681
rect 14737 4641 14749 4675
rect 14783 4672 14795 4675
rect 15654 4672 15660 4684
rect 14783 4644 15660 4672
rect 14783 4641 14795 4644
rect 14737 4635 14795 4641
rect 5629 4607 5687 4613
rect 5629 4573 5641 4607
rect 5675 4604 5687 4607
rect 7650 4604 7656 4616
rect 5675 4576 7656 4604
rect 5675 4573 5687 4576
rect 5629 4567 5687 4573
rect 7650 4564 7656 4576
rect 7708 4564 7714 4616
rect 8662 4604 8668 4616
rect 8623 4576 8668 4604
rect 8662 4564 8668 4576
rect 8720 4564 8726 4616
rect 10413 4607 10471 4613
rect 10413 4573 10425 4607
rect 10459 4604 10471 4607
rect 12618 4604 12624 4616
rect 10459 4576 12547 4604
rect 12579 4576 12624 4604
rect 10459 4573 10471 4576
rect 10413 4567 10471 4573
rect 4338 4496 4344 4548
rect 4396 4536 4402 4548
rect 6822 4536 6828 4548
rect 4396 4508 6828 4536
rect 4396 4496 4402 4508
rect 6822 4496 6828 4508
rect 6880 4496 6886 4548
rect 7190 4496 7196 4548
rect 7248 4536 7254 4548
rect 9769 4539 9827 4545
rect 9769 4536 9781 4539
rect 7248 4508 9781 4536
rect 7248 4496 7254 4508
rect 9769 4505 9781 4508
rect 9815 4536 9827 4539
rect 10686 4536 10692 4548
rect 9815 4508 10692 4536
rect 9815 4505 9827 4508
rect 9769 4499 9827 4505
rect 10686 4496 10692 4508
rect 10744 4496 10750 4548
rect 12519 4536 12547 4576
rect 12618 4564 12624 4576
rect 12676 4564 12682 4616
rect 14461 4607 14519 4613
rect 14461 4573 14473 4607
rect 14507 4604 14519 4607
rect 14752 4604 14780 4635
rect 15654 4632 15660 4644
rect 15712 4632 15718 4684
rect 17678 4672 17684 4684
rect 17639 4644 17684 4672
rect 17678 4632 17684 4644
rect 17736 4632 17742 4684
rect 22002 4632 22008 4684
rect 22060 4672 22066 4684
rect 22097 4675 22155 4681
rect 22097 4672 22109 4675
rect 22060 4644 22109 4672
rect 22060 4632 22066 4644
rect 22097 4641 22109 4644
rect 22143 4672 22155 4675
rect 22186 4672 22192 4684
rect 22143 4644 22192 4672
rect 22143 4641 22155 4644
rect 22097 4635 22155 4641
rect 22186 4632 22192 4644
rect 22244 4632 22250 4684
rect 16117 4607 16175 4613
rect 16117 4604 16129 4607
rect 14507 4576 14780 4604
rect 16040 4576 16129 4604
rect 14507 4573 14519 4576
rect 14461 4567 14519 4573
rect 16040 4548 16068 4576
rect 16117 4573 16129 4576
rect 16163 4573 16175 4607
rect 16117 4567 16175 4573
rect 16206 4564 16212 4616
rect 16264 4604 16270 4616
rect 16393 4607 16451 4613
rect 16393 4604 16405 4607
rect 16264 4576 16405 4604
rect 16264 4564 16270 4576
rect 16393 4573 16405 4576
rect 16439 4573 16451 4607
rect 19058 4604 19064 4616
rect 19019 4576 19064 4604
rect 16393 4567 16451 4573
rect 19058 4564 19064 4576
rect 19116 4564 19122 4616
rect 19426 4604 19432 4616
rect 19387 4576 19432 4604
rect 19426 4564 19432 4576
rect 19484 4564 19490 4616
rect 20714 4564 20720 4616
rect 20772 4604 20778 4616
rect 21177 4607 21235 4613
rect 21177 4604 21189 4607
rect 20772 4576 21189 4604
rect 20772 4564 20778 4576
rect 21177 4573 21189 4576
rect 21223 4604 21235 4607
rect 21358 4604 21364 4616
rect 21223 4576 21364 4604
rect 21223 4573 21235 4576
rect 21177 4567 21235 4573
rect 21358 4564 21364 4576
rect 21416 4564 21422 4616
rect 21453 4607 21511 4613
rect 21453 4573 21465 4607
rect 21499 4573 21511 4607
rect 21453 4567 21511 4573
rect 22741 4607 22799 4613
rect 22741 4573 22753 4607
rect 22787 4604 22799 4607
rect 23014 4604 23020 4616
rect 22787 4576 22876 4604
rect 22975 4576 23020 4604
rect 22787 4573 22799 4576
rect 22741 4567 22799 4573
rect 12519 4508 14964 4536
rect 9401 4471 9459 4477
rect 9401 4437 9413 4471
rect 9447 4468 9459 4471
rect 9490 4468 9496 4480
rect 9447 4440 9496 4468
rect 9447 4437 9459 4440
rect 9401 4431 9459 4437
rect 9490 4428 9496 4440
rect 9548 4428 9554 4480
rect 10042 4428 10048 4480
rect 10100 4468 10106 4480
rect 11425 4471 11483 4477
rect 11425 4468 11437 4471
rect 10100 4440 11437 4468
rect 10100 4428 10106 4440
rect 11425 4437 11437 4440
rect 11471 4437 11483 4471
rect 11425 4431 11483 4437
rect 13722 4428 13728 4480
rect 13780 4468 13786 4480
rect 14461 4471 14519 4477
rect 14461 4468 14473 4471
rect 13780 4440 14473 4468
rect 13780 4428 13786 4440
rect 14461 4437 14473 4440
rect 14507 4437 14519 4471
rect 14936 4468 14964 4508
rect 16022 4496 16028 4548
rect 16080 4496 16086 4548
rect 20898 4496 20904 4548
rect 20956 4536 20962 4548
rect 21468 4536 21496 4567
rect 20956 4508 21496 4536
rect 22848 4536 22876 4576
rect 23014 4564 23020 4576
rect 23072 4604 23078 4616
rect 23934 4604 23940 4616
rect 23072 4576 23940 4604
rect 23072 4564 23078 4576
rect 23934 4564 23940 4576
rect 23992 4564 23998 4616
rect 24581 4607 24639 4613
rect 24581 4573 24593 4607
rect 24627 4573 24639 4607
rect 24854 4604 24860 4616
rect 24815 4576 24860 4604
rect 24581 4567 24639 4573
rect 22922 4536 22928 4548
rect 22848 4508 22928 4536
rect 20956 4496 20962 4508
rect 22922 4496 22928 4508
rect 22980 4496 22986 4548
rect 23750 4536 23756 4548
rect 23663 4508 23756 4536
rect 23750 4496 23756 4508
rect 23808 4536 23814 4548
rect 24210 4536 24216 4548
rect 23808 4508 24216 4536
rect 23808 4496 23814 4508
rect 24210 4496 24216 4508
rect 24268 4496 24274 4548
rect 24596 4536 24624 4567
rect 24854 4564 24860 4576
rect 24912 4564 24918 4616
rect 25222 4536 25228 4548
rect 24596 4508 25228 4536
rect 25222 4496 25228 4508
rect 25280 4496 25286 4548
rect 16574 4468 16580 4480
rect 14936 4440 16580 4468
rect 14461 4431 14519 4437
rect 16574 4428 16580 4440
rect 16632 4428 16638 4480
rect 17494 4428 17500 4480
rect 17552 4468 17558 4480
rect 17865 4471 17923 4477
rect 17865 4468 17877 4471
rect 17552 4440 17877 4468
rect 17552 4428 17558 4440
rect 17865 4437 17877 4440
rect 17911 4437 17923 4471
rect 18782 4468 18788 4480
rect 18743 4440 18788 4468
rect 17865 4431 17923 4437
rect 18782 4428 18788 4440
rect 18840 4428 18846 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 3602 4264 3608 4276
rect 3563 4236 3608 4264
rect 3602 4224 3608 4236
rect 3660 4224 3666 4276
rect 4062 4264 4068 4276
rect 4023 4236 4068 4264
rect 4062 4224 4068 4236
rect 4120 4224 4126 4276
rect 5534 4224 5540 4276
rect 5592 4264 5598 4276
rect 7558 4264 7564 4276
rect 5592 4236 7564 4264
rect 5592 4224 5598 4236
rect 7558 4224 7564 4236
rect 7616 4224 7622 4276
rect 9033 4267 9091 4273
rect 9033 4233 9045 4267
rect 9079 4264 9091 4267
rect 9950 4264 9956 4276
rect 9079 4236 9956 4264
rect 9079 4233 9091 4236
rect 9033 4227 9091 4233
rect 9950 4224 9956 4236
rect 10008 4224 10014 4276
rect 10686 4264 10692 4276
rect 10647 4236 10692 4264
rect 10686 4224 10692 4236
rect 10744 4224 10750 4276
rect 10873 4267 10931 4273
rect 10873 4233 10885 4267
rect 10919 4264 10931 4267
rect 11146 4264 11152 4276
rect 10919 4236 11152 4264
rect 10919 4233 10931 4236
rect 10873 4227 10931 4233
rect 11146 4224 11152 4236
rect 11204 4224 11210 4276
rect 11425 4267 11483 4273
rect 11425 4233 11437 4267
rect 11471 4264 11483 4267
rect 12897 4267 12955 4273
rect 11471 4236 12801 4264
rect 11471 4233 11483 4236
rect 11425 4227 11483 4233
rect 9398 4196 9404 4208
rect 9359 4168 9404 4196
rect 9398 4156 9404 4168
rect 9456 4156 9462 4208
rect 9674 4156 9680 4208
rect 9732 4196 9738 4208
rect 9858 4196 9864 4208
rect 9732 4168 9864 4196
rect 9732 4156 9738 4168
rect 9858 4156 9864 4168
rect 9916 4196 9922 4208
rect 10321 4199 10379 4205
rect 10321 4196 10333 4199
rect 9916 4168 10333 4196
rect 9916 4156 9922 4168
rect 10321 4165 10333 4168
rect 10367 4165 10379 4199
rect 10321 4159 10379 4165
rect 11238 4156 11244 4208
rect 11296 4196 11302 4208
rect 11793 4199 11851 4205
rect 11793 4196 11805 4199
rect 11296 4168 11805 4196
rect 11296 4156 11302 4168
rect 11793 4165 11805 4168
rect 11839 4165 11851 4199
rect 12773 4196 12801 4236
rect 12897 4233 12909 4267
rect 12943 4264 12955 4267
rect 14366 4264 14372 4276
rect 12943 4236 14372 4264
rect 12943 4233 12955 4236
rect 12897 4227 12955 4233
rect 14366 4224 14372 4236
rect 14424 4224 14430 4276
rect 14645 4267 14703 4273
rect 14645 4233 14657 4267
rect 14691 4264 14703 4267
rect 16206 4264 16212 4276
rect 14691 4236 16212 4264
rect 14691 4233 14703 4236
rect 14645 4227 14703 4233
rect 16206 4224 16212 4236
rect 16264 4224 16270 4276
rect 16390 4264 16396 4276
rect 16351 4236 16396 4264
rect 16390 4224 16396 4236
rect 16448 4224 16454 4276
rect 17129 4267 17187 4273
rect 17129 4233 17141 4267
rect 17175 4264 17187 4267
rect 17310 4264 17316 4276
rect 17175 4236 17316 4264
rect 17175 4233 17187 4236
rect 17129 4227 17187 4233
rect 17310 4224 17316 4236
rect 17368 4224 17374 4276
rect 21174 4264 21180 4276
rect 21135 4236 21180 4264
rect 21174 4224 21180 4236
rect 21232 4224 21238 4276
rect 22557 4267 22615 4273
rect 22557 4233 22569 4267
rect 22603 4264 22615 4267
rect 22830 4264 22836 4276
rect 22603 4236 22836 4264
rect 22603 4233 22615 4236
rect 22557 4227 22615 4233
rect 22830 4224 22836 4236
rect 22888 4224 22894 4276
rect 25222 4224 25228 4276
rect 25280 4264 25286 4276
rect 25409 4267 25467 4273
rect 25409 4264 25421 4267
rect 25280 4236 25421 4264
rect 25280 4224 25286 4236
rect 25409 4233 25421 4236
rect 25455 4233 25467 4267
rect 25409 4227 25467 4233
rect 14458 4196 14464 4208
rect 12773 4168 14464 4196
rect 11793 4159 11851 4165
rect 14458 4156 14464 4168
rect 14516 4156 14522 4208
rect 22922 4156 22928 4208
rect 22980 4196 22986 4208
rect 24854 4196 24860 4208
rect 22980 4168 24860 4196
rect 22980 4156 22986 4168
rect 2866 4088 2872 4140
rect 2924 4128 2930 4140
rect 2961 4131 3019 4137
rect 2961 4128 2973 4131
rect 2924 4100 2973 4128
rect 2924 4088 2930 4100
rect 2961 4097 2973 4100
rect 3007 4097 3019 4131
rect 2961 4091 3019 4097
rect 2976 3992 3004 4091
rect 3326 4088 3332 4140
rect 3384 4128 3390 4140
rect 3694 4128 3700 4140
rect 3384 4100 3700 4128
rect 3384 4088 3390 4100
rect 3694 4088 3700 4100
rect 3752 4088 3758 4140
rect 5074 4088 5080 4140
rect 5132 4128 5138 4140
rect 7285 4131 7343 4137
rect 7285 4128 7297 4131
rect 5132 4100 7297 4128
rect 5132 4088 5138 4100
rect 7285 4097 7297 4100
rect 7331 4097 7343 4131
rect 7285 4091 7343 4097
rect 3212 4063 3270 4069
rect 3212 4029 3224 4063
rect 3258 4060 3270 4063
rect 3602 4060 3608 4072
rect 3258 4032 3608 4060
rect 3258 4029 3270 4032
rect 3212 4023 3270 4029
rect 3602 4020 3608 4032
rect 3660 4020 3666 4072
rect 4246 4069 4252 4072
rect 4224 4063 4252 4069
rect 4224 4060 4236 4063
rect 4159 4032 4236 4060
rect 4224 4029 4236 4032
rect 4304 4060 4310 4072
rect 4706 4060 4712 4072
rect 4304 4032 4712 4060
rect 4224 4023 4252 4029
rect 4246 4020 4252 4023
rect 4304 4020 4310 4032
rect 4706 4020 4712 4032
rect 4764 4020 4770 4072
rect 4982 4020 4988 4072
rect 5040 4060 5046 4072
rect 5169 4063 5227 4069
rect 5169 4060 5181 4063
rect 5040 4032 5181 4060
rect 5040 4020 5046 4032
rect 5169 4029 5181 4032
rect 5215 4029 5227 4063
rect 5718 4060 5724 4072
rect 5679 4032 5724 4060
rect 5169 4023 5227 4029
rect 5718 4020 5724 4032
rect 5776 4020 5782 4072
rect 7300 4060 7328 4091
rect 7558 4088 7564 4140
rect 7616 4128 7622 4140
rect 8478 4128 8484 4140
rect 7616 4100 8484 4128
rect 7616 4088 7622 4100
rect 7745 4063 7803 4069
rect 7745 4060 7757 4063
rect 7300 4032 7757 4060
rect 7745 4029 7757 4032
rect 7791 4060 7803 4063
rect 7926 4060 7932 4072
rect 7791 4032 7932 4060
rect 7791 4029 7803 4032
rect 7745 4023 7803 4029
rect 7926 4020 7932 4032
rect 7984 4020 7990 4072
rect 8220 4069 8248 4100
rect 8478 4088 8484 4100
rect 8536 4128 8542 4140
rect 8757 4131 8815 4137
rect 8757 4128 8769 4131
rect 8536 4100 8769 4128
rect 8536 4088 8542 4100
rect 8757 4097 8769 4100
rect 8803 4097 8815 4131
rect 12618 4128 12624 4140
rect 8757 4091 8815 4097
rect 9232 4100 12624 4128
rect 8205 4063 8263 4069
rect 8205 4060 8217 4063
rect 8183 4032 8217 4060
rect 8205 4029 8217 4032
rect 8251 4029 8263 4063
rect 8205 4023 8263 4029
rect 8662 4020 8668 4072
rect 8720 4060 8726 4072
rect 9232 4060 9260 4100
rect 12618 4088 12624 4100
rect 12676 4088 12682 4140
rect 13354 4128 13360 4140
rect 12728 4100 13360 4128
rect 8720 4032 9260 4060
rect 8720 4020 8726 4032
rect 9306 4020 9312 4072
rect 9364 4060 9370 4072
rect 9364 4032 9409 4060
rect 9364 4020 9370 4032
rect 9490 4020 9496 4072
rect 9548 4060 9554 4072
rect 9585 4063 9643 4069
rect 9585 4060 9597 4063
rect 9548 4032 9597 4060
rect 9548 4020 9554 4032
rect 9585 4029 9597 4032
rect 9631 4060 9643 4063
rect 9950 4060 9956 4072
rect 9631 4032 9956 4060
rect 9631 4029 9643 4032
rect 9585 4023 9643 4029
rect 9950 4020 9956 4032
rect 10008 4020 10014 4072
rect 10778 4020 10784 4072
rect 10836 4060 10842 4072
rect 10873 4063 10931 4069
rect 10873 4060 10885 4063
rect 10836 4032 10885 4060
rect 10836 4020 10842 4032
rect 10873 4029 10885 4032
rect 10919 4029 10931 4063
rect 10873 4023 10931 4029
rect 11241 4063 11299 4069
rect 11241 4029 11253 4063
rect 11287 4060 11299 4063
rect 12526 4060 12532 4072
rect 11287 4032 12532 4060
rect 11287 4029 11299 4032
rect 11241 4023 11299 4029
rect 12526 4020 12532 4032
rect 12584 4020 12590 4072
rect 12728 4069 12756 4100
rect 13354 4088 13360 4100
rect 13412 4088 13418 4140
rect 13446 4088 13452 4140
rect 13504 4128 13510 4140
rect 17773 4131 17831 4137
rect 17773 4128 17785 4131
rect 13504 4100 17785 4128
rect 13504 4088 13510 4100
rect 17773 4097 17785 4100
rect 17819 4128 17831 4131
rect 18325 4131 18383 4137
rect 18325 4128 18337 4131
rect 17819 4100 18337 4128
rect 17819 4097 17831 4100
rect 17773 4091 17831 4097
rect 18325 4097 18337 4100
rect 18371 4097 18383 4131
rect 18325 4091 18383 4097
rect 19426 4088 19432 4140
rect 19484 4128 19490 4140
rect 20441 4131 20499 4137
rect 20441 4128 20453 4131
rect 19484 4100 20453 4128
rect 19484 4088 19490 4100
rect 20441 4097 20453 4100
rect 20487 4097 20499 4131
rect 20441 4091 20499 4097
rect 21637 4131 21695 4137
rect 21637 4097 21649 4131
rect 21683 4128 21695 4131
rect 22186 4128 22192 4140
rect 21683 4100 22192 4128
rect 21683 4097 21695 4100
rect 21637 4091 21695 4097
rect 22186 4088 22192 4100
rect 22244 4088 22250 4140
rect 24780 4137 24808 4168
rect 24854 4156 24860 4168
rect 24912 4156 24918 4208
rect 24765 4131 24823 4137
rect 24765 4128 24777 4131
rect 24743 4100 24777 4128
rect 24765 4097 24777 4100
rect 24811 4097 24823 4131
rect 24765 4091 24823 4097
rect 12713 4063 12771 4069
rect 12713 4029 12725 4063
rect 12759 4029 12771 4063
rect 12713 4023 12771 4029
rect 16574 4020 16580 4072
rect 16632 4060 16638 4072
rect 16945 4063 17003 4069
rect 16945 4060 16957 4063
rect 16632 4032 16957 4060
rect 16632 4020 16638 4032
rect 16945 4029 16957 4032
rect 16991 4060 17003 4063
rect 17405 4063 17463 4069
rect 17405 4060 17417 4063
rect 16991 4032 17417 4060
rect 16991 4029 17003 4032
rect 16945 4023 17003 4029
rect 17405 4029 17417 4032
rect 17451 4029 17463 4063
rect 17405 4023 17463 4029
rect 19245 4063 19303 4069
rect 19245 4029 19257 4063
rect 19291 4060 19303 4063
rect 19291 4032 20024 4060
rect 19291 4029 19303 4032
rect 19245 4023 19303 4029
rect 5534 3992 5540 4004
rect 2976 3964 5540 3992
rect 5534 3952 5540 3964
rect 5592 3952 5598 4004
rect 5905 3995 5963 4001
rect 5905 3961 5917 3995
rect 5951 3992 5963 3995
rect 5994 3992 6000 4004
rect 5951 3964 6000 3992
rect 5951 3961 5963 3964
rect 5905 3955 5963 3961
rect 5994 3952 6000 3964
rect 6052 3952 6058 4004
rect 8481 3995 8539 4001
rect 8481 3961 8493 3995
rect 8527 3992 8539 3995
rect 12066 3992 12072 4004
rect 8527 3964 9260 3992
rect 8527 3961 8539 3964
rect 8481 3955 8539 3961
rect 3283 3927 3341 3933
rect 3283 3893 3295 3927
rect 3329 3924 3341 3927
rect 3786 3924 3792 3936
rect 3329 3896 3792 3924
rect 3329 3893 3341 3896
rect 3283 3887 3341 3893
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 4295 3927 4353 3933
rect 4295 3893 4307 3927
rect 4341 3924 4353 3927
rect 4522 3924 4528 3936
rect 4341 3896 4528 3924
rect 4341 3893 4353 3896
rect 4295 3887 4353 3893
rect 4522 3884 4528 3896
rect 4580 3884 4586 3936
rect 4706 3924 4712 3936
rect 4667 3896 4712 3924
rect 4706 3884 4712 3896
rect 4764 3884 4770 3936
rect 4982 3924 4988 3936
rect 4943 3896 4988 3924
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 6549 3927 6607 3933
rect 6549 3893 6561 3927
rect 6595 3924 6607 3927
rect 7098 3924 7104 3936
rect 6595 3896 7104 3924
rect 6595 3893 6607 3896
rect 6549 3887 6607 3893
rect 7098 3884 7104 3896
rect 7156 3884 7162 3936
rect 8294 3884 8300 3936
rect 8352 3924 8358 3936
rect 9033 3927 9091 3933
rect 9033 3924 9045 3927
rect 8352 3896 9045 3924
rect 8352 3884 8358 3896
rect 9033 3893 9045 3896
rect 9079 3924 9091 3927
rect 9125 3927 9183 3933
rect 9125 3924 9137 3927
rect 9079 3896 9137 3924
rect 9079 3893 9091 3896
rect 9033 3887 9091 3893
rect 9125 3893 9137 3896
rect 9171 3893 9183 3927
rect 9232 3924 9260 3964
rect 9646 3964 12072 3992
rect 9646 3924 9674 3964
rect 12066 3952 12072 3964
rect 12124 3952 12130 4004
rect 13909 3995 13967 4001
rect 13909 3992 13921 3995
rect 13786 3964 13921 3992
rect 9766 3924 9772 3936
rect 9232 3896 9674 3924
rect 9727 3896 9772 3924
rect 9125 3887 9183 3893
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 12253 3927 12311 3933
rect 12253 3893 12265 3927
rect 12299 3924 12311 3927
rect 12710 3924 12716 3936
rect 12299 3896 12716 3924
rect 12299 3893 12311 3896
rect 12253 3887 12311 3893
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 12894 3884 12900 3936
rect 12952 3924 12958 3936
rect 13633 3927 13691 3933
rect 13633 3924 13645 3927
rect 12952 3896 13645 3924
rect 12952 3884 12958 3896
rect 13633 3893 13645 3896
rect 13679 3924 13691 3927
rect 13786 3924 13814 3964
rect 13909 3961 13921 3964
rect 13955 3961 13967 3995
rect 13909 3955 13967 3961
rect 13998 3952 14004 4004
rect 14056 3992 14062 4004
rect 14550 3992 14556 4004
rect 14056 3964 14101 3992
rect 14511 3964 14556 3992
rect 14056 3952 14062 3964
rect 14550 3952 14556 3964
rect 14608 3992 14614 4004
rect 14645 3995 14703 4001
rect 14645 3992 14657 3995
rect 14608 3964 14657 3992
rect 14608 3952 14614 3964
rect 14645 3961 14657 3964
rect 14691 3961 14703 3995
rect 15473 3995 15531 4001
rect 15473 3992 15485 3995
rect 14645 3955 14703 3961
rect 14844 3964 15485 3992
rect 14844 3936 14872 3964
rect 15473 3961 15485 3964
rect 15519 3961 15531 3995
rect 15473 3955 15531 3961
rect 15565 3995 15623 4001
rect 15565 3961 15577 3995
rect 15611 3992 15623 3995
rect 15838 3992 15844 4004
rect 15611 3964 15844 3992
rect 15611 3961 15623 3964
rect 15565 3955 15623 3961
rect 14826 3924 14832 3936
rect 13679 3896 13814 3924
rect 14787 3896 14832 3924
rect 13679 3893 13691 3896
rect 13633 3887 13691 3893
rect 14826 3884 14832 3896
rect 14884 3884 14890 3936
rect 15286 3924 15292 3936
rect 15199 3896 15292 3924
rect 15286 3884 15292 3896
rect 15344 3924 15350 3936
rect 15580 3924 15608 3955
rect 15838 3952 15844 3964
rect 15896 3952 15902 4004
rect 16114 3992 16120 4004
rect 16075 3964 16120 3992
rect 16114 3952 16120 3964
rect 16172 3952 16178 4004
rect 15344 3896 15608 3924
rect 15344 3884 15350 3896
rect 16022 3884 16028 3936
rect 16080 3924 16086 3936
rect 16761 3927 16819 3933
rect 16761 3924 16773 3927
rect 16080 3896 16773 3924
rect 16080 3884 16086 3896
rect 16761 3893 16773 3896
rect 16807 3893 16819 3927
rect 16761 3887 16819 3893
rect 18598 3884 18604 3936
rect 18656 3924 18662 3936
rect 18693 3927 18751 3933
rect 18693 3924 18705 3927
rect 18656 3896 18705 3924
rect 18656 3884 18662 3896
rect 18693 3893 18705 3896
rect 18739 3893 18751 3927
rect 19518 3924 19524 3936
rect 19479 3896 19524 3924
rect 18693 3887 18751 3893
rect 19518 3884 19524 3896
rect 19576 3884 19582 3936
rect 19996 3933 20024 4032
rect 20916 4032 23474 4060
rect 20162 3992 20168 4004
rect 20123 3964 20168 3992
rect 20162 3952 20168 3964
rect 20220 3952 20226 4004
rect 20257 3995 20315 4001
rect 20257 3961 20269 3995
rect 20303 3961 20315 3995
rect 20257 3955 20315 3961
rect 19981 3927 20039 3933
rect 19981 3893 19993 3927
rect 20027 3924 20039 3927
rect 20272 3924 20300 3955
rect 20916 3924 20944 4032
rect 21958 3995 22016 4001
rect 21958 3961 21970 3995
rect 22004 3961 22016 3995
rect 21958 3955 22016 3961
rect 20027 3896 20944 3924
rect 20027 3893 20039 3896
rect 19981 3887 20039 3893
rect 21266 3884 21272 3936
rect 21324 3924 21330 3936
rect 21545 3927 21603 3933
rect 21545 3924 21557 3927
rect 21324 3896 21557 3924
rect 21324 3884 21330 3896
rect 21545 3893 21557 3896
rect 21591 3924 21603 3927
rect 21973 3924 22001 3955
rect 22094 3924 22100 3936
rect 21591 3896 22100 3924
rect 21591 3893 21603 3896
rect 21545 3887 21603 3893
rect 22094 3884 22100 3896
rect 22152 3884 22158 3936
rect 22922 3884 22928 3936
rect 22980 3924 22986 3936
rect 23201 3927 23259 3933
rect 23201 3924 23213 3927
rect 22980 3896 23213 3924
rect 22980 3884 22986 3896
rect 23201 3893 23213 3896
rect 23247 3893 23259 3927
rect 23446 3924 23474 4032
rect 23750 3952 23756 4004
rect 23808 3992 23814 4004
rect 24213 3995 24271 4001
rect 24213 3992 24225 3995
rect 23808 3964 24225 3992
rect 23808 3952 23814 3964
rect 24213 3961 24225 3964
rect 24259 3961 24271 3995
rect 24486 3992 24492 4004
rect 24447 3964 24492 3992
rect 24213 3955 24271 3961
rect 23937 3927 23995 3933
rect 23937 3924 23949 3927
rect 23446 3896 23949 3924
rect 23201 3887 23259 3893
rect 23937 3893 23949 3896
rect 23983 3924 23995 3927
rect 24026 3924 24032 3936
rect 23983 3896 24032 3924
rect 23983 3893 23995 3896
rect 23937 3887 23995 3893
rect 24026 3884 24032 3896
rect 24084 3884 24090 3936
rect 24228 3924 24256 3955
rect 24486 3952 24492 3964
rect 24544 3952 24550 4004
rect 24581 3995 24639 4001
rect 24581 3961 24593 3995
rect 24627 3961 24639 3995
rect 24581 3955 24639 3961
rect 24596 3924 24624 3955
rect 24228 3896 24624 3924
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 5718 3680 5724 3732
rect 5776 3720 5782 3732
rect 5905 3723 5963 3729
rect 5905 3720 5917 3723
rect 5776 3692 5917 3720
rect 5776 3680 5782 3692
rect 5905 3689 5917 3692
rect 5951 3689 5963 3723
rect 9398 3720 9404 3732
rect 9359 3692 9404 3720
rect 5905 3683 5963 3689
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 11422 3720 11428 3732
rect 11383 3692 11428 3720
rect 11422 3680 11428 3692
rect 11480 3680 11486 3732
rect 12066 3720 12072 3732
rect 12027 3692 12072 3720
rect 12066 3680 12072 3692
rect 12124 3680 12130 3732
rect 12802 3680 12808 3732
rect 12860 3720 12866 3732
rect 14642 3720 14648 3732
rect 12860 3692 14648 3720
rect 12860 3680 12866 3692
rect 14642 3680 14648 3692
rect 14700 3680 14706 3732
rect 18598 3720 18604 3732
rect 18559 3692 18604 3720
rect 18598 3680 18604 3692
rect 18656 3680 18662 3732
rect 19058 3680 19064 3732
rect 19116 3720 19122 3732
rect 19797 3723 19855 3729
rect 19797 3720 19809 3723
rect 19116 3692 19809 3720
rect 19116 3680 19122 3692
rect 19797 3689 19809 3692
rect 19843 3689 19855 3723
rect 20714 3720 20720 3732
rect 20675 3692 20720 3720
rect 19797 3683 19855 3689
rect 20714 3680 20720 3692
rect 20772 3680 20778 3732
rect 22094 3720 22100 3732
rect 22055 3692 22100 3720
rect 22094 3680 22100 3692
rect 22152 3680 22158 3732
rect 22649 3723 22707 3729
rect 22649 3689 22661 3723
rect 22695 3720 22707 3723
rect 23382 3720 23388 3732
rect 22695 3692 23388 3720
rect 22695 3689 22707 3692
rect 22649 3683 22707 3689
rect 23382 3680 23388 3692
rect 23440 3680 23446 3732
rect 24486 3680 24492 3732
rect 24544 3720 24550 3732
rect 24673 3723 24731 3729
rect 24673 3720 24685 3723
rect 24544 3692 24685 3720
rect 24544 3680 24550 3692
rect 24673 3689 24685 3692
rect 24719 3689 24731 3723
rect 24673 3683 24731 3689
rect 3099 3655 3157 3661
rect 3099 3621 3111 3655
rect 3145 3652 3157 3655
rect 8662 3652 8668 3664
rect 3145 3624 8668 3652
rect 3145 3621 3157 3624
rect 3099 3615 3157 3621
rect 8662 3612 8668 3624
rect 8720 3612 8726 3664
rect 8757 3655 8815 3661
rect 8757 3621 8769 3655
rect 8803 3652 8815 3655
rect 12615 3655 12673 3661
rect 8803 3624 11284 3652
rect 8803 3621 8815 3624
rect 8757 3615 8815 3621
rect 2016 3587 2074 3593
rect 2016 3553 2028 3587
rect 2062 3584 2074 3587
rect 2222 3584 2228 3596
rect 2062 3556 2228 3584
rect 2062 3553 2074 3556
rect 2016 3547 2074 3553
rect 2222 3544 2228 3556
rect 2280 3544 2286 3596
rect 2958 3584 2964 3596
rect 2919 3556 2964 3584
rect 2958 3544 2964 3556
rect 3016 3544 3022 3596
rect 5169 3587 5227 3593
rect 5169 3553 5181 3587
rect 5215 3584 5227 3587
rect 5258 3584 5264 3596
rect 5215 3556 5264 3584
rect 5215 3553 5227 3556
rect 5169 3547 5227 3553
rect 5258 3544 5264 3556
rect 5316 3544 5322 3596
rect 5445 3587 5503 3593
rect 5445 3553 5457 3587
rect 5491 3584 5503 3587
rect 5718 3584 5724 3596
rect 5491 3556 5724 3584
rect 5491 3553 5503 3556
rect 5445 3547 5503 3553
rect 3142 3476 3148 3528
rect 3200 3516 3206 3528
rect 3970 3516 3976 3528
rect 3200 3488 3976 3516
rect 3200 3476 3206 3488
rect 3970 3476 3976 3488
rect 4028 3516 4034 3528
rect 4801 3519 4859 3525
rect 4801 3516 4813 3519
rect 4028 3488 4813 3516
rect 4028 3476 4034 3488
rect 4801 3485 4813 3488
rect 4847 3516 4859 3519
rect 5460 3516 5488 3547
rect 5718 3544 5724 3556
rect 5776 3544 5782 3596
rect 7006 3584 7012 3596
rect 6967 3556 7012 3584
rect 7006 3544 7012 3556
rect 7064 3544 7070 3596
rect 7190 3584 7196 3596
rect 7151 3556 7196 3584
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 7285 3587 7343 3593
rect 7285 3553 7297 3587
rect 7331 3584 7343 3587
rect 8018 3584 8024 3596
rect 7331 3556 8024 3584
rect 7331 3553 7343 3556
rect 7285 3547 7343 3553
rect 8018 3544 8024 3556
rect 8076 3544 8082 3596
rect 8294 3584 8300 3596
rect 8255 3556 8300 3584
rect 8294 3544 8300 3556
rect 8352 3544 8358 3596
rect 9674 3584 9680 3596
rect 9635 3556 9680 3584
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 9950 3584 9956 3596
rect 9911 3556 9956 3584
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 11256 3593 11284 3624
rect 12615 3621 12627 3655
rect 12661 3652 12673 3655
rect 12710 3652 12716 3664
rect 12661 3624 12716 3652
rect 12661 3621 12673 3624
rect 12615 3615 12673 3621
rect 12710 3612 12716 3624
rect 12768 3612 12774 3664
rect 13909 3655 13967 3661
rect 13909 3621 13921 3655
rect 13955 3652 13967 3655
rect 13998 3652 14004 3664
rect 13955 3624 14004 3652
rect 13955 3621 13967 3624
rect 13909 3615 13967 3621
rect 13998 3612 14004 3624
rect 14056 3612 14062 3664
rect 15378 3612 15384 3664
rect 15436 3652 15442 3664
rect 15473 3655 15531 3661
rect 15473 3652 15485 3655
rect 15436 3624 15485 3652
rect 15436 3612 15442 3624
rect 15473 3621 15485 3624
rect 15519 3621 15531 3655
rect 15473 3615 15531 3621
rect 15746 3612 15752 3664
rect 15804 3652 15810 3664
rect 15804 3624 18276 3652
rect 15804 3612 15810 3624
rect 11241 3587 11299 3593
rect 11241 3553 11253 3587
rect 11287 3584 11299 3587
rect 11701 3587 11759 3593
rect 11701 3584 11713 3587
rect 11287 3556 11713 3584
rect 11287 3553 11299 3556
rect 11241 3547 11299 3553
rect 11701 3553 11713 3556
rect 11747 3553 11759 3587
rect 14090 3584 14096 3596
rect 14051 3556 14096 3584
rect 11701 3547 11759 3553
rect 14090 3544 14096 3556
rect 14148 3544 14154 3596
rect 15010 3584 15016 3596
rect 14971 3556 15016 3584
rect 15010 3544 15016 3556
rect 15068 3544 15074 3596
rect 17126 3584 17132 3596
rect 17087 3556 17132 3584
rect 17126 3544 17132 3556
rect 17184 3544 17190 3596
rect 18248 3593 18276 3624
rect 19334 3612 19340 3664
rect 19392 3652 19398 3664
rect 20162 3652 20168 3664
rect 19392 3624 20168 3652
rect 19392 3612 19398 3624
rect 20162 3612 20168 3624
rect 20220 3612 20226 3664
rect 23750 3652 23756 3664
rect 23446 3624 23756 3652
rect 18233 3587 18291 3593
rect 18233 3553 18245 3587
rect 18279 3584 18291 3587
rect 18966 3584 18972 3596
rect 18279 3556 18972 3584
rect 18279 3553 18291 3556
rect 18233 3547 18291 3553
rect 18966 3544 18972 3556
rect 19024 3544 19030 3596
rect 19150 3584 19156 3596
rect 19063 3556 19156 3584
rect 19150 3544 19156 3556
rect 19208 3584 19214 3596
rect 19518 3584 19524 3596
rect 19208 3556 19524 3584
rect 19208 3544 19214 3556
rect 19518 3544 19524 3556
rect 19576 3584 19582 3596
rect 23446 3584 23474 3624
rect 23750 3612 23756 3624
rect 23808 3652 23814 3664
rect 23845 3655 23903 3661
rect 23845 3652 23857 3655
rect 23808 3624 23857 3652
rect 23808 3612 23814 3624
rect 23845 3621 23857 3624
rect 23891 3621 23903 3655
rect 23845 3615 23903 3621
rect 24210 3612 24216 3664
rect 24268 3652 24274 3664
rect 24397 3655 24455 3661
rect 24397 3652 24409 3655
rect 24268 3624 24409 3652
rect 24268 3612 24274 3624
rect 24397 3621 24409 3624
rect 24443 3621 24455 3655
rect 24397 3615 24455 3621
rect 19576 3556 23474 3584
rect 19576 3544 19582 3556
rect 4847 3488 5488 3516
rect 5629 3519 5687 3525
rect 4847 3485 4859 3488
rect 4801 3479 4859 3485
rect 5629 3485 5641 3519
rect 5675 3516 5687 3519
rect 6270 3516 6276 3528
rect 5675 3488 6276 3516
rect 5675 3485 5687 3488
rect 5629 3479 5687 3485
rect 6270 3476 6276 3488
rect 6328 3476 6334 3528
rect 6362 3476 6368 3528
rect 6420 3516 6426 3528
rect 10137 3519 10195 3525
rect 10137 3516 10149 3519
rect 6420 3488 10149 3516
rect 6420 3476 6426 3488
rect 10137 3485 10149 3488
rect 10183 3485 10195 3519
rect 12250 3516 12256 3528
rect 12211 3488 12256 3516
rect 10137 3479 10195 3485
rect 12250 3476 12256 3488
rect 12308 3476 12314 3528
rect 12618 3476 12624 3528
rect 12676 3516 12682 3528
rect 13449 3519 13507 3525
rect 13449 3516 13461 3519
rect 12676 3488 13461 3516
rect 12676 3476 12682 3488
rect 13449 3485 13461 3488
rect 13495 3485 13507 3519
rect 15028 3516 15056 3544
rect 15381 3519 15439 3525
rect 15381 3516 15393 3519
rect 15028 3488 15393 3516
rect 13449 3479 13507 3485
rect 15381 3485 15393 3488
rect 15427 3485 15439 3519
rect 15381 3479 15439 3485
rect 15657 3519 15715 3525
rect 15657 3485 15669 3519
rect 15703 3516 15715 3519
rect 16114 3516 16120 3528
rect 15703 3488 16120 3516
rect 15703 3485 15715 3488
rect 15657 3479 15715 3485
rect 2087 3451 2145 3457
rect 2087 3417 2099 3451
rect 2133 3448 2145 3451
rect 6914 3448 6920 3460
rect 2133 3420 6920 3448
rect 2133 3417 2145 3420
rect 2087 3411 2145 3417
rect 6914 3408 6920 3420
rect 6972 3408 6978 3460
rect 7006 3408 7012 3460
rect 7064 3448 7070 3460
rect 7374 3448 7380 3460
rect 7064 3420 7380 3448
rect 7064 3408 7070 3420
rect 7374 3408 7380 3420
rect 7432 3448 7438 3460
rect 7929 3451 7987 3457
rect 7929 3448 7941 3451
rect 7432 3420 7941 3448
rect 7432 3408 7438 3420
rect 7929 3417 7941 3420
rect 7975 3448 7987 3451
rect 8113 3451 8171 3457
rect 8113 3448 8125 3451
rect 7975 3420 8125 3448
rect 7975 3417 7987 3420
rect 7929 3411 7987 3417
rect 8113 3417 8125 3420
rect 8159 3448 8171 3451
rect 9398 3448 9404 3460
rect 8159 3420 9404 3448
rect 8159 3417 8171 3420
rect 8113 3411 8171 3417
rect 9398 3408 9404 3420
rect 9456 3448 9462 3460
rect 9769 3451 9827 3457
rect 9769 3448 9781 3451
rect 9456 3420 9781 3448
rect 9456 3408 9462 3420
rect 9769 3417 9781 3420
rect 9815 3448 9827 3451
rect 9858 3448 9864 3460
rect 9815 3420 9864 3448
rect 9815 3417 9827 3420
rect 9769 3411 9827 3417
rect 9858 3408 9864 3420
rect 9916 3408 9922 3460
rect 10870 3448 10876 3460
rect 10783 3420 10876 3448
rect 10870 3408 10876 3420
rect 10928 3448 10934 3460
rect 15672 3448 15700 3479
rect 16114 3476 16120 3488
rect 16172 3476 16178 3528
rect 20806 3476 20812 3528
rect 20864 3516 20870 3528
rect 21729 3519 21787 3525
rect 21729 3516 21741 3519
rect 20864 3488 21741 3516
rect 20864 3476 20870 3488
rect 21729 3485 21741 3488
rect 21775 3485 21787 3519
rect 23750 3516 23756 3528
rect 21729 3479 21787 3485
rect 23446 3488 23756 3516
rect 10928 3420 15700 3448
rect 17313 3451 17371 3457
rect 10928 3408 10934 3420
rect 17313 3417 17325 3451
rect 17359 3448 17371 3451
rect 19058 3448 19064 3460
rect 17359 3420 19064 3448
rect 17359 3417 17371 3420
rect 17313 3411 17371 3417
rect 19058 3408 19064 3420
rect 19116 3408 19122 3460
rect 22462 3408 22468 3460
rect 22520 3448 22526 3460
rect 23446 3448 23474 3488
rect 23750 3476 23756 3488
rect 23808 3476 23814 3528
rect 23842 3476 23848 3528
rect 23900 3516 23906 3528
rect 25225 3519 25283 3525
rect 25225 3516 25237 3519
rect 23900 3488 25237 3516
rect 23900 3476 23906 3488
rect 25225 3485 25237 3488
rect 25271 3485 25283 3519
rect 25225 3479 25283 3485
rect 22520 3420 23474 3448
rect 22520 3408 22526 3420
rect 4890 3340 4896 3392
rect 4948 3380 4954 3392
rect 7285 3383 7343 3389
rect 7285 3380 7297 3383
rect 4948 3352 7297 3380
rect 4948 3340 4954 3352
rect 7285 3349 7297 3352
rect 7331 3349 7343 3383
rect 7558 3380 7564 3392
rect 7519 3352 7564 3380
rect 7285 3343 7343 3349
rect 7558 3340 7564 3352
rect 7616 3340 7622 3392
rect 12526 3340 12532 3392
rect 12584 3380 12590 3392
rect 13173 3383 13231 3389
rect 13173 3380 13185 3383
rect 12584 3352 13185 3380
rect 12584 3340 12590 3352
rect 13173 3349 13185 3352
rect 13219 3349 13231 3383
rect 14274 3380 14280 3392
rect 14235 3352 14280 3380
rect 13173 3343 13231 3349
rect 14274 3340 14280 3352
rect 14332 3340 14338 3392
rect 14642 3380 14648 3392
rect 14603 3352 14648 3380
rect 14642 3340 14648 3352
rect 14700 3340 14706 3392
rect 15654 3340 15660 3392
rect 15712 3380 15718 3392
rect 16301 3383 16359 3389
rect 16301 3380 16313 3383
rect 15712 3352 16313 3380
rect 15712 3340 15718 3352
rect 16301 3349 16313 3352
rect 16347 3349 16359 3383
rect 17678 3380 17684 3392
rect 17639 3352 17684 3380
rect 16301 3343 16359 3349
rect 17678 3340 17684 3352
rect 17736 3340 17742 3392
rect 19334 3340 19340 3392
rect 19392 3380 19398 3392
rect 19429 3383 19487 3389
rect 19429 3380 19441 3383
rect 19392 3352 19441 3380
rect 19392 3340 19398 3352
rect 19429 3349 19441 3352
rect 19475 3349 19487 3383
rect 21266 3380 21272 3392
rect 21227 3352 21272 3380
rect 19429 3343 19487 3349
rect 21266 3340 21272 3352
rect 21324 3340 21330 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 2271 3179 2329 3185
rect 2271 3145 2283 3179
rect 2317 3176 2329 3179
rect 3326 3176 3332 3188
rect 2317 3148 3332 3176
rect 2317 3145 2329 3148
rect 2271 3139 2329 3145
rect 3326 3136 3332 3148
rect 3384 3136 3390 3188
rect 3970 3176 3976 3188
rect 3931 3148 3976 3176
rect 3970 3136 3976 3148
rect 4028 3136 4034 3188
rect 4341 3179 4399 3185
rect 4341 3145 4353 3179
rect 4387 3176 4399 3179
rect 4982 3176 4988 3188
rect 4387 3148 4988 3176
rect 4387 3145 4399 3148
rect 4341 3139 4399 3145
rect 4982 3136 4988 3148
rect 5040 3136 5046 3188
rect 6273 3179 6331 3185
rect 6273 3145 6285 3179
rect 6319 3176 6331 3179
rect 6641 3179 6699 3185
rect 6641 3176 6653 3179
rect 6319 3148 6653 3176
rect 6319 3145 6331 3148
rect 6273 3139 6331 3145
rect 6641 3145 6653 3148
rect 6687 3176 6699 3179
rect 6687 3148 7420 3176
rect 6687 3145 6699 3148
rect 6641 3139 6699 3145
rect 7392 3120 7420 3148
rect 8018 3136 8024 3188
rect 8076 3176 8082 3188
rect 9122 3176 9128 3188
rect 8076 3148 9128 3176
rect 8076 3136 8082 3148
rect 9122 3136 9128 3148
rect 9180 3176 9186 3188
rect 9306 3176 9312 3188
rect 9180 3148 9312 3176
rect 9180 3136 9186 3148
rect 9306 3136 9312 3148
rect 9364 3176 9370 3188
rect 10778 3176 10784 3188
rect 9364 3148 10784 3176
rect 9364 3136 9370 3148
rect 10778 3136 10784 3148
rect 10836 3136 10842 3188
rect 14090 3176 14096 3188
rect 14051 3148 14096 3176
rect 14090 3136 14096 3148
rect 14148 3136 14154 3188
rect 15378 3176 15384 3188
rect 15339 3148 15384 3176
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 17126 3176 17132 3188
rect 17087 3148 17132 3176
rect 17126 3136 17132 3148
rect 17184 3136 17190 3188
rect 18785 3179 18843 3185
rect 18785 3176 18797 3179
rect 18156 3148 18797 3176
rect 5261 3111 5319 3117
rect 5261 3077 5273 3111
rect 5307 3108 5319 3111
rect 5718 3108 5724 3120
rect 5307 3080 5724 3108
rect 5307 3077 5319 3080
rect 5261 3071 5319 3077
rect 5718 3068 5724 3080
rect 5776 3108 5782 3120
rect 7190 3108 7196 3120
rect 5776 3080 7196 3108
rect 5776 3068 5782 3080
rect 7190 3068 7196 3080
rect 7248 3068 7254 3120
rect 7374 3108 7380 3120
rect 7335 3080 7380 3108
rect 7374 3068 7380 3080
rect 7432 3068 7438 3120
rect 11146 3068 11152 3120
rect 11204 3108 11210 3120
rect 13357 3111 13415 3117
rect 13357 3108 13369 3111
rect 11204 3080 13369 3108
rect 11204 3068 11210 3080
rect 13357 3077 13369 3080
rect 13403 3077 13415 3111
rect 13357 3071 13415 3077
rect 13998 3068 14004 3120
rect 14056 3108 14062 3120
rect 15105 3111 15163 3117
rect 15105 3108 15117 3111
rect 14056 3080 15117 3108
rect 14056 3068 14062 3080
rect 15105 3077 15117 3080
rect 15151 3108 15163 3111
rect 15194 3108 15200 3120
rect 15151 3080 15200 3108
rect 15151 3077 15163 3080
rect 15105 3071 15163 3077
rect 15194 3068 15200 3080
rect 15252 3108 15258 3120
rect 15749 3111 15807 3117
rect 15749 3108 15761 3111
rect 15252 3080 15761 3108
rect 15252 3068 15258 3080
rect 15749 3077 15761 3080
rect 15795 3077 15807 3111
rect 15749 3071 15807 3077
rect 4709 3043 4767 3049
rect 4709 3009 4721 3043
rect 4755 3040 4767 3043
rect 9766 3040 9772 3052
rect 4755 3012 9772 3040
rect 4755 3009 4767 3012
rect 4709 3003 4767 3009
rect 2200 2975 2258 2981
rect 2200 2941 2212 2975
rect 2246 2972 2258 2975
rect 4157 2975 4215 2981
rect 2246 2944 2636 2972
rect 2246 2941 2258 2944
rect 2200 2935 2258 2941
rect 2608 2848 2636 2944
rect 4157 2941 4169 2975
rect 4203 2972 4215 2975
rect 4724 2972 4752 3003
rect 9766 3000 9772 3012
rect 9824 3000 9830 3052
rect 10870 3040 10876 3052
rect 10831 3012 10876 3040
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 11517 3043 11575 3049
rect 11517 3009 11529 3043
rect 11563 3040 11575 3043
rect 11698 3040 11704 3052
rect 11563 3012 11704 3040
rect 11563 3009 11575 3012
rect 11517 3003 11575 3009
rect 11698 3000 11704 3012
rect 11756 3000 11762 3052
rect 12066 3000 12072 3052
rect 12124 3040 12130 3052
rect 12437 3043 12495 3049
rect 12437 3040 12449 3043
rect 12124 3012 12449 3040
rect 12124 3000 12130 3012
rect 12437 3009 12449 3012
rect 12483 3009 12495 3043
rect 12437 3003 12495 3009
rect 12710 3000 12716 3052
rect 12768 3000 12774 3052
rect 14185 3043 14243 3049
rect 14185 3009 14197 3043
rect 14231 3040 14243 3043
rect 14642 3040 14648 3052
rect 14231 3012 14648 3040
rect 14231 3009 14243 3012
rect 14185 3003 14243 3009
rect 14642 3000 14648 3012
rect 14700 3000 14706 3052
rect 15654 3000 15660 3052
rect 15712 3040 15718 3052
rect 16025 3043 16083 3049
rect 16025 3040 16037 3043
rect 15712 3012 16037 3040
rect 15712 3000 15718 3012
rect 16025 3009 16037 3012
rect 16071 3009 16083 3043
rect 16025 3003 16083 3009
rect 16114 3000 16120 3052
rect 16172 3040 16178 3052
rect 16301 3043 16359 3049
rect 16301 3040 16313 3043
rect 16172 3012 16313 3040
rect 16172 3000 16178 3012
rect 16301 3009 16313 3012
rect 16347 3009 16359 3043
rect 16301 3003 16359 3009
rect 4203 2944 4752 2972
rect 4203 2941 4215 2944
rect 4157 2935 4215 2941
rect 4890 2932 4896 2984
rect 4948 2972 4954 2984
rect 5169 2975 5227 2981
rect 5169 2972 5181 2975
rect 4948 2944 5181 2972
rect 4948 2932 4954 2944
rect 5169 2941 5181 2944
rect 5215 2941 5227 2975
rect 5169 2935 5227 2941
rect 5445 2975 5503 2981
rect 5445 2941 5457 2975
rect 5491 2972 5503 2975
rect 7285 2975 7343 2981
rect 5491 2944 7144 2972
rect 5491 2941 5503 2944
rect 5445 2935 5503 2941
rect 3050 2904 3056 2916
rect 3011 2876 3056 2904
rect 3050 2864 3056 2876
rect 3108 2864 3114 2916
rect 5077 2907 5135 2913
rect 5077 2873 5089 2907
rect 5123 2904 5135 2907
rect 5460 2904 5488 2935
rect 5123 2876 5488 2904
rect 5123 2873 5135 2876
rect 5077 2867 5135 2873
rect 2041 2839 2099 2845
rect 2041 2805 2053 2839
rect 2087 2836 2099 2839
rect 2222 2836 2228 2848
rect 2087 2808 2228 2836
rect 2087 2805 2099 2808
rect 2041 2799 2099 2805
rect 2222 2796 2228 2808
rect 2280 2796 2286 2848
rect 2590 2836 2596 2848
rect 2551 2808 2596 2836
rect 2590 2796 2596 2808
rect 2648 2796 2654 2848
rect 3142 2836 3148 2848
rect 3103 2808 3148 2836
rect 3142 2796 3148 2808
rect 3200 2796 3206 2848
rect 5626 2836 5632 2848
rect 5587 2808 5632 2836
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 7116 2836 7144 2944
rect 7285 2941 7297 2975
rect 7331 2941 7343 2975
rect 7558 2972 7564 2984
rect 7471 2944 7564 2972
rect 7285 2935 7343 2941
rect 7193 2907 7251 2913
rect 7193 2873 7205 2907
rect 7239 2904 7251 2907
rect 7300 2904 7328 2935
rect 7558 2932 7564 2944
rect 7616 2972 7622 2984
rect 8294 2972 8300 2984
rect 7616 2944 8300 2972
rect 7616 2932 7622 2944
rect 8294 2932 8300 2944
rect 8352 2972 8358 2984
rect 8389 2975 8447 2981
rect 8389 2972 8401 2975
rect 8352 2944 8401 2972
rect 8352 2932 8358 2944
rect 8389 2941 8401 2944
rect 8435 2972 8447 2975
rect 8754 2972 8760 2984
rect 8435 2944 8760 2972
rect 8435 2941 8447 2944
rect 8389 2935 8447 2941
rect 8754 2932 8760 2944
rect 8812 2932 8818 2984
rect 8941 2975 8999 2981
rect 8941 2941 8953 2975
rect 8987 2941 8999 2975
rect 8941 2935 8999 2941
rect 8956 2904 8984 2935
rect 9858 2932 9864 2984
rect 9916 2972 9922 2984
rect 10229 2975 10287 2981
rect 10229 2972 10241 2975
rect 9916 2944 10241 2972
rect 9916 2932 9922 2944
rect 10229 2941 10241 2944
rect 10275 2941 10287 2975
rect 10229 2935 10287 2941
rect 11885 2975 11943 2981
rect 11885 2941 11897 2975
rect 11931 2972 11943 2975
rect 12253 2975 12311 2981
rect 12253 2972 12265 2975
rect 11931 2944 12265 2972
rect 11931 2941 11943 2944
rect 11885 2935 11943 2941
rect 12253 2941 12265 2944
rect 12299 2972 12311 2975
rect 12728 2972 12756 3000
rect 18156 2981 18184 3148
rect 18785 3145 18797 3148
rect 18831 3176 18843 3179
rect 19242 3176 19248 3188
rect 18831 3148 19248 3176
rect 18831 3145 18843 3148
rect 18785 3139 18843 3145
rect 19242 3136 19248 3148
rect 19300 3136 19306 3188
rect 20806 3176 20812 3188
rect 20767 3148 20812 3176
rect 20806 3136 20812 3148
rect 20864 3136 20870 3188
rect 23750 3136 23756 3188
rect 23808 3176 23814 3188
rect 24673 3179 24731 3185
rect 24673 3176 24685 3179
rect 23808 3148 24685 3176
rect 23808 3136 23814 3148
rect 24673 3145 24685 3148
rect 24719 3145 24731 3179
rect 24673 3139 24731 3145
rect 25130 3136 25136 3188
rect 25188 3176 25194 3188
rect 25363 3179 25421 3185
rect 25363 3176 25375 3179
rect 25188 3148 25375 3176
rect 25188 3136 25194 3148
rect 25363 3145 25375 3148
rect 25409 3145 25421 3179
rect 25363 3139 25421 3145
rect 18325 3111 18383 3117
rect 18325 3077 18337 3111
rect 18371 3108 18383 3111
rect 19518 3108 19524 3120
rect 18371 3080 19524 3108
rect 18371 3077 18383 3080
rect 18325 3071 18383 3077
rect 19518 3068 19524 3080
rect 19576 3068 19582 3120
rect 18782 3000 18788 3052
rect 18840 3040 18846 3052
rect 22002 3040 22008 3052
rect 18840 3012 22008 3040
rect 18840 3000 18846 3012
rect 22002 3000 22008 3012
rect 22060 3040 22066 3052
rect 22462 3040 22468 3052
rect 22060 3012 22468 3040
rect 22060 3000 22066 3012
rect 18141 2975 18199 2981
rect 12299 2944 12842 2972
rect 12299 2941 12311 2944
rect 12253 2935 12311 2941
rect 7239 2876 8432 2904
rect 7239 2873 7251 2876
rect 7193 2867 7251 2873
rect 8404 2848 8432 2876
rect 8956 2876 9260 2904
rect 7558 2836 7564 2848
rect 7116 2808 7564 2836
rect 7558 2796 7564 2808
rect 7616 2796 7622 2848
rect 7742 2836 7748 2848
rect 7703 2808 7748 2836
rect 7742 2796 7748 2808
rect 7800 2796 7806 2848
rect 8386 2796 8392 2848
rect 8444 2836 8450 2848
rect 8665 2839 8723 2845
rect 8665 2836 8677 2839
rect 8444 2808 8677 2836
rect 8444 2796 8450 2808
rect 8665 2805 8677 2808
rect 8711 2836 8723 2839
rect 8956 2836 8984 2876
rect 8711 2808 8984 2836
rect 9232 2836 9260 2876
rect 9490 2864 9496 2916
rect 9548 2904 9554 2916
rect 9950 2904 9956 2916
rect 9548 2876 9956 2904
rect 9548 2864 9554 2876
rect 9950 2864 9956 2876
rect 10008 2904 10014 2916
rect 10597 2907 10655 2913
rect 10597 2904 10609 2907
rect 10008 2876 10609 2904
rect 10008 2864 10014 2876
rect 10597 2873 10609 2876
rect 10643 2873 10655 2907
rect 10597 2867 10655 2873
rect 10870 2864 10876 2916
rect 10928 2904 10934 2916
rect 10965 2907 11023 2913
rect 10965 2904 10977 2907
rect 10928 2876 10977 2904
rect 10928 2864 10934 2876
rect 10965 2873 10977 2876
rect 11011 2904 11023 2907
rect 12526 2904 12532 2916
rect 11011 2876 12532 2904
rect 11011 2873 11023 2876
rect 10965 2867 11023 2873
rect 12526 2864 12532 2876
rect 12584 2864 12590 2916
rect 12814 2913 12842 2944
rect 18141 2941 18153 2975
rect 18187 2941 18199 2975
rect 19242 2972 19248 2984
rect 19203 2944 19248 2972
rect 18141 2935 18199 2941
rect 19242 2932 19248 2944
rect 19300 2932 19306 2984
rect 21266 2972 21272 2984
rect 21227 2944 21272 2972
rect 21266 2932 21272 2944
rect 21324 2932 21330 2984
rect 22204 2981 22232 3012
rect 22462 3000 22468 3012
rect 22520 3040 22526 3052
rect 23017 3043 23075 3049
rect 23017 3040 23029 3043
rect 22520 3012 23029 3040
rect 22520 3000 22526 3012
rect 23017 3009 23029 3012
rect 23063 3009 23075 3043
rect 23017 3003 23075 3009
rect 23477 3043 23535 3049
rect 23477 3009 23489 3043
rect 23523 3040 23535 3043
rect 23753 3043 23811 3049
rect 23753 3040 23765 3043
rect 23523 3012 23765 3040
rect 23523 3009 23535 3012
rect 23477 3003 23535 3009
rect 23753 3009 23765 3012
rect 23799 3040 23811 3043
rect 23842 3040 23848 3052
rect 23799 3012 23848 3040
rect 23799 3009 23811 3012
rect 23753 3003 23811 3009
rect 22189 2975 22247 2981
rect 22189 2941 22201 2975
rect 22235 2941 22247 2975
rect 22189 2935 22247 2941
rect 12799 2907 12857 2913
rect 12799 2873 12811 2907
rect 12845 2904 12857 2907
rect 14506 2907 14564 2913
rect 14506 2904 14518 2907
rect 12845 2876 14518 2904
rect 12845 2873 12857 2876
rect 12799 2867 12857 2873
rect 13648 2848 13676 2876
rect 14506 2873 14518 2876
rect 14552 2904 14564 2907
rect 16114 2904 16120 2916
rect 14552 2876 15424 2904
rect 16075 2876 16120 2904
rect 14552 2873 14564 2876
rect 14506 2867 14564 2873
rect 9674 2836 9680 2848
rect 9232 2808 9680 2836
rect 8711 2805 8723 2808
rect 8665 2799 8723 2805
rect 9674 2796 9680 2808
rect 9732 2836 9738 2848
rect 9861 2839 9919 2845
rect 9861 2836 9873 2839
rect 9732 2808 9873 2836
rect 9732 2796 9738 2808
rect 9861 2805 9873 2808
rect 9907 2805 9919 2839
rect 13630 2836 13636 2848
rect 13591 2808 13636 2836
rect 9861 2799 9919 2805
rect 13630 2796 13636 2808
rect 13688 2796 13694 2848
rect 13998 2796 14004 2848
rect 14056 2836 14062 2848
rect 15286 2836 15292 2848
rect 14056 2808 15292 2836
rect 14056 2796 14062 2808
rect 15286 2796 15292 2808
rect 15344 2796 15350 2848
rect 15396 2836 15424 2876
rect 16114 2864 16120 2876
rect 16172 2864 16178 2916
rect 19566 2907 19624 2913
rect 19566 2873 19578 2907
rect 19612 2904 19624 2907
rect 21085 2907 21143 2913
rect 21085 2904 21097 2907
rect 19612 2876 21097 2904
rect 19612 2873 19624 2876
rect 19566 2867 19624 2873
rect 21085 2873 21097 2876
rect 21131 2904 21143 2907
rect 21590 2907 21648 2913
rect 21590 2904 21602 2907
rect 21131 2876 21602 2904
rect 21131 2873 21143 2876
rect 21085 2867 21143 2873
rect 21590 2873 21602 2876
rect 21636 2904 21648 2907
rect 22094 2904 22100 2916
rect 21636 2876 22100 2904
rect 21636 2873 21648 2876
rect 21590 2867 21648 2873
rect 17773 2839 17831 2845
rect 17773 2836 17785 2839
rect 15396 2808 17785 2836
rect 17773 2805 17785 2808
rect 17819 2836 17831 2839
rect 18598 2836 18604 2848
rect 17819 2808 18604 2836
rect 17819 2805 17831 2808
rect 17773 2799 17831 2805
rect 18598 2796 18604 2808
rect 18656 2836 18662 2848
rect 19061 2839 19119 2845
rect 19061 2836 19073 2839
rect 18656 2808 19073 2836
rect 18656 2796 18662 2808
rect 19061 2805 19073 2808
rect 19107 2836 19119 2839
rect 19581 2836 19609 2867
rect 22094 2864 22100 2876
rect 22152 2904 22158 2916
rect 22465 2907 22523 2913
rect 22465 2904 22477 2907
rect 22152 2876 22477 2904
rect 22152 2864 22158 2876
rect 22465 2873 22477 2876
rect 22511 2873 22523 2907
rect 23032 2904 23060 3003
rect 23842 3000 23848 3012
rect 23900 3000 23906 3052
rect 24210 3040 24216 3052
rect 24171 3012 24216 3040
rect 24210 3000 24216 3012
rect 24268 3000 24274 3052
rect 25292 2975 25350 2981
rect 25292 2941 25304 2975
rect 25338 2972 25350 2975
rect 25338 2944 25820 2972
rect 25338 2941 25350 2944
rect 25292 2935 25350 2941
rect 23845 2907 23903 2913
rect 23032 2876 23704 2904
rect 22465 2867 22523 2873
rect 19107 2808 19609 2836
rect 19107 2805 19119 2808
rect 19061 2799 19119 2805
rect 19978 2796 19984 2848
rect 20036 2836 20042 2848
rect 20165 2839 20223 2845
rect 20165 2836 20177 2839
rect 20036 2808 20177 2836
rect 20036 2796 20042 2808
rect 20165 2805 20177 2808
rect 20211 2805 20223 2839
rect 23676 2836 23704 2876
rect 23845 2873 23857 2907
rect 23891 2873 23903 2907
rect 23845 2867 23903 2873
rect 23860 2836 23888 2867
rect 25792 2848 25820 2944
rect 25774 2836 25780 2848
rect 23676 2808 23888 2836
rect 25735 2808 25780 2836
rect 20165 2799 20223 2805
rect 25774 2796 25780 2808
rect 25832 2796 25838 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 2087 2635 2145 2641
rect 2087 2601 2099 2635
rect 2133 2632 2145 2635
rect 3050 2632 3056 2644
rect 2133 2604 3056 2632
rect 2133 2601 2145 2604
rect 2087 2595 2145 2601
rect 3050 2592 3056 2604
rect 3108 2592 3114 2644
rect 4709 2635 4767 2641
rect 4709 2601 4721 2635
rect 4755 2632 4767 2635
rect 4890 2632 4896 2644
rect 4755 2604 4896 2632
rect 4755 2601 4767 2604
rect 4709 2595 4767 2601
rect 4890 2592 4896 2604
rect 4948 2592 4954 2644
rect 4985 2635 5043 2641
rect 4985 2601 4997 2635
rect 5031 2632 5043 2635
rect 5074 2632 5080 2644
rect 5031 2604 5080 2632
rect 5031 2601 5043 2604
rect 4985 2595 5043 2601
rect 5074 2592 5080 2604
rect 5132 2592 5138 2644
rect 5350 2632 5356 2644
rect 5311 2604 5356 2632
rect 5350 2592 5356 2604
rect 5408 2632 5414 2644
rect 5997 2635 6055 2641
rect 5997 2632 6009 2635
rect 5408 2604 6009 2632
rect 5408 2592 5414 2604
rect 5997 2601 6009 2604
rect 6043 2601 6055 2635
rect 6362 2632 6368 2644
rect 6323 2604 6368 2632
rect 5997 2595 6055 2601
rect 6362 2592 6368 2604
rect 6420 2592 6426 2644
rect 7653 2635 7711 2641
rect 7653 2601 7665 2635
rect 7699 2632 7711 2635
rect 7742 2632 7748 2644
rect 7699 2604 7748 2632
rect 7699 2601 7711 2604
rect 7653 2595 7711 2601
rect 5718 2564 5724 2576
rect 5679 2536 5724 2564
rect 5718 2524 5724 2536
rect 5776 2524 5782 2576
rect 2016 2499 2074 2505
rect 2016 2465 2028 2499
rect 2062 2496 2074 2499
rect 2498 2496 2504 2508
rect 2062 2468 2504 2496
rect 2062 2465 2074 2468
rect 2016 2459 2074 2465
rect 2498 2456 2504 2468
rect 2556 2456 2562 2508
rect 3028 2499 3086 2505
rect 3028 2465 3040 2499
rect 3074 2496 3086 2499
rect 3510 2496 3516 2508
rect 3074 2468 3516 2496
rect 3074 2465 3086 2468
rect 3028 2459 3086 2465
rect 3510 2456 3516 2468
rect 3568 2456 3574 2508
rect 4341 2499 4399 2505
rect 4341 2465 4353 2499
rect 4387 2496 4399 2499
rect 4801 2499 4859 2505
rect 4801 2496 4813 2499
rect 4387 2468 4813 2496
rect 4387 2465 4399 2468
rect 4341 2459 4399 2465
rect 4801 2465 4813 2468
rect 4847 2496 4859 2499
rect 5626 2496 5632 2508
rect 4847 2468 5632 2496
rect 4847 2465 4859 2468
rect 4801 2459 4859 2465
rect 5626 2456 5632 2468
rect 5684 2456 5690 2508
rect 5813 2499 5871 2505
rect 5813 2465 5825 2499
rect 5859 2496 5871 2499
rect 6380 2496 6408 2592
rect 5859 2468 6408 2496
rect 7101 2499 7159 2505
rect 5859 2465 5871 2468
rect 5813 2459 5871 2465
rect 7101 2465 7113 2499
rect 7147 2496 7159 2499
rect 7668 2496 7696 2595
rect 7742 2592 7748 2604
rect 7800 2592 7806 2644
rect 9122 2632 9128 2644
rect 9083 2604 9128 2632
rect 9122 2592 9128 2604
rect 9180 2592 9186 2644
rect 10045 2635 10103 2641
rect 10045 2601 10057 2635
rect 10091 2632 10103 2635
rect 12250 2632 12256 2644
rect 10091 2604 11928 2632
rect 12211 2604 12256 2632
rect 10091 2601 10103 2604
rect 10045 2595 10103 2601
rect 8849 2567 8907 2573
rect 8849 2533 8861 2567
rect 8895 2564 8907 2567
rect 9490 2564 9496 2576
rect 8895 2536 9496 2564
rect 8895 2533 8907 2536
rect 8849 2527 8907 2533
rect 9490 2524 9496 2536
rect 9548 2524 9554 2576
rect 9585 2567 9643 2573
rect 9585 2533 9597 2567
rect 9631 2564 9643 2567
rect 11146 2564 11152 2576
rect 9631 2536 11152 2564
rect 9631 2533 9643 2536
rect 9585 2527 9643 2533
rect 11146 2524 11152 2536
rect 11204 2524 11210 2576
rect 11698 2564 11704 2576
rect 11659 2536 11704 2564
rect 11698 2524 11704 2536
rect 11756 2524 11762 2576
rect 11900 2564 11928 2604
rect 12250 2592 12256 2604
rect 12308 2592 12314 2644
rect 16022 2632 16028 2644
rect 12360 2604 16028 2632
rect 12360 2564 12388 2604
rect 16022 2592 16028 2604
rect 16080 2592 16086 2644
rect 16850 2632 16856 2644
rect 16811 2604 16856 2632
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 18966 2632 18972 2644
rect 18927 2604 18972 2632
rect 18966 2592 18972 2604
rect 19024 2592 19030 2644
rect 21315 2635 21373 2641
rect 21315 2601 21327 2635
rect 21361 2632 21373 2635
rect 21634 2632 21640 2644
rect 21361 2604 21640 2632
rect 21361 2601 21373 2604
rect 21315 2595 21373 2601
rect 21634 2592 21640 2604
rect 21692 2592 21698 2644
rect 21729 2635 21787 2641
rect 21729 2601 21741 2635
rect 21775 2632 21787 2635
rect 24210 2632 24216 2644
rect 21775 2604 24216 2632
rect 21775 2601 21787 2604
rect 21729 2595 21787 2601
rect 11900 2536 12388 2564
rect 13725 2567 13783 2573
rect 13725 2533 13737 2567
rect 13771 2564 13783 2567
rect 13998 2564 14004 2576
rect 13771 2536 14004 2564
rect 13771 2533 13783 2536
rect 13725 2527 13783 2533
rect 13998 2524 14004 2536
rect 14056 2524 14062 2576
rect 14550 2564 14556 2576
rect 14511 2536 14556 2564
rect 14550 2524 14556 2536
rect 14608 2524 14614 2576
rect 15194 2564 15200 2576
rect 15155 2536 15200 2564
rect 15194 2524 15200 2536
rect 15252 2564 15258 2576
rect 15933 2567 15991 2573
rect 15933 2564 15945 2567
rect 15252 2536 15945 2564
rect 15252 2524 15258 2536
rect 15933 2533 15945 2536
rect 15979 2564 15991 2567
rect 16114 2564 16120 2576
rect 15979 2536 16120 2564
rect 15979 2533 15991 2536
rect 15933 2527 15991 2533
rect 16114 2524 16120 2536
rect 16172 2524 16178 2576
rect 16485 2567 16543 2573
rect 16485 2533 16497 2567
rect 16531 2564 16543 2567
rect 16758 2564 16764 2576
rect 16531 2536 16764 2564
rect 16531 2533 16543 2536
rect 16485 2527 16543 2533
rect 16758 2524 16764 2536
rect 16816 2524 16822 2576
rect 19429 2567 19487 2573
rect 19429 2533 19441 2567
rect 19475 2564 19487 2567
rect 19705 2567 19763 2573
rect 19705 2564 19717 2567
rect 19475 2536 19717 2564
rect 19475 2533 19487 2536
rect 19429 2527 19487 2533
rect 19705 2533 19717 2536
rect 19751 2564 19763 2567
rect 19978 2564 19984 2576
rect 19751 2536 19984 2564
rect 19751 2533 19763 2536
rect 19705 2527 19763 2533
rect 19978 2524 19984 2536
rect 20036 2524 20042 2576
rect 7147 2468 7696 2496
rect 8021 2499 8079 2505
rect 7147 2465 7159 2468
rect 7101 2459 7159 2465
rect 8021 2465 8033 2499
rect 8067 2496 8079 2499
rect 8754 2496 8760 2508
rect 8067 2468 8760 2496
rect 8067 2465 8079 2468
rect 8021 2459 8079 2465
rect 8754 2456 8760 2468
rect 8812 2456 8818 2508
rect 9861 2499 9919 2505
rect 9861 2465 9873 2499
rect 9907 2496 9919 2499
rect 10413 2499 10471 2505
rect 10413 2496 10425 2499
rect 9907 2468 10425 2496
rect 9907 2465 9919 2468
rect 9861 2459 9919 2465
rect 10413 2465 10425 2468
rect 10459 2465 10471 2499
rect 10870 2496 10876 2508
rect 10831 2468 10876 2496
rect 10413 2459 10471 2465
rect 4706 2388 4712 2440
rect 4764 2428 4770 2440
rect 9876 2428 9904 2459
rect 10870 2456 10876 2468
rect 10928 2456 10934 2508
rect 12710 2496 12716 2508
rect 12671 2468 12716 2496
rect 12710 2456 12716 2468
rect 12768 2496 12774 2508
rect 13265 2499 13323 2505
rect 13265 2496 13277 2499
rect 12768 2468 13277 2496
rect 12768 2456 12774 2468
rect 13265 2465 13277 2468
rect 13311 2465 13323 2499
rect 13265 2459 13323 2465
rect 18141 2499 18199 2505
rect 18141 2465 18153 2499
rect 18187 2496 18199 2499
rect 18414 2496 18420 2508
rect 18187 2468 18420 2496
rect 18187 2465 18199 2468
rect 18141 2459 18199 2465
rect 18414 2456 18420 2468
rect 18472 2456 18478 2508
rect 21244 2499 21302 2505
rect 21244 2465 21256 2499
rect 21290 2496 21302 2499
rect 21744 2496 21772 2595
rect 24210 2592 24216 2604
rect 24268 2592 24274 2644
rect 22002 2564 22008 2576
rect 21963 2536 22008 2564
rect 22002 2524 22008 2536
rect 22060 2524 22066 2576
rect 22278 2564 22284 2576
rect 22239 2536 22284 2564
rect 22278 2524 22284 2536
rect 22336 2524 22342 2576
rect 22373 2567 22431 2573
rect 22373 2533 22385 2567
rect 22419 2564 22431 2567
rect 22462 2564 22468 2576
rect 22419 2536 22468 2564
rect 22419 2533 22431 2536
rect 22373 2527 22431 2533
rect 22462 2524 22468 2536
rect 22520 2524 22526 2576
rect 22922 2564 22928 2576
rect 22883 2536 22928 2564
rect 22922 2524 22928 2536
rect 22980 2524 22986 2576
rect 23658 2564 23664 2576
rect 23619 2536 23664 2564
rect 23658 2524 23664 2536
rect 23716 2524 23722 2576
rect 24026 2524 24032 2576
rect 24084 2564 24090 2576
rect 24489 2567 24547 2573
rect 24489 2564 24501 2567
rect 24084 2536 24501 2564
rect 24084 2524 24090 2536
rect 24489 2533 24501 2536
rect 24535 2564 24547 2567
rect 25317 2567 25375 2573
rect 25317 2564 25329 2567
rect 24535 2536 25329 2564
rect 24535 2533 24547 2536
rect 24489 2527 24547 2533
rect 25317 2533 25329 2536
rect 25363 2533 25375 2567
rect 25317 2527 25375 2533
rect 21290 2468 21772 2496
rect 21290 2465 21302 2468
rect 21244 2459 21302 2465
rect 4764 2400 9904 2428
rect 11057 2431 11115 2437
rect 4764 2388 4770 2400
rect 11057 2397 11069 2431
rect 11103 2428 11115 2431
rect 11790 2428 11796 2440
rect 11103 2400 11796 2428
rect 11103 2397 11115 2400
rect 11057 2391 11115 2397
rect 11790 2388 11796 2400
rect 11848 2388 11854 2440
rect 13909 2431 13967 2437
rect 13909 2397 13921 2431
rect 13955 2397 13967 2431
rect 13909 2391 13967 2397
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2428 14979 2431
rect 15841 2431 15899 2437
rect 15841 2428 15853 2431
rect 14967 2400 15853 2428
rect 14967 2397 14979 2400
rect 14921 2391 14979 2397
rect 15841 2397 15853 2400
rect 15887 2428 15899 2431
rect 15930 2428 15936 2440
rect 15887 2400 15936 2428
rect 15887 2397 15899 2400
rect 15841 2391 15899 2397
rect 7285 2363 7343 2369
rect 7285 2329 7297 2363
rect 7331 2360 7343 2363
rect 8846 2360 8852 2372
rect 7331 2332 8852 2360
rect 7331 2329 7343 2332
rect 7285 2323 7343 2329
rect 8846 2320 8852 2332
rect 8904 2320 8910 2372
rect 13924 2360 13952 2391
rect 15930 2388 15936 2400
rect 15988 2388 15994 2440
rect 19426 2388 19432 2440
rect 19484 2428 19490 2440
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 19484 2400 19625 2428
rect 19484 2388 19490 2400
rect 19613 2397 19625 2400
rect 19659 2428 19671 2431
rect 20533 2431 20591 2437
rect 20533 2428 20545 2431
rect 19659 2400 20545 2428
rect 19659 2397 19671 2400
rect 19613 2391 19671 2397
rect 20533 2397 20545 2400
rect 20579 2397 20591 2431
rect 20533 2391 20591 2397
rect 22278 2388 22284 2440
rect 22336 2428 22342 2440
rect 23201 2431 23259 2437
rect 23201 2428 23213 2431
rect 22336 2400 23213 2428
rect 22336 2388 22342 2400
rect 23201 2397 23213 2400
rect 23247 2397 23259 2431
rect 24397 2431 24455 2437
rect 24397 2428 24409 2431
rect 23201 2391 23259 2397
rect 23446 2400 24409 2428
rect 16850 2360 16856 2372
rect 13924 2332 16856 2360
rect 16850 2320 16856 2332
rect 16908 2320 16914 2372
rect 18601 2363 18659 2369
rect 18601 2329 18613 2363
rect 18647 2360 18659 2363
rect 20162 2360 20168 2372
rect 18647 2332 19748 2360
rect 20123 2332 20168 2360
rect 18647 2329 18659 2332
rect 18601 2323 18659 2329
rect 2498 2292 2504 2304
rect 2459 2264 2504 2292
rect 2498 2252 2504 2264
rect 2556 2252 2562 2304
rect 3099 2295 3157 2301
rect 3099 2261 3111 2295
rect 3145 2292 3157 2295
rect 3326 2292 3332 2304
rect 3145 2264 3332 2292
rect 3145 2261 3157 2264
rect 3099 2255 3157 2261
rect 3326 2252 3332 2264
rect 3384 2252 3390 2304
rect 3510 2292 3516 2304
rect 3471 2264 3516 2292
rect 3510 2252 3516 2264
rect 3568 2252 3574 2304
rect 12894 2292 12900 2304
rect 12855 2264 12900 2292
rect 12894 2252 12900 2264
rect 12952 2252 12958 2304
rect 19720 2292 19748 2332
rect 20162 2320 20168 2332
rect 20220 2360 20226 2372
rect 23014 2360 23020 2372
rect 20220 2332 23020 2360
rect 20220 2320 20226 2332
rect 23014 2320 23020 2332
rect 23072 2320 23078 2372
rect 20254 2292 20260 2304
rect 19720 2264 20260 2292
rect 20254 2252 20260 2264
rect 20312 2252 20318 2304
rect 22646 2252 22652 2304
rect 22704 2292 22710 2304
rect 23446 2292 23474 2400
rect 24397 2397 24409 2400
rect 24443 2428 24455 2431
rect 25685 2431 25743 2437
rect 25685 2428 25697 2431
rect 24443 2400 25697 2428
rect 24443 2397 24455 2400
rect 24397 2391 24455 2397
rect 25685 2397 25697 2400
rect 25731 2397 25743 2431
rect 25685 2391 25743 2397
rect 24302 2320 24308 2372
rect 24360 2360 24366 2372
rect 24949 2363 25007 2369
rect 24949 2360 24961 2363
rect 24360 2332 24961 2360
rect 24360 2320 24366 2332
rect 24949 2329 24961 2332
rect 24995 2329 25007 2363
rect 24949 2323 25007 2329
rect 22704 2264 23474 2292
rect 22704 2252 22710 2264
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 4430 76 4436 128
rect 4488 116 4494 128
rect 4982 116 4988 128
rect 4488 88 4988 116
rect 4488 76 4494 88
rect 4982 76 4988 88
rect 5040 76 5046 128
rect 9582 76 9588 128
rect 9640 116 9646 128
rect 10410 116 10416 128
rect 9640 88 10416 116
rect 9640 76 9646 88
rect 10410 76 10416 88
rect 10468 76 10474 128
rect 12894 76 12900 128
rect 12952 116 12958 128
rect 15102 116 15108 128
rect 12952 88 15108 116
rect 12952 76 12958 88
rect 15102 76 15108 88
rect 15160 76 15166 128
rect 26142 76 26148 128
rect 26200 116 26206 128
rect 26786 116 26792 128
rect 26200 88 26792 116
rect 26200 76 26206 88
rect 26786 76 26792 88
rect 26844 76 26850 128
rect 14274 8 14280 60
rect 14332 48 14338 60
rect 18230 48 18236 60
rect 14332 20 18236 48
rect 14332 8 14338 20
rect 18230 8 18236 20
rect 18288 8 18294 60
rect 26234 8 26240 60
rect 26292 48 26298 60
rect 27522 48 27528 60
rect 26292 20 27528 48
rect 26292 8 26298 20
rect 27522 8 27528 20
rect 27580 8 27586 60
<< via1 >>
rect 2228 27480 2280 27532
rect 3424 27480 3476 27532
rect 14372 27480 14424 27532
rect 16212 27480 16264 27532
rect 756 26732 808 26784
rect 2780 26732 2832 26784
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 27160 24896 27212 24948
rect 24124 24692 24176 24744
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 24768 24395 24820 24404
rect 24768 24361 24777 24395
rect 24777 24361 24811 24395
rect 24811 24361 24820 24395
rect 24768 24352 24820 24361
rect 23848 24216 23900 24268
rect 24676 24216 24728 24268
rect 25596 24080 25648 24132
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 14740 23808 14792 23860
rect 17776 23808 17828 23860
rect 19340 23808 19392 23860
rect 20904 23808 20956 23860
rect 24032 23808 24084 23860
rect 24952 23808 25004 23860
rect 22468 23740 22520 23792
rect 23848 23783 23900 23792
rect 23848 23749 23857 23783
rect 23857 23749 23891 23783
rect 23891 23749 23900 23783
rect 23848 23740 23900 23749
rect 1860 23647 1912 23656
rect 1860 23613 1869 23647
rect 1869 23613 1903 23647
rect 1903 23613 1912 23647
rect 1860 23604 1912 23613
rect 12716 23604 12768 23656
rect 15384 23604 15436 23656
rect 17224 23604 17276 23656
rect 19524 23604 19576 23656
rect 22008 23647 22060 23656
rect 7104 23536 7156 23588
rect 19340 23536 19392 23588
rect 22008 23613 22017 23647
rect 22017 23613 22051 23647
rect 22051 23613 22060 23647
rect 22008 23604 22060 23613
rect 22652 23536 22704 23588
rect 24676 23536 24728 23588
rect 22744 23468 22796 23520
rect 23848 23468 23900 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 24768 23307 24820 23316
rect 24768 23273 24777 23307
rect 24777 23273 24811 23307
rect 24811 23273 24820 23307
rect 24768 23264 24820 23273
rect 24032 23128 24084 23180
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 24032 22380 24084 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 24768 22219 24820 22228
rect 24768 22185 24777 22219
rect 24777 22185 24811 22219
rect 24811 22185 24820 22219
rect 24768 22176 24820 22185
rect 7104 22108 7156 22160
rect 11980 22108 12032 22160
rect 9588 22083 9640 22092
rect 9588 22049 9597 22083
rect 9597 22049 9631 22083
rect 9631 22049 9640 22083
rect 9588 22040 9640 22049
rect 24216 22040 24268 22092
rect 18604 21836 18656 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 8944 21428 8996 21480
rect 14740 21632 14792 21684
rect 22008 21632 22060 21684
rect 8576 21360 8628 21412
rect 9588 21360 9640 21412
rect 10048 21292 10100 21344
rect 14096 21292 14148 21344
rect 24216 21292 24268 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 4896 20952 4948 21004
rect 11612 20952 11664 21004
rect 13176 20952 13228 21004
rect 10140 20884 10192 20936
rect 13636 20884 13688 20936
rect 4712 20748 4764 20800
rect 10692 20748 10744 20800
rect 13452 20748 13504 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 4896 20587 4948 20596
rect 4896 20553 4905 20587
rect 4905 20553 4939 20587
rect 4939 20553 4948 20587
rect 4896 20544 4948 20553
rect 11612 20587 11664 20596
rect 11612 20553 11621 20587
rect 11621 20553 11655 20587
rect 11655 20553 11664 20587
rect 11612 20544 11664 20553
rect 13176 20544 13228 20596
rect 10692 20451 10744 20460
rect 10692 20417 10701 20451
rect 10701 20417 10735 20451
rect 10735 20417 10744 20451
rect 10692 20408 10744 20417
rect 4436 20340 4488 20392
rect 10232 20340 10284 20392
rect 11704 20272 11756 20324
rect 9956 20204 10008 20256
rect 10692 20204 10744 20256
rect 12256 20204 12308 20256
rect 13728 20383 13780 20392
rect 13728 20349 13737 20383
rect 13737 20349 13771 20383
rect 13771 20349 13780 20383
rect 13728 20340 13780 20349
rect 15292 20340 15344 20392
rect 13820 20315 13872 20324
rect 13820 20281 13829 20315
rect 13829 20281 13863 20315
rect 13863 20281 13872 20315
rect 13820 20272 13872 20281
rect 13360 20204 13412 20256
rect 14648 20204 14700 20256
rect 15844 20247 15896 20256
rect 15844 20213 15853 20247
rect 15853 20213 15887 20247
rect 15887 20213 15896 20247
rect 15844 20204 15896 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 13452 20043 13504 20052
rect 13452 20009 13461 20043
rect 13461 20009 13495 20043
rect 13495 20009 13504 20043
rect 13452 20000 13504 20009
rect 10232 19975 10284 19984
rect 10232 19941 10241 19975
rect 10241 19941 10275 19975
rect 10275 19941 10284 19975
rect 10232 19932 10284 19941
rect 11888 19932 11940 19984
rect 25228 20000 25280 20052
rect 13820 19975 13872 19984
rect 13820 19941 13829 19975
rect 13829 19941 13863 19975
rect 13863 19941 13872 19975
rect 13820 19932 13872 19941
rect 15936 19907 15988 19916
rect 15936 19873 15945 19907
rect 15945 19873 15979 19907
rect 15979 19873 15988 19907
rect 15936 19864 15988 19873
rect 24676 19864 24728 19916
rect 11704 19839 11756 19848
rect 10048 19660 10100 19712
rect 11704 19805 11713 19839
rect 11713 19805 11747 19839
rect 11747 19805 11756 19839
rect 11704 19796 11756 19805
rect 14464 19796 14516 19848
rect 15292 19839 15344 19848
rect 15292 19805 15301 19839
rect 15301 19805 15335 19839
rect 15335 19805 15344 19839
rect 15292 19796 15344 19805
rect 12256 19771 12308 19780
rect 12256 19737 12265 19771
rect 12265 19737 12299 19771
rect 12299 19737 12308 19771
rect 12256 19728 12308 19737
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 10140 19456 10192 19508
rect 10232 19252 10284 19304
rect 10692 19320 10744 19372
rect 11704 19456 11756 19508
rect 13544 19456 13596 19508
rect 13820 19456 13872 19508
rect 15936 19499 15988 19508
rect 15936 19465 15945 19499
rect 15945 19465 15979 19499
rect 15979 19465 15988 19499
rect 15936 19456 15988 19465
rect 13636 19320 13688 19372
rect 24676 19320 24728 19372
rect 11612 19184 11664 19236
rect 13544 19227 13596 19236
rect 13544 19193 13553 19227
rect 13553 19193 13587 19227
rect 13587 19193 13596 19227
rect 13544 19184 13596 19193
rect 15016 19227 15068 19236
rect 15016 19193 15025 19227
rect 15025 19193 15059 19227
rect 15059 19193 15068 19227
rect 15016 19184 15068 19193
rect 11336 19116 11388 19168
rect 11888 19116 11940 19168
rect 13084 19116 13136 19168
rect 15292 19184 15344 19236
rect 15660 19227 15712 19236
rect 15660 19193 15669 19227
rect 15669 19193 15703 19227
rect 15703 19193 15712 19227
rect 15660 19184 15712 19193
rect 15384 19116 15436 19168
rect 16672 19116 16724 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 11612 18887 11664 18896
rect 11612 18853 11621 18887
rect 11621 18853 11655 18887
rect 11655 18853 11664 18887
rect 11612 18844 11664 18853
rect 13636 18912 13688 18964
rect 15016 18955 15068 18964
rect 15016 18921 15025 18955
rect 15025 18921 15059 18955
rect 15059 18921 15068 18955
rect 15016 18912 15068 18921
rect 15936 18912 15988 18964
rect 11796 18844 11848 18896
rect 12256 18887 12308 18896
rect 12256 18853 12265 18887
rect 12265 18853 12299 18887
rect 12299 18853 12308 18887
rect 12256 18844 12308 18853
rect 13728 18844 13780 18896
rect 13820 18887 13872 18896
rect 13820 18853 13829 18887
rect 13829 18853 13863 18887
rect 13863 18853 13872 18887
rect 15476 18887 15528 18896
rect 13820 18844 13872 18853
rect 15476 18853 15485 18887
rect 15485 18853 15519 18887
rect 15519 18853 15528 18887
rect 15476 18844 15528 18853
rect 9680 18776 9732 18828
rect 3424 18708 3476 18760
rect 4252 18708 4304 18760
rect 9956 18708 10008 18760
rect 10876 18708 10928 18760
rect 14464 18776 14516 18828
rect 11888 18708 11940 18760
rect 13728 18751 13780 18760
rect 13728 18717 13737 18751
rect 13737 18717 13771 18751
rect 13771 18717 13780 18751
rect 13728 18708 13780 18717
rect 14648 18708 14700 18760
rect 15384 18751 15436 18760
rect 15384 18717 15393 18751
rect 15393 18717 15427 18751
rect 15427 18717 15436 18751
rect 15384 18708 15436 18717
rect 15660 18751 15712 18760
rect 15660 18717 15669 18751
rect 15669 18717 15703 18751
rect 15703 18717 15712 18751
rect 15660 18708 15712 18717
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 9680 18411 9732 18420
rect 9680 18377 9689 18411
rect 9689 18377 9723 18411
rect 9723 18377 9732 18411
rect 9680 18368 9732 18377
rect 10048 18368 10100 18420
rect 10140 18368 10192 18420
rect 11796 18411 11848 18420
rect 4252 18300 4304 18352
rect 7472 18275 7524 18284
rect 7472 18241 7481 18275
rect 7481 18241 7515 18275
rect 7515 18241 7524 18275
rect 7472 18232 7524 18241
rect 8944 18275 8996 18284
rect 8944 18241 8953 18275
rect 8953 18241 8987 18275
rect 8987 18241 8996 18275
rect 8944 18232 8996 18241
rect 2044 18164 2096 18216
rect 8300 18139 8352 18148
rect 8300 18105 8309 18139
rect 8309 18105 8343 18139
rect 8343 18105 8352 18139
rect 8300 18096 8352 18105
rect 11796 18377 11805 18411
rect 11805 18377 11839 18411
rect 11839 18377 11848 18411
rect 11796 18368 11848 18377
rect 13728 18368 13780 18420
rect 15476 18368 15528 18420
rect 14832 18343 14884 18352
rect 14832 18309 14841 18343
rect 14841 18309 14875 18343
rect 14875 18309 14884 18343
rect 14832 18300 14884 18309
rect 15384 18300 15436 18352
rect 10876 18275 10928 18284
rect 10876 18241 10885 18275
rect 10885 18241 10919 18275
rect 10919 18241 10928 18275
rect 10876 18232 10928 18241
rect 11612 18232 11664 18284
rect 14096 18232 14148 18284
rect 14464 18232 14516 18284
rect 13636 18207 13688 18216
rect 13636 18173 13645 18207
rect 13645 18173 13679 18207
rect 13679 18173 13688 18207
rect 13636 18164 13688 18173
rect 16212 18164 16264 18216
rect 7196 18028 7248 18080
rect 7472 18028 7524 18080
rect 11336 18096 11388 18148
rect 14280 18096 14332 18148
rect 13820 18028 13872 18080
rect 16028 18071 16080 18080
rect 16028 18037 16037 18071
rect 16037 18037 16071 18071
rect 16071 18037 16080 18071
rect 16028 18028 16080 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 7196 17824 7248 17876
rect 11336 17867 11388 17876
rect 11336 17833 11345 17867
rect 11345 17833 11379 17867
rect 11379 17833 11388 17867
rect 11336 17824 11388 17833
rect 12532 17867 12584 17876
rect 12532 17833 12541 17867
rect 12541 17833 12575 17867
rect 12575 17833 12584 17867
rect 12532 17824 12584 17833
rect 13084 17867 13136 17876
rect 13084 17833 13093 17867
rect 13093 17833 13127 17867
rect 13127 17833 13136 17867
rect 13084 17824 13136 17833
rect 14096 17867 14148 17876
rect 14096 17833 14105 17867
rect 14105 17833 14139 17867
rect 14139 17833 14148 17867
rect 14096 17824 14148 17833
rect 14464 17867 14516 17876
rect 14464 17833 14473 17867
rect 14473 17833 14507 17867
rect 14507 17833 14516 17867
rect 14464 17824 14516 17833
rect 7380 17799 7432 17808
rect 7380 17765 7389 17799
rect 7389 17765 7423 17799
rect 7423 17765 7432 17799
rect 7380 17756 7432 17765
rect 9772 17756 9824 17808
rect 13820 17756 13872 17808
rect 15384 17799 15436 17808
rect 15384 17765 15393 17799
rect 15393 17765 15427 17799
rect 15427 17765 15436 17799
rect 15384 17756 15436 17765
rect 16028 17756 16080 17808
rect 17040 17799 17092 17808
rect 17040 17765 17049 17799
rect 17049 17765 17083 17799
rect 17083 17765 17092 17799
rect 17040 17756 17092 17765
rect 5080 17688 5132 17740
rect 13360 17688 13412 17740
rect 13912 17731 13964 17740
rect 13912 17697 13921 17731
rect 13921 17697 13955 17731
rect 13955 17697 13964 17731
rect 13912 17688 13964 17697
rect 7288 17663 7340 17672
rect 7288 17629 7297 17663
rect 7297 17629 7331 17663
rect 7331 17629 7340 17663
rect 7288 17620 7340 17629
rect 7656 17663 7708 17672
rect 7656 17629 7665 17663
rect 7665 17629 7699 17663
rect 7699 17629 7708 17663
rect 7656 17620 7708 17629
rect 8300 17620 8352 17672
rect 11428 17620 11480 17672
rect 8116 17484 8168 17536
rect 8944 17527 8996 17536
rect 8944 17493 8953 17527
rect 8953 17493 8987 17527
rect 8987 17493 8996 17527
rect 8944 17484 8996 17493
rect 11796 17484 11848 17536
rect 16764 17620 16816 17672
rect 17592 17663 17644 17672
rect 17592 17629 17601 17663
rect 17601 17629 17635 17663
rect 17635 17629 17644 17663
rect 17592 17620 17644 17629
rect 14280 17552 14332 17604
rect 16488 17552 16540 17604
rect 22744 17484 22796 17536
rect 23940 17484 23992 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 5080 17323 5132 17332
rect 5080 17289 5089 17323
rect 5089 17289 5123 17323
rect 5123 17289 5132 17323
rect 5080 17280 5132 17289
rect 6828 17280 6880 17332
rect 7288 17280 7340 17332
rect 13820 17323 13872 17332
rect 13820 17289 13829 17323
rect 13829 17289 13863 17323
rect 13863 17289 13872 17323
rect 13820 17280 13872 17289
rect 15476 17280 15528 17332
rect 16212 17323 16264 17332
rect 16212 17289 16221 17323
rect 16221 17289 16255 17323
rect 16255 17289 16264 17323
rect 16212 17280 16264 17289
rect 17040 17280 17092 17332
rect 25412 17280 25464 17332
rect 6736 17212 6788 17264
rect 16028 17212 16080 17264
rect 17776 17212 17828 17264
rect 7196 17144 7248 17196
rect 8300 17144 8352 17196
rect 8944 17187 8996 17196
rect 8944 17153 8953 17187
rect 8953 17153 8987 17187
rect 8987 17153 8996 17187
rect 8944 17144 8996 17153
rect 9036 17144 9088 17196
rect 16488 17187 16540 17196
rect 12532 17076 12584 17128
rect 7288 16940 7340 16992
rect 9220 17008 9272 17060
rect 11152 17008 11204 17060
rect 13820 17076 13872 17128
rect 16488 17153 16497 17187
rect 16497 17153 16531 17187
rect 16531 17153 16540 17187
rect 16488 17144 16540 17153
rect 16764 17187 16816 17196
rect 16764 17153 16773 17187
rect 16773 17153 16807 17187
rect 16807 17153 16816 17187
rect 16764 17144 16816 17153
rect 14648 17119 14700 17128
rect 14648 17085 14657 17119
rect 14657 17085 14691 17119
rect 14691 17085 14700 17119
rect 14648 17076 14700 17085
rect 24216 17076 24268 17128
rect 14556 17051 14608 17060
rect 14556 17017 14565 17051
rect 14565 17017 14599 17051
rect 14599 17017 14608 17051
rect 14556 17008 14608 17017
rect 8392 16983 8444 16992
rect 8392 16949 8401 16983
rect 8401 16949 8435 16983
rect 8435 16949 8444 16983
rect 8392 16940 8444 16949
rect 9772 16940 9824 16992
rect 10784 16983 10836 16992
rect 10784 16949 10793 16983
rect 10793 16949 10827 16983
rect 10827 16949 10836 16983
rect 10784 16940 10836 16949
rect 11428 16940 11480 16992
rect 11888 16983 11940 16992
rect 11888 16949 11897 16983
rect 11897 16949 11931 16983
rect 11931 16949 11940 16983
rect 11888 16940 11940 16949
rect 16212 16940 16264 16992
rect 18052 16983 18104 16992
rect 18052 16949 18061 16983
rect 18061 16949 18095 16983
rect 18095 16949 18104 16983
rect 18052 16940 18104 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 7472 16668 7524 16720
rect 7748 16711 7800 16720
rect 7748 16677 7757 16711
rect 7757 16677 7791 16711
rect 7791 16677 7800 16711
rect 7748 16668 7800 16677
rect 8300 16711 8352 16720
rect 8300 16677 8309 16711
rect 8309 16677 8343 16711
rect 8343 16677 8352 16711
rect 8300 16668 8352 16677
rect 6644 16643 6696 16652
rect 6644 16609 6653 16643
rect 6653 16609 6687 16643
rect 6687 16609 6696 16643
rect 6644 16600 6696 16609
rect 10140 16600 10192 16652
rect 10416 16643 10468 16652
rect 10416 16609 10425 16643
rect 10425 16609 10459 16643
rect 10459 16609 10468 16643
rect 10416 16600 10468 16609
rect 14648 16779 14700 16788
rect 11796 16668 11848 16720
rect 11888 16668 11940 16720
rect 12624 16668 12676 16720
rect 12808 16643 12860 16652
rect 7472 16532 7524 16584
rect 10784 16532 10836 16584
rect 12808 16609 12817 16643
rect 12817 16609 12851 16643
rect 12851 16609 12860 16643
rect 12808 16600 12860 16609
rect 14648 16745 14657 16779
rect 14657 16745 14691 16779
rect 14691 16745 14700 16779
rect 14648 16736 14700 16745
rect 15384 16736 15436 16788
rect 16764 16736 16816 16788
rect 13912 16668 13964 16720
rect 16212 16668 16264 16720
rect 17776 16668 17828 16720
rect 13636 16600 13688 16652
rect 7288 16439 7340 16448
rect 7288 16405 7297 16439
rect 7297 16405 7331 16439
rect 7331 16405 7340 16439
rect 7288 16396 7340 16405
rect 8668 16439 8720 16448
rect 8668 16405 8677 16439
rect 8677 16405 8711 16439
rect 8711 16405 8720 16439
rect 8668 16396 8720 16405
rect 11704 16396 11756 16448
rect 17040 16532 17092 16584
rect 18052 16532 18104 16584
rect 18512 16532 18564 16584
rect 17132 16464 17184 16516
rect 13452 16396 13504 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 6644 16235 6696 16244
rect 6644 16201 6653 16235
rect 6653 16201 6687 16235
rect 6687 16201 6696 16235
rect 6644 16192 6696 16201
rect 7748 16192 7800 16244
rect 9220 16235 9272 16244
rect 9220 16201 9229 16235
rect 9229 16201 9263 16235
rect 9263 16201 9272 16235
rect 9220 16192 9272 16201
rect 16212 16235 16264 16244
rect 16212 16201 16221 16235
rect 16221 16201 16255 16235
rect 16255 16201 16264 16235
rect 16212 16192 16264 16201
rect 17776 16235 17828 16244
rect 17776 16201 17785 16235
rect 17785 16201 17819 16235
rect 17819 16201 17828 16235
rect 17776 16192 17828 16201
rect 18512 16235 18564 16244
rect 18512 16201 18521 16235
rect 18521 16201 18555 16235
rect 18555 16201 18564 16235
rect 18512 16192 18564 16201
rect 24768 16235 24820 16244
rect 24768 16201 24777 16235
rect 24777 16201 24811 16235
rect 24811 16201 24820 16235
rect 24768 16192 24820 16201
rect 6092 15988 6144 16040
rect 8484 16124 8536 16176
rect 11428 16167 11480 16176
rect 11428 16133 11437 16167
rect 11437 16133 11471 16167
rect 11471 16133 11480 16167
rect 11428 16124 11480 16133
rect 13820 16167 13872 16176
rect 13820 16133 13829 16167
rect 13829 16133 13863 16167
rect 13863 16133 13872 16167
rect 13820 16124 13872 16133
rect 16948 16124 17000 16176
rect 6828 16099 6880 16108
rect 6828 16065 6837 16099
rect 6837 16065 6871 16099
rect 6871 16065 6880 16099
rect 6828 16056 6880 16065
rect 8392 15988 8444 16040
rect 8760 15988 8812 16040
rect 10140 15988 10192 16040
rect 15384 16056 15436 16108
rect 19340 16056 19392 16108
rect 7472 15920 7524 15972
rect 8208 15963 8260 15972
rect 8208 15929 8217 15963
rect 8217 15929 8251 15963
rect 8251 15929 8260 15963
rect 8208 15920 8260 15929
rect 9772 15920 9824 15972
rect 9128 15852 9180 15904
rect 10416 15920 10468 15972
rect 10784 15988 10836 16040
rect 11152 15988 11204 16040
rect 12624 16031 12676 16040
rect 12624 15997 12633 16031
rect 12633 15997 12667 16031
rect 12667 15997 12676 16031
rect 12624 15988 12676 15997
rect 12900 16031 12952 16040
rect 12900 15997 12909 16031
rect 12909 15997 12943 16031
rect 12943 15997 12952 16031
rect 12900 15988 12952 15997
rect 11704 15920 11756 15972
rect 11888 15895 11940 15904
rect 11888 15861 11897 15895
rect 11897 15861 11931 15895
rect 11931 15861 11940 15895
rect 12808 15920 12860 15972
rect 13452 15988 13504 16040
rect 14740 16031 14792 16040
rect 14740 15997 14749 16031
rect 14749 15997 14783 16031
rect 14783 15997 14792 16031
rect 14740 15988 14792 15997
rect 17592 15988 17644 16040
rect 24032 15988 24084 16040
rect 11888 15852 11940 15861
rect 12900 15852 12952 15904
rect 14556 15920 14608 15972
rect 15752 15920 15804 15972
rect 19708 15920 19760 15972
rect 16488 15895 16540 15904
rect 16488 15861 16497 15895
rect 16497 15861 16531 15895
rect 16531 15861 16540 15895
rect 16488 15852 16540 15861
rect 17040 15895 17092 15904
rect 17040 15861 17049 15895
rect 17049 15861 17083 15895
rect 17083 15861 17092 15895
rect 17040 15852 17092 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 7472 15691 7524 15700
rect 7472 15657 7481 15691
rect 7481 15657 7515 15691
rect 7515 15657 7524 15691
rect 7472 15648 7524 15657
rect 7748 15648 7800 15700
rect 8760 15648 8812 15700
rect 11704 15691 11756 15700
rect 11704 15657 11713 15691
rect 11713 15657 11747 15691
rect 11747 15657 11756 15691
rect 11704 15648 11756 15657
rect 12624 15648 12676 15700
rect 16212 15691 16264 15700
rect 16212 15657 16221 15691
rect 16221 15657 16255 15691
rect 16255 15657 16264 15691
rect 16212 15648 16264 15657
rect 17040 15648 17092 15700
rect 7288 15580 7340 15632
rect 6644 15512 6696 15564
rect 7196 15512 7248 15564
rect 8208 15580 8260 15632
rect 10140 15555 10192 15564
rect 10140 15521 10149 15555
rect 10149 15521 10183 15555
rect 10183 15521 10192 15555
rect 10140 15512 10192 15521
rect 10692 15555 10744 15564
rect 10692 15521 10701 15555
rect 10701 15521 10735 15555
rect 10735 15521 10744 15555
rect 10692 15512 10744 15521
rect 10784 15555 10836 15564
rect 10784 15521 10793 15555
rect 10793 15521 10827 15555
rect 10827 15521 10836 15555
rect 11336 15555 11388 15564
rect 10784 15512 10836 15521
rect 11336 15521 11345 15555
rect 11345 15521 11379 15555
rect 11379 15521 11388 15555
rect 11336 15512 11388 15521
rect 12440 15555 12492 15564
rect 12440 15521 12449 15555
rect 12449 15521 12483 15555
rect 12483 15521 12492 15555
rect 12440 15512 12492 15521
rect 15752 15580 15804 15632
rect 17224 15623 17276 15632
rect 17224 15589 17233 15623
rect 17233 15589 17267 15623
rect 17267 15589 17276 15623
rect 17224 15580 17276 15589
rect 12900 15512 12952 15564
rect 13084 15555 13136 15564
rect 13084 15521 13093 15555
rect 13093 15521 13127 15555
rect 13127 15521 13136 15555
rect 13084 15512 13136 15521
rect 13452 15555 13504 15564
rect 13452 15521 13461 15555
rect 13461 15521 13495 15555
rect 13495 15521 13504 15555
rect 13452 15512 13504 15521
rect 18696 15512 18748 15564
rect 8484 15444 8536 15496
rect 16120 15444 16172 15496
rect 17132 15487 17184 15496
rect 17132 15453 17141 15487
rect 17141 15453 17175 15487
rect 17175 15453 17184 15487
rect 17132 15444 17184 15453
rect 17592 15487 17644 15496
rect 17592 15453 17601 15487
rect 17601 15453 17635 15487
rect 17635 15453 17644 15487
rect 17592 15444 17644 15453
rect 9496 15351 9548 15360
rect 9496 15317 9505 15351
rect 9505 15317 9539 15351
rect 9539 15317 9548 15351
rect 9496 15308 9548 15317
rect 13912 15308 13964 15360
rect 14740 15351 14792 15360
rect 14740 15317 14749 15351
rect 14749 15317 14783 15351
rect 14783 15317 14792 15351
rect 14740 15308 14792 15317
rect 18052 15351 18104 15360
rect 18052 15317 18061 15351
rect 18061 15317 18095 15351
rect 18095 15317 18104 15351
rect 18052 15308 18104 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 6644 15147 6696 15156
rect 6644 15113 6653 15147
rect 6653 15113 6687 15147
rect 6687 15113 6696 15147
rect 6644 15104 6696 15113
rect 8024 15104 8076 15156
rect 8208 15104 8260 15156
rect 9128 15147 9180 15156
rect 9128 15113 9137 15147
rect 9137 15113 9171 15147
rect 9171 15113 9180 15147
rect 9128 15104 9180 15113
rect 16120 15147 16172 15156
rect 16120 15113 16129 15147
rect 16129 15113 16163 15147
rect 16163 15113 16172 15147
rect 16120 15104 16172 15113
rect 17132 15104 17184 15156
rect 7656 15079 7708 15088
rect 7656 15045 7665 15079
rect 7665 15045 7699 15079
rect 7699 15045 7708 15079
rect 7656 15036 7708 15045
rect 12440 15036 12492 15088
rect 13912 15011 13964 15020
rect 13912 14977 13921 15011
rect 13921 14977 13955 15011
rect 13955 14977 13964 15011
rect 13912 14968 13964 14977
rect 15292 15011 15344 15020
rect 15292 14977 15301 15011
rect 15301 14977 15335 15011
rect 15335 14977 15344 15011
rect 15292 14968 15344 14977
rect 17224 14968 17276 15020
rect 17960 14968 18012 15020
rect 9404 14900 9456 14952
rect 10140 14943 10192 14952
rect 10140 14909 10149 14943
rect 10149 14909 10183 14943
rect 10183 14909 10192 14943
rect 10140 14900 10192 14909
rect 10692 14943 10744 14952
rect 10692 14909 10701 14943
rect 10701 14909 10735 14943
rect 10735 14909 10744 14943
rect 10692 14900 10744 14909
rect 10784 14943 10836 14952
rect 10784 14909 10793 14943
rect 10793 14909 10827 14943
rect 10827 14909 10836 14943
rect 11152 14943 11204 14952
rect 10784 14900 10836 14909
rect 11152 14909 11161 14943
rect 11161 14909 11195 14943
rect 11195 14909 11204 14943
rect 11152 14900 11204 14909
rect 12440 14943 12492 14952
rect 12440 14909 12449 14943
rect 12449 14909 12483 14943
rect 12483 14909 12492 14943
rect 12440 14900 12492 14909
rect 12900 14943 12952 14952
rect 12900 14909 12909 14943
rect 12909 14909 12943 14943
rect 12943 14909 12952 14943
rect 12900 14900 12952 14909
rect 13636 14943 13688 14952
rect 7104 14875 7156 14884
rect 7104 14841 7113 14875
rect 7113 14841 7147 14875
rect 7147 14841 7156 14875
rect 7104 14832 7156 14841
rect 7196 14875 7248 14884
rect 7196 14841 7205 14875
rect 7205 14841 7239 14875
rect 7239 14841 7248 14875
rect 8484 14875 8536 14884
rect 7196 14832 7248 14841
rect 8484 14841 8493 14875
rect 8493 14841 8527 14875
rect 8527 14841 8536 14875
rect 8484 14832 8536 14841
rect 9404 14807 9456 14816
rect 9404 14773 9413 14807
rect 9413 14773 9447 14807
rect 9447 14773 9456 14807
rect 13084 14832 13136 14884
rect 13636 14909 13645 14943
rect 13645 14909 13679 14943
rect 13679 14909 13688 14943
rect 13636 14900 13688 14909
rect 16856 14943 16908 14952
rect 16856 14909 16865 14943
rect 16865 14909 16899 14943
rect 16899 14909 16908 14943
rect 16856 14900 16908 14909
rect 16948 14900 17000 14952
rect 18052 14943 18104 14952
rect 18052 14909 18096 14943
rect 18096 14909 18104 14943
rect 18052 14900 18104 14909
rect 14832 14875 14884 14884
rect 14832 14841 14841 14875
rect 14841 14841 14875 14875
rect 14875 14841 14884 14875
rect 14832 14832 14884 14841
rect 9404 14764 9456 14773
rect 14280 14764 14332 14816
rect 19708 14832 19760 14884
rect 15752 14807 15804 14816
rect 15752 14773 15761 14807
rect 15761 14773 15795 14807
rect 15795 14773 15804 14807
rect 15752 14764 15804 14773
rect 18696 14807 18748 14816
rect 18696 14773 18705 14807
rect 18705 14773 18739 14807
rect 18739 14773 18748 14807
rect 18696 14764 18748 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 10140 14560 10192 14612
rect 11704 14560 11756 14612
rect 13084 14603 13136 14612
rect 13084 14569 13093 14603
rect 13093 14569 13127 14603
rect 13127 14569 13136 14603
rect 13084 14560 13136 14569
rect 14832 14603 14884 14612
rect 14832 14569 14841 14603
rect 14841 14569 14875 14603
rect 14875 14569 14884 14603
rect 14832 14560 14884 14569
rect 16856 14560 16908 14612
rect 24768 14603 24820 14612
rect 24768 14569 24777 14603
rect 24777 14569 24811 14603
rect 24811 14569 24820 14603
rect 24768 14560 24820 14569
rect 9220 14492 9272 14544
rect 9496 14492 9548 14544
rect 11336 14492 11388 14544
rect 13636 14492 13688 14544
rect 16488 14492 16540 14544
rect 17040 14492 17092 14544
rect 6552 14424 6604 14476
rect 8852 14424 8904 14476
rect 10140 14424 10192 14476
rect 11060 14467 11112 14476
rect 11060 14433 11069 14467
rect 11069 14433 11103 14467
rect 11103 14433 11112 14467
rect 11060 14424 11112 14433
rect 11704 14424 11756 14476
rect 12900 14424 12952 14476
rect 14280 14467 14332 14476
rect 14280 14433 14289 14467
rect 14289 14433 14323 14467
rect 14323 14433 14332 14467
rect 14280 14424 14332 14433
rect 15476 14424 15528 14476
rect 17316 14424 17368 14476
rect 18144 14467 18196 14476
rect 18144 14433 18153 14467
rect 18153 14433 18187 14467
rect 18187 14433 18196 14467
rect 18144 14424 18196 14433
rect 18512 14424 18564 14476
rect 19708 14467 19760 14476
rect 19708 14433 19717 14467
rect 19717 14433 19751 14467
rect 19751 14433 19760 14467
rect 19708 14424 19760 14433
rect 24676 14424 24728 14476
rect 6368 14356 6420 14408
rect 10784 14356 10836 14408
rect 14188 14356 14240 14408
rect 14648 14356 14700 14408
rect 16948 14399 17000 14408
rect 16948 14365 16957 14399
rect 16957 14365 16991 14399
rect 16991 14365 17000 14399
rect 16948 14356 17000 14365
rect 18788 14399 18840 14408
rect 18788 14365 18797 14399
rect 18797 14365 18831 14399
rect 18831 14365 18840 14399
rect 18788 14356 18840 14365
rect 3884 14288 3936 14340
rect 7104 14331 7156 14340
rect 7104 14297 7113 14331
rect 7113 14297 7147 14331
rect 7147 14297 7156 14331
rect 7104 14288 7156 14297
rect 9588 14288 9640 14340
rect 10968 14288 11020 14340
rect 11152 14288 11204 14340
rect 13452 14331 13504 14340
rect 13452 14297 13461 14331
rect 13461 14297 13495 14331
rect 13495 14297 13504 14331
rect 13452 14288 13504 14297
rect 6552 14220 6604 14272
rect 7840 14263 7892 14272
rect 7840 14229 7849 14263
rect 7849 14229 7883 14263
rect 7883 14229 7892 14263
rect 7840 14220 7892 14229
rect 16212 14220 16264 14272
rect 20076 14220 20128 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 14280 14016 14332 14068
rect 15292 14016 15344 14068
rect 15384 14059 15436 14068
rect 15384 14025 15393 14059
rect 15393 14025 15427 14059
rect 15427 14025 15436 14059
rect 15384 14016 15436 14025
rect 18144 14016 18196 14068
rect 24676 14016 24728 14068
rect 27620 14016 27672 14068
rect 9404 13948 9456 14000
rect 10692 13948 10744 14000
rect 11244 13948 11296 14000
rect 7840 13923 7892 13932
rect 7840 13889 7849 13923
rect 7849 13889 7883 13923
rect 7883 13889 7892 13923
rect 7840 13880 7892 13889
rect 8208 13923 8260 13932
rect 8208 13889 8217 13923
rect 8217 13889 8251 13923
rect 8251 13889 8260 13923
rect 8208 13880 8260 13889
rect 9956 13880 10008 13932
rect 1860 13855 1912 13864
rect 1860 13821 1869 13855
rect 1869 13821 1903 13855
rect 1903 13821 1912 13855
rect 1860 13812 1912 13821
rect 9312 13855 9364 13864
rect 9312 13821 9321 13855
rect 9321 13821 9355 13855
rect 9355 13821 9364 13855
rect 9312 13812 9364 13821
rect 9680 13855 9732 13864
rect 9680 13821 9689 13855
rect 9689 13821 9723 13855
rect 9723 13821 9732 13855
rect 9680 13812 9732 13821
rect 11060 13812 11112 13864
rect 12072 13812 12124 13864
rect 13820 13812 13872 13864
rect 15292 13880 15344 13932
rect 16948 13880 17000 13932
rect 20076 13948 20128 14000
rect 22744 13948 22796 14000
rect 15384 13812 15436 13864
rect 18696 13880 18748 13932
rect 19708 13923 19760 13932
rect 19708 13889 19717 13923
rect 19717 13889 19751 13923
rect 19751 13889 19760 13923
rect 19708 13880 19760 13889
rect 20260 13855 20312 13864
rect 20260 13821 20278 13855
rect 20278 13821 20312 13855
rect 4160 13744 4212 13796
rect 6644 13744 6696 13796
rect 6184 13676 6236 13728
rect 8576 13744 8628 13796
rect 9772 13744 9824 13796
rect 10140 13744 10192 13796
rect 11704 13744 11756 13796
rect 13360 13744 13412 13796
rect 13912 13744 13964 13796
rect 15476 13744 15528 13796
rect 16212 13787 16264 13796
rect 16212 13753 16221 13787
rect 16221 13753 16255 13787
rect 16255 13753 16264 13787
rect 16212 13744 16264 13753
rect 17132 13744 17184 13796
rect 20260 13812 20312 13821
rect 8852 13719 8904 13728
rect 8852 13685 8861 13719
rect 8861 13685 8895 13719
rect 8895 13685 8904 13719
rect 8852 13676 8904 13685
rect 9036 13676 9088 13728
rect 9680 13676 9732 13728
rect 11336 13719 11388 13728
rect 11336 13685 11345 13719
rect 11345 13685 11379 13719
rect 11379 13685 11388 13719
rect 11336 13676 11388 13685
rect 12900 13676 12952 13728
rect 13544 13719 13596 13728
rect 13544 13685 13553 13719
rect 13553 13685 13587 13719
rect 13587 13685 13596 13719
rect 13544 13676 13596 13685
rect 14832 13676 14884 13728
rect 17040 13719 17092 13728
rect 17040 13685 17049 13719
rect 17049 13685 17083 13719
rect 17083 13685 17092 13719
rect 17040 13676 17092 13685
rect 17500 13719 17552 13728
rect 17500 13685 17509 13719
rect 17509 13685 17543 13719
rect 17543 13685 17552 13719
rect 17500 13676 17552 13685
rect 21088 13744 21140 13796
rect 21548 13744 21600 13796
rect 23388 13744 23440 13796
rect 25688 13744 25740 13796
rect 18328 13719 18380 13728
rect 18328 13685 18337 13719
rect 18337 13685 18371 13719
rect 18371 13685 18380 13719
rect 18328 13676 18380 13685
rect 18420 13676 18472 13728
rect 22284 13676 22336 13728
rect 22468 13676 22520 13728
rect 23756 13676 23808 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 9680 13472 9732 13524
rect 6552 13447 6604 13456
rect 6552 13413 6561 13447
rect 6561 13413 6595 13447
rect 6595 13413 6604 13447
rect 6552 13404 6604 13413
rect 6644 13447 6696 13456
rect 6644 13413 6653 13447
rect 6653 13413 6687 13447
rect 6687 13413 6696 13447
rect 6644 13404 6696 13413
rect 7656 13404 7708 13456
rect 9312 13404 9364 13456
rect 13820 13515 13872 13524
rect 13820 13481 13829 13515
rect 13829 13481 13863 13515
rect 13863 13481 13872 13515
rect 13820 13472 13872 13481
rect 16488 13472 16540 13524
rect 17592 13472 17644 13524
rect 20812 13472 20864 13524
rect 22652 13472 22704 13524
rect 9956 13404 10008 13456
rect 13544 13404 13596 13456
rect 15752 13404 15804 13456
rect 17040 13447 17092 13456
rect 17040 13413 17049 13447
rect 17049 13413 17083 13447
rect 17083 13413 17092 13447
rect 17040 13404 17092 13413
rect 17224 13404 17276 13456
rect 18512 13404 18564 13456
rect 8760 13336 8812 13388
rect 9496 13336 9548 13388
rect 11704 13336 11756 13388
rect 12072 13379 12124 13388
rect 12072 13345 12081 13379
rect 12081 13345 12115 13379
rect 12115 13345 12124 13379
rect 12072 13336 12124 13345
rect 12532 13379 12584 13388
rect 12532 13345 12541 13379
rect 12541 13345 12575 13379
rect 12575 13345 12584 13379
rect 12532 13336 12584 13345
rect 13268 13336 13320 13388
rect 13636 13336 13688 13388
rect 16212 13379 16264 13388
rect 16212 13345 16221 13379
rect 16221 13345 16255 13379
rect 16255 13345 16264 13379
rect 17408 13379 17460 13388
rect 16212 13336 16264 13345
rect 17408 13345 17417 13379
rect 17417 13345 17451 13379
rect 17451 13345 17460 13379
rect 17408 13336 17460 13345
rect 18880 13379 18932 13388
rect 18880 13345 18889 13379
rect 18889 13345 18923 13379
rect 18923 13345 18932 13379
rect 18880 13336 18932 13345
rect 19064 13379 19116 13388
rect 19064 13345 19073 13379
rect 19073 13345 19107 13379
rect 19107 13345 19116 13379
rect 19064 13336 19116 13345
rect 8116 13311 8168 13320
rect 8116 13277 8125 13311
rect 8125 13277 8159 13311
rect 8159 13277 8168 13311
rect 8116 13268 8168 13277
rect 8208 13268 8260 13320
rect 9956 13268 10008 13320
rect 8668 13243 8720 13252
rect 8668 13209 8677 13243
rect 8677 13209 8711 13243
rect 8711 13209 8720 13243
rect 15384 13268 15436 13320
rect 21272 13336 21324 13388
rect 22836 13336 22888 13388
rect 24216 13336 24268 13388
rect 25228 13336 25280 13388
rect 22192 13268 22244 13320
rect 8668 13200 8720 13209
rect 11060 13200 11112 13252
rect 11612 13200 11664 13252
rect 18696 13200 18748 13252
rect 7932 13175 7984 13184
rect 7932 13141 7941 13175
rect 7941 13141 7975 13175
rect 7975 13141 7984 13175
rect 7932 13132 7984 13141
rect 9036 13175 9088 13184
rect 9036 13141 9045 13175
rect 9045 13141 9079 13175
rect 9079 13141 9088 13175
rect 9036 13132 9088 13141
rect 9496 13175 9548 13184
rect 9496 13141 9505 13175
rect 9505 13141 9539 13175
rect 9539 13141 9548 13175
rect 9496 13132 9548 13141
rect 10968 13132 11020 13184
rect 11704 13132 11756 13184
rect 14280 13132 14332 13184
rect 17500 13132 17552 13184
rect 20168 13132 20220 13184
rect 24032 13132 24084 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 7656 12971 7708 12980
rect 7656 12937 7665 12971
rect 7665 12937 7699 12971
rect 7699 12937 7708 12971
rect 7656 12928 7708 12937
rect 8024 12971 8076 12980
rect 8024 12937 8033 12971
rect 8033 12937 8067 12971
rect 8067 12937 8076 12971
rect 8024 12928 8076 12937
rect 9036 12971 9088 12980
rect 9036 12937 9045 12971
rect 9045 12937 9079 12971
rect 9079 12937 9088 12971
rect 9036 12928 9088 12937
rect 11244 12928 11296 12980
rect 12532 12928 12584 12980
rect 14648 12971 14700 12980
rect 14648 12937 14657 12971
rect 14657 12937 14691 12971
rect 14691 12937 14700 12971
rect 14648 12928 14700 12937
rect 15384 12928 15436 12980
rect 17408 12971 17460 12980
rect 17408 12937 17417 12971
rect 17417 12937 17451 12971
rect 17451 12937 17460 12971
rect 17408 12928 17460 12937
rect 19064 12971 19116 12980
rect 19064 12937 19073 12971
rect 19073 12937 19107 12971
rect 19107 12937 19116 12971
rect 19064 12928 19116 12937
rect 12440 12860 12492 12912
rect 13820 12903 13872 12912
rect 13820 12869 13829 12903
rect 13829 12869 13863 12903
rect 13863 12869 13872 12903
rect 13820 12860 13872 12869
rect 14832 12860 14884 12912
rect 15752 12860 15804 12912
rect 16948 12860 17000 12912
rect 5816 12767 5868 12776
rect 5816 12733 5825 12767
rect 5825 12733 5859 12767
rect 5859 12733 5868 12767
rect 5816 12724 5868 12733
rect 7932 12724 7984 12776
rect 6644 12656 6696 12708
rect 8024 12656 8076 12708
rect 10048 12724 10100 12776
rect 10600 12767 10652 12776
rect 10600 12733 10609 12767
rect 10609 12733 10643 12767
rect 10643 12733 10652 12767
rect 10600 12724 10652 12733
rect 10784 12767 10836 12776
rect 10784 12733 10793 12767
rect 10793 12733 10827 12767
rect 10827 12733 10836 12767
rect 10784 12724 10836 12733
rect 11060 12767 11112 12776
rect 11060 12733 11069 12767
rect 11069 12733 11103 12767
rect 11103 12733 11112 12767
rect 11060 12724 11112 12733
rect 11704 12724 11756 12776
rect 15292 12835 15344 12844
rect 15292 12801 15301 12835
rect 15301 12801 15335 12835
rect 15335 12801 15344 12835
rect 15292 12792 15344 12801
rect 16488 12835 16540 12844
rect 16488 12801 16497 12835
rect 16497 12801 16531 12835
rect 16531 12801 16540 12835
rect 16488 12792 16540 12801
rect 16764 12835 16816 12844
rect 16764 12801 16773 12835
rect 16773 12801 16807 12835
rect 16807 12801 16816 12835
rect 16764 12792 16816 12801
rect 18604 12835 18656 12844
rect 18604 12801 18613 12835
rect 18613 12801 18647 12835
rect 18647 12801 18656 12835
rect 18604 12792 18656 12801
rect 19432 12860 19484 12912
rect 12532 12724 12584 12776
rect 13268 12767 13320 12776
rect 13268 12733 13277 12767
rect 13277 12733 13311 12767
rect 13311 12733 13320 12767
rect 13268 12724 13320 12733
rect 13452 12724 13504 12776
rect 20076 12724 20128 12776
rect 21364 12792 21416 12844
rect 21088 12724 21140 12776
rect 25964 12860 26016 12912
rect 25228 12835 25280 12844
rect 25228 12801 25237 12835
rect 25237 12801 25271 12835
rect 25271 12801 25280 12835
rect 25228 12792 25280 12801
rect 26332 12792 26384 12844
rect 6828 12631 6880 12640
rect 6828 12597 6837 12631
rect 6837 12597 6871 12631
rect 6871 12597 6880 12631
rect 6828 12588 6880 12597
rect 9772 12631 9824 12640
rect 9772 12597 9781 12631
rect 9781 12597 9815 12631
rect 9815 12597 9824 12631
rect 9772 12588 9824 12597
rect 14648 12656 14700 12708
rect 18144 12699 18196 12708
rect 16212 12588 16264 12640
rect 18144 12665 18153 12699
rect 18153 12665 18187 12699
rect 18187 12665 18196 12699
rect 18144 12656 18196 12665
rect 21180 12656 21232 12708
rect 25320 12656 25372 12708
rect 20536 12588 20588 12640
rect 21272 12588 21324 12640
rect 21732 12631 21784 12640
rect 21732 12597 21741 12631
rect 21741 12597 21775 12631
rect 21775 12597 21784 12631
rect 21732 12588 21784 12597
rect 22192 12588 22244 12640
rect 22836 12631 22888 12640
rect 22836 12597 22845 12631
rect 22845 12597 22879 12631
rect 22879 12597 22888 12631
rect 22836 12588 22888 12597
rect 24216 12631 24268 12640
rect 24216 12597 24225 12631
rect 24225 12597 24259 12631
rect 24259 12597 24268 12631
rect 24216 12588 24268 12597
rect 25136 12588 25188 12640
rect 25504 12631 25556 12640
rect 25504 12597 25513 12631
rect 25513 12597 25547 12631
rect 25547 12597 25556 12631
rect 25504 12588 25556 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 6828 12384 6880 12436
rect 7564 12427 7616 12436
rect 7564 12393 7573 12427
rect 7573 12393 7607 12427
rect 7607 12393 7616 12427
rect 7564 12384 7616 12393
rect 8116 12384 8168 12436
rect 5816 12316 5868 12368
rect 6184 12316 6236 12368
rect 8024 12316 8076 12368
rect 7564 12248 7616 12300
rect 7748 12248 7800 12300
rect 14832 12427 14884 12436
rect 14832 12393 14841 12427
rect 14841 12393 14875 12427
rect 14875 12393 14884 12427
rect 14832 12384 14884 12393
rect 18144 12384 18196 12436
rect 19524 12384 19576 12436
rect 21088 12384 21140 12436
rect 22560 12427 22612 12436
rect 22560 12393 22569 12427
rect 22569 12393 22603 12427
rect 22603 12393 22612 12427
rect 22560 12384 22612 12393
rect 9588 12316 9640 12368
rect 8576 12291 8628 12300
rect 8576 12257 8585 12291
rect 8585 12257 8619 12291
rect 8619 12257 8628 12291
rect 8576 12248 8628 12257
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 10048 12248 10100 12257
rect 10600 12291 10652 12300
rect 5540 12180 5592 12232
rect 9772 12180 9824 12232
rect 10600 12257 10609 12291
rect 10609 12257 10643 12291
rect 10643 12257 10652 12291
rect 10600 12248 10652 12257
rect 10784 12248 10836 12300
rect 13728 12316 13780 12368
rect 16120 12316 16172 12368
rect 16488 12359 16540 12368
rect 16488 12325 16497 12359
rect 16497 12325 16531 12359
rect 16531 12325 16540 12359
rect 16488 12316 16540 12325
rect 16580 12316 16632 12368
rect 17960 12359 18012 12368
rect 17960 12325 17969 12359
rect 17969 12325 18003 12359
rect 18003 12325 18012 12359
rect 17960 12316 18012 12325
rect 18052 12359 18104 12368
rect 18052 12325 18061 12359
rect 18061 12325 18095 12359
rect 18095 12325 18104 12359
rect 18052 12316 18104 12325
rect 13084 12248 13136 12300
rect 14648 12248 14700 12300
rect 15752 12291 15804 12300
rect 15752 12257 15761 12291
rect 15761 12257 15795 12291
rect 15795 12257 15804 12291
rect 15752 12248 15804 12257
rect 19248 12248 19300 12300
rect 20904 12291 20956 12300
rect 20904 12257 20913 12291
rect 20913 12257 20947 12291
rect 20947 12257 20956 12291
rect 20904 12248 20956 12257
rect 21364 12291 21416 12300
rect 21364 12257 21373 12291
rect 21373 12257 21407 12291
rect 21407 12257 21416 12291
rect 21364 12248 21416 12257
rect 22192 12248 22244 12300
rect 22928 12291 22980 12300
rect 22928 12257 22937 12291
rect 22937 12257 22971 12291
rect 22971 12257 22980 12291
rect 22928 12248 22980 12257
rect 23020 12248 23072 12300
rect 24676 12316 24728 12368
rect 27620 12316 27672 12368
rect 25872 12248 25924 12300
rect 10692 12180 10744 12232
rect 11980 12180 12032 12232
rect 14004 12180 14056 12232
rect 16764 12180 16816 12232
rect 17040 12223 17092 12232
rect 17040 12189 17049 12223
rect 17049 12189 17083 12223
rect 17083 12189 17092 12223
rect 17040 12180 17092 12189
rect 20076 12180 20128 12232
rect 21640 12223 21692 12232
rect 21640 12189 21649 12223
rect 21649 12189 21683 12223
rect 21683 12189 21692 12223
rect 21640 12180 21692 12189
rect 6460 12112 6512 12164
rect 9220 12112 9272 12164
rect 11060 12112 11112 12164
rect 9772 12044 9824 12096
rect 10784 12044 10836 12096
rect 13268 12112 13320 12164
rect 18604 12112 18656 12164
rect 12348 12087 12400 12096
rect 12348 12053 12357 12087
rect 12357 12053 12391 12087
rect 12391 12053 12400 12087
rect 12348 12044 12400 12053
rect 16212 12087 16264 12096
rect 16212 12053 16221 12087
rect 16221 12053 16255 12087
rect 16255 12053 16264 12087
rect 16212 12044 16264 12053
rect 16580 12044 16632 12096
rect 18880 12087 18932 12096
rect 18880 12053 18889 12087
rect 18889 12053 18923 12087
rect 18923 12053 18932 12087
rect 18880 12044 18932 12053
rect 19340 12087 19392 12096
rect 19340 12053 19349 12087
rect 19349 12053 19383 12087
rect 19383 12053 19392 12087
rect 19340 12044 19392 12053
rect 20628 12087 20680 12096
rect 20628 12053 20637 12087
rect 20637 12053 20671 12087
rect 20671 12053 20680 12087
rect 20628 12044 20680 12053
rect 23572 12044 23624 12096
rect 24768 12044 24820 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 6460 11840 6512 11892
rect 6644 11883 6696 11892
rect 6644 11849 6653 11883
rect 6653 11849 6687 11883
rect 6687 11849 6696 11883
rect 6644 11840 6696 11849
rect 8024 11840 8076 11892
rect 10048 11840 10100 11892
rect 12348 11840 12400 11892
rect 14372 11840 14424 11892
rect 16488 11883 16540 11892
rect 16488 11849 16497 11883
rect 16497 11849 16531 11883
rect 16531 11849 16540 11883
rect 16488 11840 16540 11849
rect 17960 11840 18012 11892
rect 19156 11840 19208 11892
rect 20904 11883 20956 11892
rect 20904 11849 20913 11883
rect 20913 11849 20947 11883
rect 20947 11849 20956 11883
rect 20904 11840 20956 11849
rect 21364 11840 21416 11892
rect 22928 11840 22980 11892
rect 24124 11840 24176 11892
rect 24676 11840 24728 11892
rect 6828 11772 6880 11824
rect 9404 11772 9456 11824
rect 9496 11772 9548 11824
rect 7564 11747 7616 11756
rect 7564 11713 7573 11747
rect 7573 11713 7607 11747
rect 7607 11713 7616 11747
rect 7564 11704 7616 11713
rect 8852 11704 8904 11756
rect 10600 11704 10652 11756
rect 6736 11636 6788 11688
rect 9220 11679 9272 11688
rect 9220 11645 9229 11679
rect 9229 11645 9263 11679
rect 9263 11645 9272 11679
rect 9220 11636 9272 11645
rect 10784 11679 10836 11688
rect 6644 11568 6696 11620
rect 7196 11568 7248 11620
rect 9956 11611 10008 11620
rect 9956 11577 9965 11611
rect 9965 11577 9999 11611
rect 9999 11577 10008 11611
rect 9956 11568 10008 11577
rect 4344 11500 4396 11552
rect 5540 11543 5592 11552
rect 5540 11509 5549 11543
rect 5549 11509 5583 11543
rect 5583 11509 5592 11543
rect 5540 11500 5592 11509
rect 9864 11500 9916 11552
rect 10784 11645 10793 11679
rect 10793 11645 10827 11679
rect 10827 11645 10836 11679
rect 10784 11636 10836 11645
rect 11336 11704 11388 11756
rect 17040 11772 17092 11824
rect 19248 11772 19300 11824
rect 20076 11772 20128 11824
rect 13176 11747 13228 11756
rect 13176 11713 13185 11747
rect 13185 11713 13219 11747
rect 13219 11713 13228 11747
rect 13176 11704 13228 11713
rect 14188 11704 14240 11756
rect 19340 11704 19392 11756
rect 10692 11543 10744 11552
rect 10692 11509 10701 11543
rect 10701 11509 10735 11543
rect 10735 11509 10744 11543
rect 11612 11636 11664 11688
rect 14096 11679 14148 11688
rect 14096 11645 14105 11679
rect 14105 11645 14139 11679
rect 14139 11645 14148 11679
rect 14096 11636 14148 11645
rect 16120 11636 16172 11688
rect 17960 11636 18012 11688
rect 22192 11636 22244 11688
rect 23296 11636 23348 11688
rect 24124 11636 24176 11688
rect 10692 11500 10744 11509
rect 12072 11500 12124 11552
rect 12348 11500 12400 11552
rect 15752 11568 15804 11620
rect 13820 11543 13872 11552
rect 13820 11509 13829 11543
rect 13829 11509 13863 11543
rect 13863 11509 13872 11543
rect 13820 11500 13872 11509
rect 14648 11500 14700 11552
rect 17960 11500 18012 11552
rect 19524 11568 19576 11620
rect 19432 11543 19484 11552
rect 19432 11509 19441 11543
rect 19441 11509 19475 11543
rect 19475 11509 19484 11543
rect 20628 11568 20680 11620
rect 21364 11611 21416 11620
rect 21364 11577 21373 11611
rect 21373 11577 21407 11611
rect 21407 11577 21416 11611
rect 21364 11568 21416 11577
rect 26148 11568 26200 11620
rect 19432 11500 19484 11509
rect 24952 11500 25004 11552
rect 25872 11543 25924 11552
rect 25872 11509 25881 11543
rect 25881 11509 25915 11543
rect 25915 11509 25924 11543
rect 25872 11500 25924 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 6184 11339 6236 11348
rect 6184 11305 6193 11339
rect 6193 11305 6227 11339
rect 6227 11305 6236 11339
rect 6184 11296 6236 11305
rect 7748 11339 7800 11348
rect 7748 11305 7757 11339
rect 7757 11305 7791 11339
rect 7791 11305 7800 11339
rect 7748 11296 7800 11305
rect 12532 11339 12584 11348
rect 12532 11305 12541 11339
rect 12541 11305 12575 11339
rect 12575 11305 12584 11339
rect 12532 11296 12584 11305
rect 13084 11339 13136 11348
rect 13084 11305 13093 11339
rect 13093 11305 13127 11339
rect 13127 11305 13136 11339
rect 13084 11296 13136 11305
rect 13820 11296 13872 11348
rect 14004 11339 14056 11348
rect 14004 11305 14013 11339
rect 14013 11305 14047 11339
rect 14047 11305 14056 11339
rect 14004 11296 14056 11305
rect 16120 11296 16172 11348
rect 16764 11296 16816 11348
rect 17960 11339 18012 11348
rect 17960 11305 17969 11339
rect 17969 11305 18003 11339
rect 18003 11305 18012 11339
rect 17960 11296 18012 11305
rect 18788 11296 18840 11348
rect 21180 11296 21232 11348
rect 22008 11296 22060 11348
rect 8392 11228 8444 11280
rect 9772 11228 9824 11280
rect 1584 11160 1636 11212
rect 7104 11160 7156 11212
rect 10048 11203 10100 11212
rect 10048 11169 10057 11203
rect 10057 11169 10091 11203
rect 10091 11169 10100 11203
rect 10048 11160 10100 11169
rect 10416 11160 10468 11212
rect 11888 11228 11940 11280
rect 13728 11271 13780 11280
rect 13728 11237 13737 11271
rect 13737 11237 13771 11271
rect 13771 11237 13780 11271
rect 13728 11228 13780 11237
rect 15752 11228 15804 11280
rect 17684 11228 17736 11280
rect 18972 11271 19024 11280
rect 18972 11237 18981 11271
rect 18981 11237 19015 11271
rect 19015 11237 19024 11271
rect 18972 11228 19024 11237
rect 19248 11228 19300 11280
rect 22744 11271 22796 11280
rect 22744 11237 22753 11271
rect 22753 11237 22787 11271
rect 22787 11237 22796 11271
rect 22744 11228 22796 11237
rect 23296 11271 23348 11280
rect 23296 11237 23305 11271
rect 23305 11237 23339 11271
rect 23339 11237 23348 11271
rect 23296 11228 23348 11237
rect 7288 11092 7340 11144
rect 8208 11135 8260 11144
rect 8208 11101 8217 11135
rect 8217 11101 8251 11135
rect 8251 11101 8260 11135
rect 8208 11092 8260 11101
rect 9220 11092 9272 11144
rect 14556 11160 14608 11212
rect 17592 11160 17644 11212
rect 21088 11203 21140 11212
rect 21088 11169 21097 11203
rect 21097 11169 21131 11203
rect 21131 11169 21140 11203
rect 21088 11160 21140 11169
rect 21272 11160 21324 11212
rect 24216 11203 24268 11212
rect 11796 11092 11848 11144
rect 15292 11135 15344 11144
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 18880 11135 18932 11144
rect 18880 11101 18889 11135
rect 18889 11101 18923 11135
rect 18923 11101 18932 11135
rect 18880 11092 18932 11101
rect 20076 11092 20128 11144
rect 6736 11024 6788 11076
rect 11152 11024 11204 11076
rect 11428 11024 11480 11076
rect 18052 11024 18104 11076
rect 21364 11024 21416 11076
rect 21824 11092 21876 11144
rect 22928 11092 22980 11144
rect 24216 11169 24225 11203
rect 24225 11169 24259 11203
rect 24259 11169 24268 11203
rect 24216 11160 24268 11169
rect 6000 10956 6052 11008
rect 7380 10999 7432 11008
rect 7380 10965 7389 10999
rect 7389 10965 7423 10999
rect 7423 10965 7432 10999
rect 7380 10956 7432 10965
rect 8852 10999 8904 11008
rect 8852 10965 8861 10999
rect 8861 10965 8895 10999
rect 8895 10965 8904 10999
rect 8852 10956 8904 10965
rect 9128 10956 9180 11008
rect 9772 10956 9824 11008
rect 14740 10956 14792 11008
rect 14832 10956 14884 11008
rect 18696 10956 18748 11008
rect 19524 10956 19576 11008
rect 20536 10956 20588 11008
rect 24676 11092 24728 11144
rect 23848 10956 23900 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1584 10795 1636 10804
rect 1584 10761 1593 10795
rect 1593 10761 1627 10795
rect 1627 10761 1636 10795
rect 1584 10752 1636 10761
rect 6092 10752 6144 10804
rect 9128 10752 9180 10804
rect 9680 10752 9732 10804
rect 10140 10752 10192 10804
rect 11428 10795 11480 10804
rect 11428 10761 11437 10795
rect 11437 10761 11471 10795
rect 11471 10761 11480 10795
rect 11428 10752 11480 10761
rect 11796 10795 11848 10804
rect 11796 10761 11805 10795
rect 11805 10761 11839 10795
rect 11839 10761 11848 10795
rect 11796 10752 11848 10761
rect 12532 10752 12584 10804
rect 15752 10752 15804 10804
rect 18696 10752 18748 10804
rect 18972 10795 19024 10804
rect 18972 10761 18981 10795
rect 18981 10761 19015 10795
rect 19015 10761 19024 10795
rect 18972 10752 19024 10761
rect 20628 10752 20680 10804
rect 21272 10752 21324 10804
rect 22744 10752 22796 10804
rect 24676 10795 24728 10804
rect 24676 10761 24685 10795
rect 24685 10761 24719 10795
rect 24719 10761 24728 10795
rect 24676 10752 24728 10761
rect 9312 10684 9364 10736
rect 9956 10684 10008 10736
rect 7196 10616 7248 10668
rect 8208 10616 8260 10668
rect 12808 10616 12860 10668
rect 13176 10659 13228 10668
rect 13176 10625 13185 10659
rect 13185 10625 13219 10659
rect 13219 10625 13228 10659
rect 13176 10616 13228 10625
rect 7380 10548 7432 10600
rect 8024 10480 8076 10532
rect 7104 10455 7156 10464
rect 7104 10421 7113 10455
rect 7113 10421 7147 10455
rect 7147 10421 7156 10455
rect 7104 10412 7156 10421
rect 8484 10455 8536 10464
rect 8484 10421 8493 10455
rect 8493 10421 8527 10455
rect 8527 10421 8536 10455
rect 8484 10412 8536 10421
rect 9772 10591 9824 10600
rect 9312 10480 9364 10532
rect 9772 10557 9781 10591
rect 9781 10557 9815 10591
rect 9815 10557 9824 10591
rect 9772 10548 9824 10557
rect 9956 10548 10008 10600
rect 10416 10548 10468 10600
rect 15292 10684 15344 10736
rect 17684 10727 17736 10736
rect 17684 10693 17693 10727
rect 17693 10693 17727 10727
rect 17727 10693 17736 10727
rect 17684 10684 17736 10693
rect 20076 10684 20128 10736
rect 16764 10616 16816 10668
rect 18788 10616 18840 10668
rect 10048 10480 10100 10532
rect 10140 10480 10192 10532
rect 16672 10548 16724 10600
rect 23020 10684 23072 10736
rect 21180 10659 21232 10668
rect 21180 10625 21189 10659
rect 21189 10625 21223 10659
rect 21223 10625 21232 10659
rect 21180 10616 21232 10625
rect 23848 10616 23900 10668
rect 24032 10659 24084 10668
rect 24032 10625 24041 10659
rect 24041 10625 24075 10659
rect 24075 10625 24084 10659
rect 24032 10616 24084 10625
rect 20628 10548 20680 10600
rect 22928 10591 22980 10600
rect 22928 10557 22937 10591
rect 22937 10557 22971 10591
rect 22971 10557 22980 10591
rect 22928 10548 22980 10557
rect 24860 10548 24912 10600
rect 12624 10523 12676 10532
rect 12624 10489 12633 10523
rect 12633 10489 12667 10523
rect 12667 10489 12676 10523
rect 12624 10480 12676 10489
rect 12992 10480 13044 10532
rect 13176 10480 13228 10532
rect 14832 10480 14884 10532
rect 17684 10480 17736 10532
rect 21456 10480 21508 10532
rect 23112 10480 23164 10532
rect 9772 10412 9824 10464
rect 14188 10455 14240 10464
rect 14188 10421 14197 10455
rect 14197 10421 14231 10455
rect 14231 10421 14240 10455
rect 14188 10412 14240 10421
rect 14556 10455 14608 10464
rect 14556 10421 14565 10455
rect 14565 10421 14599 10455
rect 14599 10421 14608 10455
rect 14556 10412 14608 10421
rect 16396 10455 16448 10464
rect 16396 10421 16405 10455
rect 16405 10421 16439 10455
rect 16439 10421 16448 10455
rect 16396 10412 16448 10421
rect 23940 10480 23992 10532
rect 24676 10480 24728 10532
rect 25596 10412 25648 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 7288 10251 7340 10260
rect 7288 10217 7297 10251
rect 7297 10217 7331 10251
rect 7331 10217 7340 10251
rect 7288 10208 7340 10217
rect 9312 10208 9364 10260
rect 9956 10251 10008 10260
rect 9956 10217 9965 10251
rect 9965 10217 9999 10251
rect 9999 10217 10008 10251
rect 9956 10208 10008 10217
rect 10048 10208 10100 10260
rect 12624 10208 12676 10260
rect 12808 10251 12860 10260
rect 12808 10217 12817 10251
rect 12817 10217 12851 10251
rect 12851 10217 12860 10251
rect 12808 10208 12860 10217
rect 15568 10251 15620 10260
rect 15568 10217 15577 10251
rect 15577 10217 15611 10251
rect 15611 10217 15620 10251
rect 15568 10208 15620 10217
rect 17592 10208 17644 10260
rect 7564 10183 7616 10192
rect 7564 10149 7573 10183
rect 7573 10149 7607 10183
rect 7607 10149 7616 10183
rect 7564 10140 7616 10149
rect 8208 10140 8260 10192
rect 14188 10140 14240 10192
rect 14832 10140 14884 10192
rect 112 10072 164 10124
rect 4804 10115 4856 10124
rect 4804 10081 4848 10115
rect 4848 10081 4856 10115
rect 4804 10072 4856 10081
rect 5540 10072 5592 10124
rect 6552 10072 6604 10124
rect 10140 10115 10192 10124
rect 10140 10081 10149 10115
rect 10149 10081 10183 10115
rect 10183 10081 10192 10115
rect 10140 10072 10192 10081
rect 10692 10072 10744 10124
rect 11796 10115 11848 10124
rect 11796 10081 11805 10115
rect 11805 10081 11839 10115
rect 11839 10081 11848 10115
rect 11796 10072 11848 10081
rect 13912 10115 13964 10124
rect 13912 10081 13921 10115
rect 13921 10081 13955 10115
rect 13955 10081 13964 10115
rect 13912 10072 13964 10081
rect 14280 10072 14332 10124
rect 15476 10115 15528 10124
rect 15476 10081 15485 10115
rect 15485 10081 15519 10115
rect 15519 10081 15528 10115
rect 15476 10072 15528 10081
rect 17224 10140 17276 10192
rect 18144 10140 18196 10192
rect 19432 10208 19484 10260
rect 21088 10251 21140 10260
rect 21088 10217 21097 10251
rect 21097 10217 21131 10251
rect 21131 10217 21140 10251
rect 21088 10208 21140 10217
rect 23296 10208 23348 10260
rect 18880 10140 18932 10192
rect 21456 10140 21508 10192
rect 24216 10208 24268 10260
rect 24124 10140 24176 10192
rect 24952 10140 25004 10192
rect 25228 10140 25280 10192
rect 16856 10115 16908 10124
rect 16856 10081 16865 10115
rect 16865 10081 16899 10115
rect 16899 10081 16908 10115
rect 16856 10072 16908 10081
rect 19064 10072 19116 10124
rect 19708 10072 19760 10124
rect 20720 10072 20772 10124
rect 22560 10072 22612 10124
rect 24216 10072 24268 10124
rect 6460 10047 6512 10056
rect 6460 10013 6469 10047
rect 6469 10013 6503 10047
rect 6503 10013 6512 10047
rect 6460 10004 6512 10013
rect 7472 10047 7524 10056
rect 7472 10013 7481 10047
rect 7481 10013 7515 10047
rect 7515 10013 7524 10047
rect 7472 10004 7524 10013
rect 7012 9936 7064 9988
rect 11612 10004 11664 10056
rect 14372 10047 14424 10056
rect 14372 10013 14381 10047
rect 14381 10013 14415 10047
rect 14415 10013 14424 10047
rect 14372 10004 14424 10013
rect 17500 10004 17552 10056
rect 24032 10004 24084 10056
rect 24952 10047 25004 10056
rect 24952 10013 24961 10047
rect 24961 10013 24995 10047
rect 24995 10013 25004 10047
rect 24952 10004 25004 10013
rect 9404 9936 9456 9988
rect 14464 9936 14516 9988
rect 20536 9936 20588 9988
rect 22928 9936 22980 9988
rect 4068 9868 4120 9920
rect 7196 9868 7248 9920
rect 8484 9868 8536 9920
rect 13544 9911 13596 9920
rect 13544 9877 13553 9911
rect 13553 9877 13587 9911
rect 13587 9877 13596 9911
rect 13544 9868 13596 9877
rect 15384 9868 15436 9920
rect 17224 9868 17276 9920
rect 19156 9868 19208 9920
rect 23204 9911 23256 9920
rect 23204 9877 23213 9911
rect 23213 9877 23247 9911
rect 23247 9877 23256 9911
rect 23204 9868 23256 9877
rect 23388 9868 23440 9920
rect 23664 9868 23716 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 4804 9707 4856 9716
rect 4804 9673 4813 9707
rect 4813 9673 4847 9707
rect 4847 9673 4856 9707
rect 4804 9664 4856 9673
rect 6552 9707 6604 9716
rect 6552 9673 6561 9707
rect 6561 9673 6595 9707
rect 6595 9673 6604 9707
rect 6552 9664 6604 9673
rect 12716 9664 12768 9716
rect 13360 9664 13412 9716
rect 13636 9664 13688 9716
rect 15752 9664 15804 9716
rect 17684 9664 17736 9716
rect 19708 9707 19760 9716
rect 7564 9528 7616 9580
rect 7012 9460 7064 9512
rect 7196 9503 7248 9512
rect 7196 9469 7205 9503
rect 7205 9469 7239 9503
rect 7239 9469 7248 9503
rect 7196 9460 7248 9469
rect 5540 9392 5592 9444
rect 11244 9596 11296 9648
rect 13728 9596 13780 9648
rect 16948 9596 17000 9648
rect 19708 9673 19717 9707
rect 19717 9673 19751 9707
rect 19751 9673 19760 9707
rect 19708 9664 19760 9673
rect 21456 9664 21508 9716
rect 23848 9664 23900 9716
rect 8760 9528 8812 9580
rect 6000 9324 6052 9376
rect 7840 9324 7892 9376
rect 9312 9460 9364 9512
rect 11060 9503 11112 9512
rect 11060 9469 11069 9503
rect 11069 9469 11103 9503
rect 11103 9469 11112 9503
rect 11060 9460 11112 9469
rect 11244 9503 11296 9512
rect 11244 9469 11253 9503
rect 11253 9469 11287 9503
rect 11287 9469 11296 9503
rect 11244 9460 11296 9469
rect 13544 9528 13596 9580
rect 12900 9503 12952 9512
rect 12900 9469 12909 9503
rect 12909 9469 12943 9503
rect 12943 9469 12952 9503
rect 12900 9460 12952 9469
rect 18328 9528 18380 9580
rect 10140 9392 10192 9444
rect 11520 9435 11572 9444
rect 8760 9367 8812 9376
rect 8760 9333 8769 9367
rect 8769 9333 8803 9367
rect 8803 9333 8812 9367
rect 8760 9324 8812 9333
rect 11520 9401 11529 9435
rect 11529 9401 11563 9435
rect 11563 9401 11572 9435
rect 11520 9392 11572 9401
rect 11796 9324 11848 9376
rect 12348 9324 12400 9376
rect 13084 9324 13136 9376
rect 14096 9460 14148 9512
rect 15384 9503 15436 9512
rect 15384 9469 15393 9503
rect 15393 9469 15427 9503
rect 15427 9469 15436 9503
rect 15384 9460 15436 9469
rect 16212 9460 16264 9512
rect 18052 9460 18104 9512
rect 14188 9435 14240 9444
rect 14188 9401 14197 9435
rect 14197 9401 14231 9435
rect 14231 9401 14240 9435
rect 14188 9392 14240 9401
rect 13912 9324 13964 9376
rect 15752 9392 15804 9444
rect 15844 9392 15896 9444
rect 16120 9392 16172 9444
rect 16856 9435 16908 9444
rect 16856 9401 16865 9435
rect 16865 9401 16899 9435
rect 16899 9401 16908 9435
rect 16856 9392 16908 9401
rect 20536 9596 20588 9648
rect 23112 9596 23164 9648
rect 25228 9596 25280 9648
rect 19984 9528 20036 9580
rect 20628 9571 20680 9580
rect 20628 9537 20637 9571
rect 20637 9537 20671 9571
rect 20671 9537 20680 9571
rect 20628 9528 20680 9537
rect 21732 9528 21784 9580
rect 23204 9528 23256 9580
rect 23940 9528 23992 9580
rect 24124 9571 24176 9580
rect 24124 9537 24133 9571
rect 24133 9537 24167 9571
rect 24167 9537 24176 9571
rect 24124 9528 24176 9537
rect 24676 9460 24728 9512
rect 18972 9392 19024 9444
rect 20536 9392 20588 9444
rect 21456 9392 21508 9444
rect 22192 9392 22244 9444
rect 15476 9324 15528 9376
rect 16304 9324 16356 9376
rect 17500 9367 17552 9376
rect 17500 9333 17509 9367
rect 17509 9333 17543 9367
rect 17543 9333 17552 9367
rect 17500 9324 17552 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 4068 9120 4120 9172
rect 5264 9120 5316 9172
rect 7196 9163 7248 9172
rect 7196 9129 7205 9163
rect 7205 9129 7239 9163
rect 7239 9129 7248 9163
rect 7196 9120 7248 9129
rect 9956 9120 10008 9172
rect 14280 9120 14332 9172
rect 14832 9120 14884 9172
rect 15752 9120 15804 9172
rect 15844 9120 15896 9172
rect 16396 9120 16448 9172
rect 18144 9163 18196 9172
rect 18144 9129 18153 9163
rect 18153 9129 18187 9163
rect 18187 9129 18196 9163
rect 18144 9120 18196 9129
rect 19984 9120 20036 9172
rect 20720 9163 20772 9172
rect 20720 9129 20729 9163
rect 20729 9129 20763 9163
rect 20763 9129 20772 9163
rect 20720 9120 20772 9129
rect 21732 9163 21784 9172
rect 21732 9129 21741 9163
rect 21741 9129 21775 9163
rect 21775 9129 21784 9163
rect 21732 9120 21784 9129
rect 22192 9120 22244 9172
rect 23480 9120 23532 9172
rect 4712 9052 4764 9104
rect 6184 9095 6236 9104
rect 6184 9061 6193 9095
rect 6193 9061 6227 9095
rect 6227 9061 6236 9095
rect 6184 9052 6236 9061
rect 6276 9095 6328 9104
rect 6276 9061 6285 9095
rect 6285 9061 6319 9095
rect 6319 9061 6328 9095
rect 6276 9052 6328 9061
rect 8208 9095 8260 9104
rect 8208 9061 8217 9095
rect 8217 9061 8251 9095
rect 8251 9061 8260 9095
rect 8208 9052 8260 9061
rect 12532 9052 12584 9104
rect 9404 8984 9456 9036
rect 11060 9027 11112 9036
rect 11060 8993 11069 9027
rect 11069 8993 11103 9027
rect 11103 8993 11112 9027
rect 11060 8984 11112 8993
rect 11428 8984 11480 9036
rect 15568 9027 15620 9036
rect 15568 8993 15577 9027
rect 15577 8993 15611 9027
rect 15611 8993 15620 9027
rect 15568 8984 15620 8993
rect 18972 9052 19024 9104
rect 23296 9095 23348 9104
rect 23296 9061 23305 9095
rect 23305 9061 23339 9095
rect 23339 9061 23348 9095
rect 23296 9052 23348 9061
rect 23756 9095 23808 9104
rect 23756 9061 23765 9095
rect 23765 9061 23799 9095
rect 23799 9061 23808 9095
rect 23756 9052 23808 9061
rect 24676 9120 24728 9172
rect 25228 9120 25280 9172
rect 17316 8984 17368 9036
rect 17684 8984 17736 9036
rect 20444 8984 20496 9036
rect 20904 9027 20956 9036
rect 20904 8993 20948 9027
rect 20948 8993 20956 9027
rect 20904 8984 20956 8993
rect 21640 8984 21692 9036
rect 25504 8984 25556 9036
rect 6460 8959 6512 8968
rect 6460 8925 6469 8959
rect 6469 8925 6503 8959
rect 6503 8925 6512 8959
rect 6460 8916 6512 8925
rect 9036 8916 9088 8968
rect 12716 8916 12768 8968
rect 14372 8916 14424 8968
rect 18696 8916 18748 8968
rect 24032 8959 24084 8968
rect 24032 8925 24041 8959
rect 24041 8925 24075 8959
rect 24075 8925 24084 8959
rect 24032 8916 24084 8925
rect 7472 8891 7524 8900
rect 3700 8780 3752 8832
rect 7472 8857 7481 8891
rect 7481 8857 7515 8891
rect 7515 8857 7524 8891
rect 7472 8848 7524 8857
rect 8668 8891 8720 8900
rect 8668 8857 8677 8891
rect 8677 8857 8711 8891
rect 8711 8857 8720 8891
rect 8668 8848 8720 8857
rect 8944 8848 8996 8900
rect 19800 8848 19852 8900
rect 21180 8891 21232 8900
rect 21180 8857 21189 8891
rect 21189 8857 21223 8891
rect 21223 8857 21232 8891
rect 21180 8848 21232 8857
rect 24952 8848 25004 8900
rect 25320 8848 25372 8900
rect 9312 8780 9364 8832
rect 9956 8780 10008 8832
rect 11060 8780 11112 8832
rect 12164 8780 12216 8832
rect 12532 8823 12584 8832
rect 12532 8789 12541 8823
rect 12541 8789 12575 8823
rect 12575 8789 12584 8823
rect 12532 8780 12584 8789
rect 14004 8780 14056 8832
rect 14280 8823 14332 8832
rect 14280 8789 14289 8823
rect 14289 8789 14323 8823
rect 14323 8789 14332 8823
rect 14280 8780 14332 8789
rect 17960 8780 18012 8832
rect 19432 8823 19484 8832
rect 19432 8789 19441 8823
rect 19441 8789 19475 8823
rect 19475 8789 19484 8823
rect 19432 8780 19484 8789
rect 21456 8823 21508 8832
rect 21456 8789 21465 8823
rect 21465 8789 21499 8823
rect 21499 8789 21508 8823
rect 21456 8780 21508 8789
rect 25412 8823 25464 8832
rect 25412 8789 25421 8823
rect 25421 8789 25455 8823
rect 25455 8789 25464 8823
rect 25412 8780 25464 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 6184 8576 6236 8628
rect 8024 8619 8076 8628
rect 8024 8585 8033 8619
rect 8033 8585 8067 8619
rect 8067 8585 8076 8619
rect 8024 8576 8076 8585
rect 8208 8576 8260 8628
rect 11060 8619 11112 8628
rect 11060 8585 11069 8619
rect 11069 8585 11103 8619
rect 11103 8585 11112 8619
rect 11060 8576 11112 8585
rect 11520 8576 11572 8628
rect 14004 8619 14056 8628
rect 112 8372 164 8424
rect 8944 8508 8996 8560
rect 9772 8551 9824 8560
rect 9772 8517 9781 8551
rect 9781 8517 9815 8551
rect 9815 8517 9824 8551
rect 9772 8508 9824 8517
rect 5264 8483 5316 8492
rect 5264 8449 5273 8483
rect 5273 8449 5307 8483
rect 5307 8449 5316 8483
rect 5264 8440 5316 8449
rect 6460 8440 6512 8492
rect 7748 8440 7800 8492
rect 7196 8372 7248 8424
rect 9956 8415 10008 8424
rect 9956 8381 9965 8415
rect 9965 8381 9999 8415
rect 9999 8381 10008 8415
rect 9956 8372 10008 8381
rect 14004 8585 14013 8619
rect 14013 8585 14047 8619
rect 14047 8585 14056 8619
rect 14004 8576 14056 8585
rect 15568 8576 15620 8628
rect 15844 8576 15896 8628
rect 20904 8619 20956 8628
rect 20904 8585 20913 8619
rect 20913 8585 20947 8619
rect 20947 8585 20956 8619
rect 20904 8576 20956 8585
rect 21640 8576 21692 8628
rect 23480 8619 23532 8628
rect 23480 8585 23489 8619
rect 23489 8585 23523 8619
rect 23523 8585 23532 8619
rect 23480 8576 23532 8585
rect 23756 8576 23808 8628
rect 23940 8576 23992 8628
rect 25504 8576 25556 8628
rect 12900 8508 12952 8560
rect 14280 8483 14332 8492
rect 14280 8449 14289 8483
rect 14289 8449 14323 8483
rect 14323 8449 14332 8483
rect 14280 8440 14332 8449
rect 24032 8508 24084 8560
rect 24952 8551 25004 8560
rect 24952 8517 24961 8551
rect 24961 8517 24995 8551
rect 24995 8517 25004 8551
rect 24952 8508 25004 8517
rect 17960 8440 18012 8492
rect 18880 8483 18932 8492
rect 18880 8449 18889 8483
rect 18889 8449 18923 8483
rect 18923 8449 18932 8483
rect 18880 8440 18932 8449
rect 19800 8483 19852 8492
rect 19800 8449 19809 8483
rect 19809 8449 19843 8483
rect 19843 8449 19852 8483
rect 19800 8440 19852 8449
rect 20628 8440 20680 8492
rect 21180 8440 21232 8492
rect 25412 8440 25464 8492
rect 13728 8372 13780 8424
rect 16672 8415 16724 8424
rect 16672 8381 16681 8415
rect 16681 8381 16715 8415
rect 16715 8381 16724 8415
rect 16672 8372 16724 8381
rect 5356 8347 5408 8356
rect 5356 8313 5365 8347
rect 5365 8313 5399 8347
rect 5399 8313 5408 8347
rect 5356 8304 5408 8313
rect 6276 8347 6328 8356
rect 6276 8313 6285 8347
rect 6285 8313 6319 8347
rect 6319 8313 6328 8347
rect 6276 8304 6328 8313
rect 5448 8236 5500 8288
rect 7288 8279 7340 8288
rect 7288 8245 7297 8279
rect 7297 8245 7331 8279
rect 7331 8245 7340 8279
rect 7288 8236 7340 8245
rect 8024 8304 8076 8356
rect 9404 8279 9456 8288
rect 9404 8245 9413 8279
rect 9413 8245 9447 8279
rect 9447 8245 9456 8279
rect 9404 8236 9456 8245
rect 9496 8236 9548 8288
rect 9772 8236 9824 8288
rect 10784 8236 10836 8288
rect 11428 8279 11480 8288
rect 11428 8245 11437 8279
rect 11437 8245 11471 8279
rect 11471 8245 11480 8279
rect 11428 8236 11480 8245
rect 12164 8279 12216 8288
rect 12164 8245 12173 8279
rect 12173 8245 12207 8279
rect 12207 8245 12216 8279
rect 12164 8236 12216 8245
rect 12532 8304 12584 8356
rect 14004 8304 14056 8356
rect 16488 8304 16540 8356
rect 17868 8372 17920 8424
rect 22192 8372 22244 8424
rect 17960 8304 18012 8356
rect 18052 8304 18104 8356
rect 19432 8304 19484 8356
rect 21456 8347 21508 8356
rect 13360 8279 13412 8288
rect 13360 8245 13369 8279
rect 13369 8245 13403 8279
rect 13403 8245 13412 8279
rect 13360 8236 13412 8245
rect 17684 8236 17736 8288
rect 18972 8236 19024 8288
rect 21456 8313 21465 8347
rect 21465 8313 21499 8347
rect 21499 8313 21508 8347
rect 21456 8304 21508 8313
rect 23664 8304 23716 8356
rect 24676 8304 24728 8356
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 5356 8032 5408 8084
rect 7012 8032 7064 8084
rect 7748 8075 7800 8084
rect 6184 7964 6236 8016
rect 7748 8041 7757 8075
rect 7757 8041 7791 8075
rect 7791 8041 7800 8075
rect 7748 8032 7800 8041
rect 9036 8075 9088 8084
rect 8024 7964 8076 8016
rect 9036 8041 9045 8075
rect 9045 8041 9079 8075
rect 9079 8041 9088 8075
rect 9036 8032 9088 8041
rect 12440 8075 12492 8084
rect 12440 8041 12449 8075
rect 12449 8041 12483 8075
rect 12483 8041 12492 8075
rect 12440 8032 12492 8041
rect 12716 8075 12768 8084
rect 12716 8041 12725 8075
rect 12725 8041 12759 8075
rect 12759 8041 12768 8075
rect 12716 8032 12768 8041
rect 15384 8075 15436 8084
rect 15384 8041 15393 8075
rect 15393 8041 15427 8075
rect 15427 8041 15436 8075
rect 15384 8032 15436 8041
rect 16488 8075 16540 8084
rect 16488 8041 16497 8075
rect 16497 8041 16531 8075
rect 16531 8041 16540 8075
rect 16488 8032 16540 8041
rect 18052 8075 18104 8084
rect 18052 8041 18061 8075
rect 18061 8041 18095 8075
rect 18095 8041 18104 8075
rect 18052 8032 18104 8041
rect 18696 8075 18748 8084
rect 18696 8041 18705 8075
rect 18705 8041 18739 8075
rect 18739 8041 18748 8075
rect 18696 8032 18748 8041
rect 19156 8075 19208 8084
rect 19156 8041 19165 8075
rect 19165 8041 19199 8075
rect 19199 8041 19208 8075
rect 19156 8032 19208 8041
rect 21088 8032 21140 8084
rect 23664 8075 23716 8084
rect 12164 7964 12216 8016
rect 13360 7964 13412 8016
rect 5172 7896 5224 7948
rect 7932 7896 7984 7948
rect 8760 7896 8812 7948
rect 9956 7939 10008 7948
rect 6552 7828 6604 7880
rect 7380 7828 7432 7880
rect 6644 7692 6696 7744
rect 8760 7735 8812 7744
rect 8760 7701 8769 7735
rect 8769 7701 8803 7735
rect 8803 7701 8812 7735
rect 8760 7692 8812 7701
rect 9312 7692 9364 7744
rect 9956 7905 9965 7939
rect 9965 7905 9999 7939
rect 9999 7905 10008 7939
rect 9956 7896 10008 7905
rect 10140 7896 10192 7948
rect 15292 7939 15344 7948
rect 15292 7905 15301 7939
rect 15301 7905 15335 7939
rect 15335 7905 15344 7939
rect 15292 7896 15344 7905
rect 15752 7939 15804 7948
rect 15752 7905 15761 7939
rect 15761 7905 15795 7939
rect 15795 7905 15804 7939
rect 15752 7896 15804 7905
rect 21180 7964 21232 8016
rect 21456 7964 21508 8016
rect 23664 8041 23673 8075
rect 23673 8041 23707 8075
rect 23707 8041 23716 8075
rect 23664 8032 23716 8041
rect 23388 7964 23440 8016
rect 23480 7964 23532 8016
rect 24676 7964 24728 8016
rect 24952 8007 25004 8016
rect 24952 7973 24961 8007
rect 24961 7973 24995 8007
rect 24995 7973 25004 8007
rect 24952 7964 25004 7973
rect 17132 7896 17184 7948
rect 17408 7896 17460 7948
rect 17868 7896 17920 7948
rect 19248 7939 19300 7948
rect 19248 7905 19257 7939
rect 19257 7905 19291 7939
rect 19291 7905 19300 7939
rect 19248 7896 19300 7905
rect 19800 7939 19852 7948
rect 19800 7905 19809 7939
rect 19809 7905 19843 7939
rect 19843 7905 19852 7939
rect 19800 7896 19852 7905
rect 11888 7828 11940 7880
rect 13728 7871 13780 7880
rect 13728 7837 13737 7871
rect 13737 7837 13771 7871
rect 13771 7837 13780 7871
rect 13728 7828 13780 7837
rect 17592 7871 17644 7880
rect 17592 7837 17601 7871
rect 17601 7837 17635 7871
rect 17635 7837 17644 7871
rect 17592 7828 17644 7837
rect 19984 7871 20036 7880
rect 19984 7837 19993 7871
rect 19993 7837 20027 7871
rect 20027 7837 20036 7871
rect 19984 7828 20036 7837
rect 21180 7871 21232 7880
rect 21180 7837 21189 7871
rect 21189 7837 21223 7871
rect 21223 7837 21232 7871
rect 21180 7828 21232 7837
rect 14280 7803 14332 7812
rect 14280 7769 14289 7803
rect 14289 7769 14323 7803
rect 14323 7769 14332 7803
rect 14280 7760 14332 7769
rect 14648 7760 14700 7812
rect 16672 7760 16724 7812
rect 20260 7760 20312 7812
rect 20904 7760 20956 7812
rect 23112 7828 23164 7880
rect 25044 7828 25096 7880
rect 18512 7692 18564 7744
rect 22100 7735 22152 7744
rect 22100 7701 22109 7735
rect 22109 7701 22143 7735
rect 22143 7701 22152 7735
rect 22100 7692 22152 7701
rect 22744 7692 22796 7744
rect 24124 7735 24176 7744
rect 24124 7701 24133 7735
rect 24133 7701 24167 7735
rect 24167 7701 24176 7735
rect 24124 7692 24176 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 1400 7488 1452 7540
rect 4160 7488 4212 7540
rect 3792 7420 3844 7472
rect 5172 7488 5224 7540
rect 5356 7488 5408 7540
rect 5540 7488 5592 7540
rect 6552 7531 6604 7540
rect 6552 7497 6561 7531
rect 6561 7497 6595 7531
rect 6595 7497 6604 7531
rect 6552 7488 6604 7497
rect 8024 7488 8076 7540
rect 11888 7531 11940 7540
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 12440 7488 12492 7540
rect 13728 7488 13780 7540
rect 17408 7531 17460 7540
rect 17408 7497 17417 7531
rect 17417 7497 17451 7531
rect 17451 7497 17460 7531
rect 17408 7488 17460 7497
rect 17868 7531 17920 7540
rect 17868 7497 17877 7531
rect 17877 7497 17911 7531
rect 17911 7497 17920 7531
rect 19800 7531 19852 7540
rect 17868 7488 17920 7497
rect 19800 7497 19809 7531
rect 19809 7497 19843 7531
rect 19843 7497 19852 7531
rect 19800 7488 19852 7497
rect 23388 7531 23440 7540
rect 23388 7497 23397 7531
rect 23397 7497 23431 7531
rect 23431 7497 23440 7531
rect 23388 7488 23440 7497
rect 24124 7488 24176 7540
rect 11980 7420 12032 7472
rect 14832 7463 14884 7472
rect 14832 7429 14841 7463
rect 14841 7429 14875 7463
rect 14875 7429 14884 7463
rect 14832 7420 14884 7429
rect 15844 7420 15896 7472
rect 20996 7420 21048 7472
rect 6644 7352 6696 7404
rect 8668 7352 8720 7404
rect 5540 7284 5592 7336
rect 6736 7284 6788 7336
rect 9312 7284 9364 7336
rect 14280 7395 14332 7404
rect 14280 7361 14289 7395
rect 14289 7361 14323 7395
rect 14323 7361 14332 7395
rect 14280 7352 14332 7361
rect 6092 7148 6144 7200
rect 7012 7259 7064 7268
rect 7012 7225 7021 7259
rect 7021 7225 7055 7259
rect 7055 7225 7064 7259
rect 7012 7216 7064 7225
rect 7380 7216 7432 7268
rect 8484 7259 8536 7268
rect 8484 7225 8493 7259
rect 8493 7225 8527 7259
rect 8527 7225 8536 7259
rect 8484 7216 8536 7225
rect 8116 7148 8168 7200
rect 8760 7216 8812 7268
rect 13360 7284 13412 7336
rect 15844 7327 15896 7336
rect 15844 7293 15853 7327
rect 15853 7293 15887 7327
rect 15887 7293 15896 7327
rect 15844 7284 15896 7293
rect 16948 7352 17000 7404
rect 19156 7352 19208 7404
rect 16856 7327 16908 7336
rect 16856 7293 16865 7327
rect 16865 7293 16899 7327
rect 16899 7293 16908 7327
rect 16856 7284 16908 7293
rect 17868 7284 17920 7336
rect 20260 7352 20312 7404
rect 24676 7463 24728 7472
rect 24676 7429 24685 7463
rect 24685 7429 24719 7463
rect 24719 7429 24728 7463
rect 24676 7420 24728 7429
rect 25044 7463 25096 7472
rect 25044 7429 25053 7463
rect 25053 7429 25087 7463
rect 25087 7429 25096 7463
rect 25044 7420 25096 7429
rect 24952 7352 25004 7404
rect 10692 7259 10744 7268
rect 8852 7148 8904 7200
rect 10692 7225 10701 7259
rect 10701 7225 10735 7259
rect 10735 7225 10744 7259
rect 10692 7216 10744 7225
rect 13912 7259 13964 7268
rect 13912 7225 13921 7259
rect 13921 7225 13955 7259
rect 13955 7225 13964 7259
rect 13912 7216 13964 7225
rect 10140 7148 10192 7200
rect 12164 7148 12216 7200
rect 12716 7148 12768 7200
rect 13360 7191 13412 7200
rect 13360 7157 13369 7191
rect 13369 7157 13403 7191
rect 13403 7157 13412 7191
rect 13360 7148 13412 7157
rect 18420 7216 18472 7268
rect 18512 7259 18564 7268
rect 18512 7225 18521 7259
rect 18521 7225 18555 7259
rect 18555 7225 18564 7259
rect 18512 7216 18564 7225
rect 19248 7216 19300 7268
rect 20444 7259 20496 7268
rect 20444 7225 20453 7259
rect 20453 7225 20487 7259
rect 20487 7225 20496 7259
rect 20444 7216 20496 7225
rect 14832 7148 14884 7200
rect 15292 7148 15344 7200
rect 21640 7216 21692 7268
rect 22100 7259 22152 7268
rect 22100 7225 22109 7259
rect 22109 7225 22143 7259
rect 22143 7225 22152 7259
rect 22100 7216 22152 7225
rect 22744 7259 22796 7268
rect 21088 7148 21140 7200
rect 21456 7191 21508 7200
rect 21456 7157 21465 7191
rect 21465 7157 21499 7191
rect 21499 7157 21508 7191
rect 21456 7148 21508 7157
rect 21732 7148 21784 7200
rect 22744 7225 22753 7259
rect 22753 7225 22787 7259
rect 22787 7225 22796 7259
rect 22744 7216 22796 7225
rect 23112 7191 23164 7200
rect 23112 7157 23121 7191
rect 23121 7157 23155 7191
rect 23155 7157 23164 7191
rect 23112 7148 23164 7157
rect 23664 7148 23716 7200
rect 25964 7148 26016 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 664 6944 716 6996
rect 5540 6944 5592 6996
rect 6276 6987 6328 6996
rect 6276 6953 6285 6987
rect 6285 6953 6319 6987
rect 6319 6953 6328 6987
rect 6276 6944 6328 6953
rect 4712 6808 4764 6860
rect 5448 6876 5500 6928
rect 6092 6876 6144 6928
rect 8484 6944 8536 6996
rect 11980 6987 12032 6996
rect 11980 6953 11989 6987
rect 11989 6953 12023 6987
rect 12023 6953 12032 6987
rect 11980 6944 12032 6953
rect 13452 6987 13504 6996
rect 13452 6953 13461 6987
rect 13461 6953 13495 6987
rect 13495 6953 13504 6987
rect 13452 6944 13504 6953
rect 13912 6944 13964 6996
rect 14740 6944 14792 6996
rect 15384 6944 15436 6996
rect 17500 6944 17552 6996
rect 21180 6987 21232 6996
rect 21180 6953 21189 6987
rect 21189 6953 21223 6987
rect 21223 6953 21232 6987
rect 21180 6944 21232 6953
rect 21456 6944 21508 6996
rect 23480 6944 23532 6996
rect 7012 6876 7064 6928
rect 7380 6919 7432 6928
rect 7380 6885 7389 6919
rect 7389 6885 7423 6919
rect 7423 6885 7432 6919
rect 7380 6876 7432 6885
rect 7932 6919 7984 6928
rect 7932 6885 7941 6919
rect 7941 6885 7975 6919
rect 7975 6885 7984 6919
rect 7932 6876 7984 6885
rect 8116 6876 8168 6928
rect 5540 6808 5592 6860
rect 10048 6876 10100 6928
rect 11428 6876 11480 6928
rect 13544 6876 13596 6928
rect 17684 6876 17736 6928
rect 18972 6876 19024 6928
rect 22100 6919 22152 6928
rect 22100 6885 22109 6919
rect 22109 6885 22143 6919
rect 22143 6885 22152 6919
rect 22100 6876 22152 6885
rect 23848 6919 23900 6928
rect 23848 6885 23857 6919
rect 23857 6885 23891 6919
rect 23891 6885 23900 6919
rect 23848 6876 23900 6885
rect 8300 6740 8352 6792
rect 4804 6672 4856 6724
rect 5080 6672 5132 6724
rect 9312 6672 9364 6724
rect 10692 6740 10744 6792
rect 11612 6851 11664 6860
rect 11612 6817 11621 6851
rect 11621 6817 11655 6851
rect 11655 6817 11664 6851
rect 11796 6851 11848 6860
rect 11612 6808 11664 6817
rect 11796 6817 11805 6851
rect 11805 6817 11839 6851
rect 11839 6817 11848 6851
rect 11796 6808 11848 6817
rect 16304 6851 16356 6860
rect 16304 6817 16313 6851
rect 16313 6817 16347 6851
rect 16347 6817 16356 6851
rect 16304 6808 16356 6817
rect 13176 6783 13228 6792
rect 12348 6672 12400 6724
rect 13176 6749 13185 6783
rect 13185 6749 13219 6783
rect 13219 6749 13228 6783
rect 13176 6740 13228 6749
rect 16856 6808 16908 6860
rect 17592 6851 17644 6860
rect 17592 6817 17601 6851
rect 17601 6817 17635 6851
rect 17635 6817 17644 6851
rect 17592 6808 17644 6817
rect 19432 6808 19484 6860
rect 21824 6851 21876 6860
rect 21824 6817 21833 6851
rect 21833 6817 21867 6851
rect 21867 6817 21876 6851
rect 21824 6808 21876 6817
rect 25780 6808 25832 6860
rect 18052 6740 18104 6792
rect 23204 6740 23256 6792
rect 24032 6783 24084 6792
rect 24032 6749 24041 6783
rect 24041 6749 24075 6783
rect 24075 6749 24084 6783
rect 24032 6740 24084 6749
rect 14280 6715 14332 6724
rect 14280 6681 14289 6715
rect 14289 6681 14323 6715
rect 14323 6681 14332 6715
rect 14280 6672 14332 6681
rect 20444 6715 20496 6724
rect 20444 6681 20453 6715
rect 20453 6681 20487 6715
rect 20487 6681 20496 6715
rect 20444 6672 20496 6681
rect 9220 6647 9272 6656
rect 9220 6613 9229 6647
rect 9229 6613 9263 6647
rect 9263 6613 9272 6647
rect 9220 6604 9272 6613
rect 9588 6604 9640 6656
rect 13360 6604 13412 6656
rect 18512 6647 18564 6656
rect 18512 6613 18521 6647
rect 18521 6613 18555 6647
rect 18555 6613 18564 6647
rect 18512 6604 18564 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 4712 6443 4764 6452
rect 4712 6409 4721 6443
rect 4721 6409 4755 6443
rect 4755 6409 4764 6443
rect 4712 6400 4764 6409
rect 5080 6443 5132 6452
rect 5080 6409 5089 6443
rect 5089 6409 5123 6443
rect 5123 6409 5132 6443
rect 5080 6400 5132 6409
rect 7932 6400 7984 6452
rect 8300 6443 8352 6452
rect 8300 6409 8309 6443
rect 8309 6409 8343 6443
rect 8343 6409 8352 6443
rect 8300 6400 8352 6409
rect 11612 6400 11664 6452
rect 13176 6400 13228 6452
rect 17040 6443 17092 6452
rect 6000 6332 6052 6384
rect 7380 6332 7432 6384
rect 7472 6332 7524 6384
rect 9220 6332 9272 6384
rect 3976 6103 4028 6112
rect 3976 6069 3985 6103
rect 3985 6069 4019 6103
rect 4019 6069 4028 6103
rect 4896 6196 4948 6248
rect 6368 6264 6420 6316
rect 6460 6264 6512 6316
rect 7564 6264 7616 6316
rect 9588 6264 9640 6316
rect 5540 6196 5592 6248
rect 11612 6264 11664 6316
rect 13360 6332 13412 6384
rect 16120 6332 16172 6384
rect 16304 6375 16356 6384
rect 16304 6341 16313 6375
rect 16313 6341 16347 6375
rect 16347 6341 16356 6375
rect 16304 6332 16356 6341
rect 16764 6375 16816 6384
rect 16764 6341 16773 6375
rect 16773 6341 16807 6375
rect 16807 6341 16816 6375
rect 16764 6332 16816 6341
rect 15384 6307 15436 6316
rect 15384 6273 15393 6307
rect 15393 6273 15427 6307
rect 15427 6273 15436 6307
rect 15384 6264 15436 6273
rect 6460 6128 6512 6180
rect 6920 6171 6972 6180
rect 3976 6060 4028 6069
rect 4528 6060 4580 6112
rect 5080 6060 5132 6112
rect 6920 6137 6929 6171
rect 6929 6137 6963 6171
rect 6963 6137 6972 6171
rect 6920 6128 6972 6137
rect 7012 6171 7064 6180
rect 7012 6137 7021 6171
rect 7021 6137 7055 6171
rect 7055 6137 7064 6171
rect 7012 6128 7064 6137
rect 7564 6128 7616 6180
rect 8668 6103 8720 6112
rect 8668 6069 8677 6103
rect 8677 6069 8711 6103
rect 8711 6069 8720 6103
rect 8668 6060 8720 6069
rect 9036 6103 9088 6112
rect 9036 6069 9045 6103
rect 9045 6069 9079 6103
rect 9079 6069 9088 6103
rect 11796 6196 11848 6248
rect 11244 6128 11296 6180
rect 9036 6060 9088 6069
rect 10048 6060 10100 6112
rect 12716 6060 12768 6112
rect 13176 6060 13228 6112
rect 13268 6060 13320 6112
rect 13820 6196 13872 6248
rect 14096 6239 14148 6248
rect 14096 6205 14105 6239
rect 14105 6205 14139 6239
rect 14139 6205 14148 6239
rect 17040 6409 17049 6443
rect 17049 6409 17083 6443
rect 17083 6409 17092 6443
rect 17040 6400 17092 6409
rect 23848 6400 23900 6452
rect 25044 6400 25096 6452
rect 25872 6400 25924 6452
rect 19432 6375 19484 6384
rect 19432 6341 19441 6375
rect 19441 6341 19475 6375
rect 19475 6341 19484 6375
rect 19432 6332 19484 6341
rect 23480 6332 23532 6384
rect 23572 6332 23624 6384
rect 18052 6307 18104 6316
rect 18052 6273 18061 6307
rect 18061 6273 18095 6307
rect 18095 6273 18104 6307
rect 18052 6264 18104 6273
rect 18420 6264 18472 6316
rect 19524 6264 19576 6316
rect 14096 6196 14148 6205
rect 17960 6196 18012 6248
rect 22192 6264 22244 6316
rect 23848 6264 23900 6316
rect 24032 6264 24084 6316
rect 15200 6128 15252 6180
rect 15476 6171 15528 6180
rect 15476 6137 15485 6171
rect 15485 6137 15519 6171
rect 15519 6137 15528 6171
rect 15476 6128 15528 6137
rect 16764 6128 16816 6180
rect 14832 6060 14884 6112
rect 15292 6060 15344 6112
rect 15660 6060 15712 6112
rect 17684 6103 17736 6112
rect 17684 6069 17693 6103
rect 17693 6069 17727 6103
rect 17727 6069 17736 6103
rect 17684 6060 17736 6069
rect 18236 6060 18288 6112
rect 21732 6128 21784 6180
rect 25872 6196 25924 6248
rect 23572 6128 23624 6180
rect 20720 6103 20772 6112
rect 20720 6069 20729 6103
rect 20729 6069 20763 6103
rect 20763 6069 20772 6103
rect 20720 6060 20772 6069
rect 21272 6103 21324 6112
rect 21272 6069 21281 6103
rect 21281 6069 21315 6103
rect 21315 6069 21324 6103
rect 21272 6060 21324 6069
rect 22100 6060 22152 6112
rect 22560 6060 22612 6112
rect 23204 6060 23256 6112
rect 23756 6060 23808 6112
rect 25780 6103 25832 6112
rect 25780 6069 25789 6103
rect 25789 6069 25823 6103
rect 25823 6069 25832 6103
rect 25780 6060 25832 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 3240 5788 3292 5840
rect 8668 5856 8720 5908
rect 4528 5788 4580 5840
rect 6920 5788 6972 5840
rect 7196 5831 7248 5840
rect 7196 5797 7205 5831
rect 7205 5797 7239 5831
rect 7239 5797 7248 5831
rect 7196 5788 7248 5797
rect 7564 5831 7616 5840
rect 7564 5797 7573 5831
rect 7573 5797 7607 5831
rect 7607 5797 7616 5831
rect 7564 5788 7616 5797
rect 7932 5831 7984 5840
rect 7932 5797 7941 5831
rect 7941 5797 7975 5831
rect 7975 5797 7984 5831
rect 7932 5788 7984 5797
rect 4620 5720 4672 5772
rect 5172 5763 5224 5772
rect 5172 5729 5181 5763
rect 5181 5729 5215 5763
rect 5215 5729 5224 5763
rect 5172 5720 5224 5729
rect 6368 5720 6420 5772
rect 6460 5763 6512 5772
rect 6460 5729 6469 5763
rect 6469 5729 6503 5763
rect 6503 5729 6512 5763
rect 6460 5720 6512 5729
rect 8024 5763 8076 5772
rect 4712 5652 4764 5704
rect 6644 5652 6696 5704
rect 8024 5729 8033 5763
rect 8033 5729 8067 5763
rect 8067 5729 8076 5763
rect 8024 5720 8076 5729
rect 8392 5720 8444 5772
rect 9404 5856 9456 5908
rect 10692 5899 10744 5908
rect 10692 5865 10701 5899
rect 10701 5865 10735 5899
rect 10735 5865 10744 5899
rect 10692 5856 10744 5865
rect 11428 5856 11480 5908
rect 13544 5899 13596 5908
rect 13544 5865 13553 5899
rect 13553 5865 13587 5899
rect 13587 5865 13596 5899
rect 13544 5856 13596 5865
rect 15660 5899 15712 5908
rect 15660 5865 15669 5899
rect 15669 5865 15703 5899
rect 15703 5865 15712 5899
rect 15660 5856 15712 5865
rect 17592 5899 17644 5908
rect 17592 5865 17601 5899
rect 17601 5865 17635 5899
rect 17635 5865 17644 5899
rect 17592 5856 17644 5865
rect 18144 5856 18196 5908
rect 19340 5899 19392 5908
rect 19340 5865 19349 5899
rect 19349 5865 19383 5899
rect 19383 5865 19392 5899
rect 19340 5856 19392 5865
rect 19524 5856 19576 5908
rect 20260 5899 20312 5908
rect 20260 5865 20269 5899
rect 20269 5865 20303 5899
rect 20303 5865 20312 5899
rect 20260 5856 20312 5865
rect 21272 5899 21324 5908
rect 21272 5865 21281 5899
rect 21281 5865 21315 5899
rect 21315 5865 21324 5899
rect 21272 5856 21324 5865
rect 21824 5856 21876 5908
rect 22192 5856 22244 5908
rect 23112 5899 23164 5908
rect 23112 5865 23121 5899
rect 23121 5865 23155 5899
rect 23155 5865 23164 5899
rect 23112 5856 23164 5865
rect 23756 5899 23808 5908
rect 23756 5865 23765 5899
rect 23765 5865 23799 5899
rect 23799 5865 23808 5899
rect 23756 5856 23808 5865
rect 13820 5831 13872 5840
rect 13820 5797 13829 5831
rect 13829 5797 13863 5831
rect 13863 5797 13872 5831
rect 13820 5788 13872 5797
rect 17224 5788 17276 5840
rect 17776 5788 17828 5840
rect 18236 5788 18288 5840
rect 24216 5831 24268 5840
rect 24216 5797 24225 5831
rect 24225 5797 24259 5831
rect 24259 5797 24268 5831
rect 24216 5788 24268 5797
rect 24676 5788 24728 5840
rect 9036 5652 9088 5704
rect 11336 5720 11388 5772
rect 12164 5720 12216 5772
rect 13544 5720 13596 5772
rect 15200 5720 15252 5772
rect 12808 5695 12860 5704
rect 4988 5627 5040 5636
rect 4988 5593 4997 5627
rect 4997 5593 5031 5627
rect 5031 5593 5040 5627
rect 4988 5584 5040 5593
rect 6552 5627 6604 5636
rect 6552 5593 6561 5627
rect 6561 5593 6595 5627
rect 6595 5593 6604 5627
rect 6552 5584 6604 5593
rect 7380 5584 7432 5636
rect 7932 5584 7984 5636
rect 12808 5661 12817 5695
rect 12817 5661 12851 5695
rect 12851 5661 12860 5695
rect 12808 5652 12860 5661
rect 13728 5695 13780 5704
rect 13728 5661 13737 5695
rect 13737 5661 13771 5695
rect 13771 5661 13780 5695
rect 13728 5652 13780 5661
rect 19708 5720 19760 5772
rect 19984 5720 20036 5772
rect 21088 5720 21140 5772
rect 21824 5763 21876 5772
rect 21824 5729 21833 5763
rect 21833 5729 21867 5763
rect 21867 5729 21876 5763
rect 21824 5720 21876 5729
rect 22100 5720 22152 5772
rect 9772 5627 9824 5636
rect 9772 5593 9781 5627
rect 9781 5593 9815 5627
rect 9815 5593 9824 5627
rect 9772 5584 9824 5593
rect 11704 5584 11756 5636
rect 21364 5652 21416 5704
rect 22744 5652 22796 5704
rect 16120 5584 16172 5636
rect 5540 5516 5592 5568
rect 9404 5559 9456 5568
rect 9404 5525 9413 5559
rect 9413 5525 9447 5559
rect 9447 5525 9456 5559
rect 9404 5516 9456 5525
rect 13084 5559 13136 5568
rect 13084 5525 13093 5559
rect 13093 5525 13127 5559
rect 13127 5525 13136 5559
rect 13084 5516 13136 5525
rect 16212 5559 16264 5568
rect 16212 5525 16221 5559
rect 16221 5525 16255 5559
rect 16255 5525 16264 5559
rect 16212 5516 16264 5525
rect 19340 5516 19392 5568
rect 23572 5516 23624 5568
rect 25504 5516 25556 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 1676 5355 1728 5364
rect 1676 5321 1685 5355
rect 1685 5321 1719 5355
rect 1719 5321 1728 5355
rect 1676 5312 1728 5321
rect 3240 5355 3292 5364
rect 3240 5321 3249 5355
rect 3249 5321 3283 5355
rect 3283 5321 3292 5355
rect 3240 5312 3292 5321
rect 3884 5312 3936 5364
rect 5172 5312 5224 5364
rect 9404 5312 9456 5364
rect 11336 5312 11388 5364
rect 14464 5312 14516 5364
rect 15384 5312 15436 5364
rect 17776 5355 17828 5364
rect 17776 5321 17785 5355
rect 17785 5321 17819 5355
rect 17819 5321 17828 5355
rect 17776 5312 17828 5321
rect 18236 5355 18288 5364
rect 18236 5321 18245 5355
rect 18245 5321 18279 5355
rect 18279 5321 18288 5355
rect 18236 5312 18288 5321
rect 19708 5355 19760 5364
rect 19708 5321 19717 5355
rect 19717 5321 19751 5355
rect 19751 5321 19760 5355
rect 19708 5312 19760 5321
rect 19984 5312 20036 5364
rect 21824 5355 21876 5364
rect 21824 5321 21833 5355
rect 21833 5321 21867 5355
rect 21867 5321 21876 5355
rect 21824 5312 21876 5321
rect 23204 5312 23256 5364
rect 25596 5312 25648 5364
rect 3148 5244 3200 5296
rect 204 5108 256 5160
rect 5080 5244 5132 5296
rect 6644 5244 6696 5296
rect 8024 5244 8076 5296
rect 8852 5244 8904 5296
rect 12532 5244 12584 5296
rect 19340 5244 19392 5296
rect 20260 5244 20312 5296
rect 20904 5287 20956 5296
rect 4712 5151 4764 5160
rect 4712 5117 4721 5151
rect 4721 5117 4755 5151
rect 4755 5117 4764 5151
rect 4712 5108 4764 5117
rect 5264 5151 5316 5160
rect 5264 5117 5273 5151
rect 5273 5117 5307 5151
rect 5307 5117 5316 5151
rect 5264 5108 5316 5117
rect 6920 5176 6972 5228
rect 7472 5151 7524 5160
rect 7472 5117 7481 5151
rect 7481 5117 7515 5151
rect 7515 5117 7524 5151
rect 7472 5108 7524 5117
rect 6184 5040 6236 5092
rect 6552 5040 6604 5092
rect 9036 5108 9088 5160
rect 9588 5151 9640 5160
rect 9588 5117 9597 5151
rect 9597 5117 9631 5151
rect 9631 5117 9640 5151
rect 9588 5108 9640 5117
rect 10692 5108 10744 5160
rect 12164 5108 12216 5160
rect 13084 5108 13136 5160
rect 14188 5176 14240 5228
rect 16120 5219 16172 5228
rect 16120 5185 16129 5219
rect 16129 5185 16163 5219
rect 16163 5185 16172 5219
rect 16120 5176 16172 5185
rect 19248 5176 19300 5228
rect 20904 5253 20913 5287
rect 20913 5253 20947 5287
rect 20947 5253 20956 5287
rect 20904 5244 20956 5253
rect 24676 5287 24728 5296
rect 24676 5253 24685 5287
rect 24685 5253 24719 5287
rect 24719 5253 24728 5287
rect 24676 5244 24728 5253
rect 21180 5176 21232 5228
rect 23848 5176 23900 5228
rect 23940 5176 23992 5228
rect 15752 5108 15804 5160
rect 25596 5108 25648 5160
rect 9772 5040 9824 5092
rect 11060 5040 11112 5092
rect 12256 5040 12308 5092
rect 4896 5015 4948 5024
rect 4896 4981 4905 5015
rect 4905 4981 4939 5015
rect 4939 4981 4948 5015
rect 4896 4972 4948 4981
rect 6368 4972 6420 5024
rect 9864 4972 9916 5024
rect 10048 4972 10100 5024
rect 10692 5015 10744 5024
rect 10692 4981 10701 5015
rect 10701 4981 10735 5015
rect 10735 4981 10744 5015
rect 10692 4972 10744 4981
rect 12716 4972 12768 5024
rect 15660 5040 15712 5092
rect 16212 5083 16264 5092
rect 16212 5049 16221 5083
rect 16221 5049 16255 5083
rect 16255 5049 16264 5083
rect 16764 5083 16816 5092
rect 16212 5040 16264 5049
rect 16764 5049 16773 5083
rect 16773 5049 16807 5083
rect 16807 5049 16816 5083
rect 16764 5040 16816 5049
rect 18880 5083 18932 5092
rect 18880 5049 18889 5083
rect 18889 5049 18923 5083
rect 18923 5049 18932 5083
rect 19432 5083 19484 5092
rect 18880 5040 18932 5049
rect 19432 5049 19441 5083
rect 19441 5049 19475 5083
rect 19475 5049 19484 5083
rect 19432 5040 19484 5049
rect 20720 5040 20772 5092
rect 22100 5083 22152 5092
rect 22100 5049 22109 5083
rect 22109 5049 22143 5083
rect 22143 5049 22152 5083
rect 22100 5040 22152 5049
rect 23756 5083 23808 5092
rect 15844 5015 15896 5024
rect 15844 4981 15853 5015
rect 15853 4981 15887 5015
rect 15887 4981 15896 5015
rect 21272 5015 21324 5024
rect 15844 4972 15896 4981
rect 21272 4981 21281 5015
rect 21281 4981 21315 5015
rect 21315 4981 21324 5015
rect 21272 4972 21324 4981
rect 21824 4972 21876 5024
rect 23756 5049 23765 5083
rect 23765 5049 23799 5083
rect 23799 5049 23808 5083
rect 23756 5040 23808 5049
rect 23388 5015 23440 5024
rect 23388 4981 23397 5015
rect 23397 4981 23431 5015
rect 23431 4981 23440 5015
rect 23388 4972 23440 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 4344 4768 4396 4820
rect 4620 4768 4672 4820
rect 4988 4768 5040 4820
rect 7472 4768 7524 4820
rect 7932 4811 7984 4820
rect 7932 4777 7941 4811
rect 7941 4777 7975 4811
rect 7975 4777 7984 4811
rect 7932 4768 7984 4777
rect 6460 4743 6512 4752
rect 6460 4709 6469 4743
rect 6469 4709 6503 4743
rect 6503 4709 6512 4743
rect 6460 4700 6512 4709
rect 2872 4632 2924 4684
rect 4068 4632 4120 4684
rect 4896 4675 4948 4684
rect 4896 4641 4905 4675
rect 4905 4641 4939 4675
rect 4939 4641 4948 4675
rect 4896 4632 4948 4641
rect 5448 4675 5500 4684
rect 5448 4641 5457 4675
rect 5457 4641 5491 4675
rect 5491 4641 5500 4675
rect 5448 4632 5500 4641
rect 6920 4632 6972 4684
rect 7104 4675 7156 4684
rect 7104 4641 7113 4675
rect 7113 4641 7147 4675
rect 7147 4641 7156 4675
rect 7104 4632 7156 4641
rect 10784 4768 10836 4820
rect 12164 4811 12216 4820
rect 12164 4777 12173 4811
rect 12173 4777 12207 4811
rect 12207 4777 12216 4811
rect 12164 4768 12216 4777
rect 12532 4811 12584 4820
rect 12532 4777 12541 4811
rect 12541 4777 12575 4811
rect 12575 4777 12584 4811
rect 12532 4768 12584 4777
rect 13820 4811 13872 4820
rect 13820 4777 13829 4811
rect 13829 4777 13863 4811
rect 13863 4777 13872 4811
rect 13820 4768 13872 4777
rect 14188 4768 14240 4820
rect 15292 4768 15344 4820
rect 15660 4768 15712 4820
rect 16764 4768 16816 4820
rect 17684 4768 17736 4820
rect 19524 4768 19576 4820
rect 20168 4768 20220 4820
rect 20720 4768 20772 4820
rect 22100 4768 22152 4820
rect 23572 4768 23624 4820
rect 24216 4811 24268 4820
rect 24216 4777 24225 4811
rect 24225 4777 24259 4811
rect 24259 4777 24268 4811
rect 24216 4768 24268 4777
rect 8484 4632 8536 4684
rect 12716 4700 12768 4752
rect 15384 4700 15436 4752
rect 16396 4700 16448 4752
rect 19156 4743 19208 4752
rect 19156 4709 19165 4743
rect 19165 4709 19199 4743
rect 19199 4709 19208 4743
rect 19156 4700 19208 4709
rect 21180 4700 21232 4752
rect 22560 4700 22612 4752
rect 22836 4743 22888 4752
rect 22836 4709 22845 4743
rect 22845 4709 22879 4743
rect 22879 4709 22888 4743
rect 22836 4700 22888 4709
rect 24032 4700 24084 4752
rect 9680 4675 9732 4684
rect 9680 4641 9689 4675
rect 9689 4641 9723 4675
rect 9723 4641 9732 4675
rect 9680 4632 9732 4641
rect 9956 4675 10008 4684
rect 9956 4641 9965 4675
rect 9965 4641 9999 4675
rect 9999 4641 10008 4675
rect 9956 4632 10008 4641
rect 11244 4675 11296 4684
rect 11244 4641 11253 4675
rect 11253 4641 11287 4675
rect 11287 4641 11296 4675
rect 11244 4632 11296 4641
rect 11796 4675 11848 4684
rect 11796 4641 11805 4675
rect 11805 4641 11839 4675
rect 11839 4641 11848 4675
rect 11796 4632 11848 4641
rect 14556 4632 14608 4684
rect 7656 4564 7708 4616
rect 8668 4607 8720 4616
rect 8668 4573 8677 4607
rect 8677 4573 8711 4607
rect 8711 4573 8720 4607
rect 8668 4564 8720 4573
rect 12624 4607 12676 4616
rect 4344 4496 4396 4548
rect 6828 4496 6880 4548
rect 7196 4496 7248 4548
rect 10692 4496 10744 4548
rect 12624 4573 12633 4607
rect 12633 4573 12667 4607
rect 12667 4573 12676 4607
rect 12624 4564 12676 4573
rect 15660 4632 15712 4684
rect 17684 4675 17736 4684
rect 17684 4641 17693 4675
rect 17693 4641 17727 4675
rect 17727 4641 17736 4675
rect 17684 4632 17736 4641
rect 22008 4632 22060 4684
rect 22192 4632 22244 4684
rect 16212 4564 16264 4616
rect 19064 4607 19116 4616
rect 19064 4573 19073 4607
rect 19073 4573 19107 4607
rect 19107 4573 19116 4607
rect 19064 4564 19116 4573
rect 19432 4607 19484 4616
rect 19432 4573 19441 4607
rect 19441 4573 19475 4607
rect 19475 4573 19484 4607
rect 19432 4564 19484 4573
rect 20720 4564 20772 4616
rect 21364 4564 21416 4616
rect 23020 4607 23072 4616
rect 9496 4428 9548 4480
rect 10048 4428 10100 4480
rect 13728 4428 13780 4480
rect 16028 4496 16080 4548
rect 20904 4496 20956 4548
rect 23020 4573 23029 4607
rect 23029 4573 23063 4607
rect 23063 4573 23072 4607
rect 23020 4564 23072 4573
rect 23940 4564 23992 4616
rect 24860 4607 24912 4616
rect 22928 4496 22980 4548
rect 23756 4539 23808 4548
rect 23756 4505 23765 4539
rect 23765 4505 23799 4539
rect 23799 4505 23808 4539
rect 23756 4496 23808 4505
rect 24216 4496 24268 4548
rect 24860 4573 24869 4607
rect 24869 4573 24903 4607
rect 24903 4573 24912 4607
rect 24860 4564 24912 4573
rect 25228 4496 25280 4548
rect 16580 4428 16632 4480
rect 17500 4428 17552 4480
rect 18788 4471 18840 4480
rect 18788 4437 18797 4471
rect 18797 4437 18831 4471
rect 18831 4437 18840 4471
rect 18788 4428 18840 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 3608 4267 3660 4276
rect 3608 4233 3617 4267
rect 3617 4233 3651 4267
rect 3651 4233 3660 4267
rect 3608 4224 3660 4233
rect 4068 4267 4120 4276
rect 4068 4233 4077 4267
rect 4077 4233 4111 4267
rect 4111 4233 4120 4267
rect 4068 4224 4120 4233
rect 5540 4224 5592 4276
rect 7564 4267 7616 4276
rect 7564 4233 7573 4267
rect 7573 4233 7607 4267
rect 7607 4233 7616 4267
rect 7564 4224 7616 4233
rect 9956 4224 10008 4276
rect 10692 4267 10744 4276
rect 10692 4233 10701 4267
rect 10701 4233 10735 4267
rect 10735 4233 10744 4267
rect 10692 4224 10744 4233
rect 11152 4267 11204 4276
rect 11152 4233 11161 4267
rect 11161 4233 11195 4267
rect 11195 4233 11204 4267
rect 11152 4224 11204 4233
rect 9404 4199 9456 4208
rect 9404 4165 9413 4199
rect 9413 4165 9447 4199
rect 9447 4165 9456 4199
rect 9404 4156 9456 4165
rect 9680 4156 9732 4208
rect 9864 4156 9916 4208
rect 11244 4156 11296 4208
rect 14372 4224 14424 4276
rect 16212 4224 16264 4276
rect 16396 4267 16448 4276
rect 16396 4233 16405 4267
rect 16405 4233 16439 4267
rect 16439 4233 16448 4267
rect 16396 4224 16448 4233
rect 17316 4224 17368 4276
rect 21180 4267 21232 4276
rect 21180 4233 21189 4267
rect 21189 4233 21223 4267
rect 21223 4233 21232 4267
rect 21180 4224 21232 4233
rect 22836 4267 22888 4276
rect 22836 4233 22845 4267
rect 22845 4233 22879 4267
rect 22879 4233 22888 4267
rect 22836 4224 22888 4233
rect 25228 4224 25280 4276
rect 14464 4156 14516 4208
rect 22928 4156 22980 4208
rect 2872 4088 2924 4140
rect 3332 4088 3384 4140
rect 3700 4088 3752 4140
rect 5080 4088 5132 4140
rect 3608 4020 3660 4072
rect 4252 4063 4304 4072
rect 4252 4029 4270 4063
rect 4270 4029 4304 4063
rect 4252 4020 4304 4029
rect 4712 4020 4764 4072
rect 4988 4020 5040 4072
rect 5724 4063 5776 4072
rect 5724 4029 5733 4063
rect 5733 4029 5767 4063
rect 5767 4029 5776 4063
rect 5724 4020 5776 4029
rect 7564 4088 7616 4140
rect 7932 4020 7984 4072
rect 8484 4088 8536 4140
rect 8668 4020 8720 4072
rect 12624 4088 12676 4140
rect 13360 4131 13412 4140
rect 9312 4063 9364 4072
rect 9312 4029 9321 4063
rect 9321 4029 9355 4063
rect 9355 4029 9364 4063
rect 9312 4020 9364 4029
rect 9496 4020 9548 4072
rect 9956 4020 10008 4072
rect 10784 4020 10836 4072
rect 12532 4020 12584 4072
rect 13360 4097 13369 4131
rect 13369 4097 13403 4131
rect 13403 4097 13412 4131
rect 13360 4088 13412 4097
rect 13452 4088 13504 4140
rect 19432 4088 19484 4140
rect 22192 4088 22244 4140
rect 24860 4156 24912 4208
rect 16580 4020 16632 4072
rect 5540 3952 5592 4004
rect 6000 3952 6052 4004
rect 3792 3884 3844 3936
rect 4528 3884 4580 3936
rect 4712 3927 4764 3936
rect 4712 3893 4721 3927
rect 4721 3893 4755 3927
rect 4755 3893 4764 3927
rect 4712 3884 4764 3893
rect 4988 3927 5040 3936
rect 4988 3893 4997 3927
rect 4997 3893 5031 3927
rect 5031 3893 5040 3927
rect 4988 3884 5040 3893
rect 7104 3884 7156 3936
rect 8300 3884 8352 3936
rect 12072 3952 12124 4004
rect 9772 3927 9824 3936
rect 9772 3893 9781 3927
rect 9781 3893 9815 3927
rect 9815 3893 9824 3927
rect 9772 3884 9824 3893
rect 12716 3884 12768 3936
rect 12900 3884 12952 3936
rect 14004 3995 14056 4004
rect 14004 3961 14013 3995
rect 14013 3961 14047 3995
rect 14047 3961 14056 3995
rect 14556 3995 14608 4004
rect 14004 3952 14056 3961
rect 14556 3961 14565 3995
rect 14565 3961 14599 3995
rect 14599 3961 14608 3995
rect 14556 3952 14608 3961
rect 14832 3927 14884 3936
rect 14832 3893 14841 3927
rect 14841 3893 14875 3927
rect 14875 3893 14884 3927
rect 14832 3884 14884 3893
rect 15292 3927 15344 3936
rect 15292 3893 15301 3927
rect 15301 3893 15335 3927
rect 15335 3893 15344 3927
rect 15844 3952 15896 4004
rect 16120 3995 16172 4004
rect 16120 3961 16129 3995
rect 16129 3961 16163 3995
rect 16163 3961 16172 3995
rect 16120 3952 16172 3961
rect 15292 3884 15344 3893
rect 16028 3884 16080 3936
rect 18604 3884 18656 3936
rect 19524 3927 19576 3936
rect 19524 3893 19533 3927
rect 19533 3893 19567 3927
rect 19567 3893 19576 3927
rect 19524 3884 19576 3893
rect 20168 3995 20220 4004
rect 20168 3961 20177 3995
rect 20177 3961 20211 3995
rect 20211 3961 20220 3995
rect 20168 3952 20220 3961
rect 21272 3884 21324 3936
rect 22100 3884 22152 3936
rect 22928 3884 22980 3936
rect 23756 3952 23808 4004
rect 24492 3995 24544 4004
rect 24032 3884 24084 3936
rect 24492 3961 24501 3995
rect 24501 3961 24535 3995
rect 24535 3961 24544 3995
rect 24492 3952 24544 3961
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 5724 3680 5776 3732
rect 9404 3723 9456 3732
rect 9404 3689 9413 3723
rect 9413 3689 9447 3723
rect 9447 3689 9456 3723
rect 9404 3680 9456 3689
rect 11428 3723 11480 3732
rect 11428 3689 11437 3723
rect 11437 3689 11471 3723
rect 11471 3689 11480 3723
rect 11428 3680 11480 3689
rect 12072 3723 12124 3732
rect 12072 3689 12081 3723
rect 12081 3689 12115 3723
rect 12115 3689 12124 3723
rect 12072 3680 12124 3689
rect 12808 3680 12860 3732
rect 14648 3680 14700 3732
rect 18604 3723 18656 3732
rect 18604 3689 18613 3723
rect 18613 3689 18647 3723
rect 18647 3689 18656 3723
rect 18604 3680 18656 3689
rect 19064 3680 19116 3732
rect 20720 3723 20772 3732
rect 20720 3689 20729 3723
rect 20729 3689 20763 3723
rect 20763 3689 20772 3723
rect 20720 3680 20772 3689
rect 22100 3723 22152 3732
rect 22100 3689 22109 3723
rect 22109 3689 22143 3723
rect 22143 3689 22152 3723
rect 22100 3680 22152 3689
rect 23388 3680 23440 3732
rect 24492 3680 24544 3732
rect 8668 3612 8720 3664
rect 2228 3544 2280 3596
rect 2964 3587 3016 3596
rect 2964 3553 2973 3587
rect 2973 3553 3007 3587
rect 3007 3553 3016 3587
rect 2964 3544 3016 3553
rect 5264 3544 5316 3596
rect 3148 3476 3200 3528
rect 3976 3476 4028 3528
rect 5724 3544 5776 3596
rect 7012 3587 7064 3596
rect 7012 3553 7021 3587
rect 7021 3553 7055 3587
rect 7055 3553 7064 3587
rect 7012 3544 7064 3553
rect 7196 3587 7248 3596
rect 7196 3553 7205 3587
rect 7205 3553 7239 3587
rect 7239 3553 7248 3587
rect 7196 3544 7248 3553
rect 8024 3587 8076 3596
rect 8024 3553 8033 3587
rect 8033 3553 8067 3587
rect 8067 3553 8076 3587
rect 8024 3544 8076 3553
rect 8300 3587 8352 3596
rect 8300 3553 8309 3587
rect 8309 3553 8343 3587
rect 8343 3553 8352 3587
rect 8300 3544 8352 3553
rect 9680 3587 9732 3596
rect 9680 3553 9689 3587
rect 9689 3553 9723 3587
rect 9723 3553 9732 3587
rect 9680 3544 9732 3553
rect 9956 3587 10008 3596
rect 9956 3553 9965 3587
rect 9965 3553 9999 3587
rect 9999 3553 10008 3587
rect 9956 3544 10008 3553
rect 12716 3612 12768 3664
rect 14004 3612 14056 3664
rect 15384 3612 15436 3664
rect 15752 3612 15804 3664
rect 14096 3587 14148 3596
rect 14096 3553 14105 3587
rect 14105 3553 14139 3587
rect 14139 3553 14148 3587
rect 14096 3544 14148 3553
rect 15016 3587 15068 3596
rect 15016 3553 15025 3587
rect 15025 3553 15059 3587
rect 15059 3553 15068 3587
rect 15016 3544 15068 3553
rect 17132 3587 17184 3596
rect 17132 3553 17141 3587
rect 17141 3553 17175 3587
rect 17175 3553 17184 3587
rect 17132 3544 17184 3553
rect 19340 3612 19392 3664
rect 20168 3655 20220 3664
rect 20168 3621 20177 3655
rect 20177 3621 20211 3655
rect 20211 3621 20220 3655
rect 20168 3612 20220 3621
rect 18972 3544 19024 3596
rect 19156 3587 19208 3596
rect 19156 3553 19165 3587
rect 19165 3553 19199 3587
rect 19199 3553 19208 3587
rect 19156 3544 19208 3553
rect 19524 3544 19576 3596
rect 23756 3612 23808 3664
rect 24216 3612 24268 3664
rect 6276 3476 6328 3528
rect 6368 3476 6420 3528
rect 12256 3519 12308 3528
rect 12256 3485 12265 3519
rect 12265 3485 12299 3519
rect 12299 3485 12308 3519
rect 12256 3476 12308 3485
rect 12624 3476 12676 3528
rect 6920 3408 6972 3460
rect 7012 3408 7064 3460
rect 7380 3408 7432 3460
rect 9404 3408 9456 3460
rect 9864 3408 9916 3460
rect 10876 3451 10928 3460
rect 10876 3417 10885 3451
rect 10885 3417 10919 3451
rect 10919 3417 10928 3451
rect 16120 3476 16172 3528
rect 20812 3476 20864 3528
rect 23756 3519 23808 3528
rect 10876 3408 10928 3417
rect 19064 3408 19116 3460
rect 22468 3408 22520 3460
rect 23756 3485 23765 3519
rect 23765 3485 23799 3519
rect 23799 3485 23808 3519
rect 23756 3476 23808 3485
rect 23848 3476 23900 3528
rect 4896 3340 4948 3392
rect 7564 3383 7616 3392
rect 7564 3349 7573 3383
rect 7573 3349 7607 3383
rect 7607 3349 7616 3383
rect 7564 3340 7616 3349
rect 12532 3340 12584 3392
rect 14280 3383 14332 3392
rect 14280 3349 14289 3383
rect 14289 3349 14323 3383
rect 14323 3349 14332 3383
rect 14280 3340 14332 3349
rect 14648 3383 14700 3392
rect 14648 3349 14657 3383
rect 14657 3349 14691 3383
rect 14691 3349 14700 3383
rect 14648 3340 14700 3349
rect 15660 3340 15712 3392
rect 17684 3383 17736 3392
rect 17684 3349 17693 3383
rect 17693 3349 17727 3383
rect 17727 3349 17736 3383
rect 17684 3340 17736 3349
rect 19340 3340 19392 3392
rect 21272 3383 21324 3392
rect 21272 3349 21281 3383
rect 21281 3349 21315 3383
rect 21315 3349 21324 3383
rect 21272 3340 21324 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 3332 3136 3384 3188
rect 3976 3179 4028 3188
rect 3976 3145 3985 3179
rect 3985 3145 4019 3179
rect 4019 3145 4028 3179
rect 3976 3136 4028 3145
rect 4988 3136 5040 3188
rect 8024 3136 8076 3188
rect 9128 3179 9180 3188
rect 9128 3145 9137 3179
rect 9137 3145 9171 3179
rect 9171 3145 9180 3179
rect 9128 3136 9180 3145
rect 9312 3136 9364 3188
rect 10784 3136 10836 3188
rect 14096 3179 14148 3188
rect 14096 3145 14105 3179
rect 14105 3145 14139 3179
rect 14139 3145 14148 3179
rect 14096 3136 14148 3145
rect 15384 3179 15436 3188
rect 15384 3145 15393 3179
rect 15393 3145 15427 3179
rect 15427 3145 15436 3179
rect 15384 3136 15436 3145
rect 17132 3179 17184 3188
rect 17132 3145 17141 3179
rect 17141 3145 17175 3179
rect 17175 3145 17184 3179
rect 17132 3136 17184 3145
rect 5724 3068 5776 3120
rect 7196 3068 7248 3120
rect 7380 3111 7432 3120
rect 7380 3077 7389 3111
rect 7389 3077 7423 3111
rect 7423 3077 7432 3111
rect 7380 3068 7432 3077
rect 11152 3068 11204 3120
rect 14004 3068 14056 3120
rect 15200 3068 15252 3120
rect 9772 3000 9824 3052
rect 10876 3043 10928 3052
rect 10876 3009 10885 3043
rect 10885 3009 10919 3043
rect 10919 3009 10928 3043
rect 10876 3000 10928 3009
rect 11704 3000 11756 3052
rect 12072 3000 12124 3052
rect 12716 3000 12768 3052
rect 14648 3000 14700 3052
rect 15660 3000 15712 3052
rect 16120 3000 16172 3052
rect 4896 2932 4948 2984
rect 3056 2907 3108 2916
rect 3056 2873 3065 2907
rect 3065 2873 3099 2907
rect 3099 2873 3108 2907
rect 3056 2864 3108 2873
rect 2228 2796 2280 2848
rect 2596 2839 2648 2848
rect 2596 2805 2605 2839
rect 2605 2805 2639 2839
rect 2639 2805 2648 2839
rect 2596 2796 2648 2805
rect 3148 2839 3200 2848
rect 3148 2805 3157 2839
rect 3157 2805 3191 2839
rect 3191 2805 3200 2839
rect 3148 2796 3200 2805
rect 5632 2839 5684 2848
rect 5632 2805 5641 2839
rect 5641 2805 5675 2839
rect 5675 2805 5684 2839
rect 5632 2796 5684 2805
rect 7564 2975 7616 2984
rect 7564 2941 7573 2975
rect 7573 2941 7607 2975
rect 7607 2941 7616 2975
rect 7564 2932 7616 2941
rect 8300 2932 8352 2984
rect 8760 2932 8812 2984
rect 9864 2932 9916 2984
rect 19248 3136 19300 3188
rect 20812 3179 20864 3188
rect 20812 3145 20821 3179
rect 20821 3145 20855 3179
rect 20855 3145 20864 3179
rect 20812 3136 20864 3145
rect 23756 3136 23808 3188
rect 25136 3136 25188 3188
rect 19524 3068 19576 3120
rect 18788 3000 18840 3052
rect 22008 3000 22060 3052
rect 7564 2796 7616 2848
rect 7748 2839 7800 2848
rect 7748 2805 7757 2839
rect 7757 2805 7791 2839
rect 7791 2805 7800 2839
rect 7748 2796 7800 2805
rect 8392 2796 8444 2848
rect 9496 2864 9548 2916
rect 9956 2864 10008 2916
rect 10876 2864 10928 2916
rect 12532 2864 12584 2916
rect 19248 2975 19300 2984
rect 19248 2941 19257 2975
rect 19257 2941 19291 2975
rect 19291 2941 19300 2975
rect 19248 2932 19300 2941
rect 21272 2975 21324 2984
rect 21272 2941 21281 2975
rect 21281 2941 21315 2975
rect 21315 2941 21324 2975
rect 21272 2932 21324 2941
rect 22468 3000 22520 3052
rect 16120 2907 16172 2916
rect 9680 2796 9732 2848
rect 13636 2839 13688 2848
rect 13636 2805 13645 2839
rect 13645 2805 13679 2839
rect 13679 2805 13688 2839
rect 13636 2796 13688 2805
rect 14004 2796 14056 2848
rect 15292 2796 15344 2848
rect 16120 2873 16129 2907
rect 16129 2873 16163 2907
rect 16163 2873 16172 2907
rect 16120 2864 16172 2873
rect 18604 2796 18656 2848
rect 22100 2864 22152 2916
rect 23848 3000 23900 3052
rect 24216 3043 24268 3052
rect 24216 3009 24225 3043
rect 24225 3009 24259 3043
rect 24259 3009 24268 3043
rect 24216 3000 24268 3009
rect 19984 2796 20036 2848
rect 25780 2839 25832 2848
rect 25780 2805 25789 2839
rect 25789 2805 25823 2839
rect 25823 2805 25832 2839
rect 25780 2796 25832 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 3056 2592 3108 2644
rect 4896 2592 4948 2644
rect 5080 2592 5132 2644
rect 5356 2635 5408 2644
rect 5356 2601 5365 2635
rect 5365 2601 5399 2635
rect 5399 2601 5408 2635
rect 5356 2592 5408 2601
rect 6368 2635 6420 2644
rect 6368 2601 6377 2635
rect 6377 2601 6411 2635
rect 6411 2601 6420 2635
rect 6368 2592 6420 2601
rect 5724 2567 5776 2576
rect 5724 2533 5733 2567
rect 5733 2533 5767 2567
rect 5767 2533 5776 2567
rect 5724 2524 5776 2533
rect 2504 2456 2556 2508
rect 3516 2456 3568 2508
rect 5632 2456 5684 2508
rect 7748 2592 7800 2644
rect 9128 2635 9180 2644
rect 9128 2601 9137 2635
rect 9137 2601 9171 2635
rect 9171 2601 9180 2635
rect 9128 2592 9180 2601
rect 12256 2635 12308 2644
rect 9496 2524 9548 2576
rect 11152 2567 11204 2576
rect 11152 2533 11161 2567
rect 11161 2533 11195 2567
rect 11195 2533 11204 2567
rect 11152 2524 11204 2533
rect 11704 2567 11756 2576
rect 11704 2533 11713 2567
rect 11713 2533 11747 2567
rect 11747 2533 11756 2567
rect 11704 2524 11756 2533
rect 12256 2601 12265 2635
rect 12265 2601 12299 2635
rect 12299 2601 12308 2635
rect 12256 2592 12308 2601
rect 16028 2592 16080 2644
rect 16856 2635 16908 2644
rect 16856 2601 16865 2635
rect 16865 2601 16899 2635
rect 16899 2601 16908 2635
rect 16856 2592 16908 2601
rect 18972 2635 19024 2644
rect 18972 2601 18981 2635
rect 18981 2601 19015 2635
rect 19015 2601 19024 2635
rect 18972 2592 19024 2601
rect 21640 2592 21692 2644
rect 14004 2567 14056 2576
rect 14004 2533 14013 2567
rect 14013 2533 14047 2567
rect 14047 2533 14056 2567
rect 14004 2524 14056 2533
rect 14556 2567 14608 2576
rect 14556 2533 14565 2567
rect 14565 2533 14599 2567
rect 14599 2533 14608 2567
rect 14556 2524 14608 2533
rect 15200 2567 15252 2576
rect 15200 2533 15209 2567
rect 15209 2533 15243 2567
rect 15243 2533 15252 2567
rect 15200 2524 15252 2533
rect 16120 2524 16172 2576
rect 16764 2524 16816 2576
rect 19984 2524 20036 2576
rect 8760 2499 8812 2508
rect 8760 2465 8769 2499
rect 8769 2465 8803 2499
rect 8803 2465 8812 2499
rect 8760 2456 8812 2465
rect 10876 2499 10928 2508
rect 4712 2388 4764 2440
rect 10876 2465 10885 2499
rect 10885 2465 10919 2499
rect 10919 2465 10928 2499
rect 10876 2456 10928 2465
rect 12716 2499 12768 2508
rect 12716 2465 12725 2499
rect 12725 2465 12759 2499
rect 12759 2465 12768 2499
rect 12716 2456 12768 2465
rect 18420 2499 18472 2508
rect 18420 2465 18429 2499
rect 18429 2465 18463 2499
rect 18463 2465 18472 2499
rect 18420 2456 18472 2465
rect 24216 2592 24268 2644
rect 22008 2567 22060 2576
rect 22008 2533 22017 2567
rect 22017 2533 22051 2567
rect 22051 2533 22060 2567
rect 22008 2524 22060 2533
rect 22284 2567 22336 2576
rect 22284 2533 22293 2567
rect 22293 2533 22327 2567
rect 22327 2533 22336 2567
rect 22284 2524 22336 2533
rect 22468 2524 22520 2576
rect 22928 2567 22980 2576
rect 22928 2533 22937 2567
rect 22937 2533 22971 2567
rect 22971 2533 22980 2567
rect 22928 2524 22980 2533
rect 23664 2567 23716 2576
rect 23664 2533 23673 2567
rect 23673 2533 23707 2567
rect 23707 2533 23716 2567
rect 23664 2524 23716 2533
rect 24032 2524 24084 2576
rect 11796 2388 11848 2440
rect 8852 2320 8904 2372
rect 15936 2388 15988 2440
rect 19432 2388 19484 2440
rect 22284 2388 22336 2440
rect 16856 2320 16908 2372
rect 20168 2363 20220 2372
rect 2504 2295 2556 2304
rect 2504 2261 2513 2295
rect 2513 2261 2547 2295
rect 2547 2261 2556 2295
rect 2504 2252 2556 2261
rect 3332 2252 3384 2304
rect 3516 2295 3568 2304
rect 3516 2261 3525 2295
rect 3525 2261 3559 2295
rect 3559 2261 3568 2295
rect 3516 2252 3568 2261
rect 12900 2295 12952 2304
rect 12900 2261 12909 2295
rect 12909 2261 12943 2295
rect 12943 2261 12952 2295
rect 12900 2252 12952 2261
rect 20168 2329 20177 2363
rect 20177 2329 20211 2363
rect 20211 2329 20220 2363
rect 20168 2320 20220 2329
rect 23020 2320 23072 2372
rect 20260 2252 20312 2304
rect 22652 2252 22704 2304
rect 24308 2320 24360 2372
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 4436 76 4488 128
rect 4988 76 5040 128
rect 9588 76 9640 128
rect 10416 76 10468 128
rect 12900 76 12952 128
rect 15108 76 15160 128
rect 26148 76 26200 128
rect 26792 76 26844 128
rect 14280 8 14332 60
rect 18236 8 18288 60
rect 26240 8 26292 60
rect 27528 8 27580 60
<< metal2 >>
rect 754 27520 810 28000
rect 2226 27532 2282 28000
rect 2226 27520 2228 27532
rect 768 26790 796 27520
rect 2280 27520 2282 27532
rect 3424 27532 3476 27538
rect 2228 27474 2280 27480
rect 3790 27520 3846 28000
rect 5092 27526 5304 27554
rect 3424 27474 3476 27480
rect 2240 27443 2268 27474
rect 756 26784 808 26790
rect 756 26726 808 26732
rect 2780 26784 2832 26790
rect 2780 26726 2832 26732
rect 1858 25664 1914 25673
rect 1858 25599 1914 25608
rect 1872 23662 1900 25599
rect 1860 23656 1912 23662
rect 1860 23598 1912 23604
rect 1582 18592 1638 18601
rect 1582 18527 1638 18536
rect 110 12200 166 12209
rect 110 12135 166 12144
rect 124 10130 152 12135
rect 1596 11218 1624 18527
rect 2044 18216 2096 18222
rect 2044 18158 2096 18164
rect 1858 15192 1914 15201
rect 1858 15127 1914 15136
rect 1872 13870 1900 15127
rect 1860 13864 1912 13870
rect 1860 13806 1912 13812
rect 1584 11212 1636 11218
rect 1584 11154 1636 11160
rect 1596 10810 1624 11154
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 112 10124 164 10130
rect 112 10066 164 10072
rect 110 8664 166 8673
rect 110 8599 166 8608
rect 124 8430 152 8599
rect 112 8424 164 8430
rect 112 8366 164 8372
rect 1674 8392 1730 8401
rect 1674 8327 1730 8336
rect 1400 7540 1452 7546
rect 1400 7482 1452 7488
rect 664 6996 716 7002
rect 664 6938 716 6944
rect 204 5160 256 5166
rect 110 5128 166 5137
rect 166 5108 204 5114
rect 166 5102 256 5108
rect 166 5086 244 5102
rect 110 5063 166 5072
rect 386 82 442 480
rect 676 82 704 6938
rect 386 54 704 82
rect 1122 82 1178 480
rect 1412 82 1440 7482
rect 1688 5370 1716 8327
rect 1676 5364 1728 5370
rect 1676 5306 1728 5312
rect 1122 54 1440 82
rect 1858 82 1914 480
rect 2056 82 2084 18158
rect 2792 17785 2820 26726
rect 3436 18766 3464 27474
rect 3804 21593 3832 27520
rect 4894 22128 4950 22137
rect 4894 22063 4950 22072
rect 3790 21584 3846 21593
rect 3790 21519 3846 21528
rect 4908 21010 4936 22063
rect 4896 21004 4948 21010
rect 4896 20946 4948 20952
rect 4712 20800 4764 20806
rect 4712 20742 4764 20748
rect 4436 20392 4488 20398
rect 4436 20334 4488 20340
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 4252 18760 4304 18766
rect 4252 18702 4304 18708
rect 4264 18358 4292 18702
rect 4252 18352 4304 18358
rect 4252 18294 4304 18300
rect 2778 17776 2834 17785
rect 2778 17711 2834 17720
rect 3054 17776 3110 17785
rect 3054 17711 3110 17720
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 2884 4146 2912 4626
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 2964 3596 3016 3602
rect 3068 3584 3096 17711
rect 3884 14340 3936 14346
rect 3884 14282 3936 14288
rect 3606 13560 3662 13569
rect 3606 13495 3662 13504
rect 3240 5840 3292 5846
rect 3240 5782 3292 5788
rect 3252 5370 3280 5782
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3148 5296 3200 5302
rect 3148 5238 3200 5244
rect 3016 3556 3096 3584
rect 2964 3538 3016 3544
rect 2240 2854 2268 3538
rect 3068 2922 3096 3556
rect 3160 3534 3188 5238
rect 3620 4282 3648 13495
rect 3700 8832 3752 8838
rect 3700 8774 3752 8780
rect 3608 4276 3660 4282
rect 3608 4218 3660 4224
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3148 3528 3200 3534
rect 3148 3470 3200 3476
rect 3344 3194 3372 4082
rect 3620 4078 3648 4218
rect 3712 4146 3740 8774
rect 3792 7472 3844 7478
rect 3792 7414 3844 7420
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 3608 4072 3660 4078
rect 3804 4026 3832 7414
rect 3896 5370 3924 14282
rect 4160 13796 4212 13802
rect 4160 13738 4212 13744
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 4080 9178 4108 9862
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4172 7546 4200 13738
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 3988 4154 4016 6054
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 4080 4282 4108 4626
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 3608 4014 3660 4020
rect 3712 3998 3832 4026
rect 3896 4126 4016 4154
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3056 2916 3108 2922
rect 3056 2858 3108 2864
rect 2228 2848 2280 2854
rect 2228 2790 2280 2796
rect 2596 2848 2648 2854
rect 3068 2825 3096 2858
rect 3148 2848 3200 2854
rect 2596 2790 2648 2796
rect 3054 2816 3110 2825
rect 2240 2009 2268 2790
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 2516 2310 2544 2450
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 2226 2000 2282 2009
rect 2226 1935 2282 1944
rect 2516 1057 2544 2246
rect 2502 1048 2558 1057
rect 2502 983 2558 992
rect 1858 54 2084 82
rect 2608 82 2636 2790
rect 3148 2790 3200 2796
rect 3054 2751 3110 2760
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 3068 2417 3096 2586
rect 3160 2553 3188 2790
rect 3146 2544 3202 2553
rect 3146 2479 3202 2488
rect 3516 2508 3568 2514
rect 3516 2450 3568 2456
rect 3054 2408 3110 2417
rect 3054 2343 3110 2352
rect 3528 2310 3556 2450
rect 3332 2304 3384 2310
rect 3332 2246 3384 2252
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 3344 1601 3372 2246
rect 3528 1737 3556 2246
rect 3514 1728 3570 1737
rect 3514 1663 3570 1672
rect 3330 1592 3386 1601
rect 3330 1527 3386 1536
rect 2686 82 2742 480
rect 2608 54 2742 82
rect 386 0 442 54
rect 1122 0 1178 54
rect 1858 0 1914 54
rect 2686 0 2742 54
rect 3422 82 3478 480
rect 3712 82 3740 3998
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3804 3097 3832 3878
rect 3790 3088 3846 3097
rect 3790 3023 3846 3032
rect 3896 2281 3924 4126
rect 4264 4078 4292 18294
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4356 4826 4384 11494
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 4344 4548 4396 4554
rect 4344 4490 4396 4496
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3988 3194 4016 3470
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 3882 2272 3938 2281
rect 3882 2207 3938 2216
rect 3422 54 3740 82
rect 4250 82 4306 480
rect 4356 82 4384 4490
rect 4448 134 4476 20334
rect 4724 9110 4752 20742
rect 4908 20602 4936 20946
rect 4896 20596 4948 20602
rect 4896 20538 4948 20544
rect 5092 17746 5120 27526
rect 5276 27418 5304 27526
rect 5354 27520 5410 28000
rect 6918 27520 6974 28000
rect 8482 27520 8538 28000
rect 10046 27568 10102 28000
rect 5368 27418 5396 27520
rect 5276 27390 5396 27418
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5080 17740 5132 17746
rect 5080 17682 5132 17688
rect 5092 17338 5120 17682
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6736 17264 6788 17270
rect 6656 17224 6736 17252
rect 6656 16658 6684 17224
rect 6736 17206 6788 17212
rect 6644 16652 6696 16658
rect 6644 16594 6696 16600
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6656 16250 6684 16594
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 6840 16114 6868 17274
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 6092 16040 6144 16046
rect 6092 15982 6144 15988
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5170 13288 5226 13297
rect 5170 13223 5226 13232
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4816 9722 4844 10066
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 5184 7954 5212 13223
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5816 12776 5868 12782
rect 5816 12718 5868 12724
rect 5828 12374 5856 12718
rect 5816 12368 5868 12374
rect 5816 12310 5868 12316
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5552 11558 5580 12174
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 6104 10962 6132 15982
rect 6644 15564 6696 15570
rect 6644 15506 6696 15512
rect 6656 15162 6684 15506
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 6552 14476 6604 14482
rect 6604 14436 6684 14464
rect 6552 14418 6604 14424
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6196 12753 6224 13670
rect 6182 12744 6238 12753
rect 6182 12679 6238 12688
rect 6184 12368 6236 12374
rect 6184 12310 6236 12316
rect 6196 11354 6224 12310
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 6012 10713 6040 10950
rect 6104 10934 6224 10962
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 5998 10704 6054 10713
rect 5998 10639 6054 10648
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5552 9450 5580 10066
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5276 8498 5304 9114
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5368 8090 5396 8298
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5184 7546 5212 7890
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 4710 7440 4766 7449
rect 4710 7375 4766 7384
rect 4724 6866 4752 7375
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4724 6458 4752 6802
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 5080 6724 5132 6730
rect 5080 6666 5132 6672
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4540 5846 4568 6054
rect 4528 5840 4580 5846
rect 4528 5782 4580 5788
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 4632 4826 4660 5714
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4724 5166 4752 5646
rect 4712 5160 4764 5166
rect 4816 5137 4844 6666
rect 5092 6458 5120 6666
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 4712 5102 4764 5108
rect 4802 5128 4858 5137
rect 4802 5063 4858 5072
rect 4908 5030 4936 6190
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 4988 5636 5040 5642
rect 4988 5578 5040 5584
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 5000 4826 5028 5578
rect 5092 5302 5120 6054
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 5184 5370 5212 5714
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 5080 5296 5132 5302
rect 5080 5238 5132 5244
rect 5262 5264 5318 5273
rect 5262 5199 5318 5208
rect 5276 5166 5304 5199
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4986 4720 5042 4729
rect 4896 4684 4948 4690
rect 4986 4655 5042 4664
rect 4896 4626 4948 4632
rect 4908 4593 4936 4626
rect 4894 4584 4950 4593
rect 4894 4519 4950 4528
rect 5000 4078 5028 4655
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4988 4072 5040 4078
rect 4988 4014 5040 4020
rect 4724 3942 4752 4014
rect 5000 3942 5028 4014
rect 4528 3936 4580 3942
rect 4528 3878 4580 3884
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 4540 1465 4568 3878
rect 4724 2446 4752 3878
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4908 2990 4936 3334
rect 5000 3194 5028 3878
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 4896 2984 4948 2990
rect 4896 2926 4948 2932
rect 4908 2650 4936 2926
rect 5092 2650 5120 4082
rect 5264 3596 5316 3602
rect 5368 3584 5396 7482
rect 5460 6934 5488 8230
rect 5552 7546 5580 9386
rect 6000 9376 6052 9382
rect 6104 9364 6132 10746
rect 6052 9336 6132 9364
rect 6000 9318 6052 9324
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5552 7002 5580 7278
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5448 6928 5500 6934
rect 5448 6870 5500 6876
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5552 6254 5580 6802
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6012 6390 6040 9318
rect 6196 9194 6224 10934
rect 6104 9166 6224 9194
rect 6104 7290 6132 9166
rect 6184 9104 6236 9110
rect 6184 9046 6236 9052
rect 6276 9104 6328 9110
rect 6276 9046 6328 9052
rect 6196 8634 6224 9046
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6288 8362 6316 9046
rect 6276 8356 6328 8362
rect 6276 8298 6328 8304
rect 6184 8016 6236 8022
rect 6288 8004 6316 8298
rect 6236 7976 6316 8004
rect 6184 7958 6236 7964
rect 6104 7262 6224 7290
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 6104 6934 6132 7142
rect 6092 6928 6144 6934
rect 6092 6870 6144 6876
rect 6000 6384 6052 6390
rect 6000 6326 6052 6332
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5448 4684 5500 4690
rect 5448 4626 5500 4632
rect 5460 4154 5488 4626
rect 5552 4282 5580 5510
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6196 5273 6224 7262
rect 6288 7002 6316 7976
rect 6276 6996 6328 7002
rect 6276 6938 6328 6944
rect 6380 6322 6408 14350
rect 6552 14272 6604 14278
rect 6552 14214 6604 14220
rect 6564 13462 6592 14214
rect 6656 13802 6684 14436
rect 6644 13796 6696 13802
rect 6644 13738 6696 13744
rect 6932 13569 6960 27520
rect 7104 23588 7156 23594
rect 7104 23530 7156 23536
rect 7116 22166 7144 23530
rect 7104 22160 7156 22166
rect 7104 22102 7156 22108
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 7484 18193 7512 18226
rect 7470 18184 7526 18193
rect 7470 18119 7526 18128
rect 8300 18148 8352 18154
rect 8300 18090 8352 18096
rect 7196 18080 7248 18086
rect 7196 18022 7248 18028
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7208 17882 7236 18022
rect 7196 17876 7248 17882
rect 7196 17818 7248 17824
rect 7208 17202 7236 17818
rect 7380 17808 7432 17814
rect 7380 17750 7432 17756
rect 7288 17672 7340 17678
rect 7288 17614 7340 17620
rect 7300 17338 7328 17614
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7288 16992 7340 16998
rect 7392 16980 7420 17750
rect 7340 16952 7420 16980
rect 7288 16934 7340 16940
rect 7300 16454 7328 16934
rect 7484 16726 7512 18022
rect 8312 17678 8340 18090
rect 7656 17672 7708 17678
rect 8300 17672 8352 17678
rect 7656 17614 7708 17620
rect 8114 17640 8170 17649
rect 7472 16720 7524 16726
rect 7472 16662 7524 16668
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 7300 15638 7328 16390
rect 7484 15978 7512 16526
rect 7472 15972 7524 15978
rect 7472 15914 7524 15920
rect 7484 15706 7512 15914
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7288 15632 7340 15638
rect 7288 15574 7340 15580
rect 7196 15564 7248 15570
rect 7196 15506 7248 15512
rect 7208 14890 7236 15506
rect 7668 15094 7696 17614
rect 8300 17614 8352 17620
rect 8114 17575 8170 17584
rect 8128 17542 8156 17575
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 8312 16726 8340 17138
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 7748 16720 7800 16726
rect 7748 16662 7800 16668
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 7760 16250 7788 16662
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 7760 15706 7788 16186
rect 8404 16046 8432 16934
rect 8496 16182 8524 27520
rect 11610 27520 11666 28000
rect 13174 27520 13230 28000
rect 14372 27532 14424 27538
rect 10046 27503 10102 27512
rect 10060 27443 10088 27503
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 9588 22092 9640 22098
rect 9588 22034 9640 22040
rect 8944 21480 8996 21486
rect 8944 21422 8996 21428
rect 8576 21412 8628 21418
rect 8576 21354 8628 21360
rect 8484 16176 8536 16182
rect 8484 16118 8536 16124
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 8208 15972 8260 15978
rect 8208 15914 8260 15920
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 8220 15638 8248 15914
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 8220 15162 8248 15574
rect 8484 15496 8536 15502
rect 8588 15484 8616 21354
rect 8956 18290 8984 21422
rect 9600 21418 9628 22034
rect 9588 21412 9640 21418
rect 9588 21354 9640 21360
rect 10048 21344 10100 21350
rect 10048 21286 10100 21292
rect 10060 20369 10088 21286
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 11624 21010 11652 27520
rect 12716 23656 12768 23662
rect 12716 23598 12768 23604
rect 11980 22160 12032 22166
rect 11980 22102 12032 22108
rect 11612 21004 11664 21010
rect 11612 20946 11664 20952
rect 10140 20936 10192 20942
rect 10140 20878 10192 20884
rect 10046 20360 10102 20369
rect 10046 20295 10102 20304
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9692 18426 9720 18770
rect 9968 18766 9996 20198
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 10060 18426 10088 19654
rect 10152 19514 10180 20878
rect 10692 20800 10744 20806
rect 10692 20742 10744 20748
rect 10230 20496 10286 20505
rect 10704 20466 10732 20742
rect 11624 20602 11652 20946
rect 11612 20596 11664 20602
rect 11612 20538 11664 20544
rect 10230 20431 10286 20440
rect 10692 20460 10744 20466
rect 10244 20398 10272 20431
rect 10692 20402 10744 20408
rect 10232 20392 10284 20398
rect 10232 20334 10284 20340
rect 11704 20324 11756 20330
rect 11704 20266 11756 20272
rect 10692 20256 10744 20262
rect 10692 20198 10744 20204
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10232 19984 10284 19990
rect 10232 19926 10284 19932
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 10244 19310 10272 19926
rect 10704 19378 10732 20198
rect 11716 19854 11744 20266
rect 11888 19984 11940 19990
rect 11888 19926 11940 19932
rect 11704 19848 11756 19854
rect 11704 19790 11756 19796
rect 11716 19514 11744 19790
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10232 19304 10284 19310
rect 10152 19264 10232 19292
rect 10152 18426 10180 19264
rect 10232 19246 10284 19252
rect 11612 19236 11664 19242
rect 11612 19178 11664 19184
rect 11336 19168 11388 19174
rect 11336 19110 11388 19116
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10876 18760 10928 18766
rect 10876 18702 10928 18708
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 10048 18420 10100 18426
rect 10048 18362 10100 18368
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 10888 18290 10916 18702
rect 8944 18284 8996 18290
rect 10876 18284 10928 18290
rect 8996 18244 9076 18272
rect 8944 18226 8996 18232
rect 8944 17536 8996 17542
rect 8944 17478 8996 17484
rect 8956 17202 8984 17478
rect 9048 17202 9076 18244
rect 10876 18226 10928 18232
rect 11348 18154 11376 19110
rect 11624 18902 11652 19178
rect 11900 19174 11928 19926
rect 11888 19168 11940 19174
rect 11888 19110 11940 19116
rect 11612 18896 11664 18902
rect 11612 18838 11664 18844
rect 11796 18896 11848 18902
rect 11796 18838 11848 18844
rect 11624 18290 11652 18838
rect 11808 18426 11836 18838
rect 11900 18766 11928 19110
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 11796 18420 11848 18426
rect 11796 18362 11848 18368
rect 11612 18284 11664 18290
rect 11612 18226 11664 18232
rect 11336 18148 11388 18154
rect 11336 18090 11388 18096
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 11348 17882 11376 18090
rect 11336 17876 11388 17882
rect 11336 17818 11388 17824
rect 9772 17808 9824 17814
rect 9772 17750 9824 17756
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 9036 17196 9088 17202
rect 9036 17138 9088 17144
rect 9220 17060 9272 17066
rect 9220 17002 9272 17008
rect 8668 16448 8720 16454
rect 8668 16390 8720 16396
rect 8680 15586 8708 16390
rect 9232 16250 9260 17002
rect 9784 16998 9812 17750
rect 11428 17672 11480 17678
rect 11428 17614 11480 17620
rect 11152 17060 11204 17066
rect 11152 17002 11204 17008
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 8760 16040 8812 16046
rect 8760 15982 8812 15988
rect 8772 15706 8800 15982
rect 9784 15978 9812 16934
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10140 16652 10192 16658
rect 10140 16594 10192 16600
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 10152 16046 10180 16594
rect 10140 16040 10192 16046
rect 10140 15982 10192 15988
rect 9772 15972 9824 15978
rect 9772 15914 9824 15920
rect 9128 15904 9180 15910
rect 9128 15846 9180 15852
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8680 15558 8800 15586
rect 8588 15456 8708 15484
rect 8484 15438 8536 15444
rect 8024 15156 8076 15162
rect 8024 15098 8076 15104
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 7656 15088 7708 15094
rect 7656 15030 7708 15036
rect 7104 14884 7156 14890
rect 7104 14826 7156 14832
rect 7196 14884 7248 14890
rect 7196 14826 7248 14832
rect 7116 14346 7144 14826
rect 7104 14340 7156 14346
rect 7104 14282 7156 14288
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7852 13938 7880 14214
rect 7840 13932 7892 13938
rect 7840 13874 7892 13880
rect 6918 13560 6974 13569
rect 6918 13495 6974 13504
rect 6552 13456 6604 13462
rect 6552 13398 6604 13404
rect 6644 13456 6696 13462
rect 6644 13398 6696 13404
rect 7656 13456 7708 13462
rect 7656 13398 7708 13404
rect 6656 12714 6684 13398
rect 7668 12986 7696 13398
rect 7932 13184 7984 13190
rect 7932 13126 7984 13132
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 7944 12782 7972 13126
rect 8036 12986 8064 15098
rect 8496 14890 8524 15438
rect 8484 14884 8536 14890
rect 8484 14826 8536 14832
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8220 13326 8248 13874
rect 8576 13796 8628 13802
rect 8576 13738 8628 13744
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 7932 12776 7984 12782
rect 7932 12718 7984 12724
rect 8036 12714 8064 12922
rect 6644 12708 6696 12714
rect 6644 12650 6696 12656
rect 8024 12708 8076 12714
rect 8024 12650 8076 12656
rect 6460 12164 6512 12170
rect 6460 12106 6512 12112
rect 6472 11898 6500 12106
rect 6656 11898 6684 12650
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6840 12442 6868 12582
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6656 11626 6684 11834
rect 6840 11830 6868 12378
rect 7576 12306 7604 12378
rect 8036 12374 8064 12650
rect 8128 12442 8156 13262
rect 8116 12436 8168 12442
rect 8116 12378 8168 12384
rect 8024 12368 8076 12374
rect 8024 12310 8076 12316
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 6828 11824 6880 11830
rect 6828 11766 6880 11772
rect 7576 11762 7604 12242
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6644 11620 6696 11626
rect 6644 11562 6696 11568
rect 6748 11082 6776 11630
rect 7196 11620 7248 11626
rect 7196 11562 7248 11568
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 6736 11076 6788 11082
rect 6736 11018 6788 11024
rect 6826 10568 6882 10577
rect 6826 10503 6882 10512
rect 6458 10160 6514 10169
rect 6458 10095 6514 10104
rect 6552 10124 6604 10130
rect 6472 10062 6500 10095
rect 6552 10066 6604 10072
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6564 9761 6592 10066
rect 6734 9888 6790 9897
rect 6734 9823 6790 9832
rect 6550 9752 6606 9761
rect 6550 9687 6552 9696
rect 6604 9687 6606 9696
rect 6552 9658 6604 9664
rect 6564 9627 6592 9658
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6472 8498 6500 8910
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6472 6322 6500 8434
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6564 7546 6592 7822
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6656 7410 6684 7686
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6748 7342 6776 9823
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6380 5778 6408 6258
rect 6460 6180 6512 6186
rect 6460 6122 6512 6128
rect 6472 5778 6500 6122
rect 6368 5772 6420 5778
rect 6368 5714 6420 5720
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6182 5264 6238 5273
rect 6182 5199 6238 5208
rect 6184 5092 6236 5098
rect 6184 5034 6236 5040
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5460 4126 5764 4154
rect 5736 4078 5764 4126
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 5316 3556 5396 3584
rect 5264 3538 5316 3544
rect 5368 2650 5396 3556
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 4526 1456 4582 1465
rect 4526 1391 4582 1400
rect 4250 54 4384 82
rect 4436 128 4488 134
rect 4436 70 4488 76
rect 4986 128 5042 480
rect 4986 76 4988 128
rect 5040 76 5042 128
rect 3422 0 3478 54
rect 4250 0 4306 54
rect 4986 0 5042 76
rect 5552 82 5580 3946
rect 5736 3738 5764 4014
rect 6000 4004 6052 4010
rect 6000 3946 6052 3952
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5736 3602 5764 3674
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5724 3120 5776 3126
rect 5724 3062 5776 3068
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5644 2514 5672 2790
rect 5736 2582 5764 3062
rect 5724 2576 5776 2582
rect 5724 2518 5776 2524
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6012 1329 6040 3946
rect 5998 1320 6054 1329
rect 5998 1255 6054 1264
rect 5814 82 5870 480
rect 5552 54 5870 82
rect 6196 82 6224 5034
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6380 3777 6408 4966
rect 6472 4758 6500 5714
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6552 5636 6604 5642
rect 6552 5578 6604 5584
rect 6564 5098 6592 5578
rect 6656 5302 6684 5646
rect 6644 5296 6696 5302
rect 6644 5238 6696 5244
rect 6552 5092 6604 5098
rect 6552 5034 6604 5040
rect 6460 4752 6512 4758
rect 6460 4694 6512 4700
rect 6840 4554 6868 10503
rect 7116 10470 7144 11154
rect 7208 10674 7236 11562
rect 7760 11354 7788 12242
rect 8036 11898 8064 12310
rect 8588 12306 8616 13738
rect 8680 13258 8708 15456
rect 8772 13394 8800 15558
rect 9140 15162 9168 15846
rect 10152 15570 10180 15982
rect 10428 15978 10456 16594
rect 10796 16590 10824 16934
rect 10784 16584 10836 16590
rect 10784 16526 10836 16532
rect 10796 16046 10824 16526
rect 11164 16046 11192 17002
rect 11440 16998 11468 17614
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11440 16182 11468 16934
rect 11808 16726 11836 17478
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11900 16726 11928 16934
rect 11796 16720 11848 16726
rect 11796 16662 11848 16668
rect 11888 16720 11940 16726
rect 11888 16662 11940 16668
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11428 16176 11480 16182
rect 11428 16118 11480 16124
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 10416 15972 10468 15978
rect 10416 15914 10468 15920
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10140 15564 10192 15570
rect 10140 15506 10192 15512
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10784 15564 10836 15570
rect 10784 15506 10836 15512
rect 9496 15360 9548 15366
rect 9496 15302 9548 15308
rect 9128 15156 9180 15162
rect 9128 15098 9180 15104
rect 9404 14952 9456 14958
rect 9404 14894 9456 14900
rect 9416 14822 9444 14894
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9220 14544 9272 14550
rect 9220 14486 9272 14492
rect 8852 14476 8904 14482
rect 8852 14418 8904 14424
rect 8864 13734 8892 14418
rect 8852 13728 8904 13734
rect 8850 13696 8852 13705
rect 9036 13728 9088 13734
rect 8904 13696 8906 13705
rect 9036 13670 9088 13676
rect 8850 13631 8906 13640
rect 8864 13605 8892 13631
rect 8760 13388 8812 13394
rect 8760 13330 8812 13336
rect 8668 13252 8720 13258
rect 8668 13194 8720 13200
rect 9048 13190 9076 13670
rect 9036 13184 9088 13190
rect 9036 13126 9088 13132
rect 9048 12986 9076 13126
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 9232 12170 9260 14486
rect 9416 14006 9444 14758
rect 9508 14550 9536 15302
rect 10152 14958 10180 15506
rect 10704 14958 10732 15506
rect 10796 14958 10824 15506
rect 11164 14958 11192 15982
rect 11716 15978 11744 16390
rect 11704 15972 11756 15978
rect 11704 15914 11756 15920
rect 11716 15706 11744 15914
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 11152 14952 11204 14958
rect 11152 14894 11204 14900
rect 10152 14618 10180 14894
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 9496 14544 9548 14550
rect 9496 14486 9548 14492
rect 10140 14476 10192 14482
rect 10140 14418 10192 14424
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 9404 14000 9456 14006
rect 9404 13942 9456 13948
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 9324 13462 9352 13806
rect 9312 13456 9364 13462
rect 9312 13398 9364 13404
rect 9220 12164 9272 12170
rect 9220 12106 9272 12112
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 7024 9518 7052 9930
rect 7116 9897 7144 10406
rect 7300 10266 7328 11086
rect 7380 11008 7432 11014
rect 7380 10950 7432 10956
rect 7392 10606 7420 10950
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 8036 10538 8064 11834
rect 9416 11830 9444 13942
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 9508 13190 9536 13330
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9508 11830 9536 13126
rect 9600 12374 9628 14282
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9680 13864 9732 13870
rect 9680 13806 9732 13812
rect 9692 13734 9720 13806
rect 9772 13796 9824 13802
rect 9772 13738 9824 13744
rect 9680 13728 9732 13734
rect 9680 13670 9732 13676
rect 9692 13530 9720 13670
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9784 13161 9812 13738
rect 9968 13569 9996 13874
rect 10152 13802 10180 14418
rect 10704 14006 10732 14894
rect 10796 14414 10824 14894
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10968 14340 11020 14346
rect 10968 14282 11020 14288
rect 10692 14000 10744 14006
rect 10692 13942 10744 13948
rect 10140 13796 10192 13802
rect 10140 13738 10192 13744
rect 9954 13560 10010 13569
rect 9954 13495 10010 13504
rect 9956 13456 10008 13462
rect 9956 13398 10008 13404
rect 9968 13326 9996 13398
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 9770 13152 9826 13161
rect 9770 13087 9826 13096
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9588 12368 9640 12374
rect 9588 12310 9640 12316
rect 9784 12238 9812 12582
rect 10060 12306 10088 12718
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9784 12102 9812 12174
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9404 11824 9456 11830
rect 9404 11766 9456 11772
rect 9496 11824 9548 11830
rect 9496 11766 9548 11772
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8392 11280 8444 11286
rect 8444 11240 8524 11268
rect 8392 11222 8444 11228
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 8220 10674 8248 11086
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7564 10192 7616 10198
rect 7564 10134 7616 10140
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7196 9920 7248 9926
rect 7102 9888 7158 9897
rect 7196 9862 7248 9868
rect 7102 9823 7158 9832
rect 7208 9518 7236 9862
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7208 9178 7236 9454
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7484 8906 7512 9998
rect 7576 9586 7604 10134
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7472 8900 7524 8906
rect 7472 8842 7524 8848
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 7024 7274 7052 8026
rect 7012 7268 7064 7274
rect 7012 7210 7064 7216
rect 7012 6928 7064 6934
rect 7012 6870 7064 6876
rect 7024 6186 7052 6870
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 6932 5846 6960 6122
rect 7208 5846 7236 8366
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7300 7993 7328 8230
rect 7760 8090 7788 8434
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7286 7984 7342 7993
rect 7286 7919 7342 7928
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7392 7274 7420 7822
rect 7852 7721 7880 9318
rect 8036 8634 8064 10474
rect 8220 10198 8248 10610
rect 8496 10470 8524 11240
rect 8864 11014 8892 11698
rect 9220 11688 9272 11694
rect 9220 11630 9272 11636
rect 9232 11150 9260 11630
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 8852 11008 8904 11014
rect 8852 10950 8904 10956
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8496 9926 8524 10406
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8760 9580 8812 9586
rect 8680 9540 8760 9568
rect 8208 9104 8260 9110
rect 8208 9046 8260 9052
rect 8220 8634 8248 9046
rect 8680 8906 8708 9540
rect 8760 9522 8812 9528
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8668 8900 8720 8906
rect 8668 8842 8720 8848
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8036 8362 8064 8570
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 8036 8022 8064 8298
rect 8024 8016 8076 8022
rect 8024 7958 8076 7964
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 7838 7712 7894 7721
rect 7838 7647 7894 7656
rect 7380 7268 7432 7274
rect 7380 7210 7432 7216
rect 7392 6934 7420 7210
rect 7380 6928 7432 6934
rect 7380 6870 7432 6876
rect 7380 6384 7432 6390
rect 7380 6326 7432 6332
rect 7472 6384 7524 6390
rect 7472 6326 7524 6332
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 7196 5840 7248 5846
rect 7196 5782 7248 5788
rect 7392 5642 7420 6326
rect 7380 5636 7432 5642
rect 7380 5578 7432 5584
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6932 4690 6960 5170
rect 7484 5166 7512 6326
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7576 6186 7604 6258
rect 7564 6180 7616 6186
rect 7564 6122 7616 6128
rect 7576 5846 7604 6122
rect 7564 5840 7616 5846
rect 7564 5782 7616 5788
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7484 4826 7512 5102
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 6828 4548 6880 4554
rect 6828 4490 6880 4496
rect 7116 3942 7144 4626
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7196 4548 7248 4554
rect 7196 4490 7248 4496
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 6366 3768 6422 3777
rect 6366 3703 6422 3712
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 6288 1873 6316 3470
rect 6380 2650 6408 3470
rect 7024 3466 7052 3538
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 7012 3460 7064 3466
rect 7012 3402 7064 3408
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 6274 1864 6330 1873
rect 6274 1799 6330 1808
rect 6932 1193 6960 3402
rect 6918 1184 6974 1193
rect 6918 1119 6974 1128
rect 6550 82 6606 480
rect 6196 54 6606 82
rect 7116 82 7144 3878
rect 7208 3602 7236 4490
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7576 4146 7604 4218
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7668 4049 7696 4558
rect 7852 4154 7880 7647
rect 7944 6934 7972 7890
rect 8036 7546 8064 7958
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 8680 7410 8708 8842
rect 8772 7954 8800 9318
rect 8864 7993 8892 10950
rect 9140 10810 9168 10950
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 9312 10736 9364 10742
rect 9312 10678 9364 10684
rect 9324 10538 9352 10678
rect 9312 10532 9364 10538
rect 9312 10474 9364 10480
rect 9324 10266 9352 10474
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9416 9994 9444 11766
rect 9784 11286 9812 12038
rect 10060 11898 10088 12242
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 9956 11620 10008 11626
rect 9956 11562 10008 11568
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9772 11280 9824 11286
rect 9772 11222 9824 11228
rect 9784 11014 9812 11222
rect 9772 11008 9824 11014
rect 9772 10950 9824 10956
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9404 9988 9456 9994
rect 9404 9930 9456 9936
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 8944 8900 8996 8906
rect 8944 8842 8996 8848
rect 8956 8566 8984 8842
rect 8944 8560 8996 8566
rect 8944 8502 8996 8508
rect 9048 8090 9076 8910
rect 9324 8838 9352 9454
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 8850 7984 8906 7993
rect 8760 7948 8812 7954
rect 8850 7919 8906 7928
rect 8760 7890 8812 7896
rect 9324 7750 9352 8774
rect 9416 8294 9444 8978
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8772 7274 8800 7686
rect 9324 7342 9352 7686
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 8484 7268 8536 7274
rect 8484 7210 8536 7216
rect 8760 7268 8812 7274
rect 8760 7210 8812 7216
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8128 6934 8156 7142
rect 8496 7002 8524 7210
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 7932 6928 7984 6934
rect 7932 6870 7984 6876
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 8390 6896 8446 6905
rect 8390 6831 8446 6840
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8312 6458 8340 6734
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 7944 5846 7972 6394
rect 7932 5840 7984 5846
rect 7932 5782 7984 5788
rect 8404 5778 8432 6831
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8680 5914 8708 6054
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8024 5772 8076 5778
rect 8024 5714 8076 5720
rect 8392 5772 8444 5778
rect 8392 5714 8444 5720
rect 7932 5636 7984 5642
rect 7932 5578 7984 5584
rect 7944 4826 7972 5578
rect 8036 5302 8064 5714
rect 8864 5302 8892 7142
rect 9324 6730 9352 7278
rect 9312 6724 9364 6730
rect 9312 6666 9364 6672
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9232 6390 9260 6598
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 9036 6112 9088 6118
rect 9036 6054 9088 6060
rect 9048 5710 9076 6054
rect 9416 5914 9444 8230
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 8024 5296 8076 5302
rect 8024 5238 8076 5244
rect 8852 5296 8904 5302
rect 8852 5238 8904 5244
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 7852 4126 7972 4154
rect 8496 4146 8524 4626
rect 8668 4616 8720 4622
rect 8668 4558 8720 4564
rect 7944 4078 7972 4126
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8680 4078 8708 4558
rect 7932 4072 7984 4078
rect 7654 4040 7710 4049
rect 7932 4014 7984 4020
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 7654 3975 7710 3984
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8312 3602 8340 3878
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 7208 3126 7236 3538
rect 7380 3460 7432 3466
rect 7380 3402 7432 3408
rect 7392 3126 7420 3402
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7196 3120 7248 3126
rect 7196 3062 7248 3068
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 7576 2990 7604 3334
rect 8036 3194 8064 3538
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8312 2990 8340 3538
rect 8680 3505 8708 3606
rect 8666 3496 8722 3505
rect 8666 3431 8722 3440
rect 7564 2984 7616 2990
rect 7564 2926 7616 2932
rect 8300 2984 8352 2990
rect 8300 2926 8352 2932
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 7576 2854 7604 2926
rect 7564 2848 7616 2854
rect 7564 2790 7616 2796
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 7760 2650 7788 2790
rect 7748 2644 7800 2650
rect 7748 2586 7800 2592
rect 7378 82 7434 480
rect 7116 54 7434 82
rect 5814 0 5870 54
rect 6550 0 6606 54
rect 7378 0 7434 54
rect 8114 82 8170 480
rect 8404 82 8432 2790
rect 8772 2514 8800 2926
rect 8760 2508 8812 2514
rect 8760 2450 8812 2456
rect 8114 54 8432 82
rect 8772 82 8800 2450
rect 8864 2378 8892 5238
rect 9048 5166 9076 5646
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9416 5370 9444 5510
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9036 5160 9088 5166
rect 9036 5102 9088 5108
rect 9508 4729 9536 8230
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9600 6322 9628 6598
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9494 4720 9550 4729
rect 9494 4655 9550 4664
rect 9496 4480 9548 4486
rect 9496 4422 9548 4428
rect 9404 4208 9456 4214
rect 9404 4150 9456 4156
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9324 3194 9352 4014
rect 9416 3738 9444 4150
rect 9508 4078 9536 4422
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9416 3466 9444 3674
rect 9404 3460 9456 3466
rect 9404 3402 9456 3408
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9140 2650 9168 3130
rect 9496 2916 9548 2922
rect 9496 2858 9548 2864
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 9508 2582 9536 2858
rect 9496 2576 9548 2582
rect 9496 2518 9548 2524
rect 8852 2372 8904 2378
rect 8852 2314 8904 2320
rect 8850 82 8906 480
rect 9600 134 9628 5102
rect 9692 4690 9720 10746
rect 9784 10606 9812 10950
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9784 10470 9812 10542
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9772 8560 9824 8566
rect 9772 8502 9824 8508
rect 9784 8294 9812 8502
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9772 5636 9824 5642
rect 9772 5578 9824 5584
rect 9784 5098 9812 5578
rect 9772 5092 9824 5098
rect 9772 5034 9824 5040
rect 9876 5030 9904 11494
rect 9968 10742 9996 11562
rect 10060 11218 10088 11834
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 9956 10736 10008 10742
rect 9956 10678 10008 10684
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9968 10266 9996 10542
rect 10060 10538 10088 11154
rect 10152 10810 10180 13738
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10980 13190 11008 14282
rect 11072 13870 11100 14418
rect 11164 14346 11192 14894
rect 11348 14550 11376 15506
rect 11716 14618 11744 15642
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 11336 14544 11388 14550
rect 11336 14486 11388 14492
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11152 14340 11204 14346
rect 11152 14282 11204 14288
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11060 13252 11112 13258
rect 11060 13194 11112 13200
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 11072 12782 11100 13194
rect 11256 12986 11284 13942
rect 11716 13802 11744 14418
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 10600 12776 10652 12782
rect 10784 12776 10836 12782
rect 10652 12736 10732 12764
rect 10600 12718 10652 12724
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 10612 11762 10640 12242
rect 10704 12238 10732 12736
rect 10784 12718 10836 12724
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 10796 12306 10824 12718
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 11072 12170 11100 12718
rect 11060 12164 11112 12170
rect 11060 12106 11112 12112
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10796 11694 10824 12038
rect 11348 11762 11376 13670
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11612 13252 11664 13258
rect 11612 13194 11664 13200
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 11624 11694 11652 13194
rect 11716 13190 11744 13330
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11716 12782 11744 13126
rect 11704 12776 11756 12782
rect 11704 12718 11756 12724
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10152 10538 10180 10746
rect 10428 10606 10456 11154
rect 10416 10600 10468 10606
rect 10416 10542 10468 10548
rect 10048 10532 10100 10538
rect 10048 10474 10100 10480
rect 10140 10532 10192 10538
rect 10140 10474 10192 10480
rect 10060 10266 10088 10474
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 9968 9178 9996 10202
rect 10704 10130 10732 11494
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 11428 11076 11480 11082
rect 11428 11018 11480 11024
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10152 9450 10180 10066
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 10140 9444 10192 9450
rect 10140 9386 10192 9392
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 11072 9042 11100 9454
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 11072 8838 11100 8978
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 9968 8430 9996 8774
rect 11072 8634 11100 8774
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9968 7954 9996 8366
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 10140 7948 10192 7954
rect 10140 7890 10192 7896
rect 10152 7206 10180 7890
rect 10692 7268 10744 7274
rect 10692 7210 10744 7216
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10048 6928 10100 6934
rect 10048 6870 10100 6876
rect 10060 6118 10088 6870
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9692 4214 9720 4626
rect 9968 4282 9996 4626
rect 10060 4486 10088 4966
rect 10152 4593 10180 7142
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10704 6798 10732 7210
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10704 5914 10732 6734
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10704 5030 10732 5102
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10704 4729 10732 4966
rect 10796 4826 10824 8230
rect 11060 5092 11112 5098
rect 11060 5034 11112 5040
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10690 4720 10746 4729
rect 10690 4655 10746 4664
rect 10138 4584 10194 4593
rect 10138 4519 10194 4528
rect 10692 4548 10744 4554
rect 10692 4490 10744 4496
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 10704 4282 10732 4490
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 9680 4208 9732 4214
rect 9680 4150 9732 4156
rect 9864 4208 9916 4214
rect 9864 4150 9916 4156
rect 9876 4060 9904 4150
rect 9692 4032 9904 4060
rect 9956 4072 10008 4078
rect 9692 3602 9720 4032
rect 9956 4014 10008 4020
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9692 2854 9720 3538
rect 9784 3058 9812 3878
rect 9968 3602 9996 4014
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9864 3460 9916 3466
rect 9864 3402 9916 3408
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9876 2990 9904 3402
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 8772 54 8906 82
rect 9588 128 9640 134
rect 9588 70 9640 76
rect 9678 82 9734 480
rect 9876 82 9904 2926
rect 9968 2922 9996 3538
rect 10796 3194 10824 4014
rect 10876 3460 10928 3466
rect 10876 3402 10928 3408
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 10888 3058 10916 3402
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 9956 2916 10008 2922
rect 9956 2858 10008 2864
rect 10876 2916 10928 2922
rect 10876 2858 10928 2864
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10888 2514 10916 2858
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 8114 0 8170 54
rect 8850 0 8906 54
rect 9678 54 9904 82
rect 10414 128 10470 480
rect 10414 76 10416 128
rect 10468 76 10470 128
rect 9678 0 9734 54
rect 10414 0 10470 76
rect 11072 82 11100 5034
rect 11164 4282 11192 11018
rect 11440 10810 11468 11018
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 11256 9518 11284 9590
rect 11244 9512 11296 9518
rect 11296 9472 11376 9500
rect 11244 9454 11296 9460
rect 11348 7177 11376 9472
rect 11520 9444 11572 9450
rect 11520 9386 11572 9392
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 11440 8294 11468 8978
rect 11532 8634 11560 9386
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 11426 7984 11482 7993
rect 11426 7919 11482 7928
rect 11334 7168 11390 7177
rect 11334 7103 11390 7112
rect 11244 6180 11296 6186
rect 11244 6122 11296 6128
rect 11256 4690 11284 6122
rect 11348 5778 11376 7103
rect 11440 6934 11468 7919
rect 11428 6928 11480 6934
rect 11428 6870 11480 6876
rect 11440 5914 11468 6870
rect 11624 6866 11652 9998
rect 11612 6860 11664 6866
rect 11716 6848 11744 12718
rect 11900 11286 11928 15846
rect 11992 12238 12020 22102
rect 12256 20256 12308 20262
rect 12256 20198 12308 20204
rect 12268 19786 12296 20198
rect 12256 19780 12308 19786
rect 12256 19722 12308 19728
rect 12268 18902 12296 19722
rect 12256 18896 12308 18902
rect 12256 18838 12308 18844
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12544 17134 12572 17818
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 12624 16720 12676 16726
rect 12624 16662 12676 16668
rect 12636 16046 12664 16662
rect 12624 16040 12676 16046
rect 12624 15982 12676 15988
rect 12636 15706 12664 15982
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12452 15094 12480 15506
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 12452 14958 12480 15030
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 12084 13394 12112 13806
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 12452 12918 12480 14894
rect 12532 13388 12584 13394
rect 12532 13330 12584 13336
rect 12544 12986 12572 13330
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 12544 12782 12572 12922
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12360 11898 12388 12038
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12360 11558 12388 11834
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 11888 11280 11940 11286
rect 11888 11222 11940 11228
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11808 10810 11836 11086
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11796 10124 11848 10130
rect 11796 10066 11848 10072
rect 11808 9382 11836 10066
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11900 7546 11928 7822
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11980 7472 12032 7478
rect 11980 7414 12032 7420
rect 11992 7002 12020 7414
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 12084 6905 12112 11494
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12544 10810 12572 11290
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12636 10266 12664 10474
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12728 9722 12756 23598
rect 13188 21010 13216 27520
rect 14738 27520 14794 28000
rect 16210 27532 16266 28000
rect 16210 27520 16212 27532
rect 14372 27474 14424 27480
rect 14096 21344 14148 21350
rect 14096 21286 14148 21292
rect 13176 21004 13228 21010
rect 13176 20946 13228 20952
rect 13188 20602 13216 20946
rect 13636 20936 13688 20942
rect 13636 20878 13688 20884
rect 13452 20800 13504 20806
rect 13452 20742 13504 20748
rect 13176 20596 13228 20602
rect 13176 20538 13228 20544
rect 13360 20256 13412 20262
rect 13360 20198 13412 20204
rect 13084 19168 13136 19174
rect 13084 19110 13136 19116
rect 13096 17882 13124 19110
rect 13084 17876 13136 17882
rect 13084 17818 13136 17824
rect 13372 17746 13400 20198
rect 13464 20058 13492 20742
rect 13452 20052 13504 20058
rect 13452 19994 13504 20000
rect 13544 19508 13596 19514
rect 13544 19450 13596 19456
rect 13556 19242 13584 19450
rect 13648 19378 13676 20878
rect 13728 20392 13780 20398
rect 13728 20334 13780 20340
rect 13636 19372 13688 19378
rect 13636 19314 13688 19320
rect 13544 19236 13596 19242
rect 13544 19178 13596 19184
rect 13648 18970 13676 19314
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 13740 18902 13768 20334
rect 13820 20324 13872 20330
rect 13820 20266 13872 20272
rect 13832 19990 13860 20266
rect 13820 19984 13872 19990
rect 13820 19926 13872 19932
rect 13832 19514 13860 19926
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13728 18896 13780 18902
rect 13728 18838 13780 18844
rect 13820 18896 13872 18902
rect 13820 18838 13872 18844
rect 13728 18760 13780 18766
rect 13728 18702 13780 18708
rect 13740 18426 13768 18702
rect 13728 18420 13780 18426
rect 13728 18362 13780 18368
rect 13636 18216 13688 18222
rect 13636 18158 13688 18164
rect 13648 17785 13676 18158
rect 13832 18086 13860 18838
rect 14108 18290 14136 21286
rect 14096 18284 14148 18290
rect 14096 18226 14148 18232
rect 14280 18148 14332 18154
rect 14280 18090 14332 18096
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13832 17814 13860 18022
rect 14096 17876 14148 17882
rect 14096 17818 14148 17824
rect 13820 17808 13872 17814
rect 13634 17776 13690 17785
rect 13360 17740 13412 17746
rect 14108 17785 14136 17818
rect 13820 17750 13872 17756
rect 14094 17776 14150 17785
rect 13634 17711 13690 17720
rect 13360 17682 13412 17688
rect 13832 17338 13860 17750
rect 13912 17740 13964 17746
rect 14094 17711 14150 17720
rect 13912 17682 13964 17688
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 12820 15978 12848 16594
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13464 16046 13492 16390
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 13452 16040 13504 16046
rect 13452 15982 13504 15988
rect 12808 15972 12860 15978
rect 12808 15914 12860 15920
rect 12912 15910 12940 15982
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 12912 15570 12940 15846
rect 13464 15570 13492 15982
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 13084 15564 13136 15570
rect 13084 15506 13136 15512
rect 13452 15564 13504 15570
rect 13452 15506 13504 15512
rect 12912 14958 12940 15506
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 13096 14890 13124 15506
rect 13084 14884 13136 14890
rect 13084 14826 13136 14832
rect 13096 14618 13124 14826
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 12912 13734 12940 14418
rect 13464 14346 13492 15506
rect 13648 14958 13676 16594
rect 13832 16182 13860 17070
rect 13924 16726 13952 17682
rect 14292 17610 14320 18090
rect 14280 17604 14332 17610
rect 14280 17546 14332 17552
rect 13912 16720 13964 16726
rect 13912 16662 13964 16668
rect 13820 16176 13872 16182
rect 13820 16118 13872 16124
rect 13912 15360 13964 15366
rect 13912 15302 13964 15308
rect 13924 15026 13952 15302
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 13648 14550 13676 14894
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13452 14340 13504 14346
rect 13452 14282 13504 14288
rect 13360 13796 13412 13802
rect 13360 13738 13412 13744
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12820 10266 12848 10610
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 12912 9761 12940 13670
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 13280 12782 13308 13330
rect 13268 12776 13320 12782
rect 13268 12718 13320 12724
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 13096 11354 13124 12242
rect 13280 12170 13308 12718
rect 13268 12164 13320 12170
rect 13268 12106 13320 12112
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 13188 11665 13216 11698
rect 13174 11656 13230 11665
rect 13174 11591 13230 11600
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 12992 10532 13044 10538
rect 13096 10520 13124 11290
rect 13188 10674 13216 11591
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 13044 10492 13124 10520
rect 13176 10532 13228 10538
rect 12992 10474 13044 10480
rect 13176 10474 13228 10480
rect 12898 9752 12954 9761
rect 12716 9716 12768 9722
rect 12898 9687 12954 9696
rect 12716 9658 12768 9664
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12176 8294 12204 8774
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 12176 8022 12204 8230
rect 12164 8016 12216 8022
rect 12164 7958 12216 7964
rect 12176 7206 12204 7958
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12070 6896 12126 6905
rect 11796 6860 11848 6866
rect 11716 6820 11796 6848
rect 11612 6802 11664 6808
rect 12070 6831 12126 6840
rect 11796 6802 11848 6808
rect 11624 6458 11652 6802
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11428 5908 11480 5914
rect 11428 5850 11480 5856
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 11348 5370 11376 5714
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11256 4214 11284 4626
rect 11426 4584 11482 4593
rect 11426 4519 11482 4528
rect 11244 4208 11296 4214
rect 11244 4150 11296 4156
rect 11440 3738 11468 4519
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 11152 3120 11204 3126
rect 11152 3062 11204 3068
rect 11164 2582 11192 3062
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 11242 82 11298 480
rect 11072 54 11298 82
rect 11624 82 11652 6258
rect 11808 6254 11836 6802
rect 12360 6730 12388 9318
rect 12532 9104 12584 9110
rect 12532 9046 12584 9052
rect 12544 8838 12572 9046
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12544 8362 12572 8774
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12728 8090 12756 8910
rect 12912 8566 12940 9454
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12452 7546 12480 8026
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12716 7200 12768 7206
rect 12716 7142 12768 7148
rect 12348 6724 12400 6730
rect 12348 6666 12400 6672
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 12164 5772 12216 5778
rect 12164 5714 12216 5720
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 11716 3058 11744 5578
rect 12176 5166 12204 5714
rect 12164 5160 12216 5166
rect 12164 5102 12216 5108
rect 12176 4826 12204 5102
rect 12256 5092 12308 5098
rect 12256 5034 12308 5040
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11716 2582 11744 2994
rect 11704 2576 11756 2582
rect 11704 2518 11756 2524
rect 11808 2446 11836 4626
rect 12072 4004 12124 4010
rect 12072 3946 12124 3952
rect 12084 3738 12112 3946
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 12084 3058 12112 3674
rect 12268 3534 12296 5034
rect 12256 3528 12308 3534
rect 12256 3470 12308 3476
rect 12072 3052 12124 3058
rect 12072 2994 12124 3000
rect 12268 2650 12296 3470
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 11978 82 12034 480
rect 12360 116 12388 6666
rect 12728 6118 12756 7142
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12532 5296 12584 5302
rect 12532 5238 12584 5244
rect 12544 4826 12572 5238
rect 12728 5030 12756 6054
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12544 4078 12572 4762
rect 12728 4758 12756 4966
rect 12716 4752 12768 4758
rect 12716 4694 12768 4700
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12636 4146 12664 4558
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12532 4072 12584 4078
rect 12532 4014 12584 4020
rect 12636 3534 12664 4082
rect 12728 3942 12756 4694
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12728 3670 12756 3878
rect 12820 3738 12848 5646
rect 13096 5574 13124 9318
rect 13188 8401 13216 10474
rect 13372 9722 13400 13738
rect 13464 12782 13492 14282
rect 13544 13728 13596 13734
rect 13544 13670 13596 13676
rect 13556 13462 13584 13670
rect 13544 13456 13596 13462
rect 13544 13398 13596 13404
rect 13648 13394 13676 14486
rect 14292 14482 14320 14758
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14188 14408 14240 14414
rect 14188 14350 14240 14356
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13832 13530 13860 13806
rect 13912 13796 13964 13802
rect 13912 13738 13964 13744
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 13832 12918 13860 13466
rect 13820 12912 13872 12918
rect 13820 12854 13872 12860
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 13740 11286 13768 12310
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13832 11354 13860 11494
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13728 11280 13780 11286
rect 13924 11234 13952 13738
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 14016 11354 14044 12174
rect 14200 11762 14228 14350
rect 14292 14074 14320 14418
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14096 11688 14148 11694
rect 14096 11630 14148 11636
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 13728 11222 13780 11228
rect 13832 11206 13952 11234
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13360 9716 13412 9722
rect 13360 9658 13412 9664
rect 13556 9586 13584 9862
rect 13636 9716 13688 9722
rect 13688 9664 13768 9674
rect 13636 9658 13768 9664
rect 13648 9654 13768 9658
rect 13648 9648 13780 9654
rect 13648 9646 13728 9648
rect 13728 9590 13780 9596
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13740 8430 13768 9590
rect 13728 8424 13780 8430
rect 13174 8392 13230 8401
rect 13728 8366 13780 8372
rect 13174 8327 13230 8336
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 13372 8022 13400 8230
rect 13360 8016 13412 8022
rect 13360 7958 13412 7964
rect 13372 7426 13400 7958
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13740 7546 13768 7822
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13372 7398 13492 7426
rect 13360 7336 13412 7342
rect 13358 7304 13360 7313
rect 13412 7304 13414 7313
rect 13358 7239 13414 7248
rect 13372 7206 13400 7239
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 13464 7002 13492 7398
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13544 6928 13596 6934
rect 13544 6870 13596 6876
rect 13832 6882 13860 11206
rect 13912 10124 13964 10130
rect 13912 10066 13964 10072
rect 13924 9382 13952 10066
rect 14108 9897 14136 11630
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14200 10198 14228 10406
rect 14188 10192 14240 10198
rect 14188 10134 14240 10140
rect 14094 9888 14150 9897
rect 14094 9823 14150 9832
rect 14200 9761 14228 10134
rect 14292 10130 14320 13126
rect 14384 11898 14412 27474
rect 14752 23866 14780 27520
rect 16264 27520 16266 27532
rect 17774 27520 17830 28000
rect 19338 27520 19394 28000
rect 20902 27520 20958 28000
rect 22466 27520 22522 28000
rect 24030 27520 24086 28000
rect 25594 27520 25650 28000
rect 27158 27520 27214 28000
rect 16212 27474 16264 27480
rect 16224 27443 16252 27474
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 17788 23866 17816 27520
rect 19352 23866 19380 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20916 23866 20944 27520
rect 14740 23860 14792 23866
rect 14740 23802 14792 23808
rect 17776 23860 17828 23866
rect 17776 23802 17828 23808
rect 19340 23860 19392 23866
rect 19340 23802 19392 23808
rect 20904 23860 20956 23866
rect 20904 23802 20956 23808
rect 22480 23798 22508 27520
rect 23848 24268 23900 24274
rect 23848 24210 23900 24216
rect 23860 23798 23888 24210
rect 24044 23866 24072 27520
rect 24950 26752 25006 26761
rect 24950 26687 25006 26696
rect 24766 25392 24822 25401
rect 24766 25327 24822 25336
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24124 24744 24176 24750
rect 24124 24686 24176 24692
rect 24032 23860 24084 23866
rect 24032 23802 24084 23808
rect 22468 23792 22520 23798
rect 22468 23734 22520 23740
rect 23848 23792 23900 23798
rect 23848 23734 23900 23740
rect 15384 23656 15436 23662
rect 15384 23598 15436 23604
rect 17224 23656 17276 23662
rect 17224 23598 17276 23604
rect 19524 23656 19576 23662
rect 19524 23598 19576 23604
rect 22008 23656 22060 23662
rect 22008 23598 22060 23604
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14740 21684 14792 21690
rect 14740 21626 14792 21632
rect 14648 20256 14700 20262
rect 14648 20198 14700 20204
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 14476 18834 14504 19790
rect 14464 18828 14516 18834
rect 14464 18770 14516 18776
rect 14660 18766 14688 20198
rect 14648 18760 14700 18766
rect 14648 18702 14700 18708
rect 14464 18284 14516 18290
rect 14464 18226 14516 18232
rect 14476 17882 14504 18226
rect 14464 17876 14516 17882
rect 14464 17818 14516 17824
rect 14648 17128 14700 17134
rect 14648 17070 14700 17076
rect 14556 17060 14608 17066
rect 14556 17002 14608 17008
rect 14568 15978 14596 17002
rect 14660 16794 14688 17070
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 14752 16130 14780 21626
rect 15290 21584 15346 21593
rect 15290 21519 15346 21528
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15304 20398 15332 21519
rect 15292 20392 15344 20398
rect 15292 20334 15344 20340
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15304 19242 15332 19790
rect 15016 19236 15068 19242
rect 15016 19178 15068 19184
rect 15292 19236 15344 19242
rect 15292 19178 15344 19184
rect 15028 18970 15056 19178
rect 15396 19174 15424 23598
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 15660 19236 15712 19242
rect 15660 19178 15712 19184
rect 15384 19168 15436 19174
rect 15384 19110 15436 19116
rect 15016 18964 15068 18970
rect 14844 18924 15016 18952
rect 14844 18358 14872 18924
rect 15016 18906 15068 18912
rect 15476 18896 15528 18902
rect 15476 18838 15528 18844
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15396 18358 15424 18702
rect 15488 18426 15516 18838
rect 15672 18766 15700 19178
rect 15660 18760 15712 18766
rect 15660 18702 15712 18708
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 14832 18352 14884 18358
rect 14832 18294 14884 18300
rect 15384 18352 15436 18358
rect 15384 18294 15436 18300
rect 15384 17808 15436 17814
rect 15384 17750 15436 17756
rect 15396 17649 15424 17750
rect 15382 17640 15438 17649
rect 15382 17575 15438 17584
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15396 16794 15424 17575
rect 15488 17338 15516 18362
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 15384 16788 15436 16794
rect 15384 16730 15436 16736
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14660 16102 14780 16130
rect 15384 16108 15436 16114
rect 14556 15972 14608 15978
rect 14556 15914 14608 15920
rect 14660 15178 14688 16102
rect 15384 16050 15436 16056
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 14752 15366 14780 15982
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14660 15150 14780 15178
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 14660 12986 14688 14350
rect 14648 12980 14700 12986
rect 14648 12922 14700 12928
rect 14660 12714 14688 12922
rect 14648 12708 14700 12714
rect 14648 12650 14700 12656
rect 14648 12300 14700 12306
rect 14752 12288 14780 15150
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 14832 14884 14884 14890
rect 14832 14826 14884 14832
rect 14844 14618 14872 14826
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15304 14074 15332 14962
rect 15396 14074 15424 16050
rect 15752 15972 15804 15978
rect 15752 15914 15804 15920
rect 15764 15638 15792 15914
rect 15752 15632 15804 15638
rect 15752 15574 15804 15580
rect 15764 14822 15792 15574
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15384 14068 15436 14074
rect 15384 14010 15436 14016
rect 15304 13938 15332 14010
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 14832 13728 14884 13734
rect 14832 13670 14884 13676
rect 14844 12918 14872 13670
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14832 12912 14884 12918
rect 14832 12854 14884 12860
rect 14844 12442 14872 12854
rect 15304 12850 15332 13874
rect 15396 13870 15424 14010
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15396 13433 15424 13806
rect 15488 13802 15516 14418
rect 15476 13796 15528 13802
rect 15476 13738 15528 13744
rect 15764 13462 15792 14758
rect 15752 13456 15804 13462
rect 15382 13424 15438 13433
rect 15752 13398 15804 13404
rect 15382 13359 15438 13368
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 15396 12986 15424 13262
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15764 12918 15792 13398
rect 15752 12912 15804 12918
rect 15752 12854 15804 12860
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 14832 12436 14884 12442
rect 14832 12378 14884 12384
rect 15764 12306 15792 12854
rect 14700 12260 14780 12288
rect 15752 12300 15804 12306
rect 14648 12242 14700 12248
rect 15752 12242 15804 12248
rect 14372 11892 14424 11898
rect 14372 11834 14424 11840
rect 14660 11558 14688 12242
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15764 11626 15792 12242
rect 15752 11620 15804 11626
rect 15752 11562 15804 11568
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14568 10470 14596 11154
rect 14660 10577 14688 11494
rect 15764 11286 15792 11562
rect 15752 11280 15804 11286
rect 15752 11222 15804 11228
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 14832 11008 14884 11014
rect 14832 10950 14884 10956
rect 14646 10568 14702 10577
rect 14646 10503 14702 10512
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14186 9752 14242 9761
rect 14186 9687 14242 9696
rect 14096 9512 14148 9518
rect 14096 9454 14148 9460
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 14004 8832 14056 8838
rect 14004 8774 14056 8780
rect 14016 8634 14044 8774
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 14016 8362 14044 8570
rect 14004 8356 14056 8362
rect 14004 8298 14056 8304
rect 13912 7268 13964 7274
rect 13912 7210 13964 7216
rect 13924 7002 13952 7210
rect 13912 6996 13964 7002
rect 13912 6938 13964 6944
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 13188 6458 13216 6734
rect 13360 6656 13412 6662
rect 13556 6644 13584 6870
rect 13832 6854 14044 6882
rect 13412 6616 13584 6644
rect 13360 6598 13412 6604
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13360 6384 13412 6390
rect 13360 6326 13412 6332
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 13268 6112 13320 6118
rect 13268 6054 13320 6060
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 13096 5166 13124 5510
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 12716 3664 12768 3670
rect 12716 3606 12768 3612
rect 12624 3528 12676 3534
rect 12624 3470 12676 3476
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12544 2922 12572 3334
rect 12728 3058 12756 3606
rect 12716 3052 12768 3058
rect 12716 2994 12768 3000
rect 12714 2952 12770 2961
rect 12532 2916 12584 2922
rect 12714 2887 12770 2896
rect 12532 2858 12584 2864
rect 12728 2514 12756 2887
rect 12912 2553 12940 3878
rect 13188 2961 13216 6054
rect 13280 4593 13308 6054
rect 13266 4584 13322 4593
rect 13266 4519 13322 4528
rect 13372 4146 13400 6326
rect 13556 5914 13584 6616
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13832 5930 13860 6190
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13648 5902 13860 5930
rect 13544 5772 13596 5778
rect 13648 5760 13676 5902
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 13596 5732 13676 5760
rect 13544 5714 13596 5720
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13740 4486 13768 5646
rect 13832 4826 13860 5782
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13728 4480 13780 4486
rect 13728 4422 13780 4428
rect 14016 4154 14044 6854
rect 14108 6254 14136 9454
rect 14188 9444 14240 9450
rect 14188 9386 14240 9392
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 14200 5234 14228 9386
rect 14292 9178 14320 10066
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 14384 8974 14412 9998
rect 14464 9988 14516 9994
rect 14464 9930 14516 9936
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 14292 8498 14320 8774
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14292 7818 14320 8434
rect 14280 7812 14332 7818
rect 14280 7754 14332 7760
rect 14292 7410 14320 7754
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14292 6730 14320 7346
rect 14280 6724 14332 6730
rect 14280 6666 14332 6672
rect 14476 5370 14504 9930
rect 14568 7313 14596 10406
rect 14648 7812 14700 7818
rect 14648 7754 14700 7760
rect 14660 7721 14688 7754
rect 14646 7712 14702 7721
rect 14646 7647 14702 7656
rect 14554 7304 14610 7313
rect 14554 7239 14610 7248
rect 14752 7002 14780 10950
rect 14844 10538 14872 10950
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15304 10742 15332 11086
rect 15764 10810 15792 11222
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 15292 10736 15344 10742
rect 15292 10678 15344 10684
rect 14832 10532 14884 10538
rect 14832 10474 14884 10480
rect 14832 10192 14884 10198
rect 15304 10169 15332 10678
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 14832 10134 14884 10140
rect 15290 10160 15346 10169
rect 14844 9178 14872 10134
rect 15290 10095 15346 10104
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15396 9518 15424 9862
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 14832 9172 14884 9178
rect 14832 9114 14884 9120
rect 14844 7478 14872 9114
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15396 8090 15424 9454
rect 15488 9382 15516 10066
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15580 9042 15608 10202
rect 15764 9722 15792 10746
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15764 9450 15792 9658
rect 15856 9450 15884 20198
rect 15936 19916 15988 19922
rect 15936 19858 15988 19864
rect 15948 19514 15976 19858
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 15948 18970 15976 19450
rect 16672 19168 16724 19174
rect 16672 19110 16724 19116
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 16212 18216 16264 18222
rect 16212 18158 16264 18164
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 16040 17814 16068 18022
rect 16028 17808 16080 17814
rect 16028 17750 16080 17756
rect 16040 17270 16068 17750
rect 16224 17338 16252 18158
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 16028 17264 16080 17270
rect 16028 17206 16080 17212
rect 16224 16998 16252 17274
rect 16500 17202 16528 17546
rect 16488 17196 16540 17202
rect 16488 17138 16540 17144
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 16224 16726 16252 16934
rect 16212 16720 16264 16726
rect 16212 16662 16264 16668
rect 16224 16250 16252 16662
rect 16212 16244 16264 16250
rect 16212 16186 16264 16192
rect 16224 15706 16252 16186
rect 16488 15904 16540 15910
rect 16488 15846 16540 15852
rect 16212 15700 16264 15706
rect 16212 15642 16264 15648
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 16132 15162 16160 15438
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 16500 14550 16528 15846
rect 16488 14544 16540 14550
rect 16488 14486 16540 14492
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 16224 13802 16252 14214
rect 16212 13796 16264 13802
rect 16212 13738 16264 13744
rect 16224 13394 16252 13738
rect 16500 13530 16528 14486
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16212 13388 16264 13394
rect 16212 13330 16264 13336
rect 16684 13297 16712 19110
rect 17236 18193 17264 23598
rect 19340 23588 19392 23594
rect 19340 23530 19392 23536
rect 18604 21888 18656 21894
rect 18604 21830 18656 21836
rect 18616 21049 18644 21830
rect 18602 21040 18658 21049
rect 18602 20975 18658 20984
rect 17222 18184 17278 18193
rect 17222 18119 17278 18128
rect 17040 17808 17092 17814
rect 17040 17750 17092 17756
rect 16764 17672 16816 17678
rect 16764 17614 16816 17620
rect 16776 17202 16804 17614
rect 17052 17338 17080 17750
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17040 17332 17092 17338
rect 16960 17292 17040 17320
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 16776 16794 16804 17138
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 16960 16182 16988 17292
rect 17040 17274 17092 17280
rect 17040 16584 17092 16590
rect 17040 16526 17092 16532
rect 16948 16176 17000 16182
rect 16868 16136 16948 16164
rect 16868 14958 16896 16136
rect 16948 16118 17000 16124
rect 17052 15910 17080 16526
rect 17132 16516 17184 16522
rect 17132 16458 17184 16464
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 17052 15706 17080 15846
rect 17040 15700 17092 15706
rect 17040 15642 17092 15648
rect 17144 15502 17172 16458
rect 17604 16046 17632 17614
rect 17776 17264 17828 17270
rect 17776 17206 17828 17212
rect 17788 16726 17816 17206
rect 18052 16992 18104 16998
rect 18052 16934 18104 16940
rect 17776 16720 17828 16726
rect 17776 16662 17828 16668
rect 17788 16250 17816 16662
rect 18064 16590 18092 16934
rect 18052 16584 18104 16590
rect 18052 16526 18104 16532
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 18524 16250 18552 16526
rect 17776 16244 17828 16250
rect 17776 16186 17828 16192
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 19352 16114 19380 23530
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17224 15632 17276 15638
rect 17224 15574 17276 15580
rect 17132 15496 17184 15502
rect 17132 15438 17184 15444
rect 17144 15162 17172 15438
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 17236 15026 17264 15574
rect 17604 15502 17632 15982
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 17592 15496 17644 15502
rect 17592 15438 17644 15444
rect 18052 15360 18104 15366
rect 18052 15302 18104 15308
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16868 14618 16896 14894
rect 16856 14612 16908 14618
rect 16856 14554 16908 14560
rect 16960 14414 16988 14894
rect 17040 14544 17092 14550
rect 17040 14486 17092 14492
rect 16948 14408 17000 14414
rect 16948 14350 17000 14356
rect 16960 13938 16988 14350
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 17052 13734 17080 14486
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 17132 13796 17184 13802
rect 17132 13738 17184 13744
rect 17040 13728 17092 13734
rect 17040 13670 17092 13676
rect 17052 13462 17080 13670
rect 17040 13456 17092 13462
rect 17040 13398 17092 13404
rect 16670 13288 16726 13297
rect 16670 13223 16726 13232
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 16500 12753 16528 12786
rect 16486 12744 16542 12753
rect 16542 12702 16620 12730
rect 16486 12679 16542 12688
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16120 12368 16172 12374
rect 16120 12310 16172 12316
rect 15934 12200 15990 12209
rect 15934 12135 15990 12144
rect 15752 9444 15804 9450
rect 15752 9386 15804 9392
rect 15844 9444 15896 9450
rect 15844 9386 15896 9392
rect 15764 9330 15792 9386
rect 15764 9302 15884 9330
rect 15856 9178 15884 9302
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15844 9172 15896 9178
rect 15844 9114 15896 9120
rect 15568 9036 15620 9042
rect 15568 8978 15620 8984
rect 15580 8634 15608 8978
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15764 7954 15792 9114
rect 15856 8634 15884 9114
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14832 7472 14884 7478
rect 14832 7414 14884 7420
rect 15304 7206 15332 7890
rect 15844 7472 15896 7478
rect 15842 7440 15844 7449
rect 15896 7440 15898 7449
rect 15842 7375 15898 7384
rect 15856 7342 15884 7375
rect 15844 7336 15896 7342
rect 15844 7278 15896 7284
rect 14832 7200 14884 7206
rect 14832 7142 14884 7148
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 14740 6996 14792 7002
rect 14740 6938 14792 6944
rect 14844 6118 14872 7142
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15396 6322 15424 6938
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 15200 6180 15252 6186
rect 15476 6180 15528 6186
rect 15200 6122 15252 6128
rect 15396 6140 15476 6168
rect 14832 6112 14884 6118
rect 14832 6054 14884 6060
rect 15212 5778 15240 6122
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15304 5828 15332 6054
rect 15396 5828 15424 6140
rect 15476 6122 15528 6128
rect 15660 6112 15712 6118
rect 15660 6054 15712 6060
rect 15672 5914 15700 6054
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15304 5800 15424 5828
rect 15200 5772 15252 5778
rect 15252 5732 15332 5760
rect 15200 5714 15252 5720
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 14200 4826 14228 5170
rect 15304 4826 15332 5732
rect 15396 5370 15424 5800
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15396 4758 15424 5306
rect 15672 5098 15700 5850
rect 15752 5160 15804 5166
rect 15752 5102 15804 5108
rect 15660 5092 15712 5098
rect 15660 5034 15712 5040
rect 15660 4820 15712 4826
rect 15660 4762 15712 4768
rect 15384 4752 15436 4758
rect 15384 4694 15436 4700
rect 14556 4684 14608 4690
rect 14556 4626 14608 4632
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 14384 4185 14412 4218
rect 14464 4208 14516 4214
rect 14370 4176 14426 4185
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 13452 4140 13504 4146
rect 14016 4126 14136 4154
rect 13452 4082 13504 4088
rect 13464 4049 13492 4082
rect 13450 4040 13506 4049
rect 13450 3975 13506 3984
rect 14004 4004 14056 4010
rect 14004 3946 14056 3952
rect 14016 3670 14044 3946
rect 14004 3664 14056 3670
rect 14004 3606 14056 3612
rect 14016 3126 14044 3606
rect 14108 3602 14136 4126
rect 14464 4150 14516 4156
rect 14370 4111 14426 4120
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 14108 3194 14136 3538
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 14096 3188 14148 3194
rect 14096 3130 14148 3136
rect 14004 3120 14056 3126
rect 14004 3062 14056 3068
rect 13174 2952 13230 2961
rect 13174 2887 13230 2896
rect 12898 2544 12954 2553
rect 12716 2508 12768 2514
rect 12898 2479 12954 2488
rect 12716 2450 12768 2456
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 12360 88 12480 116
rect 11624 54 12034 82
rect 12452 82 12480 88
rect 12806 82 12862 480
rect 12912 134 12940 2246
rect 13188 1737 13216 2887
rect 13636 2848 13688 2854
rect 13636 2790 13688 2796
rect 14004 2848 14056 2854
rect 14004 2790 14056 2796
rect 13174 1728 13230 1737
rect 13174 1663 13230 1672
rect 12452 54 12862 82
rect 12900 128 12952 134
rect 12900 70 12952 76
rect 13542 82 13598 480
rect 13648 82 13676 2790
rect 14016 2582 14044 2790
rect 14004 2576 14056 2582
rect 14004 2518 14056 2524
rect 11242 0 11298 54
rect 11978 0 12034 54
rect 12806 0 12862 54
rect 13542 54 13676 82
rect 14292 66 14320 3334
rect 14370 82 14426 480
rect 14476 82 14504 4150
rect 14568 4010 14596 4626
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14556 4004 14608 4010
rect 14556 3946 14608 3952
rect 14568 2582 14596 3946
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14660 3398 14688 3674
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 14660 3058 14688 3334
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 14556 2576 14608 2582
rect 14556 2518 14608 2524
rect 14844 2417 14872 3878
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 15028 3505 15056 3538
rect 15014 3496 15070 3505
rect 15014 3431 15070 3440
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15200 3120 15252 3126
rect 15200 3062 15252 3068
rect 15212 2582 15240 3062
rect 15304 2854 15332 3878
rect 15396 3670 15424 4694
rect 15672 4690 15700 4762
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15764 3670 15792 5102
rect 15844 5024 15896 5030
rect 15844 4966 15896 4972
rect 15856 4010 15884 4966
rect 15844 4004 15896 4010
rect 15844 3946 15896 3952
rect 15384 3664 15436 3670
rect 15384 3606 15436 3612
rect 15752 3664 15804 3670
rect 15752 3606 15804 3612
rect 15396 3194 15424 3606
rect 15660 3392 15712 3398
rect 15660 3334 15712 3340
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15672 3058 15700 3334
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 15200 2576 15252 2582
rect 15200 2518 15252 2524
rect 14830 2408 14886 2417
rect 14830 2343 14886 2352
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15672 1601 15700 2994
rect 15948 2446 15976 12135
rect 16132 11694 16160 12310
rect 16224 12102 16252 12582
rect 16592 12374 16620 12702
rect 16488 12368 16540 12374
rect 16488 12310 16540 12316
rect 16580 12368 16632 12374
rect 16580 12310 16632 12316
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 16132 11354 16160 11630
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16224 9518 16252 12038
rect 16500 11898 16528 12310
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16212 9512 16264 9518
rect 16212 9454 16264 9460
rect 16120 9444 16172 9450
rect 16120 9386 16172 9392
rect 16132 6390 16160 9386
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16316 6866 16344 9318
rect 16408 9178 16436 10406
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16592 8412 16620 12038
rect 16684 10606 16712 13223
rect 16948 12912 17000 12918
rect 16948 12854 17000 12860
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 16776 12238 16804 12786
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16776 11354 16804 12174
rect 16764 11348 16816 11354
rect 16764 11290 16816 11296
rect 16776 10674 16804 11290
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16868 9450 16896 10066
rect 16960 9654 16988 12854
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 17052 11830 17080 12174
rect 17040 11824 17092 11830
rect 17040 11766 17092 11772
rect 16948 9648 17000 9654
rect 16948 9590 17000 9596
rect 16856 9444 16908 9450
rect 16856 9386 16908 9392
rect 16672 8424 16724 8430
rect 16592 8384 16672 8412
rect 16672 8366 16724 8372
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 16500 8090 16528 8298
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16684 7818 16712 8366
rect 16672 7812 16724 7818
rect 16672 7754 16724 7760
rect 16960 7410 16988 9590
rect 17144 7954 17172 13738
rect 17224 13456 17276 13462
rect 17224 13398 17276 13404
rect 17236 10198 17264 13398
rect 17224 10192 17276 10198
rect 17224 10134 17276 10140
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 17132 7948 17184 7954
rect 17132 7890 17184 7896
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16868 6866 16896 7278
rect 17038 6896 17094 6905
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 16856 6860 16908 6866
rect 17038 6831 17094 6840
rect 16856 6802 16908 6808
rect 16316 6390 16344 6802
rect 16120 6384 16172 6390
rect 16120 6326 16172 6332
rect 16304 6384 16356 6390
rect 16304 6326 16356 6332
rect 16764 6384 16816 6390
rect 16868 6372 16896 6802
rect 17052 6458 17080 6831
rect 17040 6452 17092 6458
rect 17040 6394 17092 6400
rect 16816 6344 16896 6372
rect 16764 6326 16816 6332
rect 16764 6180 16816 6186
rect 16764 6122 16816 6128
rect 16120 5636 16172 5642
rect 16120 5578 16172 5584
rect 16132 5234 16160 5578
rect 16212 5568 16264 5574
rect 16212 5510 16264 5516
rect 16120 5228 16172 5234
rect 16120 5170 16172 5176
rect 16132 5137 16160 5170
rect 16118 5128 16174 5137
rect 16224 5098 16252 5510
rect 16776 5098 16804 6122
rect 17236 5846 17264 9862
rect 17328 9042 17356 14418
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 17420 12986 17448 13330
rect 17512 13190 17540 13670
rect 17592 13524 17644 13530
rect 17592 13466 17644 13472
rect 17500 13184 17552 13190
rect 17500 13126 17552 13132
rect 17408 12980 17460 12986
rect 17408 12922 17460 12928
rect 17604 11218 17632 13466
rect 17972 12374 18000 14962
rect 18064 14958 18092 15302
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 18708 14822 18736 15506
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 18144 14476 18196 14482
rect 18144 14418 18196 14424
rect 18512 14476 18564 14482
rect 18512 14418 18564 14424
rect 18156 14074 18184 14418
rect 18144 14068 18196 14074
rect 18144 14010 18196 14016
rect 18328 13728 18380 13734
rect 18328 13670 18380 13676
rect 18420 13728 18472 13734
rect 18420 13670 18472 13676
rect 18144 12708 18196 12714
rect 18144 12650 18196 12656
rect 18156 12442 18184 12650
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 17960 12368 18012 12374
rect 17960 12310 18012 12316
rect 18052 12368 18104 12374
rect 18052 12310 18104 12316
rect 17972 11898 18000 12310
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 17960 11688 18012 11694
rect 18064 11676 18092 12310
rect 18012 11648 18092 11676
rect 17960 11630 18012 11636
rect 17960 11552 18012 11558
rect 17960 11494 18012 11500
rect 17972 11354 18000 11494
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 17684 11280 17736 11286
rect 17684 11222 17736 11228
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17604 10266 17632 11154
rect 17696 10742 17724 11222
rect 18064 11082 18092 11648
rect 18052 11076 18104 11082
rect 18052 11018 18104 11024
rect 17684 10736 17736 10742
rect 17684 10678 17736 10684
rect 17696 10538 17724 10678
rect 17684 10532 17736 10538
rect 17684 10474 17736 10480
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 17500 10056 17552 10062
rect 17500 9998 17552 10004
rect 17512 9382 17540 9998
rect 17696 9722 17724 10474
rect 18144 10192 18196 10198
rect 18144 10134 18196 10140
rect 17684 9716 17736 9722
rect 17684 9658 17736 9664
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17316 9036 17368 9042
rect 17316 8978 17368 8984
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 17130 5264 17186 5273
rect 17130 5199 17186 5208
rect 16118 5063 16174 5072
rect 16212 5092 16264 5098
rect 16212 5034 16264 5040
rect 16764 5092 16816 5098
rect 16764 5034 16816 5040
rect 16776 4826 16804 5034
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 16396 4752 16448 4758
rect 16396 4694 16448 4700
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 16028 4548 16080 4554
rect 16028 4490 16080 4496
rect 16040 3942 16068 4490
rect 16224 4282 16252 4558
rect 16408 4282 16436 4694
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 16212 4276 16264 4282
rect 16212 4218 16264 4224
rect 16396 4276 16448 4282
rect 16396 4218 16448 4224
rect 16486 4176 16542 4185
rect 16486 4111 16542 4120
rect 16120 4004 16172 4010
rect 16120 3946 16172 3952
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 16040 2825 16068 3878
rect 16132 3534 16160 3946
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 16132 3058 16160 3470
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 16120 2916 16172 2922
rect 16120 2858 16172 2864
rect 16026 2816 16082 2825
rect 16026 2751 16082 2760
rect 16028 2644 16080 2650
rect 16028 2586 16080 2592
rect 15936 2440 15988 2446
rect 15936 2382 15988 2388
rect 15658 1592 15714 1601
rect 15658 1527 15714 1536
rect 14280 60 14332 66
rect 13542 0 13598 54
rect 14280 2 14332 8
rect 14370 54 14504 82
rect 15106 128 15162 480
rect 15106 76 15108 128
rect 15160 76 15162 128
rect 14370 0 14426 54
rect 15106 0 15162 76
rect 15842 82 15898 480
rect 16040 82 16068 2586
rect 16132 2582 16160 2858
rect 16120 2576 16172 2582
rect 16120 2518 16172 2524
rect 15842 54 16068 82
rect 16500 82 16528 4111
rect 16592 4078 16620 4422
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16776 2582 16804 4762
rect 16854 4040 16910 4049
rect 16854 3975 16910 3984
rect 16868 2650 16896 3975
rect 17144 3602 17172 5199
rect 17328 4282 17356 8978
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 17420 7546 17448 7890
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 17512 7002 17540 9318
rect 17684 9036 17736 9042
rect 17684 8978 17736 8984
rect 17696 8294 17724 8978
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 17972 8498 18000 8774
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 17684 8288 17736 8294
rect 17684 8230 17736 8236
rect 17592 7880 17644 7886
rect 17696 7857 17724 8230
rect 17880 7954 17908 8366
rect 18064 8362 18092 9454
rect 18156 9178 18184 10134
rect 18340 9586 18368 13670
rect 18328 9580 18380 9586
rect 18328 9522 18380 9528
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 18052 8356 18104 8362
rect 18052 8298 18104 8304
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 17592 7822 17644 7828
rect 17682 7848 17738 7857
rect 17500 6996 17552 7002
rect 17500 6938 17552 6944
rect 17604 6866 17632 7822
rect 17682 7783 17738 7792
rect 17880 7546 17908 7890
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17880 7342 17908 7482
rect 17868 7336 17920 7342
rect 17868 7278 17920 7284
rect 17684 6928 17736 6934
rect 17684 6870 17736 6876
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17604 5914 17632 6802
rect 17696 6118 17724 6870
rect 17972 6254 18000 8298
rect 18064 8090 18092 8298
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 18432 7392 18460 13670
rect 18524 13462 18552 14418
rect 18708 14385 18736 14758
rect 18788 14408 18840 14414
rect 18694 14376 18750 14385
rect 18788 14350 18840 14356
rect 18694 14311 18750 14320
rect 18696 13932 18748 13938
rect 18696 13874 18748 13880
rect 18512 13456 18564 13462
rect 18512 13398 18564 13404
rect 18708 13258 18736 13874
rect 18696 13252 18748 13258
rect 18696 13194 18748 13200
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18616 12170 18644 12786
rect 18604 12164 18656 12170
rect 18604 12106 18656 12112
rect 18800 11354 18828 14350
rect 18880 13388 18932 13394
rect 18880 13330 18932 13336
rect 19064 13388 19116 13394
rect 19064 13330 19116 13336
rect 18892 12102 18920 13330
rect 19076 12986 19104 13330
rect 19064 12980 19116 12986
rect 19064 12922 19116 12928
rect 19432 12912 19484 12918
rect 19062 12880 19118 12889
rect 19432 12854 19484 12860
rect 19062 12815 19118 12824
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18696 11008 18748 11014
rect 18696 10950 18748 10956
rect 18708 10810 18736 10950
rect 18696 10804 18748 10810
rect 18696 10746 18748 10752
rect 18800 10674 18828 11290
rect 18972 11280 19024 11286
rect 18972 11222 19024 11228
rect 18880 11144 18932 11150
rect 18880 11086 18932 11092
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 18892 10198 18920 11086
rect 18984 10810 19012 11222
rect 18972 10804 19024 10810
rect 18972 10746 19024 10752
rect 18880 10192 18932 10198
rect 18880 10134 18932 10140
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18708 8090 18736 8910
rect 18892 8498 18920 10134
rect 19076 10130 19104 12815
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19156 11892 19208 11898
rect 19156 11834 19208 11840
rect 19168 11132 19196 11834
rect 19260 11830 19288 12242
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 19248 11824 19300 11830
rect 19248 11766 19300 11772
rect 19260 11286 19288 11766
rect 19352 11762 19380 12038
rect 19340 11756 19392 11762
rect 19340 11698 19392 11704
rect 19444 11642 19472 12854
rect 19536 12442 19564 23598
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 22020 21690 22048 23598
rect 22652 23588 22704 23594
rect 22652 23530 22704 23536
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 20442 18184 20498 18193
rect 20442 18119 20498 18128
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19798 16008 19854 16017
rect 19720 15978 19798 15994
rect 19708 15972 19798 15978
rect 19760 15966 19798 15972
rect 19798 15943 19854 15952
rect 19708 15914 19760 15920
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19798 14920 19854 14929
rect 19720 14890 19798 14906
rect 19708 14884 19798 14890
rect 19760 14878 19798 14884
rect 19798 14855 19854 14864
rect 19708 14826 19760 14832
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19708 14476 19760 14482
rect 19708 14418 19760 14424
rect 19720 13938 19748 14418
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 20088 14006 20116 14214
rect 20076 14000 20128 14006
rect 20076 13942 20128 13948
rect 19708 13932 19760 13938
rect 19708 13874 19760 13880
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 20088 12782 20116 13942
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 20168 13184 20220 13190
rect 20168 13126 20220 13132
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19524 12436 19576 12442
rect 19524 12378 19576 12384
rect 20088 12238 20116 12718
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 20076 11824 20128 11830
rect 20076 11766 20128 11772
rect 19352 11614 19472 11642
rect 19524 11620 19576 11626
rect 19248 11280 19300 11286
rect 19248 11222 19300 11228
rect 19168 11104 19288 11132
rect 19064 10124 19116 10130
rect 19064 10066 19116 10072
rect 18972 9444 19024 9450
rect 18972 9386 19024 9392
rect 18984 9110 19012 9386
rect 18972 9104 19024 9110
rect 18972 9046 19024 9052
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18984 8294 19012 9046
rect 18972 8288 19024 8294
rect 18972 8230 19024 8236
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18340 7364 18460 7392
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 18064 6322 18092 6734
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 17960 6248 18012 6254
rect 17960 6190 18012 6196
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17592 5908 17644 5914
rect 17592 5850 17644 5856
rect 17696 4826 17724 6054
rect 18064 5896 18092 6258
rect 18340 6202 18368 7364
rect 18524 7274 18552 7686
rect 18420 7268 18472 7274
rect 18420 7210 18472 7216
rect 18512 7268 18564 7274
rect 18512 7210 18564 7216
rect 18432 6322 18460 7210
rect 18524 6662 18552 7210
rect 18984 6934 19012 8230
rect 18972 6928 19024 6934
rect 18972 6870 19024 6876
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 18524 6225 18552 6598
rect 18510 6216 18566 6225
rect 18340 6174 18460 6202
rect 18236 6112 18288 6118
rect 18236 6054 18288 6060
rect 18144 5908 18196 5914
rect 18064 5868 18144 5896
rect 18144 5850 18196 5856
rect 18248 5846 18276 6054
rect 17776 5840 17828 5846
rect 17776 5782 17828 5788
rect 18236 5840 18288 5846
rect 18236 5782 18288 5788
rect 17788 5370 17816 5782
rect 18248 5370 18276 5782
rect 17776 5364 17828 5370
rect 17776 5306 17828 5312
rect 18236 5364 18288 5370
rect 18236 5306 18288 5312
rect 17684 4820 17736 4826
rect 17684 4762 17736 4768
rect 17684 4684 17736 4690
rect 17684 4626 17736 4632
rect 17500 4480 17552 4486
rect 17500 4422 17552 4428
rect 17316 4276 17368 4282
rect 17316 4218 17368 4224
rect 17132 3596 17184 3602
rect 17132 3538 17184 3544
rect 17144 3194 17172 3538
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 16764 2576 16816 2582
rect 16764 2518 16816 2524
rect 16868 2378 16896 2586
rect 16856 2372 16908 2378
rect 16856 2314 16908 2320
rect 16670 82 16726 480
rect 16500 54 16726 82
rect 15842 0 15898 54
rect 16670 0 16726 54
rect 17406 82 17462 480
rect 17512 82 17540 4422
rect 17696 3398 17724 4626
rect 17684 3392 17736 3398
rect 17684 3334 17736 3340
rect 17696 1193 17724 3334
rect 18432 2514 18460 6174
rect 18510 6151 18566 6160
rect 19076 5114 19104 10066
rect 19156 9920 19208 9926
rect 19156 9862 19208 9868
rect 19168 8090 19196 9862
rect 19156 8084 19208 8090
rect 19156 8026 19208 8032
rect 19168 7410 19196 8026
rect 19260 7954 19288 11104
rect 19248 7948 19300 7954
rect 19248 7890 19300 7896
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19260 7274 19288 7890
rect 19248 7268 19300 7274
rect 19248 7210 19300 7216
rect 19260 7177 19288 7210
rect 19246 7168 19302 7177
rect 19246 7103 19302 7112
rect 19352 5914 19380 11614
rect 19524 11562 19576 11568
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19444 10266 19472 11494
rect 19536 11014 19564 11562
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 20088 11150 20116 11766
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 19524 11008 19576 11014
rect 19524 10950 19576 10956
rect 20088 10742 20116 11086
rect 20076 10736 20128 10742
rect 19982 10704 20038 10713
rect 20076 10678 20128 10684
rect 19982 10639 20038 10648
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19432 10260 19484 10266
rect 19432 10202 19484 10208
rect 19708 10124 19760 10130
rect 19708 10066 19760 10072
rect 19720 9722 19748 10066
rect 19708 9716 19760 9722
rect 19708 9658 19760 9664
rect 19996 9586 20024 10639
rect 19984 9580 20036 9586
rect 19984 9522 20036 9528
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19996 9178 20024 9522
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 19800 8900 19852 8906
rect 19800 8842 19852 8848
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 19444 8362 19472 8774
rect 19812 8498 19840 8842
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 19432 8356 19484 8362
rect 19432 8298 19484 8304
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19800 7948 19852 7954
rect 19800 7890 19852 7896
rect 19812 7546 19840 7890
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19444 6390 19472 6802
rect 19432 6384 19484 6390
rect 19432 6326 19484 6332
rect 19524 6316 19576 6322
rect 19524 6258 19576 6264
rect 19536 5914 19564 6258
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19340 5908 19392 5914
rect 19260 5868 19340 5896
rect 19260 5234 19288 5868
rect 19340 5850 19392 5856
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19996 5778 20024 7822
rect 19708 5772 19760 5778
rect 19708 5714 19760 5720
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19352 5302 19380 5510
rect 19720 5370 19748 5714
rect 19996 5370 20024 5714
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 19248 5228 19300 5234
rect 19248 5170 19300 5176
rect 18880 5092 18932 5098
rect 18800 5052 18880 5080
rect 18800 4486 18828 5052
rect 19076 5086 19288 5114
rect 18880 5034 18932 5040
rect 19156 4752 19208 4758
rect 19156 4694 19208 4700
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18604 3936 18656 3942
rect 18604 3878 18656 3884
rect 18616 3738 18644 3878
rect 18604 3732 18656 3738
rect 18604 3674 18656 3680
rect 18616 2854 18644 3674
rect 18800 3058 18828 4422
rect 19076 3738 19104 4558
rect 19064 3732 19116 3738
rect 19064 3674 19116 3680
rect 19076 3641 19104 3674
rect 19062 3632 19118 3641
rect 18972 3596 19024 3602
rect 19168 3602 19196 4694
rect 19062 3567 19118 3576
rect 19156 3596 19208 3602
rect 18972 3538 19024 3544
rect 19156 3538 19208 3544
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 18604 2848 18656 2854
rect 18604 2790 18656 2796
rect 18984 2650 19012 3538
rect 19064 3460 19116 3466
rect 19064 3402 19116 3408
rect 18972 2644 19024 2650
rect 18972 2586 19024 2592
rect 18420 2508 18472 2514
rect 18420 2450 18472 2456
rect 17682 1184 17738 1193
rect 17682 1119 17738 1128
rect 17406 54 17540 82
rect 18234 60 18290 480
rect 17406 0 17462 54
rect 18234 8 18236 60
rect 18288 8 18290 60
rect 18234 0 18290 8
rect 18970 82 19026 480
rect 19076 82 19104 3402
rect 19260 3194 19288 5086
rect 19432 5092 19484 5098
rect 19432 5034 19484 5040
rect 19444 4622 19472 5034
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 20180 4826 20208 13126
rect 20272 7818 20300 13806
rect 20456 9042 20484 18119
rect 21088 13796 21140 13802
rect 21088 13738 21140 13744
rect 21548 13796 21600 13802
rect 21548 13738 21600 13744
rect 20812 13524 20864 13530
rect 20812 13466 20864 13472
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20548 11014 20576 12582
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20640 11626 20668 12038
rect 20628 11620 20680 11626
rect 20628 11562 20680 11568
rect 20536 11008 20588 11014
rect 20536 10950 20588 10956
rect 20548 9994 20576 10950
rect 20640 10810 20668 11562
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 20628 10600 20680 10606
rect 20628 10542 20680 10548
rect 20536 9988 20588 9994
rect 20536 9930 20588 9936
rect 20536 9648 20588 9654
rect 20536 9590 20588 9596
rect 20548 9450 20576 9590
rect 20640 9586 20668 10542
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20536 9444 20588 9450
rect 20536 9386 20588 9392
rect 20444 9036 20496 9042
rect 20444 8978 20496 8984
rect 20640 8498 20668 9522
rect 20732 9178 20760 10066
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20260 7812 20312 7818
rect 20260 7754 20312 7760
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 20272 5914 20300 7346
rect 20444 7268 20496 7274
rect 20444 7210 20496 7216
rect 20456 6730 20484 7210
rect 20444 6724 20496 6730
rect 20444 6666 20496 6672
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 20272 5302 20300 5850
rect 20260 5296 20312 5302
rect 20260 5238 20312 5244
rect 20732 5098 20760 6054
rect 20720 5092 20772 5098
rect 20720 5034 20772 5040
rect 20732 4826 20760 5034
rect 19524 4820 19576 4826
rect 19524 4762 19576 4768
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19444 4146 19472 4558
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19338 3768 19394 3777
rect 19338 3703 19394 3712
rect 19352 3670 19380 3703
rect 19340 3664 19392 3670
rect 19340 3606 19392 3612
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19248 3188 19300 3194
rect 19248 3130 19300 3136
rect 19248 2984 19300 2990
rect 19352 2972 19380 3334
rect 19300 2944 19380 2972
rect 19248 2926 19300 2932
rect 19260 1329 19288 2926
rect 19444 2446 19472 4082
rect 19536 4049 19564 4762
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 19522 4040 19578 4049
rect 19522 3975 19578 3984
rect 20168 4004 20220 4010
rect 20168 3946 20220 3952
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 19536 3602 19564 3878
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 20180 3670 20208 3946
rect 20732 3738 20760 4558
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20168 3664 20220 3670
rect 20168 3606 20220 3612
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 20824 3534 20852 13466
rect 21100 12782 21128 13738
rect 21272 13388 21324 13394
rect 21272 13330 21324 13336
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 21100 12442 21128 12718
rect 21180 12708 21232 12714
rect 21180 12650 21232 12656
rect 21088 12436 21140 12442
rect 21088 12378 21140 12384
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20916 11898 20944 12242
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 21100 11218 21128 12378
rect 21192 11354 21220 12650
rect 21284 12646 21312 13330
rect 21364 12844 21416 12850
rect 21364 12786 21416 12792
rect 21272 12640 21324 12646
rect 21272 12582 21324 12588
rect 21376 12306 21404 12786
rect 21364 12300 21416 12306
rect 21364 12242 21416 12248
rect 21376 11898 21404 12242
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 21364 11620 21416 11626
rect 21364 11562 21416 11568
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21088 11212 21140 11218
rect 21088 11154 21140 11160
rect 20994 10704 21050 10713
rect 20994 10639 21050 10648
rect 20904 9036 20956 9042
rect 20904 8978 20956 8984
rect 20916 8634 20944 8978
rect 20904 8628 20956 8634
rect 20904 8570 20956 8576
rect 20904 7812 20956 7818
rect 20904 7754 20956 7760
rect 20916 5302 20944 7754
rect 21008 7478 21036 10639
rect 21100 10266 21128 11154
rect 21192 10674 21220 11290
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 21284 10810 21312 11154
rect 21376 11082 21404 11562
rect 21364 11076 21416 11082
rect 21364 11018 21416 11024
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 21180 10668 21232 10674
rect 21180 10610 21232 10616
rect 21088 10260 21140 10266
rect 21088 10202 21140 10208
rect 21180 8900 21232 8906
rect 21180 8842 21232 8848
rect 21192 8498 21220 8842
rect 21180 8492 21232 8498
rect 21180 8434 21232 8440
rect 21088 8084 21140 8090
rect 21088 8026 21140 8032
rect 20996 7472 21048 7478
rect 20996 7414 21048 7420
rect 21100 7206 21128 8026
rect 21180 8016 21232 8022
rect 21284 8004 21312 10746
rect 21456 10532 21508 10538
rect 21456 10474 21508 10480
rect 21468 10198 21496 10474
rect 21456 10192 21508 10198
rect 21456 10134 21508 10140
rect 21468 9722 21496 10134
rect 21456 9716 21508 9722
rect 21456 9658 21508 9664
rect 21468 9450 21496 9658
rect 21456 9444 21508 9450
rect 21456 9386 21508 9392
rect 21456 8832 21508 8838
rect 21456 8774 21508 8780
rect 21468 8362 21496 8774
rect 21456 8356 21508 8362
rect 21456 8298 21508 8304
rect 21232 7976 21312 8004
rect 21456 8016 21508 8022
rect 21180 7958 21232 7964
rect 21456 7958 21508 7964
rect 21180 7880 21232 7886
rect 21180 7822 21232 7828
rect 21088 7200 21140 7206
rect 21088 7142 21140 7148
rect 21100 5778 21128 7142
rect 21192 7002 21220 7822
rect 21468 7206 21496 7958
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 21468 7002 21496 7142
rect 21180 6996 21232 7002
rect 21180 6938 21232 6944
rect 21456 6996 21508 7002
rect 21456 6938 21508 6944
rect 21088 5772 21140 5778
rect 21088 5714 21140 5720
rect 20904 5296 20956 5302
rect 20904 5238 20956 5244
rect 20916 4554 20944 5238
rect 21192 5234 21220 6938
rect 21272 6112 21324 6118
rect 21272 6054 21324 6060
rect 21284 5914 21312 6054
rect 21272 5908 21324 5914
rect 21272 5850 21324 5856
rect 21180 5228 21232 5234
rect 21180 5170 21232 5176
rect 21284 5030 21312 5850
rect 21364 5704 21416 5710
rect 21364 5646 21416 5652
rect 21272 5024 21324 5030
rect 21272 4966 21324 4972
rect 21180 4752 21232 4758
rect 21180 4694 21232 4700
rect 20904 4548 20956 4554
rect 20904 4490 20956 4496
rect 21192 4282 21220 4694
rect 21180 4276 21232 4282
rect 21180 4218 21232 4224
rect 21284 3942 21312 4966
rect 21376 4622 21404 5646
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 21560 4154 21588 13738
rect 22284 13728 22336 13734
rect 22284 13670 22336 13676
rect 22468 13728 22520 13734
rect 22468 13670 22520 13676
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 22204 12646 22232 13262
rect 21732 12640 21784 12646
rect 21732 12582 21784 12588
rect 22192 12640 22244 12646
rect 22192 12582 22244 12588
rect 21640 12232 21692 12238
rect 21640 12174 21692 12180
rect 21652 9042 21680 12174
rect 21744 9586 21772 12582
rect 22204 12306 22232 12582
rect 22192 12300 22244 12306
rect 22192 12242 22244 12248
rect 22204 11694 22232 12242
rect 22192 11688 22244 11694
rect 22192 11630 22244 11636
rect 22008 11348 22060 11354
rect 22008 11290 22060 11296
rect 21824 11144 21876 11150
rect 21824 11086 21876 11092
rect 21732 9580 21784 9586
rect 21732 9522 21784 9528
rect 21744 9178 21772 9522
rect 21732 9172 21784 9178
rect 21732 9114 21784 9120
rect 21640 9036 21692 9042
rect 21640 8978 21692 8984
rect 21652 8634 21680 8978
rect 21640 8628 21692 8634
rect 21640 8570 21692 8576
rect 21640 7268 21692 7274
rect 21640 7210 21692 7216
rect 21468 4126 21588 4154
rect 21272 3936 21324 3942
rect 21272 3878 21324 3884
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 20824 3194 20852 3470
rect 21272 3392 21324 3398
rect 21272 3334 21324 3340
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 19524 3120 19576 3126
rect 19524 3062 19576 3068
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19246 1320 19302 1329
rect 19246 1255 19302 1264
rect 18970 54 19104 82
rect 19536 82 19564 3062
rect 21284 2990 21312 3334
rect 21272 2984 21324 2990
rect 21272 2926 21324 2932
rect 19984 2848 20036 2854
rect 19984 2790 20036 2796
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19996 2582 20024 2790
rect 19984 2576 20036 2582
rect 19984 2518 20036 2524
rect 20168 2372 20220 2378
rect 20168 2314 20220 2320
rect 20180 2009 20208 2314
rect 20260 2304 20312 2310
rect 20260 2246 20312 2252
rect 20166 2000 20222 2009
rect 20166 1935 20222 1944
rect 19798 82 19854 480
rect 19536 54 19854 82
rect 20272 82 20300 2246
rect 21284 1873 21312 2926
rect 21270 1864 21326 1873
rect 21270 1799 21326 1808
rect 20534 82 20590 480
rect 20272 54 20590 82
rect 18970 0 19026 54
rect 19798 0 19854 54
rect 20534 0 20590 54
rect 21362 82 21418 480
rect 21468 82 21496 4126
rect 21652 2650 21680 7210
rect 21732 7200 21784 7206
rect 21732 7142 21784 7148
rect 21744 6186 21772 7142
rect 21836 6866 21864 11086
rect 21824 6860 21876 6866
rect 21824 6802 21876 6808
rect 21732 6180 21784 6186
rect 21732 6122 21784 6128
rect 21836 5914 21864 6802
rect 21824 5908 21876 5914
rect 21824 5850 21876 5856
rect 21824 5772 21876 5778
rect 21824 5714 21876 5720
rect 21836 5370 21864 5714
rect 21824 5364 21876 5370
rect 21824 5306 21876 5312
rect 21836 5030 21864 5306
rect 21824 5024 21876 5030
rect 21824 4966 21876 4972
rect 22020 4690 22048 11290
rect 22192 9444 22244 9450
rect 22192 9386 22244 9392
rect 22204 9178 22232 9386
rect 22192 9172 22244 9178
rect 22192 9114 22244 9120
rect 22204 8430 22232 9114
rect 22192 8424 22244 8430
rect 22192 8366 22244 8372
rect 22100 7744 22152 7750
rect 22100 7686 22152 7692
rect 22112 7274 22140 7686
rect 22100 7268 22152 7274
rect 22100 7210 22152 7216
rect 22100 6928 22152 6934
rect 22100 6870 22152 6876
rect 22112 6118 22140 6870
rect 22192 6316 22244 6322
rect 22192 6258 22244 6264
rect 22100 6112 22152 6118
rect 22100 6054 22152 6060
rect 22112 5778 22140 6054
rect 22204 5914 22232 6258
rect 22192 5908 22244 5914
rect 22192 5850 22244 5856
rect 22100 5772 22152 5778
rect 22100 5714 22152 5720
rect 22100 5092 22152 5098
rect 22100 5034 22152 5040
rect 22112 4826 22140 5034
rect 22100 4820 22152 4826
rect 22100 4762 22152 4768
rect 22008 4684 22060 4690
rect 22008 4626 22060 4632
rect 22192 4684 22244 4690
rect 22192 4626 22244 4632
rect 22204 4146 22232 4626
rect 22192 4140 22244 4146
rect 22192 4082 22244 4088
rect 22100 3936 22152 3942
rect 22100 3878 22152 3884
rect 22112 3738 22140 3878
rect 22100 3732 22152 3738
rect 22100 3674 22152 3680
rect 22008 3052 22060 3058
rect 22008 2994 22060 3000
rect 21640 2644 21692 2650
rect 21640 2586 21692 2592
rect 22020 2582 22048 2994
rect 22112 2922 22140 3674
rect 22100 2916 22152 2922
rect 22100 2858 22152 2864
rect 22296 2582 22324 13670
rect 22374 9344 22430 9353
rect 22374 9279 22430 9288
rect 22008 2576 22060 2582
rect 22008 2518 22060 2524
rect 22284 2576 22336 2582
rect 22284 2518 22336 2524
rect 22296 2446 22324 2518
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 21362 54 21496 82
rect 22098 82 22154 480
rect 22388 82 22416 9279
rect 22480 3466 22508 13670
rect 22664 13530 22692 23530
rect 23860 23526 23888 23734
rect 22744 23520 22796 23526
rect 22744 23462 22796 23468
rect 23848 23520 23900 23526
rect 23848 23462 23900 23468
rect 22756 20505 22784 23462
rect 24032 23180 24084 23186
rect 24032 23122 24084 23128
rect 24044 22438 24072 23122
rect 24032 22432 24084 22438
rect 24032 22374 24084 22380
rect 24044 21049 24072 22374
rect 24030 21040 24086 21049
rect 24030 20975 24086 20984
rect 22742 20496 22798 20505
rect 22742 20431 22798 20440
rect 22756 17542 22784 20431
rect 23478 18728 23534 18737
rect 23478 18663 23534 18672
rect 23492 17785 23520 18663
rect 23478 17776 23534 17785
rect 23478 17711 23534 17720
rect 22744 17536 22796 17542
rect 22744 17478 22796 17484
rect 23940 17536 23992 17542
rect 23940 17478 23992 17484
rect 22744 14000 22796 14006
rect 22744 13942 22796 13948
rect 22652 13524 22704 13530
rect 22652 13466 22704 13472
rect 22560 12436 22612 12442
rect 22560 12378 22612 12384
rect 22572 10130 22600 12378
rect 22756 11370 22784 13942
rect 23388 13796 23440 13802
rect 23388 13738 23440 13744
rect 22836 13388 22888 13394
rect 22836 13330 22888 13336
rect 22848 12646 22876 13330
rect 22836 12640 22888 12646
rect 22836 12582 22888 12588
rect 22848 11665 22876 12582
rect 22928 12300 22980 12306
rect 22928 12242 22980 12248
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 22940 11898 22968 12242
rect 22928 11892 22980 11898
rect 22928 11834 22980 11840
rect 22834 11656 22890 11665
rect 22834 11591 22890 11600
rect 22664 11342 22784 11370
rect 22560 10124 22612 10130
rect 22560 10066 22612 10072
rect 22560 6112 22612 6118
rect 22560 6054 22612 6060
rect 22572 4758 22600 6054
rect 22560 4752 22612 4758
rect 22560 4694 22612 4700
rect 22468 3460 22520 3466
rect 22468 3402 22520 3408
rect 22468 3052 22520 3058
rect 22468 2994 22520 3000
rect 22480 2582 22508 2994
rect 22468 2576 22520 2582
rect 22468 2518 22520 2524
rect 22664 2310 22692 11342
rect 22744 11280 22796 11286
rect 22744 11222 22796 11228
rect 22756 10810 22784 11222
rect 22928 11144 22980 11150
rect 22928 11086 22980 11092
rect 22744 10804 22796 10810
rect 22744 10746 22796 10752
rect 22940 10606 22968 11086
rect 23032 10742 23060 12242
rect 23296 11688 23348 11694
rect 23296 11630 23348 11636
rect 23308 11286 23336 11630
rect 23296 11280 23348 11286
rect 23296 11222 23348 11228
rect 23020 10736 23072 10742
rect 23020 10678 23072 10684
rect 22928 10600 22980 10606
rect 22928 10542 22980 10548
rect 22940 9994 22968 10542
rect 23112 10532 23164 10538
rect 23112 10474 23164 10480
rect 22928 9988 22980 9994
rect 22928 9930 22980 9936
rect 23124 9654 23152 10474
rect 23296 10260 23348 10266
rect 23296 10202 23348 10208
rect 23204 9920 23256 9926
rect 23204 9862 23256 9868
rect 23112 9648 23164 9654
rect 23112 9590 23164 9596
rect 23124 8514 23152 9590
rect 23216 9586 23244 9862
rect 23204 9580 23256 9586
rect 23204 9522 23256 9528
rect 23308 9110 23336 10202
rect 23400 9926 23428 13738
rect 23756 13728 23808 13734
rect 23756 13670 23808 13676
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 23388 9920 23440 9926
rect 23388 9862 23440 9868
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 23296 9104 23348 9110
rect 23296 9046 23348 9052
rect 23492 8634 23520 9114
rect 23480 8628 23532 8634
rect 23480 8570 23532 8576
rect 23124 8486 23520 8514
rect 23492 8022 23520 8486
rect 23388 8016 23440 8022
rect 23388 7958 23440 7964
rect 23480 8016 23532 8022
rect 23480 7958 23532 7964
rect 23112 7880 23164 7886
rect 23112 7822 23164 7828
rect 22744 7744 22796 7750
rect 22744 7686 22796 7692
rect 22756 7274 22784 7686
rect 22744 7268 22796 7274
rect 22744 7210 22796 7216
rect 22756 5710 22784 7210
rect 23124 7206 23152 7822
rect 23400 7546 23428 7958
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 23112 7200 23164 7206
rect 23112 7142 23164 7148
rect 23124 5914 23152 7142
rect 23480 6996 23532 7002
rect 23480 6938 23532 6944
rect 23204 6792 23256 6798
rect 23204 6734 23256 6740
rect 23216 6118 23244 6734
rect 23492 6390 23520 6938
rect 23584 6390 23612 12038
rect 23664 9920 23716 9926
rect 23664 9862 23716 9868
rect 23676 8514 23704 9862
rect 23768 9110 23796 13670
rect 23848 11008 23900 11014
rect 23848 10950 23900 10956
rect 23860 10674 23888 10950
rect 23848 10668 23900 10674
rect 23848 10610 23900 10616
rect 23860 9722 23888 10610
rect 23952 10538 23980 17478
rect 24032 16040 24084 16046
rect 24032 15982 24084 15988
rect 24044 14929 24072 15982
rect 24030 14920 24086 14929
rect 24030 14855 24086 14864
rect 24032 13184 24084 13190
rect 24032 13126 24084 13132
rect 24044 12209 24072 13126
rect 24030 12200 24086 12209
rect 24030 12135 24086 12144
rect 24136 11898 24164 24686
rect 24780 24410 24808 25327
rect 24768 24404 24820 24410
rect 24768 24346 24820 24352
rect 24676 24268 24728 24274
rect 24676 24210 24728 24216
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24688 23594 24716 24210
rect 24766 24168 24822 24177
rect 24766 24103 24822 24112
rect 24676 23588 24728 23594
rect 24676 23530 24728 23536
rect 24780 23322 24808 24103
rect 24964 23866 24992 26687
rect 25608 24138 25636 27520
rect 27172 24954 27200 27520
rect 27160 24948 27212 24954
rect 27160 24890 27212 24896
rect 25596 24132 25648 24138
rect 25596 24074 25648 24080
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 24768 23316 24820 23322
rect 24768 23258 24820 23264
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24766 22672 24822 22681
rect 24766 22607 24822 22616
rect 24780 22234 24808 22607
rect 24768 22228 24820 22234
rect 24768 22170 24820 22176
rect 24216 22092 24268 22098
rect 24216 22034 24268 22040
rect 24228 21350 24256 22034
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24216 21344 24268 21350
rect 24216 21286 24268 21292
rect 24766 21312 24822 21321
rect 24228 20369 24256 21286
rect 24766 21247 24822 21256
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24214 20360 24270 20369
rect 24214 20295 24270 20304
rect 24676 19916 24728 19922
rect 24676 19858 24728 19864
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24688 19378 24716 19858
rect 24676 19372 24728 19378
rect 24676 19314 24728 19320
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24216 17128 24268 17134
rect 24216 17070 24268 17076
rect 24228 16017 24256 17070
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24780 16250 24808 21247
rect 25226 20224 25282 20233
rect 25226 20159 25282 20168
rect 25240 20058 25268 20159
rect 25228 20052 25280 20058
rect 25228 19994 25280 20000
rect 25410 17504 25466 17513
rect 25410 17439 25466 17448
rect 25424 17338 25452 17439
rect 25412 17332 25464 17338
rect 25412 17274 25464 17280
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 24214 16008 24270 16017
rect 24214 15943 24270 15952
rect 24766 16008 24822 16017
rect 24766 15943 24822 15952
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24780 14618 24808 15943
rect 24768 14612 24820 14618
rect 24768 14554 24820 14560
rect 24676 14476 24728 14482
rect 24676 14418 24728 14424
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24688 14074 24716 14418
rect 24676 14068 24728 14074
rect 24676 14010 24728 14016
rect 27620 14068 27672 14074
rect 27620 14010 27672 14016
rect 27632 13977 27660 14010
rect 27618 13968 27674 13977
rect 27618 13903 27674 13912
rect 25688 13796 25740 13802
rect 25688 13738 25740 13744
rect 24216 13388 24268 13394
rect 24216 13330 24268 13336
rect 25228 13388 25280 13394
rect 25228 13330 25280 13336
rect 24228 12646 24256 13330
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 25240 12850 25268 13330
rect 25228 12844 25280 12850
rect 25228 12786 25280 12792
rect 25320 12708 25372 12714
rect 25320 12650 25372 12656
rect 24216 12640 24268 12646
rect 24216 12582 24268 12588
rect 25136 12640 25188 12646
rect 25136 12582 25188 12588
rect 24676 12368 24728 12374
rect 24676 12310 24728 12316
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24688 11898 24716 12310
rect 24768 12096 24820 12102
rect 24768 12038 24820 12044
rect 24124 11892 24176 11898
rect 24124 11834 24176 11840
rect 24676 11892 24728 11898
rect 24676 11834 24728 11840
rect 24124 11688 24176 11694
rect 24124 11630 24176 11636
rect 24032 10668 24084 10674
rect 24032 10610 24084 10616
rect 23940 10532 23992 10538
rect 23940 10474 23992 10480
rect 24044 10062 24072 10610
rect 24136 10198 24164 11630
rect 24216 11212 24268 11218
rect 24216 11154 24268 11160
rect 24228 10266 24256 11154
rect 24676 11144 24728 11150
rect 24676 11086 24728 11092
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24688 10810 24716 11086
rect 24676 10804 24728 10810
rect 24676 10746 24728 10752
rect 24676 10532 24728 10538
rect 24676 10474 24728 10480
rect 24216 10260 24268 10266
rect 24216 10202 24268 10208
rect 24124 10192 24176 10198
rect 24124 10134 24176 10140
rect 24032 10056 24084 10062
rect 24032 9998 24084 10004
rect 23848 9716 23900 9722
rect 23848 9658 23900 9664
rect 23940 9580 23992 9586
rect 23940 9522 23992 9528
rect 23756 9104 23808 9110
rect 23756 9046 23808 9052
rect 23768 8634 23796 9046
rect 23952 8634 23980 9522
rect 24044 8974 24072 9998
rect 24136 9586 24164 10134
rect 24216 10124 24268 10130
rect 24216 10066 24268 10072
rect 24124 9580 24176 9586
rect 24124 9522 24176 9528
rect 24032 8968 24084 8974
rect 24032 8910 24084 8916
rect 23756 8628 23808 8634
rect 23756 8570 23808 8576
rect 23940 8628 23992 8634
rect 23940 8570 23992 8576
rect 24044 8566 24072 8910
rect 24032 8560 24084 8566
rect 23676 8486 23796 8514
rect 24032 8502 24084 8508
rect 23664 8356 23716 8362
rect 23664 8298 23716 8304
rect 23676 8090 23704 8298
rect 23664 8084 23716 8090
rect 23664 8026 23716 8032
rect 23676 7206 23704 8026
rect 23664 7200 23716 7206
rect 23664 7142 23716 7148
rect 23768 7018 23796 8486
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 24136 7546 24164 7686
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 23676 6990 23796 7018
rect 23480 6384 23532 6390
rect 23480 6326 23532 6332
rect 23572 6384 23624 6390
rect 23572 6326 23624 6332
rect 23584 6186 23612 6326
rect 23572 6180 23624 6186
rect 23572 6122 23624 6128
rect 23204 6112 23256 6118
rect 23204 6054 23256 6060
rect 23112 5908 23164 5914
rect 23112 5850 23164 5856
rect 22744 5704 22796 5710
rect 22744 5646 22796 5652
rect 23216 5370 23244 6054
rect 23572 5568 23624 5574
rect 23572 5510 23624 5516
rect 23204 5364 23256 5370
rect 23204 5306 23256 5312
rect 23388 5024 23440 5030
rect 23388 4966 23440 4972
rect 22836 4752 22888 4758
rect 22836 4694 22888 4700
rect 22848 4282 22876 4694
rect 23020 4616 23072 4622
rect 23020 4558 23072 4564
rect 22928 4548 22980 4554
rect 22928 4490 22980 4496
rect 22836 4276 22888 4282
rect 22836 4218 22888 4224
rect 22940 4214 22968 4490
rect 22928 4208 22980 4214
rect 22928 4150 22980 4156
rect 22940 3942 22968 4150
rect 22928 3936 22980 3942
rect 22928 3878 22980 3884
rect 22940 2582 22968 3878
rect 22928 2576 22980 2582
rect 22928 2518 22980 2524
rect 23032 2378 23060 4558
rect 23400 3738 23428 4966
rect 23584 4826 23612 5510
rect 23572 4820 23624 4826
rect 23572 4762 23624 4768
rect 23676 4154 23704 6990
rect 23848 6928 23900 6934
rect 23848 6870 23900 6876
rect 23860 6458 23888 6870
rect 24032 6792 24084 6798
rect 24032 6734 24084 6740
rect 23848 6452 23900 6458
rect 23848 6394 23900 6400
rect 24044 6322 24072 6734
rect 23848 6316 23900 6322
rect 23848 6258 23900 6264
rect 24032 6316 24084 6322
rect 24032 6258 24084 6264
rect 23754 6216 23810 6225
rect 23754 6151 23810 6160
rect 23768 6118 23796 6151
rect 23756 6112 23808 6118
rect 23756 6054 23808 6060
rect 23768 5914 23796 6054
rect 23756 5908 23808 5914
rect 23756 5850 23808 5856
rect 23860 5234 23888 6258
rect 24228 5846 24256 10066
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24688 9518 24716 10474
rect 24676 9512 24728 9518
rect 24676 9454 24728 9460
rect 24676 9172 24728 9178
rect 24676 9114 24728 9120
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24688 8362 24716 9114
rect 24676 8356 24728 8362
rect 24676 8298 24728 8304
rect 24676 8016 24728 8022
rect 24676 7958 24728 7964
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24688 7478 24716 7958
rect 24676 7472 24728 7478
rect 24676 7414 24728 7420
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24216 5840 24268 5846
rect 24216 5782 24268 5788
rect 24676 5840 24728 5846
rect 24676 5782 24728 5788
rect 23848 5228 23900 5234
rect 23848 5170 23900 5176
rect 23940 5228 23992 5234
rect 23940 5170 23992 5176
rect 23756 5092 23808 5098
rect 23756 5034 23808 5040
rect 23768 4554 23796 5034
rect 23952 4622 23980 5170
rect 24228 4826 24256 5782
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24688 5302 24716 5782
rect 24676 5296 24728 5302
rect 24676 5238 24728 5244
rect 24216 4820 24268 4826
rect 24216 4762 24268 4768
rect 24032 4752 24084 4758
rect 24032 4694 24084 4700
rect 23940 4616 23992 4622
rect 23940 4558 23992 4564
rect 23756 4548 23808 4554
rect 23756 4490 23808 4496
rect 23676 4126 23980 4154
rect 23756 4004 23808 4010
rect 23756 3946 23808 3952
rect 23388 3732 23440 3738
rect 23388 3674 23440 3680
rect 23768 3670 23796 3946
rect 23756 3664 23808 3670
rect 23676 3624 23756 3652
rect 23676 2582 23704 3624
rect 23756 3606 23808 3612
rect 23756 3528 23808 3534
rect 23756 3470 23808 3476
rect 23848 3528 23900 3534
rect 23848 3470 23900 3476
rect 23768 3194 23796 3470
rect 23756 3188 23808 3194
rect 23756 3130 23808 3136
rect 23860 3058 23888 3470
rect 23848 3052 23900 3058
rect 23848 2994 23900 3000
rect 23664 2576 23716 2582
rect 23664 2518 23716 2524
rect 23020 2372 23072 2378
rect 23020 2314 23072 2320
rect 22652 2304 22704 2310
rect 22652 2246 22704 2252
rect 22926 1048 22982 1057
rect 22926 983 22982 992
rect 22098 54 22416 82
rect 22834 82 22890 480
rect 22940 82 22968 983
rect 22834 54 22968 82
rect 23662 82 23718 480
rect 23952 82 23980 4126
rect 24044 3942 24072 4694
rect 24216 4548 24268 4554
rect 24216 4490 24268 4496
rect 24032 3936 24084 3942
rect 24032 3878 24084 3884
rect 24044 2582 24072 3878
rect 24228 3670 24256 4490
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24780 4154 24808 12038
rect 24952 11552 25004 11558
rect 24952 11494 25004 11500
rect 24860 10600 24912 10606
rect 24860 10542 24912 10548
rect 24872 9353 24900 10542
rect 24964 10198 24992 11494
rect 24952 10192 25004 10198
rect 24952 10134 25004 10140
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 24858 9344 24914 9353
rect 24858 9279 24914 9288
rect 24964 8906 24992 9998
rect 24952 8900 25004 8906
rect 24952 8842 25004 8848
rect 24952 8560 25004 8566
rect 24952 8502 25004 8508
rect 24964 8022 24992 8502
rect 24952 8016 25004 8022
rect 24952 7958 25004 7964
rect 24964 7410 24992 7958
rect 25044 7880 25096 7886
rect 25044 7822 25096 7828
rect 25056 7478 25084 7822
rect 25044 7472 25096 7478
rect 25044 7414 25096 7420
rect 24952 7404 25004 7410
rect 24952 7346 25004 7352
rect 25056 6458 25084 7414
rect 25044 6452 25096 6458
rect 25044 6394 25096 6400
rect 25148 6338 25176 12582
rect 25228 10192 25280 10198
rect 25228 10134 25280 10140
rect 25240 9654 25268 10134
rect 25228 9648 25280 9654
rect 25228 9590 25280 9596
rect 25240 9178 25268 9590
rect 25228 9172 25280 9178
rect 25228 9114 25280 9120
rect 25332 9058 25360 12650
rect 25504 12640 25556 12646
rect 25504 12582 25556 12588
rect 25516 9353 25544 12582
rect 25596 10464 25648 10470
rect 25596 10406 25648 10412
rect 25502 9344 25558 9353
rect 25502 9279 25558 9288
rect 24964 6310 25176 6338
rect 25240 9030 25360 9058
rect 25516 9042 25544 9279
rect 25504 9036 25556 9042
rect 24860 4616 24912 4622
rect 24860 4558 24912 4564
rect 24872 4214 24900 4558
rect 24504 4126 24808 4154
rect 24860 4208 24912 4214
rect 24860 4150 24912 4156
rect 24504 4010 24532 4126
rect 24492 4004 24544 4010
rect 24492 3946 24544 3952
rect 24504 3738 24532 3946
rect 24492 3732 24544 3738
rect 24492 3674 24544 3680
rect 24216 3664 24268 3670
rect 24216 3606 24268 3612
rect 24228 3058 24256 3606
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24216 3052 24268 3058
rect 24268 3012 24348 3040
rect 24216 2994 24268 3000
rect 24216 2644 24268 2650
rect 24216 2586 24268 2592
rect 24032 2576 24084 2582
rect 24032 2518 24084 2524
rect 23662 54 23980 82
rect 24228 82 24256 2586
rect 24320 2378 24348 3012
rect 24308 2372 24360 2378
rect 24308 2314 24360 2320
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24398 82 24454 480
rect 24228 54 24454 82
rect 24964 82 24992 6310
rect 25240 4554 25268 9030
rect 25504 8978 25556 8984
rect 25320 8900 25372 8906
rect 25320 8842 25372 8848
rect 25228 4548 25280 4554
rect 25228 4490 25280 4496
rect 25240 4282 25268 4490
rect 25228 4276 25280 4282
rect 25228 4218 25280 4224
rect 25332 4154 25360 8842
rect 25412 8832 25464 8838
rect 25412 8774 25464 8780
rect 25424 8498 25452 8774
rect 25516 8634 25544 8978
rect 25504 8628 25556 8634
rect 25504 8570 25556 8576
rect 25412 8492 25464 8498
rect 25412 8434 25464 8440
rect 25608 7970 25636 10406
rect 25516 7942 25636 7970
rect 25516 5574 25544 7942
rect 25594 7848 25650 7857
rect 25594 7783 25650 7792
rect 25504 5568 25556 5574
rect 25504 5510 25556 5516
rect 25608 5370 25636 7783
rect 25596 5364 25648 5370
rect 25596 5306 25648 5312
rect 25608 5166 25636 5306
rect 25596 5160 25648 5166
rect 25596 5102 25648 5108
rect 25148 4126 25360 4154
rect 25148 3194 25176 4126
rect 25136 3188 25188 3194
rect 25136 3130 25188 3136
rect 25226 82 25282 480
rect 24964 54 25282 82
rect 25700 82 25728 13738
rect 25964 12912 26016 12918
rect 25964 12854 26016 12860
rect 25872 12300 25924 12306
rect 25872 12242 25924 12248
rect 25884 11558 25912 12242
rect 25872 11552 25924 11558
rect 25872 11494 25924 11500
rect 25780 6860 25832 6866
rect 25780 6802 25832 6808
rect 25792 6118 25820 6802
rect 25884 6458 25912 11494
rect 25976 7206 26004 12854
rect 26332 12844 26384 12850
rect 26332 12786 26384 12792
rect 26148 11620 26200 11626
rect 26148 11562 26200 11568
rect 25964 7200 26016 7206
rect 25964 7142 26016 7148
rect 25872 6452 25924 6458
rect 25872 6394 25924 6400
rect 25884 6254 25912 6394
rect 25872 6248 25924 6254
rect 25870 6216 25872 6225
rect 25924 6216 25926 6225
rect 25870 6151 25926 6160
rect 25780 6112 25832 6118
rect 25780 6054 25832 6060
rect 25792 5137 25820 6054
rect 25778 5128 25834 5137
rect 25778 5063 25834 5072
rect 25976 4154 26004 7142
rect 25884 4126 26004 4154
rect 25780 2848 25832 2854
rect 25780 2790 25832 2796
rect 25792 1193 25820 2790
rect 25884 2145 25912 4126
rect 25870 2136 25926 2145
rect 25870 2071 25926 2080
rect 25778 1184 25834 1193
rect 25778 1119 25834 1128
rect 25962 82 26018 480
rect 26160 134 26188 11562
rect 26344 4154 26372 12786
rect 27618 12608 27674 12617
rect 27618 12543 27674 12552
rect 27632 12374 27660 12543
rect 27620 12368 27672 12374
rect 27620 12310 27672 12316
rect 26252 4126 26372 4154
rect 25700 54 26018 82
rect 26148 128 26200 134
rect 26148 70 26200 76
rect 26252 66 26280 4126
rect 26790 128 26846 480
rect 26790 76 26792 128
rect 26844 76 26846 128
rect 21362 0 21418 54
rect 22098 0 22154 54
rect 22834 0 22890 54
rect 23662 0 23718 54
rect 24398 0 24454 54
rect 25226 0 25282 54
rect 25962 0 26018 54
rect 26240 60 26292 66
rect 26240 2 26292 8
rect 26790 0 26846 76
rect 27526 60 27582 480
rect 27526 8 27528 60
rect 27580 8 27582 60
rect 27526 0 27582 8
<< via2 >>
rect 1858 25608 1914 25664
rect 1582 18536 1638 18592
rect 110 12144 166 12200
rect 1858 15136 1914 15192
rect 110 8608 166 8664
rect 1674 8336 1730 8392
rect 110 5072 166 5128
rect 4894 22072 4950 22128
rect 3790 21528 3846 21584
rect 2778 17720 2834 17776
rect 3054 17720 3110 17776
rect 3606 13504 3662 13560
rect 2226 1944 2282 2000
rect 2502 992 2558 1048
rect 3054 2760 3110 2816
rect 3146 2488 3202 2544
rect 3054 2352 3110 2408
rect 3514 1672 3570 1728
rect 3330 1536 3386 1592
rect 3790 3032 3846 3088
rect 3882 2216 3938 2272
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5170 13232 5226 13288
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 6182 12688 6238 12744
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5998 10648 6054 10704
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 4710 7384 4766 7440
rect 4802 5072 4858 5128
rect 5262 5208 5318 5264
rect 4986 4664 5042 4720
rect 4894 4528 4950 4584
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 7470 18128 7526 18184
rect 8114 17584 8170 17640
rect 10046 27512 10102 27568
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10046 20304 10102 20360
rect 10230 20440 10286 20496
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 6918 13504 6974 13560
rect 6826 10512 6882 10568
rect 6458 10104 6514 10160
rect 6734 9832 6790 9888
rect 6550 9716 6606 9752
rect 6550 9696 6552 9716
rect 6552 9696 6604 9716
rect 6604 9696 6606 9716
rect 6182 5208 6238 5264
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 4526 1400 4582 1456
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 5998 1264 6054 1320
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 8850 13676 8852 13696
rect 8852 13676 8904 13696
rect 8904 13676 8906 13696
rect 8850 13640 8906 13676
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 9954 13504 10010 13560
rect 9770 13096 9826 13152
rect 7102 9832 7158 9888
rect 7286 7928 7342 7984
rect 7838 7656 7894 7712
rect 6366 3712 6422 3768
rect 6274 1808 6330 1864
rect 6918 1128 6974 1184
rect 8850 7928 8906 7984
rect 8390 6840 8446 6896
rect 7654 3984 7710 4040
rect 8666 3440 8722 3496
rect 9494 4664 9550 4720
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10690 4664 10746 4720
rect 10138 4528 10194 4584
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 11426 7928 11482 7984
rect 11334 7112 11390 7168
rect 13634 17720 13690 17776
rect 14094 17720 14150 17776
rect 13174 11600 13230 11656
rect 12898 9696 12954 9752
rect 12070 6840 12126 6896
rect 11426 4528 11482 4584
rect 13174 8336 13230 8392
rect 13358 7284 13360 7304
rect 13360 7284 13412 7304
rect 13412 7284 13414 7304
rect 13358 7248 13414 7284
rect 14094 9832 14150 9888
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 24950 26696 25006 26752
rect 24766 25336 24822 25392
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 15290 21528 15346 21584
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 15382 17584 15438 17640
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 15382 13368 15438 13424
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14646 10512 14702 10568
rect 14186 9696 14242 9752
rect 12714 2896 12770 2952
rect 13266 4528 13322 4584
rect 14646 7656 14702 7712
rect 14554 7248 14610 7304
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 15290 10104 15346 10160
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 18602 20984 18658 21040
rect 17222 18128 17278 18184
rect 16670 13232 16726 13288
rect 16486 12688 16542 12744
rect 15934 12144 15990 12200
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 15842 7420 15844 7440
rect 15844 7420 15896 7440
rect 15896 7420 15898 7440
rect 15842 7384 15898 7420
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 13450 3984 13506 4040
rect 14370 4120 14426 4176
rect 13174 2896 13230 2952
rect 12898 2488 12954 2544
rect 13174 1672 13230 1728
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15014 3440 15070 3496
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14830 2352 14886 2408
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 17038 6840 17094 6896
rect 16118 5072 16174 5128
rect 17130 5208 17186 5264
rect 16486 4120 16542 4176
rect 16026 2760 16082 2816
rect 15658 1536 15714 1592
rect 16854 3984 16910 4040
rect 17682 7792 17738 7848
rect 18694 14320 18750 14376
rect 19062 12824 19118 12880
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 20442 18128 20498 18184
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19798 15952 19854 16008
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19798 14864 19854 14920
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 18510 6160 18566 6216
rect 19246 7112 19302 7168
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19982 10648 20038 10704
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19062 3576 19118 3632
rect 17682 1128 17738 1184
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19338 3712 19394 3768
rect 19522 3984 19578 4040
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 20994 10648 21050 10704
rect 19246 1264 19302 1320
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20166 1944 20222 2000
rect 21270 1808 21326 1864
rect 22374 9288 22430 9344
rect 24030 20984 24086 21040
rect 22742 20440 22798 20496
rect 23478 18672 23534 18728
rect 23478 17720 23534 17776
rect 22834 11600 22890 11656
rect 24030 14864 24086 14920
rect 24030 12144 24086 12200
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24766 24112 24822 24168
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24766 22616 24822 22672
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24766 21256 24822 21312
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24214 20304 24270 20360
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 25226 20168 25282 20224
rect 25410 17448 25466 17504
rect 24214 15952 24270 16008
rect 24766 15952 24822 16008
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 27618 13912 27674 13968
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 23754 6160 23810 6216
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 22926 992 22982 1048
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24858 9288 24914 9344
rect 25502 9288 25558 9344
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 25594 7792 25650 7848
rect 25870 6196 25872 6216
rect 25872 6196 25924 6216
rect 25924 6196 25926 6216
rect 25870 6160 25926 6196
rect 25778 5072 25834 5128
rect 25870 2080 25926 2136
rect 25778 1128 25834 1184
rect 27618 12552 27674 12608
<< metal3 >>
rect 9806 27508 9812 27572
rect 9876 27570 9882 27572
rect 10041 27570 10107 27573
rect 9876 27568 10107 27570
rect 9876 27512 10046 27568
rect 10102 27512 10107 27568
rect 9876 27510 10107 27512
rect 9876 27508 9882 27510
rect 10041 27507 10107 27510
rect 27520 27208 28000 27328
rect 24945 26754 25011 26757
rect 27662 26754 27722 27208
rect 24945 26752 27722 26754
rect 24945 26696 24950 26752
rect 25006 26696 27722 26752
rect 24945 26694 27722 26696
rect 24945 26691 25011 26694
rect 0 26120 480 26240
rect 62 25666 122 26120
rect 27520 25848 28000 25968
rect 1853 25666 1919 25669
rect 62 25664 1919 25666
rect 62 25608 1858 25664
rect 1914 25608 1919 25664
rect 62 25606 1919 25608
rect 1853 25603 1919 25606
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 24761 25394 24827 25397
rect 27662 25394 27722 25848
rect 24761 25392 27722 25394
rect 24761 25336 24766 25392
rect 24822 25336 27722 25392
rect 24761 25334 27722 25336
rect 24761 25331 24827 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 27520 24488 28000 24608
rect 19610 24447 19930 24448
rect 24761 24170 24827 24173
rect 27662 24170 27722 24488
rect 24761 24168 27722 24170
rect 24761 24112 24766 24168
rect 24822 24112 27722 24168
rect 24761 24110 27722 24112
rect 24761 24107 24827 24110
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 27520 23128 28000 23248
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 0 22584 480 22704
rect 24761 22674 24827 22677
rect 27662 22674 27722 23128
rect 24761 22672 27722 22674
rect 24761 22616 24766 22672
rect 24822 22616 27722 22672
rect 24761 22614 27722 22616
rect 24761 22611 24827 22614
rect 62 22130 122 22584
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 4889 22130 4955 22133
rect 62 22128 4955 22130
rect 62 22072 4894 22128
rect 4950 22072 4955 22128
rect 62 22070 4955 22072
rect 4889 22067 4955 22070
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 27520 21768 28000 21888
rect 24277 21727 24597 21728
rect 3785 21586 3851 21589
rect 15285 21586 15351 21589
rect 3785 21584 15351 21586
rect 3785 21528 3790 21584
rect 3846 21528 15290 21584
rect 15346 21528 15351 21584
rect 3785 21526 15351 21528
rect 3785 21523 3851 21526
rect 15285 21523 15351 21526
rect 24761 21314 24827 21317
rect 27662 21314 27722 21768
rect 24761 21312 27722 21314
rect 24761 21256 24766 21312
rect 24822 21256 27722 21312
rect 24761 21254 27722 21256
rect 24761 21251 24827 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 18597 21042 18663 21045
rect 24025 21042 24091 21045
rect 18597 21040 24091 21042
rect 18597 20984 18602 21040
rect 18658 20984 24030 21040
rect 24086 20984 24091 21040
rect 18597 20982 24091 20984
rect 18597 20979 18663 20982
rect 24025 20979 24091 20982
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 27520 20544 28000 20664
rect 10225 20498 10291 20501
rect 22737 20498 22803 20501
rect 10225 20496 22803 20498
rect 10225 20440 10230 20496
rect 10286 20440 22742 20496
rect 22798 20440 22803 20496
rect 10225 20438 22803 20440
rect 10225 20435 10291 20438
rect 22737 20435 22803 20438
rect 10041 20362 10107 20365
rect 24209 20362 24275 20365
rect 10041 20360 24275 20362
rect 10041 20304 10046 20360
rect 10102 20304 24214 20360
rect 24270 20304 24275 20360
rect 10041 20302 24275 20304
rect 10041 20299 10107 20302
rect 24209 20299 24275 20302
rect 25221 20226 25287 20229
rect 27662 20226 27722 20544
rect 25221 20224 27722 20226
rect 25221 20168 25226 20224
rect 25282 20168 27722 20224
rect 25221 20166 27722 20168
rect 25221 20163 25287 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 27520 19184 28000 19304
rect 0 19048 480 19168
rect 10277 19072 10597 19073
rect 62 18594 122 19048
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 23473 18730 23539 18733
rect 27662 18730 27722 19184
rect 23473 18728 27722 18730
rect 23473 18672 23478 18728
rect 23534 18672 27722 18728
rect 23473 18670 27722 18672
rect 23473 18667 23539 18670
rect 1577 18594 1643 18597
rect 62 18592 1643 18594
rect 62 18536 1582 18592
rect 1638 18536 1643 18592
rect 62 18534 1643 18536
rect 1577 18531 1643 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 7465 18186 7531 18189
rect 17217 18186 17283 18189
rect 20437 18186 20503 18189
rect 7465 18184 20503 18186
rect 7465 18128 7470 18184
rect 7526 18128 17222 18184
rect 17278 18128 20442 18184
rect 20498 18128 20503 18184
rect 7465 18126 20503 18128
rect 7465 18123 7531 18126
rect 17217 18123 17283 18126
rect 20437 18123 20503 18126
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 27520 17824 28000 17944
rect 2773 17778 2839 17781
rect 3049 17778 3115 17781
rect 13629 17778 13695 17781
rect 2773 17776 13695 17778
rect 2773 17720 2778 17776
rect 2834 17720 3054 17776
rect 3110 17720 13634 17776
rect 13690 17720 13695 17776
rect 2773 17718 13695 17720
rect 2773 17715 2839 17718
rect 3049 17715 3115 17718
rect 13629 17715 13695 17718
rect 14089 17778 14155 17781
rect 23473 17778 23539 17781
rect 14089 17776 23539 17778
rect 14089 17720 14094 17776
rect 14150 17720 23478 17776
rect 23534 17720 23539 17776
rect 14089 17718 23539 17720
rect 14089 17715 14155 17718
rect 23473 17715 23539 17718
rect 8109 17642 8175 17645
rect 15377 17642 15443 17645
rect 8109 17640 15443 17642
rect 8109 17584 8114 17640
rect 8170 17584 15382 17640
rect 15438 17584 15443 17640
rect 8109 17582 15443 17584
rect 8109 17579 8175 17582
rect 15377 17579 15443 17582
rect 25405 17506 25471 17509
rect 27662 17506 27722 17824
rect 25405 17504 27722 17506
rect 25405 17448 25410 17504
rect 25466 17448 27722 17504
rect 25405 17446 27722 17448
rect 25405 17443 25471 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 27520 16464 28000 16584
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 19793 16010 19859 16013
rect 24209 16010 24275 16013
rect 19793 16008 24275 16010
rect 19793 15952 19798 16008
rect 19854 15952 24214 16008
rect 24270 15952 24275 16008
rect 19793 15950 24275 15952
rect 19793 15947 19859 15950
rect 24209 15947 24275 15950
rect 24761 16010 24827 16013
rect 27662 16010 27722 16464
rect 24761 16008 27722 16010
rect 24761 15952 24766 16008
rect 24822 15952 27722 16008
rect 24761 15950 27722 15952
rect 24761 15947 24827 15950
rect 10277 15808 10597 15809
rect 0 15648 480 15768
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 62 15194 122 15648
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 1853 15194 1919 15197
rect 62 15192 1919 15194
rect 62 15136 1858 15192
rect 1914 15136 1919 15192
rect 62 15134 1919 15136
rect 1853 15131 1919 15134
rect 27520 15104 28000 15224
rect 19793 14922 19859 14925
rect 24025 14922 24091 14925
rect 19793 14920 24091 14922
rect 19793 14864 19798 14920
rect 19854 14864 24030 14920
rect 24086 14864 24091 14920
rect 19793 14862 24091 14864
rect 19793 14859 19859 14862
rect 24025 14859 24091 14862
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 18689 14378 18755 14381
rect 27662 14378 27722 15104
rect 18689 14376 27722 14378
rect 18689 14320 18694 14376
rect 18750 14320 27722 14376
rect 18689 14318 27722 14320
rect 18689 14315 18755 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 27520 13968 28000 14000
rect 27520 13912 27618 13968
rect 27674 13912 28000 13968
rect 27520 13880 28000 13912
rect 8845 13698 8911 13701
rect 9806 13698 9812 13700
rect 8845 13696 9812 13698
rect 8845 13640 8850 13696
rect 8906 13640 9812 13696
rect 8845 13638 9812 13640
rect 8845 13635 8911 13638
rect 9806 13636 9812 13638
rect 9876 13636 9882 13700
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 3601 13562 3667 13565
rect 6913 13562 6979 13565
rect 9949 13562 10015 13565
rect 3601 13560 10015 13562
rect 3601 13504 3606 13560
rect 3662 13504 6918 13560
rect 6974 13504 9954 13560
rect 10010 13504 10015 13560
rect 3601 13502 10015 13504
rect 3601 13499 3667 13502
rect 6913 13499 6979 13502
rect 9949 13499 10015 13502
rect 15377 13426 15443 13429
rect 11470 13424 15443 13426
rect 11470 13368 15382 13424
rect 15438 13368 15443 13424
rect 11470 13366 15443 13368
rect 5165 13290 5231 13293
rect 11470 13290 11530 13366
rect 15377 13363 15443 13366
rect 16665 13290 16731 13293
rect 5165 13288 11530 13290
rect 5165 13232 5170 13288
rect 5226 13232 11530 13288
rect 5165 13230 11530 13232
rect 13770 13288 16731 13290
rect 13770 13232 16670 13288
rect 16726 13232 16731 13288
rect 13770 13230 16731 13232
rect 5165 13227 5231 13230
rect 9765 13154 9831 13157
rect 13770 13154 13830 13230
rect 16665 13227 16731 13230
rect 9765 13152 13830 13154
rect 9765 13096 9770 13152
rect 9826 13096 13830 13152
rect 9765 13094 13830 13096
rect 9765 13091 9831 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 9806 12820 9812 12884
rect 9876 12882 9882 12884
rect 19057 12882 19123 12885
rect 9876 12880 19123 12882
rect 9876 12824 19062 12880
rect 19118 12824 19123 12880
rect 9876 12822 19123 12824
rect 9876 12820 9882 12822
rect 19057 12819 19123 12822
rect 6177 12746 6243 12749
rect 16481 12746 16547 12749
rect 6177 12744 16547 12746
rect 6177 12688 6182 12744
rect 6238 12688 16486 12744
rect 16542 12688 16547 12744
rect 6177 12686 16547 12688
rect 6177 12683 6243 12686
rect 16481 12683 16547 12686
rect 27520 12608 28000 12640
rect 27520 12552 27618 12608
rect 27674 12552 28000 12608
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 27520 12520 28000 12552
rect 19610 12479 19930 12480
rect 0 12200 480 12232
rect 0 12144 110 12200
rect 166 12144 480 12200
rect 0 12112 480 12144
rect 15929 12202 15995 12205
rect 24025 12202 24091 12205
rect 15929 12200 24091 12202
rect 15929 12144 15934 12200
rect 15990 12144 24030 12200
rect 24086 12144 24091 12200
rect 15929 12142 24091 12144
rect 15929 12139 15995 12142
rect 24025 12139 24091 12142
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 13169 11658 13235 11661
rect 22829 11658 22895 11661
rect 13169 11656 22895 11658
rect 13169 11600 13174 11656
rect 13230 11600 22834 11656
rect 22890 11600 22895 11656
rect 13169 11598 22895 11600
rect 13169 11595 13235 11598
rect 22829 11595 22895 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 27520 11160 28000 11280
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 5993 10706 6059 10709
rect 19977 10706 20043 10709
rect 5993 10704 20043 10706
rect 5993 10648 5998 10704
rect 6054 10648 19982 10704
rect 20038 10648 20043 10704
rect 5993 10646 20043 10648
rect 5993 10643 6059 10646
rect 19977 10643 20043 10646
rect 20989 10706 21055 10709
rect 27662 10706 27722 11160
rect 20989 10704 27722 10706
rect 20989 10648 20994 10704
rect 21050 10648 27722 10704
rect 20989 10646 27722 10648
rect 20989 10643 21055 10646
rect 6821 10570 6887 10573
rect 14641 10570 14707 10573
rect 6821 10568 14707 10570
rect 6821 10512 6826 10568
rect 6882 10512 14646 10568
rect 14702 10512 14707 10568
rect 6821 10510 14707 10512
rect 6821 10507 6887 10510
rect 14641 10507 14707 10510
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 6453 10162 6519 10165
rect 15285 10162 15351 10165
rect 6453 10160 15351 10162
rect 6453 10104 6458 10160
rect 6514 10104 15290 10160
rect 15346 10104 15351 10160
rect 6453 10102 15351 10104
rect 6453 10099 6519 10102
rect 15285 10099 15351 10102
rect 6729 9890 6795 9893
rect 7097 9890 7163 9893
rect 14089 9890 14155 9893
rect 6729 9888 14155 9890
rect 6729 9832 6734 9888
rect 6790 9832 7102 9888
rect 7158 9832 14094 9888
rect 14150 9832 14155 9888
rect 6729 9830 14155 9832
rect 6729 9827 6795 9830
rect 7097 9827 7163 9830
rect 14089 9827 14155 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 27520 9800 28000 9920
rect 24277 9759 24597 9760
rect 6545 9754 6611 9757
rect 12893 9754 12959 9757
rect 14181 9754 14247 9757
rect 6545 9752 14247 9754
rect 6545 9696 6550 9752
rect 6606 9696 12898 9752
rect 12954 9696 14186 9752
rect 14242 9696 14247 9752
rect 6545 9694 14247 9696
rect 6545 9691 6611 9694
rect 12893 9691 12959 9694
rect 14181 9691 14247 9694
rect 22369 9346 22435 9349
rect 24853 9346 24919 9349
rect 22369 9344 24919 9346
rect 22369 9288 22374 9344
rect 22430 9288 24858 9344
rect 24914 9288 24919 9344
rect 22369 9286 24919 9288
rect 22369 9283 22435 9286
rect 24853 9283 24919 9286
rect 25497 9346 25563 9349
rect 27662 9346 27722 9800
rect 25497 9344 27722 9346
rect 25497 9288 25502 9344
rect 25558 9288 27722 9344
rect 25497 9286 27722 9288
rect 25497 9283 25563 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 5610 8736 5930 8737
rect 0 8664 480 8696
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 0 8608 110 8664
rect 166 8608 480 8664
rect 0 8576 480 8608
rect 27520 8440 28000 8560
rect 1669 8394 1735 8397
rect 13169 8394 13235 8397
rect 1669 8392 13235 8394
rect 1669 8336 1674 8392
rect 1730 8336 13174 8392
rect 13230 8336 13235 8392
rect 1669 8334 13235 8336
rect 1669 8331 1735 8334
rect 13169 8331 13235 8334
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 7281 7986 7347 7989
rect 8845 7986 8911 7989
rect 11421 7986 11487 7989
rect 7281 7984 11487 7986
rect 7281 7928 7286 7984
rect 7342 7928 8850 7984
rect 8906 7928 11426 7984
rect 11482 7928 11487 7984
rect 7281 7926 11487 7928
rect 7281 7923 7347 7926
rect 8845 7923 8911 7926
rect 11421 7923 11487 7926
rect 17677 7850 17743 7853
rect 25589 7850 25655 7853
rect 27662 7850 27722 8440
rect 17677 7848 27722 7850
rect 17677 7792 17682 7848
rect 17738 7792 25594 7848
rect 25650 7792 27722 7848
rect 17677 7790 27722 7792
rect 17677 7787 17743 7790
rect 25589 7787 25655 7790
rect 7833 7714 7899 7717
rect 14641 7714 14707 7717
rect 7833 7712 14707 7714
rect 7833 7656 7838 7712
rect 7894 7656 14646 7712
rect 14702 7656 14707 7712
rect 7833 7654 14707 7656
rect 7833 7651 7899 7654
rect 14641 7651 14707 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 4705 7442 4771 7445
rect 15837 7442 15903 7445
rect 4705 7440 15903 7442
rect 4705 7384 4710 7440
rect 4766 7384 15842 7440
rect 15898 7384 15903 7440
rect 4705 7382 15903 7384
rect 4705 7379 4771 7382
rect 15837 7379 15903 7382
rect 13353 7306 13419 7309
rect 14549 7306 14615 7309
rect 27520 7308 28000 7336
rect 13353 7304 27354 7306
rect 13353 7248 13358 7304
rect 13414 7248 14554 7304
rect 14610 7248 27354 7304
rect 13353 7246 27354 7248
rect 13353 7243 13419 7246
rect 14549 7243 14615 7246
rect 11329 7170 11395 7173
rect 19241 7170 19307 7173
rect 11329 7168 19307 7170
rect 11329 7112 11334 7168
rect 11390 7112 19246 7168
rect 19302 7112 19307 7168
rect 11329 7110 19307 7112
rect 11329 7107 11395 7110
rect 19241 7107 19307 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 27294 7034 27354 7246
rect 27520 7244 27660 7308
rect 27724 7244 28000 7308
rect 27520 7216 28000 7244
rect 27654 7034 27660 7036
rect 27294 6974 27660 7034
rect 27654 6972 27660 6974
rect 27724 6972 27730 7036
rect 8385 6898 8451 6901
rect 12065 6898 12131 6901
rect 17033 6898 17099 6901
rect 8385 6896 17099 6898
rect 8385 6840 8390 6896
rect 8446 6840 12070 6896
rect 12126 6840 17038 6896
rect 17094 6840 17099 6896
rect 8385 6838 17099 6840
rect 8385 6835 8451 6838
rect 12065 6835 12131 6838
rect 17033 6835 17099 6838
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 18505 6218 18571 6221
rect 23749 6218 23815 6221
rect 18505 6216 23815 6218
rect 18505 6160 18510 6216
rect 18566 6160 23754 6216
rect 23810 6160 23815 6216
rect 18505 6158 23815 6160
rect 18505 6155 18571 6158
rect 23749 6155 23815 6158
rect 25865 6218 25931 6221
rect 27654 6218 27660 6220
rect 25865 6216 27660 6218
rect 25865 6160 25870 6216
rect 25926 6160 27660 6216
rect 25865 6158 27660 6160
rect 25865 6155 25931 6158
rect 27654 6156 27660 6158
rect 27724 6156 27730 6220
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 27520 5948 28000 5976
rect 27520 5884 27660 5948
rect 27724 5884 28000 5948
rect 27520 5856 28000 5884
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 5257 5266 5323 5269
rect 6177 5266 6243 5269
rect 17125 5266 17191 5269
rect 5257 5264 17191 5266
rect 5257 5208 5262 5264
rect 5318 5208 6182 5264
rect 6238 5208 17130 5264
rect 17186 5208 17191 5264
rect 5257 5206 17191 5208
rect 5257 5203 5323 5206
rect 6177 5203 6243 5206
rect 17125 5203 17191 5206
rect 0 5128 480 5160
rect 0 5072 110 5128
rect 166 5072 480 5128
rect 0 5040 480 5072
rect 4797 5130 4863 5133
rect 16113 5130 16179 5133
rect 4797 5128 16179 5130
rect 4797 5072 4802 5128
rect 4858 5072 16118 5128
rect 16174 5072 16179 5128
rect 4797 5070 16179 5072
rect 4797 5067 4863 5070
rect 16113 5067 16179 5070
rect 25773 5130 25839 5133
rect 25773 5128 27722 5130
rect 25773 5072 25778 5128
rect 25834 5072 27722 5128
rect 25773 5070 27722 5072
rect 25773 5067 25839 5070
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 4981 4722 5047 4725
rect 9489 4722 9555 4725
rect 10685 4722 10751 4725
rect 4981 4720 10751 4722
rect 4981 4664 4986 4720
rect 5042 4664 9494 4720
rect 9550 4664 10690 4720
rect 10746 4664 10751 4720
rect 4981 4662 10751 4664
rect 4981 4659 5047 4662
rect 9489 4659 9555 4662
rect 10685 4659 10751 4662
rect 27662 4616 27722 5070
rect 4889 4586 4955 4589
rect 10133 4586 10199 4589
rect 11421 4586 11487 4589
rect 13261 4586 13327 4589
rect 4889 4584 13327 4586
rect 4889 4528 4894 4584
rect 4950 4528 10138 4584
rect 10194 4528 11426 4584
rect 11482 4528 13266 4584
rect 13322 4528 13327 4584
rect 4889 4526 13327 4528
rect 4889 4523 4955 4526
rect 10133 4523 10199 4526
rect 11421 4523 11487 4526
rect 13261 4523 13327 4526
rect 27520 4496 28000 4616
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 14365 4178 14431 4181
rect 16481 4178 16547 4181
rect 14365 4176 16547 4178
rect 14365 4120 14370 4176
rect 14426 4120 16486 4176
rect 16542 4120 16547 4176
rect 14365 4118 16547 4120
rect 14365 4115 14431 4118
rect 16481 4115 16547 4118
rect 7649 4042 7715 4045
rect 13445 4042 13511 4045
rect 7649 4040 13511 4042
rect 7649 3984 7654 4040
rect 7710 3984 13450 4040
rect 13506 3984 13511 4040
rect 7649 3982 13511 3984
rect 7649 3979 7715 3982
rect 13445 3979 13511 3982
rect 16849 4042 16915 4045
rect 19517 4042 19583 4045
rect 16849 4040 19583 4042
rect 16849 3984 16854 4040
rect 16910 3984 19522 4040
rect 19578 3984 19583 4040
rect 16849 3982 19583 3984
rect 16849 3979 16915 3982
rect 19517 3979 19583 3982
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 6361 3770 6427 3773
rect 6494 3770 6500 3772
rect 6361 3768 6500 3770
rect 6361 3712 6366 3768
rect 6422 3712 6500 3768
rect 6361 3710 6500 3712
rect 6361 3707 6427 3710
rect 6494 3708 6500 3710
rect 6564 3708 6570 3772
rect 19190 3708 19196 3772
rect 19260 3770 19266 3772
rect 19333 3770 19399 3773
rect 19260 3768 19399 3770
rect 19260 3712 19338 3768
rect 19394 3712 19399 3768
rect 19260 3710 19399 3712
rect 19260 3708 19266 3710
rect 19333 3707 19399 3710
rect 17902 3572 17908 3636
rect 17972 3634 17978 3636
rect 19057 3634 19123 3637
rect 17972 3632 19123 3634
rect 17972 3576 19062 3632
rect 19118 3576 19123 3632
rect 17972 3574 19123 3576
rect 17972 3572 17978 3574
rect 19057 3571 19123 3574
rect 8661 3498 8727 3501
rect 15009 3498 15075 3501
rect 8661 3496 15075 3498
rect 8661 3440 8666 3496
rect 8722 3440 15014 3496
rect 15070 3440 15075 3496
rect 8661 3438 15075 3440
rect 8661 3435 8727 3438
rect 15009 3435 15075 3438
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 27520 3136 28000 3256
rect 3785 3090 3851 3093
rect 4102 3090 4108 3092
rect 3785 3088 4108 3090
rect 3785 3032 3790 3088
rect 3846 3032 4108 3088
rect 3785 3030 4108 3032
rect 3785 3027 3851 3030
rect 4102 3028 4108 3030
rect 4172 3028 4178 3092
rect 12709 2954 12775 2957
rect 4110 2952 12775 2954
rect 4110 2896 12714 2952
rect 12770 2896 12775 2952
rect 4110 2894 12775 2896
rect 3049 2818 3115 2821
rect 4110 2818 4170 2894
rect 12709 2891 12775 2894
rect 13169 2954 13235 2957
rect 27662 2954 27722 3136
rect 13169 2952 27722 2954
rect 13169 2896 13174 2952
rect 13230 2896 27722 2952
rect 13169 2894 27722 2896
rect 13169 2891 13235 2894
rect 16021 2818 16087 2821
rect 3049 2816 4170 2818
rect 3049 2760 3054 2816
rect 3110 2760 4170 2816
rect 3049 2758 4170 2760
rect 13770 2816 16087 2818
rect 13770 2760 16026 2816
rect 16082 2760 16087 2816
rect 13770 2758 16087 2760
rect 3049 2755 3115 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 3141 2546 3207 2549
rect 12893 2546 12959 2549
rect 3141 2544 12959 2546
rect 3141 2488 3146 2544
rect 3202 2488 12898 2544
rect 12954 2488 12959 2544
rect 3141 2486 12959 2488
rect 3141 2483 3207 2486
rect 12893 2483 12959 2486
rect 3049 2410 3115 2413
rect 13770 2410 13830 2758
rect 16021 2755 16087 2758
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 3049 2408 13830 2410
rect 3049 2352 3054 2408
rect 3110 2352 13830 2408
rect 3049 2350 13830 2352
rect 3049 2347 3115 2350
rect 14590 2348 14596 2412
rect 14660 2410 14666 2412
rect 14825 2410 14891 2413
rect 14660 2408 14891 2410
rect 14660 2352 14830 2408
rect 14886 2352 14891 2408
rect 14660 2350 14891 2352
rect 14660 2348 14666 2350
rect 14825 2347 14891 2350
rect 3877 2274 3943 2277
rect 62 2272 3943 2274
rect 62 2216 3882 2272
rect 3938 2216 3943 2272
rect 62 2214 3943 2216
rect 62 1760 122 2214
rect 3877 2211 3943 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 25865 2138 25931 2141
rect 25865 2136 27722 2138
rect 25865 2080 25870 2136
rect 25926 2080 27722 2136
rect 25865 2078 27722 2080
rect 25865 2075 25931 2078
rect 2221 2002 2287 2005
rect 20161 2002 20227 2005
rect 2221 2000 20227 2002
rect 2221 1944 2226 2000
rect 2282 1944 20166 2000
rect 20222 1944 20227 2000
rect 2221 1942 20227 1944
rect 2221 1939 2287 1942
rect 20161 1939 20227 1942
rect 27662 1896 27722 2078
rect 6269 1866 6335 1869
rect 21265 1866 21331 1869
rect 6269 1864 21331 1866
rect 6269 1808 6274 1864
rect 6330 1808 21270 1864
rect 21326 1808 21331 1864
rect 6269 1806 21331 1808
rect 6269 1803 6335 1806
rect 21265 1803 21331 1806
rect 27520 1776 28000 1896
rect 0 1640 480 1760
rect 3509 1730 3575 1733
rect 13169 1730 13235 1733
rect 3509 1728 13235 1730
rect 3509 1672 3514 1728
rect 3570 1672 13174 1728
rect 13230 1672 13235 1728
rect 3509 1670 13235 1672
rect 3509 1667 3575 1670
rect 13169 1667 13235 1670
rect 3325 1594 3391 1597
rect 15653 1594 15719 1597
rect 3325 1592 15719 1594
rect 3325 1536 3330 1592
rect 3386 1536 15658 1592
rect 15714 1536 15719 1592
rect 3325 1534 15719 1536
rect 3325 1531 3391 1534
rect 15653 1531 15719 1534
rect 4521 1458 4587 1461
rect 12382 1458 12388 1460
rect 4521 1456 12388 1458
rect 4521 1400 4526 1456
rect 4582 1400 12388 1456
rect 4521 1398 12388 1400
rect 4521 1395 4587 1398
rect 12382 1396 12388 1398
rect 12452 1396 12458 1460
rect 5993 1322 6059 1325
rect 19241 1322 19307 1325
rect 5993 1320 19307 1322
rect 5993 1264 5998 1320
rect 6054 1264 19246 1320
rect 19302 1264 19307 1320
rect 5993 1262 19307 1264
rect 5993 1259 6059 1262
rect 19241 1259 19307 1262
rect 6913 1186 6979 1189
rect 17677 1186 17743 1189
rect 6913 1184 17743 1186
rect 6913 1128 6918 1184
rect 6974 1128 17682 1184
rect 17738 1128 17743 1184
rect 6913 1126 17743 1128
rect 6913 1123 6979 1126
rect 17677 1123 17743 1126
rect 25773 1186 25839 1189
rect 25773 1184 27722 1186
rect 25773 1128 25778 1184
rect 25834 1128 27722 1184
rect 25773 1126 27722 1128
rect 25773 1123 25839 1126
rect 2497 1050 2563 1053
rect 22921 1050 22987 1053
rect 2497 1048 22987 1050
rect 2497 992 2502 1048
rect 2558 992 22926 1048
rect 22982 992 22987 1048
rect 2497 990 22987 992
rect 2497 987 2563 990
rect 22921 987 22987 990
rect 27662 672 27722 1126
rect 27520 552 28000 672
<< via3 >>
rect 9812 27508 9876 27572
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 9812 13636 9876 13700
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 9812 12820 9876 12884
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 27660 7244 27724 7308
rect 27660 6972 27724 7036
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 27660 6156 27724 6220
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 27660 5884 27724 5948
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 6500 3708 6564 3772
rect 19196 3708 19260 3772
rect 17908 3572 17972 3636
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 4108 3028 4172 3092
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 14596 2348 14660 2412
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 12388 1396 12452 1460
<< metal4 >>
rect 9811 27572 9877 27573
rect 9811 27508 9812 27572
rect 9876 27508 9877 27572
rect 9811 27507 9877 27508
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 9814 13701 9874 27507
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 9811 13700 9877 13701
rect 9811 13636 9812 13700
rect 9876 13636 9877 13700
rect 9811 13635 9877 13636
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 9814 12885 9874 13635
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 9811 12884 9877 12885
rect 9811 12820 9812 12884
rect 9876 12820 9877 12884
rect 9811 12819 9877 12820
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 4107 3092 4173 3093
rect 4107 3028 4108 3092
rect 4172 3028 4173 3092
rect 4107 3027 4173 3028
rect 4110 2498 4170 3027
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 17907 3636 17973 3637
rect 17907 3572 17908 3636
rect 17972 3572 17973 3636
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 17907 3571 17973 3572
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 12387 1460 12453 1461
rect 12387 1396 12388 1460
rect 12452 1396 12453 1460
rect 12387 1395 12453 1396
rect 12390 1138 12450 1395
rect 17910 1138 17970 3571
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 27659 7308 27725 7309
rect 27659 7244 27660 7308
rect 27724 7244 27725 7308
rect 27659 7243 27725 7244
rect 27662 7037 27722 7243
rect 27659 7036 27725 7037
rect 27659 6972 27660 7036
rect 27724 6972 27725 7036
rect 27659 6971 27725 6972
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 27659 6220 27725 6221
rect 27659 6156 27660 6220
rect 27724 6156 27725 6220
rect 27659 6155 27725 6156
rect 27662 5949 27722 6155
rect 27659 5948 27725 5949
rect 27659 5884 27660 5948
rect 27724 5884 27725 5948
rect 27659 5883 27725 5884
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 6414 3772 6650 3858
rect 6414 3708 6500 3772
rect 6500 3708 6564 3772
rect 6564 3708 6650 3772
rect 6414 3622 6650 3708
rect 4022 2262 4258 2498
rect 19110 3772 19346 3858
rect 19110 3708 19196 3772
rect 19196 3708 19260 3772
rect 19260 3708 19346 3772
rect 19110 3622 19346 3708
rect 14510 2412 14746 2498
rect 14510 2348 14596 2412
rect 14596 2348 14660 2412
rect 14660 2348 14746 2412
rect 14510 2262 14746 2348
rect 12302 902 12538 1138
rect 17822 902 18058 1138
<< metal5 >>
rect 6372 3858 19388 3900
rect 6372 3622 6414 3858
rect 6650 3622 19110 3858
rect 19346 3622 19388 3858
rect 6372 3580 19388 3622
rect 3980 2498 14788 2540
rect 3980 2262 4022 2498
rect 4258 2262 14510 2498
rect 14746 2262 14788 2498
rect 3980 2220 14788 2262
rect 12260 1138 18100 1180
rect 12260 902 12302 1138
rect 12538 902 17822 1138
rect 18058 902 18100 1138
rect 12260 860 18100 902
use scs8hd_decap_6  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 590 592
use scs8hd_decap_6  FILLER_0_3
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_12 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1932 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_14
timestamp 1586364061
transform 1 0 2392 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_16 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2576 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2576 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_18
timestamp 1586364061
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 2720
box -38 -48 314 592
use scs8hd_conb_1  _187_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3128 0 1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_1_25
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 590 592
use scs8hd_decap_4  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 4232 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_1  _091_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_40
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_36
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_43
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_36
timestamp 1586364061
transform 1 0 4416 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__C
timestamp 1586364061
transform 1 0 4600 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _078_
timestamp 1586364061
transform 1 0 4784 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_47
timestamp 1586364061
transform 1 0 5428 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 5612 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_1  _094_
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 314 592
use scs8hd_or3_4  _077_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use scs8hd_decap_3  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_68
timestamp 1586364061
transform 1 0 7360 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__C
timestamp 1586364061
transform 1 0 7084 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 7084 0 -1 2720
box -38 -48 314 592
use scs8hd_or3_4  _099_
timestamp 1586364061
transform 1 0 7268 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_80
timestamp 1586364061
transform 1 0 8464 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_76
timestamp 1586364061
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__C
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _089_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _076_
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_97
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_93
timestamp 1586364061
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_94 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__C
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _215_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9844 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_101
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_99
timestamp 1586364061
transform 1 0 10212 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__215__A
timestamp 1586364061
transform 1 0 10396 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_123
timestamp 1586364061
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12236 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_5_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_0_130
timestamp 1586364061
transform 1 0 13064 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__216__A
timestamp 1586364061
transform 1 0 13248 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _216_
timestamp 1586364061
transform 1 0 12696 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_138
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_134
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__212__A
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_157
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_153
timestamp 1586364061
transform 1 0 15180 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__211__A
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_172 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16928 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_170
timestamp 1586364061
transform 1 0 16744 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_176
timestamp 1586364061
transform 1 0 17296 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_180
timestamp 1586364061
transform 1 0 17664 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _210_
timestamp 1586364061
transform 1 0 18124 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _209_
timestamp 1586364061
transform 1 0 18400 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_189
timestamp 1586364061
transform 1 0 18492 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_192
timestamp 1586364061
transform 1 0 18768 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__210__A
timestamp 1586364061
transform 1 0 18676 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18952 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20700 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_209
timestamp 1586364061
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_212
timestamp 1586364061
transform 1 0 20608 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_215
timestamp 1586364061
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_221
timestamp 1586364061
transform 1 0 21436 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_230
timestamp 1586364061
transform 1 0 22264 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_225
timestamp 1586364061
transform 1 0 21804 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22172 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 21252 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_234
timestamp 1586364061
transform 1 0 22632 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_238
timestamp 1586364061
transform 1 0 23000 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_247
timestamp 1586364061
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23644 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_258
timestamp 1586364061
transform 1 0 24840 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_254
timestamp 1586364061
transform 1 0 24472 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_265
timestamp 1586364061
transform 1 0 25484 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_265
timestamp 1586364061
transform 1 0 25484 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25668 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25300 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24288 0 -1 2720
box -38 -48 866 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_0_269 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25852 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_8  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1932 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_6  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_8  FILLER_2_12
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_6  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 590 592
use scs8hd_nor2_4  _142_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 4692 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 5888 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_38
timestamp 1586364061
transform 1 0 4600 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_50
timestamp 1586364061
transform 1 0 5704 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _075_
timestamp 1586364061
transform 1 0 6440 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_54
timestamp 1586364061
transform 1 0 6072 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_67
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_71
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_or3_4  _096_
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 9292 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 130 592
use scs8hd_or3_4  _093_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_91
timestamp 1586364061
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_107
timestamp 1586364061
transform 1 0 10948 0 -1 3808
box -38 -48 314 592
use scs8hd_buf_1  _097_
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12236 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 11684 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12052 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_113
timestamp 1586364061
transform 1 0 11500 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _212_
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13432 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_132
timestamp 1586364061
transform 1 0 13248 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_136
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_140
timestamp 1586364061
transform 1 0 13984 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _211_
timestamp 1586364061
transform 1 0 17112 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_167
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_173
timestamp 1586364061
transform 1 0 17020 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18216 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__213__A
timestamp 1586364061
transform 1 0 17664 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_182
timestamp 1586364061
transform 1 0 17848 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19412 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_197
timestamp 1586364061
transform 1 0 19228 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_201
timestamp 1586364061
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_205
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_209
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 21712 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21252 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  FILLER_2_221
timestamp 1586364061
transform 1 0 21436 0 -1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_8  FILLER_2_235
timestamp 1586364061
transform 1 0 22724 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_2_243
timestamp 1586364061
transform 1 0 23460 0 -1 3808
box -38 -48 222 592
use scs8hd_conb_1  _189_
timestamp 1586364061
transform 1 0 25208 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_254
timestamp 1586364061
transform 1 0 24472 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_258
timestamp 1586364061
transform 1 0 24840 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_265
timestamp 1586364061
transform 1 0 25484 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_273
timestamp 1586364061
transform 1 0 26220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3128 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_25
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_29
timestamp 1586364061
transform 1 0 3772 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_36
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_40
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 6440 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_60
timestamp 1586364061
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_68
timestamp 1586364061
transform 1 0 7360 0 1 3808
box -38 -48 222 592
use scs8hd_or3_4  _090_
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 866 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 7728 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 8740 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_81
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_85
timestamp 1586364061
transform 1 0 8924 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__C
timestamp 1586364061
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 10672 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_102
timestamp 1586364061
transform 1 0 10488 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_106
timestamp 1586364061
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _217_
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__C
timestamp 1586364061
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use scs8hd_buf_2  _214_
timestamp 1586364061
transform 1 0 12696 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__214__A
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_130
timestamp 1586364061
transform 1 0 13064 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_134
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_151
timestamp 1586364061
transform 1 0 14996 0 1 3808
box -38 -48 222 592
use scs8hd_buf_1  _087_
timestamp 1586364061
transform 1 0 16928 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_164
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_168
timestamp 1586364061
transform 1 0 16560 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18308 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20056 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19504 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19872 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_198
timestamp 1586364061
transform 1 0 19320 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_202
timestamp 1586364061
transform 1 0 19688 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 21620 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_215
timestamp 1586364061
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_219
timestamp 1586364061
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23828 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_234
timestamp 1586364061
transform 1 0 22632 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_238
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_242
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_249
timestamp 1586364061
transform 1 0 24012 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24380 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24196 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25392 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_262
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_266
timestamp 1586364061
transform 1 0 25576 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_274
timestamp 1586364061
transform 1 0 26312 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__C
timestamp 1586364061
transform 1 0 4324 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_19
timestamp 1586364061
transform 1 0 2852 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 314 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 4692 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_37
timestamp 1586364061
transform 1 0 4508 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_50
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 590 592
use scs8hd_inv_8  _080_
timestamp 1586364061
transform 1 0 6440 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__081__C
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_67
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_71
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 9292 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 130 592
use scs8hd_or3_4  _086_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_91
timestamp 1586364061
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_107
timestamp 1586364061
transform 1 0 10948 0 -1 4896
box -38 -48 314 592
use scs8hd_buf_1  _116_
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__217__A
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_113
timestamp 1586364061
transform 1 0 11500 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_121
timestamp 1586364061
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_136
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_140
timestamp 1586364061
transform 1 0 13984 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_158
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_171
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 774 592
use scs8hd_buf_2  _213_
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18952 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 18308 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18676 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_179
timestamp 1586364061
transform 1 0 17572 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_184
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_189
timestamp 1586364061
transform 1 0 18492 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_193
timestamp 1586364061
transform 1 0 18860 0 -1 4896
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_203
timestamp 1586364061
transform 1 0 19780 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_207
timestamp 1586364061
transform 1 0 20148 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22080 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_226
timestamp 1586364061
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_230
timestamp 1586364061
transform 1 0 22264 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22448 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_243
timestamp 1586364061
transform 1 0 23460 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_247
timestamp 1586364061
transform 1 0 23828 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24472 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24104 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_252
timestamp 1586364061
transform 1 0 24288 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_buf_1  _138_
timestamp 1586364061
transform 1 0 2668 0 1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_6
timestamp 1586364061
transform 1 0 1656 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_10
timestamp 1586364061
transform 1 0 2024 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_16
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3680 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4140 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 3128 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 3496 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_20
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_24
timestamp 1586364061
transform 1 0 3312 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_31
timestamp 1586364061
transform 1 0 3956 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_35
timestamp 1586364061
transform 1 0 4324 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _136_
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 4508 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_42
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_46
timestamp 1586364061
transform 1 0 5336 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 406 592
use scs8hd_inv_8  _114_
timestamp 1586364061
transform 1 0 7452 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 6440 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 7268 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_60
timestamp 1586364061
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_66
timestamp 1586364061
transform 1 0 7176 0 1 4896
box -38 -48 130 592
use scs8hd_inv_8  _103_
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__C
timestamp 1586364061
transform 1 0 8464 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_78
timestamp 1586364061
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_82
timestamp 1586364061
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_95
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_99
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_121
timestamp 1586364061
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 12696 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14076 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_139
timestamp 1586364061
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_154
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_158
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18216 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_188
timestamp 1586364061
transform 1 0 18400 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20056 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19688 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_200
timestamp 1586364061
transform 1 0 19504 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_204
timestamp 1586364061
transform 1 0 19872 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 21252 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_217
timestamp 1586364061
transform 1 0 21068 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_221
timestamp 1586364061
transform 1 0 21436 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_265
timestamp 1586364061
transform 1 0 25484 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_buf_1  _128_
timestamp 1586364061
transform 1 0 2944 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_19
timestamp 1586364061
transform 1 0 2852 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_6  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_4  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_40
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_36
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_38
timestamp 1586364061
transform 1 0 4600 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 4692 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_50
timestamp 1586364061
transform 1 0 5704 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__C
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 222 592
use scs8hd_or3_4  _137_
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use scs8hd_or3_4  _135_
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_54
timestamp 1586364061
transform 1 0 6072 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_71
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_67
timestamp 1586364061
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_or3_4  _081_
timestamp 1586364061
transform 1 0 6440 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_80
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_84
timestamp 1586364061
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 8648 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use scs8hd_or3_4  _127_
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use scs8hd_or3_4  _115_
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_97
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_101
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _145_
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 866 592
use scs8hd_or3_4  _104_
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_115
timestamp 1586364061
transform 1 0 11684 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_112
timestamp 1586364061
transform 1 0 11408 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__146__C
timestamp 1586364061
transform 1 0 11500 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12512 0 1 5984
box -38 -48 314 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 12052 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_131
timestamp 1586364061
transform 1 0 13156 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_127
timestamp 1586364061
transform 1 0 12788 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_132
timestamp 1586364061
transform 1 0 13248 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_128
timestamp 1586364061
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 13064 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 13340 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12972 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 14536 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15088 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_144
timestamp 1586364061
transform 1 0 14352 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_148
timestamp 1586364061
transform 1 0 14720 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_167
timestamp 1586364061
transform 1 0 16468 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_163
timestamp 1586364061
transform 1 0 16100 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_169
timestamp 1586364061
transform 1 0 16652 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_165
timestamp 1586364061
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 16652 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 16284 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_178
timestamp 1586364061
transform 1 0 17480 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_174
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_177
timestamp 1586364061
transform 1 0 17388 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 17296 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _079_
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_182
timestamp 1586364061
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_181
timestamp 1586364061
transform 1 0 17756 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17572 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17664 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_195
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_195
timestamp 1586364061
transform 1 0 19044 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_191
timestamp 1586364061
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18860 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17848 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_7_200
timestamp 1586364061
transform 1 0 19504 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19872 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19320 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_214
timestamp 1586364061
transform 1 0 20792 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_6_210
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 19780 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 21252 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22080 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_226
timestamp 1586364061
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_230
timestamp 1586364061
transform 1 0 22264 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_218
timestamp 1586364061
transform 1 0 21160 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_221
timestamp 1586364061
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_238
timestamp 1586364061
transform 1 0 23000 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_234
timestamp 1586364061
transform 1 0 22632 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 222 592
use scs8hd_conb_1  _188_
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_248
timestamp 1586364061
transform 1 0 23920 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_242
timestamp 1586364061
transform 1 0 23368 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23736 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23736 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25300 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_259
timestamp 1586364061
transform 1 0 24932 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_255
timestamp 1586364061
transform 1 0 24564 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_259
timestamp 1586364061
transform 1 0 24932 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_266
timestamp 1586364061
transform 1 0 25576 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25760 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26128 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_271
timestamp 1586364061
transform 1 0 26036 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_270
timestamp 1586364061
transform 1 0 25944 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_274
timestamp 1586364061
transform 1 0 26312 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_35
timestamp 1586364061
transform 1 0 4324 0 -1 7072
box -38 -48 222 592
use scs8hd_or3_4  _083_
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 4508 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_39
timestamp 1586364061
transform 1 0 4692 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_52
timestamp 1586364061
transform 1 0 5888 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6624 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_58
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_69
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 406 592
use scs8hd_buf_1  _084_
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_75
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_79
timestamp 1586364061
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_90
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_104
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use scs8hd_or3_4  _146_
timestamp 1586364061
transform 1 0 11500 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_4  FILLER_8_108
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_112
timestamp 1586364061
transform 1 0 11408 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_122
timestamp 1586364061
transform 1 0 12328 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_132
timestamp 1586364061
transform 1 0 13248 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_149
timestamp 1586364061
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_158
timestamp 1586364061
transform 1 0 15640 0 -1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 16008 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_171
timestamp 1586364061
transform 1 0 16836 0 -1 7072
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17572 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18768 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_194
timestamp 1586364061
transform 1 0 18952 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19320 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19780 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20332 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_201
timestamp 1586364061
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_205
timestamp 1586364061
transform 1 0 19964 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  FILLER_8_211
timestamp 1586364061
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 21804 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21068 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_219
timestamp 1586364061
transform 1 0 21252 0 -1 7072
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_236
timestamp 1586364061
transform 1 0 22816 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_244
timestamp 1586364061
transform 1 0 23552 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_254
timestamp 1586364061
transform 1 0 24472 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_8  FILLER_8_265
timestamp 1586364061
transform 1 0 25484 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_273
timestamp 1586364061
transform 1 0 26220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _147_
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5244 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_42
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_47
timestamp 1586364061
transform 1 0 5428 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_88
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 10948 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_92
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_105
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11868 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_109
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_115
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_119
timestamp 1586364061
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_130
timestamp 1586364061
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_134
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_151
timestamp 1586364061
transform 1 0 14996 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_158
timestamp 1586364061
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_162
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20332 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 19320 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 19688 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20148 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_200
timestamp 1586364061
transform 1 0 19504 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_204
timestamp 1586364061
transform 1 0 19872 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_218
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_222
timestamp 1586364061
transform 1 0 21528 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_236
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_240
timestamp 1586364061
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_254
timestamp 1586364061
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_265
timestamp 1586364061
transform 1 0 25484 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_conb_1  _197_
timestamp 1586364061
transform 1 0 4232 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_37
timestamp 1586364061
transform 1 0 4508 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_6  FILLER_10_48
timestamp 1586364061
transform 1 0 5520 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_65
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_69
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _098_
timestamp 1586364061
transform 1 0 9936 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11500 0 -1 8160
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_10_124
timestamp 1586364061
transform 1 0 12512 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12696 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_128
timestamp 1586364061
transform 1 0 12880 0 -1 8160
box -38 -48 590 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 16928 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 16744 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_168
timestamp 1586364061
transform 1 0 16560 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18676 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17940 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_181
timestamp 1586364061
transform 1 0 17756 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_185
timestamp 1586364061
transform 1 0 18124 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_189
timestamp 1586364061
transform 1 0 18492 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_193
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_226
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_230
timestamp 1586364061
transform 1 0 22264 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24012 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_243
timestamp 1586364061
transform 1 0 23460 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_247
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_12  FILLER_10_260
timestamp 1586364061
transform 1 0 25024 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_272
timestamp 1586364061
transform 1 0 26128 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_6
timestamp 1586364061
transform 1 0 1656 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_10
timestamp 1586364061
transform 1 0 2024 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_22
timestamp 1586364061
transform 1 0 3128 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_34
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_buf_1  _082_
timestamp 1586364061
transform 1 0 7084 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 7544 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_68
timestamp 1586364061
transform 1 0 7360 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 8096 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_72
timestamp 1586364061
transform 1 0 7728 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_87
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _092_
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_91
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_104
timestamp 1586364061
transform 1 0 10672 0 1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_134
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15180 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_151
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_155
timestamp 1586364061
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17480 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_163
timestamp 1586364061
transform 1 0 16100 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_180
timestamp 1586364061
transform 1 0 17664 0 1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_194
timestamp 1586364061
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19688 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_198
timestamp 1586364061
transform 1 0 19320 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_211
timestamp 1586364061
transform 1 0 20516 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21252 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 22264 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_217
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_228
timestamp 1586364061
transform 1 0 22080 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_236
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_240
timestamp 1586364061
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23828 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_11_249
timestamp 1586364061
transform 1 0 24012 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24288 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25300 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25668 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_261
timestamp 1586364061
transform 1 0 25116 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_265
timestamp 1586364061
transform 1 0 25484 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_46
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6072 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 7084 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_63
timestamp 1586364061
transform 1 0 6900 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_67
timestamp 1586364061
transform 1 0 7268 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_71
timestamp 1586364061
transform 1 0 7636 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use scs8hd_buf_1  _105_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 10120 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_96
timestamp 1586364061
transform 1 0 9936 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_100
timestamp 1586364061
transform 1 0 10304 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_104
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_107
timestamp 1586364061
transform 1 0 10948 0 -1 9248
box -38 -48 130 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_136
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_140
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15548 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_144
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_150
timestamp 1586364061
transform 1 0 14904 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_168
timestamp 1586364061
transform 1 0 16560 0 -1 9248
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18492 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_181
timestamp 1586364061
transform 1 0 17756 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_200
timestamp 1586364061
transform 1 0 19504 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_204
timestamp 1586364061
transform 1 0 19872 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 21896 0 -1 9248
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_218
timestamp 1586364061
transform 1 0 21160 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_222
timestamp 1586364061
transform 1 0 21528 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23276 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_237
timestamp 1586364061
transform 1 0 22908 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_243
timestamp 1586364061
transform 1 0 23460 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_254
timestamp 1586364061
transform 1 0 24472 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_258
timestamp 1586364061
transform 1 0 24840 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_265
timestamp 1586364061
transform 1 0 25484 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_273
timestamp 1586364061
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 774 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 5796 0 -1 10336
box -38 -48 866 592
use scs8hd_buf_1  _126_
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4784 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_13_42
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_43
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_8  _186_
timestamp 1586364061
transform 1 0 7084 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_14_60
timestamp 1586364061
transform 1 0 6624 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_77
timestamp 1586364061
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_78
timestamp 1586364061
transform 1 0 8280 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 8464 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_87
timestamp 1586364061
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_81
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 8924 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__C
timestamp 1586364061
transform 1 0 9292 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 8648 0 1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_14_97
timestamp 1586364061
transform 1 0 10028 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_91
timestamp 1586364061
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_97
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_13_91
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__171__C
timestamp 1586364061
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_1  _102_
timestamp 1586364061
transform 1 0 10120 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_101
timestamp 1586364061
transform 1 0 10396 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_100
timestamp 1586364061
transform 1 0 10304 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 10580 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use scs8hd_inv_8  _125_
timestamp 1586364061
transform 1 0 11132 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 406 592
use scs8hd_decap_4  FILLER_14_118
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_122
timestamp 1586364061
transform 1 0 12328 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_133
timestamp 1586364061
transform 1 0 13340 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_130
timestamp 1586364061
transform 1 0 13064 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_126
timestamp 1586364061
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_6  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_151
timestamp 1586364061
transform 1 0 14996 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_143
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 14812 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15364 0 1 9248
box -38 -48 1050 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_4  FILLER_13_166
timestamp 1586364061
transform 1 0 16376 0 1 9248
box -38 -48 406 592
use scs8hd_decap_6  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_174
timestamp 1586364061
transform 1 0 17112 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_173
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_170
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17296 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18492 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 18308 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_193
timestamp 1586364061
transform 1 0 18860 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19688 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20056 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_200
timestamp 1586364061
transform 1 0 19504 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_204
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_204
timestamp 1586364061
transform 1 0 19872 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_212
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 21804 0 1 9248
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 21528 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 21528 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 21068 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_221
timestamp 1586364061
transform 1 0 21436 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_224
timestamp 1586364061
transform 1 0 21712 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_219
timestamp 1586364061
transform 1 0 21252 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_237
timestamp 1586364061
transform 1 0 22908 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_233
timestamp 1586364061
transform 1 0 22540 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_236
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22724 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23276 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 866 592
use scs8hd_decap_4  FILLER_14_254
timestamp 1586364061
transform 1 0 24472 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_250
timestamp 1586364061
transform 1 0 24104 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_254
timestamp 1586364061
transform 1 0 24472 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 24288 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_267
timestamp 1586364061
transform 1 0 25668 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_265
timestamp 1586364061
transform 1 0 25484 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_260
timestamp 1586364061
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_19
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_31
timestamp 1586364061
transform 1 0 3956 0 1 10336
box -38 -48 1142 592
use scs8hd_buf_1  _154_
timestamp 1586364061
transform 1 0 5704 0 1 10336
box -38 -48 314 592
use scs8hd_decap_6  FILLER_15_43
timestamp 1586364061
transform 1 0 5060 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_49
timestamp 1586364061
transform 1 0 5612 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7544 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6992 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7360 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_66
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 222 592
use scs8hd_nor4_4  _172_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__172__D
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_81
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_85
timestamp 1586364061
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_106
timestamp 1586364061
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__D
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _107_
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_151
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_163
timestamp 1586364061
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_167
timestamp 1586364061
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_174
timestamp 1586364061
transform 1 0 17112 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_178
timestamp 1586364061
transform 1 0 17480 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 17664 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_182
timestamp 1586364061
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_195
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 20608 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_199
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_206
timestamp 1586364061
transform 1 0 20056 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_210
timestamp 1586364061
transform 1 0 20424 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_214
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 21160 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 20976 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_229
timestamp 1586364061
transform 1 0 22172 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22540 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22908 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_235
timestamp 1586364061
transform 1 0 22724 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_239
timestamp 1586364061
transform 1 0 23092 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 24656 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_254
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_258
timestamp 1586364061
transform 1 0 24840 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_265
timestamp 1586364061
transform 1 0 25484 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_18
timestamp 1586364061
transform 1 0 2760 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_30
timestamp 1586364061
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_52
timestamp 1586364061
transform 1 0 5888 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6072 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_2  FILLER_16_65
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_69
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__106__C
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_82
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_86
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use scs8hd_nor4_4  _171_
timestamp 1586364061
transform 1 0 9844 0 -1 11424
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_90
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12144 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_16_112
timestamp 1586364061
transform 1 0 11408 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_131
timestamp 1586364061
transform 1 0 13156 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_135
timestamp 1586364061
transform 1 0 13524 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_138
timestamp 1586364061
transform 1 0 13800 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 17020 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_165
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_169
timestamp 1586364061
transform 1 0 16652 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18768 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_184
timestamp 1586364061
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_188
timestamp 1586364061
transform 1 0 18400 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20148 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_201
timestamp 1586364061
transform 1 0 19596 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_205
timestamp 1586364061
transform 1 0 19964 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_209
timestamp 1586364061
transform 1 0 20332 0 -1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_224
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_228
timestamp 1586364061
transform 1 0 22080 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22540 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_232
timestamp 1586364061
transform 1 0 22448 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_242
timestamp 1586364061
transform 1 0 23368 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_247
timestamp 1586364061
transform 1 0 23828 0 -1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 24104 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_12  FILLER_16_259
timestamp 1586364061
transform 1 0 24932 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_271
timestamp 1586364061
transform 1 0 26036 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_buf_1  _156_
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_17_47
timestamp 1586364061
transform 1 0 5428 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_71
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use scs8hd_or3_4  _106_
timestamp 1586364061
transform 1 0 9200 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_80
timestamp 1586364061
transform 1 0 8464 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_84
timestamp 1586364061
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use scs8hd_or3_4  _117_
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__C
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_97
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_101
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _225_
timestamp 1586364061
transform 1 0 14076 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_136
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_140
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__225__A
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15088 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_145
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_149
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_165
timestamp 1586364061
transform 1 0 16284 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_169
timestamp 1586364061
transform 1 0 16652 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_173
timestamp 1586364061
transform 1 0 17020 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_193
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_197
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_210
timestamp 1586364061
transform 1 0 20424 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_214
timestamp 1586364061
transform 1 0 20792 0 1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 22172 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_217
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_227
timestamp 1586364061
transform 1 0 21988 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_231
timestamp 1586364061
transform 1 0 22356 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23920 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 22540 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 22908 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_235
timestamp 1586364061
transform 1 0 22724 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_239
timestamp 1586364061
transform 1 0 23092 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_243
timestamp 1586364061
transform 1 0 23460 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24932 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24380 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_251
timestamp 1586364061
transform 1 0 24196 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_255
timestamp 1586364061
transform 1 0 24564 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_262
timestamp 1586364061
transform 1 0 25208 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_266
timestamp 1586364061
transform 1 0 25576 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25760 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_270
timestamp 1586364061
transform 1 0 25944 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_276
timestamp 1586364061
transform 1 0 26496 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_52
timestamp 1586364061
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7636 0 -1 12512
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6072 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_63
timestamp 1586364061
transform 1 0 6900 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_67
timestamp 1586364061
transform 1 0 7268 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__D
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_82
timestamp 1586364061
transform 1 0 8648 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use scs8hd_nor4_4  _168_
timestamp 1586364061
transform 1 0 9752 0 -1 12512
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 130 592
use scs8hd_inv_8  _185_
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__169__C
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__D
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_111
timestamp 1586364061
transform 1 0 11316 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_115
timestamp 1586364061
transform 1 0 11684 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_128
timestamp 1586364061
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_132
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15732 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_151
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_157
timestamp 1586364061
transform 1 0 15548 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_161
timestamp 1586364061
transform 1 0 15916 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_174
timestamp 1586364061
transform 1 0 17112 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17848 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 18860 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_191
timestamp 1586364061
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_195
timestamp 1586364061
transform 1 0 19044 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 19872 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 590 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 21896 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_224
timestamp 1586364061
transform 1 0 21712 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_228
timestamp 1586364061
transform 1 0 22080 0 -1 12512
box -38 -48 406 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 22448 0 -1 12512
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24012 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_241
timestamp 1586364061
transform 1 0 23276 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25024 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_252
timestamp 1586364061
transform 1 0 24288 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_8  _182_
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_19_60
timestamp 1586364061
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6440 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_conb_1  _191_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_20_67
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_69
timestamp 1586364061
transform 1 0 7452 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_65
timestamp 1586364061
transform 1 0 7084 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_72
timestamp 1586364061
transform 1 0 7728 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_87
timestamp 1586364061
transform 1 0 9108 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 9292 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8096 0 1 12512
box -38 -48 1050 592
use scs8hd_nor4_4  _167_
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 1602 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__D
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__C
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_91
timestamp 1586364061
transform 1 0 9476 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_115
timestamp 1586364061
transform 1 0 11684 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_110
timestamp 1586364061
transform 1 0 11224 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_19_112
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__D
timestamp 1586364061
transform 1 0 11500 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_nor4_4  _170_
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1602 592
use scs8hd_nor4_4  _169_
timestamp 1586364061
transform 1 0 12052 0 -1 13600
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13800 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_140
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_136
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_140
timestamp 1586364061
transform 1 0 13984 0 -1 13600
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14812 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_144
timestamp 1586364061
transform 1 0 14352 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_158
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_152
timestamp 1586364061
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_8  _183_
timestamp 1586364061
transform 1 0 17020 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_162
timestamp 1586364061
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_165
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_170
timestamp 1586364061
transform 1 0 16744 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_182
timestamp 1586364061
transform 1 0 17848 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 18124 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_193
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _108_
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 19872 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 19688 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_197
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_201
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_213
timestamp 1586364061
transform 1 0 20700 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 314 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 21436 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 21252 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_217
timestamp 1586364061
transform 1 0 21068 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_230
timestamp 1586364061
transform 1 0 22264 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_224
timestamp 1586364061
transform 1 0 21712 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_8  FILLER_20_236
timestamp 1586364061
transform 1 0 22816 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_232
timestamp 1586364061
transform 1 0 22448 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_238
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_234
timestamp 1586364061
transform 1 0 22632 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_247
timestamp 1586364061
transform 1 0 23828 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_248
timestamp 1586364061
transform 1 0 23920 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_252
timestamp 1586364061
transform 1 0 24288 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_19_267
timestamp 1586364061
transform 1 0 25668 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_263
timestamp 1586364061
transform 1 0 25300 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_259
timestamp 1586364061
transform 1 0 24932 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25484 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_258
timestamp 1586364061
transform 1 0 24840 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_275
timestamp 1586364061
transform 1 0 26404 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_270
timestamp 1586364061
transform 1 0 25944 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_274
timestamp 1586364061
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_6
timestamp 1586364061
transform 1 0 1656 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_10
timestamp 1586364061
transform 1 0 2024 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_22
timestamp 1586364061
transform 1 0 3128 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_34
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_46
timestamp 1586364061
transform 1 0 5336 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6992 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7544 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_58
timestamp 1586364061
transform 1 0 6440 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_66
timestamp 1586364061
transform 1 0 7176 0 1 13600
box -38 -48 406 592
use scs8hd_inv_8  _181_
timestamp 1586364061
transform 1 0 9292 0 1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_81
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_85
timestamp 1586364061
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 10304 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_98
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_102
timestamp 1586364061
transform 1 0 10488 0 1 13600
box -38 -48 590 592
use scs8hd_conb_1  _192_
timestamp 1586364061
transform 1 0 11316 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 12052 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_21_121
timestamp 1586364061
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13156 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12972 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 12604 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_127
timestamp 1586364061
transform 1 0 12788 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_142
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14904 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15364 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14720 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_146
timestamp 1586364061
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_153
timestamp 1586364061
transform 1 0 15180 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_157
timestamp 1586364061
transform 1 0 15548 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17020 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_161
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_193
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20148 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 19688 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20608 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_197
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_201
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_21_204
timestamp 1586364061
transform 1 0 19872 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_210
timestamp 1586364061
transform 1 0 20424 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_214
timestamp 1586364061
transform 1 0 20792 0 1 13600
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_221
timestamp 1586364061
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_225
timestamp 1586364061
transform 1 0 21804 0 1 13600
box -38 -48 774 592
use scs8hd_conb_1  _198_
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_236
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_240
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 406 592
use scs8hd_decap_6  FILLER_21_248
timestamp 1586364061
transform 1 0 23920 0 1 13600
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 24472 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_259
timestamp 1586364061
transform 1 0 24932 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_263
timestamp 1586364061
transform 1 0 25300 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_275
timestamp 1586364061
transform 1 0 26404 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6624 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_63
timestamp 1586364061
transform 1 0 6900 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_67
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_71
timestamp 1586364061
transform 1 0 7636 0 -1 14688
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7728 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_74
timestamp 1586364061
transform 1 0 7912 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_79
timestamp 1586364061
transform 1 0 8372 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_85
timestamp 1586364061
transform 1 0 8924 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_buf_1  _158_
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__D
timestamp 1586364061
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_100
timestamp 1586364061
transform 1 0 10304 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_104
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _110_
timestamp 1586364061
transform 1 0 12052 0 -1 14688
box -38 -48 866 592
use scs8hd_buf_1  _160_
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__D
timestamp 1586364061
transform 1 0 11500 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_111
timestamp 1586364061
transform 1 0 11316 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_115
timestamp 1586364061
transform 1 0 11684 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_8  _184_
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 13064 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__D
timestamp 1586364061
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_128
timestamp 1586364061
transform 1 0 12880 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_132
timestamp 1586364061
transform 1 0 13248 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14720 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_150
timestamp 1586364061
transform 1 0 14904 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_22_157
timestamp 1586364061
transform 1 0 15548 0 -1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16560 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 16284 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_167
timestamp 1586364061
transform 1 0 16468 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_177
timestamp 1586364061
transform 1 0 17388 0 -1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 18124 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_194
timestamp 1586364061
transform 1 0 18952 0 -1 14688
box -38 -48 774 592
use scs8hd_buf_1  _118_
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_205
timestamp 1586364061
transform 1 0 19964 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_213
timestamp 1586364061
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use scs8hd_buf_2  _208_
timestamp 1586364061
transform 1 0 24564 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_4  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_259
timestamp 1586364061
transform 1 0 24932 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_271
timestamp 1586364061
transform 1 0 26036 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 6072 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_56
timestamp 1586364061
transform 1 0 6256 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 8924 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_73
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_77
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_81
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_88
timestamp 1586364061
transform 1 0 9200 0 1 14688
box -38 -48 222 592
use scs8hd_nor4_4  _166_
timestamp 1586364061
transform 1 0 9936 0 1 14688
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 9752 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_92
timestamp 1586364061
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use scs8hd_nor4_4  _157_
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__165__C
timestamp 1586364061
transform 1 0 11684 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__C
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_113
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_117
timestamp 1586364061
transform 1 0 11868 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 14168 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_140
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14720 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_144
timestamp 1586364061
transform 1 0 14352 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_157
timestamp 1586364061
transform 1 0 15548 0 1 14688
box -38 -48 222 592
use scs8hd_inv_8  _173_
timestamp 1586364061
transform 1 0 16284 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17296 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_161
timestamp 1586364061
transform 1 0 15916 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_174
timestamp 1586364061
transform 1 0 17112 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_178
timestamp 1586364061
transform 1 0 17480 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _199_
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18584 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_182
timestamp 1586364061
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_23_187
timestamp 1586364061
transform 1 0 18308 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_192
timestamp 1586364061
transform 1 0 18768 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_198
timestamp 1586364061
transform 1 0 19320 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_210
timestamp 1586364061
transform 1 0 20424 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_222
timestamp 1586364061
transform 1 0 21528 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_23_234
timestamp 1586364061
transform 1 0 22632 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_242
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_52
timestamp 1586364061
transform 1 0 5888 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_8  _180_
timestamp 1586364061
transform 1 0 6072 0 -1 15776
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7636 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_63
timestamp 1586364061
transform 1 0 6900 0 -1 15776
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_82
timestamp 1586364061
transform 1 0 8648 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use scs8hd_nor4_4  _165_
timestamp 1586364061
transform 1 0 9936 0 -1 15776
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__D
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use scs8hd_nor4_4  _159_
timestamp 1586364061
transform 1 0 12236 0 -1 15776
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 12052 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 11684 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_113
timestamp 1586364061
transform 1 0 11500 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_117
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 13984 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_138
timestamp 1586364061
transform 1 0 13800 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_142
timestamp 1586364061
transform 1 0 14168 0 -1 15776
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14720 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_150
timestamp 1586364061
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_165
timestamp 1586364061
transform 1 0 16284 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_182
timestamp 1586364061
transform 1 0 17848 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_186
timestamp 1586364061
transform 1 0 18216 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_193
timestamp 1586364061
transform 1 0 18860 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_205
timestamp 1586364061
transform 1 0 19964 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_24_213
timestamp 1586364061
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_25_47
timestamp 1586364061
transform 1 0 5428 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _190_
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7544 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_65
timestamp 1586364061
transform 1 0 7084 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_69
timestamp 1586364061
transform 1 0 7452 0 1 15776
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8280 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8096 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_72
timestamp 1586364061
transform 1 0 7728 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_89
timestamp 1586364061
transform 1 0 9292 0 1 15776
box -38 -48 222 592
use scs8hd_nor4_4  _162_
timestamp 1586364061
transform 1 0 10028 0 1 15776
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 9476 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_93
timestamp 1586364061
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use scs8hd_nor4_4  _164_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__164__C
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 14168 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_140
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14720 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14536 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_144
timestamp 1586364061
transform 1 0 14352 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 406 592
use scs8hd_conb_1  _196_
timestamp 1586364061
transform 1 0 16468 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_165
timestamp 1586364061
transform 1 0 16284 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_170
timestamp 1586364061
transform 1 0 16744 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_174
timestamp 1586364061
transform 1 0 17112 0 1 15776
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17664 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_182
timestamp 1586364061
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_187
timestamp 1586364061
transform 1 0 18308 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_191
timestamp 1586364061
transform 1 0 18676 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_195
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_207
timestamp 1586364061
transform 1 0 20148 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_219
timestamp 1586364061
transform 1 0 21252 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_231
timestamp 1586364061
transform 1 0 22356 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_243
timestamp 1586364061
transform 1 0 23460 0 1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 774 592
use scs8hd_buf_2  _204_
timestamp 1586364061
transform 1 0 24564 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 25116 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_253
timestamp 1586364061
transform 1 0 24380 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_259
timestamp 1586364061
transform 1 0 24932 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_263
timestamp 1586364061
transform 1 0 25300 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_275
timestamp 1586364061
transform 1 0 26404 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_inv_8  _179_
timestamp 1586364061
transform 1 0 5980 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_26_52
timestamp 1586364061
transform 1 0 5888 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_44
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_56
timestamp 1586364061
transform 1 0 6256 0 1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_26_62
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_69
timestamp 1586364061
transform 1 0 7452 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_66
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_80
timestamp 1586364061
transform 1 0 8464 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_76
timestamp 1586364061
transform 1 0 8096 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_79
timestamp 1586364061
transform 1 0 8372 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8280 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_88
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__C
timestamp 1586364061
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8832 0 1 16864
box -38 -48 866 592
use scs8hd_decap_4  FILLER_27_93
timestamp 1586364061
transform 1 0 9660 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__D
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_107
timestamp 1586364061
transform 1 0 10948 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_103
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_99
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__C
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_nor4_4  _161_
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1602 592
use scs8hd_fill_1  FILLER_27_115
timestamp 1586364061
transform 1 0 11684 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_111
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_114
timestamp 1586364061
transform 1 0 11592 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_110
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 11408 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 11776 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_nor4_4  _163_
timestamp 1586364061
transform 1 0 11960 0 -1 16864
box -38 -48 1602 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12880 0 1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12696 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__D
timestamp 1586364061
transform 1 0 13708 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14076 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_135
timestamp 1586364061
transform 1 0 13524 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_139
timestamp 1586364061
transform 1 0 13892 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_139
timestamp 1586364061
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_143
timestamp 1586364061
transform 1 0 14260 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_149
timestamp 1586364061
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_26_143
timestamp 1586364061
transform 1 0 14260 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14444 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_158
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_158
timestamp 1586364061
transform 1 0 15640 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_27_162
timestamp 1586364061
transform 1 0 16008 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_162
timestamp 1586364061
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_175
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_176
timestamp 1586364061
transform 1 0 17296 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_172
timestamp 1586364061
transform 1 0 16928 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 16864
box -38 -48 866 592
use scs8hd_conb_1  _193_
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17664 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_189
timestamp 1586364061
transform 1 0 18492 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_27_187
timestamp 1586364061
transform 1 0 18308 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_201
timestamp 1586364061
transform 1 0 19596 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_26_213
timestamp 1586364061
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_199
timestamp 1586364061
transform 1 0 19412 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_211
timestamp 1586364061
transform 1 0 20516 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_223
timestamp 1586364061
transform 1 0 21620 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_235
timestamp 1586364061
transform 1 0 22724 0 1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_243
timestamp 1586364061
transform 1 0 23460 0 1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 774 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 24564 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 25116 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_253
timestamp 1586364061
transform 1 0 24380 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_259
timestamp 1586364061
transform 1 0 24932 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_263
timestamp 1586364061
transform 1 0 25300 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_275
timestamp 1586364061
transform 1 0 26404 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_8  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4968 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_40
timestamp 1586364061
transform 1 0 4784 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_45
timestamp 1586364061
transform 1 0 5244 0 -1 17952
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_57
timestamp 1586364061
transform 1 0 6348 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_63
timestamp 1586364061
transform 1 0 6900 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_75
timestamp 1586364061
transform 1 0 8004 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_79
timestamp 1586364061
transform 1 0 8372 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_83
timestamp 1586364061
transform 1 0 8740 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_28_86
timestamp 1586364061
transform 1 0 9016 0 -1 17952
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10396 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12144 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11960 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_112
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 590 592
use scs8hd_buf_2  _206_
timestamp 1586364061
transform 1 0 13892 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_131
timestamp 1586364061
transform 1 0 13156 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_135
timestamp 1586364061
transform 1 0 13524 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_138
timestamp 1586364061
transform 1 0 13800 0 -1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_143
timestamp 1586364061
transform 1 0 14260 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_147
timestamp 1586364061
transform 1 0 14628 0 -1 17952
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_163
timestamp 1586364061
transform 1 0 16100 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_168
timestamp 1586364061
transform 1 0 16560 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_180
timestamp 1586364061
transform 1 0 17664 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_192
timestamp 1586364061
transform 1 0 18768 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_204
timestamp 1586364061
transform 1 0 19872 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_212
timestamp 1586364061
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_66
timestamp 1586364061
transform 1 0 7176 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_70
timestamp 1586364061
transform 1 0 7544 0 1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8188 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 9568 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_97
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_101
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13156 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_134
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_138
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_inv_8  _174_
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 15548 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_151
timestamp 1586364061
transform 1 0 14996 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_155
timestamp 1586364061
transform 1 0 15364 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_168
timestamp 1586364061
transform 1 0 16560 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_172
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_180
timestamp 1586364061
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_8  _175_
timestamp 1586364061
transform 1 0 9936 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10948 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_4  FILLER_30_109
timestamp 1586364061
transform 1 0 11132 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_8  FILLER_30_122
timestamp 1586364061
transform 1 0 12328 0 -1 19040
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_130
timestamp 1586364061
transform 1 0 13064 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_30_135
timestamp 1586364061
transform 1 0 13524 0 -1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_149
timestamp 1586364061
transform 1 0 14812 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_152
timestamp 1586364061
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_163
timestamp 1586364061
transform 1 0 16100 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_175
timestamp 1586364061
transform 1 0 17204 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_187
timestamp 1586364061
transform 1 0 18308 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_199
timestamp 1586364061
transform 1 0 19412 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_30_211
timestamp 1586364061
transform 1 0 20516 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_inv_8  _176_
timestamp 1586364061
transform 1 0 9200 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_97
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_101
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13156 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_127
timestamp 1586364061
transform 1 0 12788 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_142
timestamp 1586364061
transform 1 0 14168 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14904 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14352 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14720 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_146
timestamp 1586364061
transform 1 0 14536 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16468 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_163
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_170
timestamp 1586364061
transform 1 0 16744 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_174
timestamp 1586364061
transform 1 0 17112 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_182
timestamp 1586364061
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 24564 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_253
timestamp 1586364061
transform 1 0 24380 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_106
timestamp 1586364061
transform 1 0 10856 0 -1 20128
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11592 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_8  FILLER_32_123
timestamp 1586364061
transform 1 0 12420 0 -1 20128
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_131
timestamp 1586364061
transform 1 0 13156 0 -1 20128
box -38 -48 314 592
use scs8hd_inv_8  _177_
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_32_163
timestamp 1586364061
transform 1 0 16100 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_175
timestamp 1586364061
transform 1 0 17204 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_187
timestamp 1586364061
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_199
timestamp 1586364061
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_32_211
timestamp 1586364061
transform 1 0 20516 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_buf_2  _205_
timestamp 1586364061
transform 1 0 24564 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_4  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_259
timestamp 1586364061
transform 1 0 24932 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_271
timestamp 1586364061
transform 1 0 26036 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_8  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4876 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4876 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_43
timestamp 1586364061
transform 1 0 5060 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_40
timestamp 1586364061
transform 1 0 4784 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_6  FILLER_33_55
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_95
timestamp 1586364061
transform 1 0 9844 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9568 0 1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_34_107
timestamp 1586364061
transform 1 0 10948 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_103
timestamp 1586364061
transform 1 0 10580 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_99
timestamp 1586364061
transform 1 0 10212 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_99
timestamp 1586364061
transform 1 0 10212 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 20128
box -38 -48 222 592
use scs8hd_conb_1  _194_
timestamp 1586364061
transform 1 0 10304 0 -1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 20128
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_112
timestamp 1586364061
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_116
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_114
timestamp 1586364061
transform 1 0 11592 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_130
timestamp 1586364061
transform 1 0 13064 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_126
timestamp 1586364061
transform 1 0 12696 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_130
timestamp 1586364061
transform 1 0 13064 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 -1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_138
timestamp 1586364061
transform 1 0 13800 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_134
timestamp 1586364061
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use scs8hd_conb_1  _195_
timestamp 1586364061
transform 1 0 13984 0 -1 21216
box -38 -48 314 592
use scs8hd_inv_8  _178_
timestamp 1586364061
transform 1 0 13800 0 1 20128
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15824 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_158
timestamp 1586364061
transform 1 0 15640 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_143
timestamp 1586364061
transform 1 0 14260 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_151
timestamp 1586364061
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_162
timestamp 1586364061
transform 1 0 16008 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_174
timestamp 1586364061
transform 1 0 17112 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_182
timestamp 1586364061
transform 1 0 17848 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9292 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_92
timestamp 1586364061
transform 1 0 9568 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_96
timestamp 1586364061
transform 1 0 9936 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_100
timestamp 1586364061
transform 1 0 10304 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_35_112
timestamp 1586364061
transform 1 0 11408 0 1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_35_120
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13800 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_141
timestamp 1586364061
transform 1 0 14076 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14260 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_145
timestamp 1586364061
transform 1 0 14444 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_157
timestamp 1586364061
transform 1 0 15548 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_169
timestamp 1586364061
transform 1 0 16652 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_181
timestamp 1586364061
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 24564 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_253
timestamp 1586364061
transform 1 0 24380 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_96
timestamp 1586364061
transform 1 0 9936 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_108
timestamp 1586364061
transform 1 0 11040 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_120
timestamp 1586364061
transform 1 0 12144 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_132
timestamp 1586364061
transform 1 0 13248 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_144
timestamp 1586364061
transform 1 0 14352 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_36_152
timestamp 1586364061
transform 1 0 15088 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_buf_2  _203_
timestamp 1586364061
transform 1 0 24564 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_4  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_259
timestamp 1586364061
transform 1 0 24932 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_271
timestamp 1586364061
transform 1 0 26036 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_171
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 24564 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_253
timestamp 1586364061
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 24564 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_259
timestamp 1586364061
transform 1 0 24932 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_271
timestamp 1586364061
transform 1 0 26036 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_22
timestamp 1586364061
transform 1 0 3128 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_34
timestamp 1586364061
transform 1 0 4232 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_46
timestamp 1586364061
transform 1 0 5336 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_58
timestamp 1586364061
transform 1 0 6440 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 13800 0 1 23392
box -38 -48 406 592
use scs8hd_decap_3  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_142
timestamp 1586364061
transform 1 0 14168 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 14352 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_146
timestamp 1586364061
transform 1 0 14536 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_158
timestamp 1586364061
transform 1 0 15640 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _224_
timestamp 1586364061
transform 1 0 16376 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__224__A
timestamp 1586364061
transform 1 0 16928 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_170
timestamp 1586364061
transform 1 0 16744 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_174
timestamp 1586364061
transform 1 0 17112 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _223_
timestamp 1586364061
transform 1 0 18124 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__223__A
timestamp 1586364061
transform 1 0 18676 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_182
timestamp 1586364061
transform 1 0 17848 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_189
timestamp 1586364061
transform 1 0 18492 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_193
timestamp 1586364061
transform 1 0 18860 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _221_
timestamp 1586364061
transform 1 0 20424 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _222_
timestamp 1586364061
transform 1 0 19228 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__222__A
timestamp 1586364061
transform 1 0 19780 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_201
timestamp 1586364061
transform 1 0 19596 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_205
timestamp 1586364061
transform 1 0 19964 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_209
timestamp 1586364061
transform 1 0 20332 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_214
timestamp 1586364061
transform 1 0 20792 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _220_
timestamp 1586364061
transform 1 0 21988 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__221__A
timestamp 1586364061
transform 1 0 20976 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_218
timestamp 1586364061
transform 1 0 21160 0 1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_39_226
timestamp 1586364061
transform 1 0 21896 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_231
timestamp 1586364061
transform 1 0 22356 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_8  FILLER_39_235
timestamp 1586364061
transform 1 0 22724 0 1 23392
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__220__A
timestamp 1586364061
transform 1 0 22540 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_247
timestamp 1586364061
transform 1 0 23828 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_6  FILLER_39_249
timestamp 1586364061
transform 1 0 24012 0 1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_243
timestamp 1586364061
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__219__A
timestamp 1586364061
transform 1 0 23828 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_buf_2  _219_
timestamp 1586364061
transform 1 0 23460 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _200_
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _201_
timestamp 1586364061
transform 1 0 24564 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_259
timestamp 1586364061
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_263
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_259
timestamp 1586364061
transform 1 0 24932 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_275
timestamp 1586364061
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_271
timestamp 1586364061
transform 1 0 26036 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 774 592
use scs8hd_buf_2  _218_
timestamp 1586364061
transform 1 0 24564 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__218__A
timestamp 1586364061
transform 1 0 25116 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_253
timestamp 1586364061
transform 1 0 24380 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_259
timestamp 1586364061
transform 1 0 24932 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_263
timestamp 1586364061
transform 1 0 25300 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_275
timestamp 1586364061
transform 1 0 26404 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 8114 0 8170 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 8850 0 8906 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 9678 0 9734 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 10414 0 10470 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 11242 0 11298 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 11978 0 12034 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 12806 0 12862 480 6 address[6]
port 6 nsew default input
rlabel metal2 s 25226 0 25282 480 6 bottom_left_grid_pin_11_
port 7 nsew default input
rlabel metal2 s 25962 0 26018 480 6 bottom_left_grid_pin_13_
port 8 nsew default input
rlabel metal2 s 26790 0 26846 480 6 bottom_left_grid_pin_15_
port 9 nsew default input
rlabel metal2 s 21362 0 21418 480 6 bottom_left_grid_pin_1_
port 10 nsew default input
rlabel metal2 s 22098 0 22154 480 6 bottom_left_grid_pin_3_
port 11 nsew default input
rlabel metal2 s 22834 0 22890 480 6 bottom_left_grid_pin_5_
port 12 nsew default input
rlabel metal2 s 23662 0 23718 480 6 bottom_left_grid_pin_7_
port 13 nsew default input
rlabel metal2 s 24398 0 24454 480 6 bottom_left_grid_pin_9_
port 14 nsew default input
rlabel metal2 s 27526 0 27582 480 6 bottom_right_grid_pin_11_
port 15 nsew default input
rlabel metal3 s 27520 1776 28000 1896 6 chanx_right_in[0]
port 16 nsew default input
rlabel metal3 s 27520 3136 28000 3256 6 chanx_right_in[1]
port 17 nsew default input
rlabel metal3 s 27520 4496 28000 4616 6 chanx_right_in[2]
port 18 nsew default input
rlabel metal3 s 27520 5856 28000 5976 6 chanx_right_in[3]
port 19 nsew default input
rlabel metal3 s 27520 7216 28000 7336 6 chanx_right_in[4]
port 20 nsew default input
rlabel metal3 s 27520 8440 28000 8560 6 chanx_right_in[5]
port 21 nsew default input
rlabel metal3 s 27520 9800 28000 9920 6 chanx_right_in[6]
port 22 nsew default input
rlabel metal3 s 27520 11160 28000 11280 6 chanx_right_in[7]
port 23 nsew default input
rlabel metal3 s 27520 12520 28000 12640 6 chanx_right_in[8]
port 24 nsew default input
rlabel metal3 s 27520 16464 28000 16584 6 chanx_right_out[0]
port 25 nsew default tristate
rlabel metal3 s 27520 17824 28000 17944 6 chanx_right_out[1]
port 26 nsew default tristate
rlabel metal3 s 27520 19184 28000 19304 6 chanx_right_out[2]
port 27 nsew default tristate
rlabel metal3 s 27520 20544 28000 20664 6 chanx_right_out[3]
port 28 nsew default tristate
rlabel metal3 s 27520 21768 28000 21888 6 chanx_right_out[4]
port 29 nsew default tristate
rlabel metal3 s 27520 23128 28000 23248 6 chanx_right_out[5]
port 30 nsew default tristate
rlabel metal3 s 27520 24488 28000 24608 6 chanx_right_out[6]
port 31 nsew default tristate
rlabel metal3 s 27520 25848 28000 25968 6 chanx_right_out[7]
port 32 nsew default tristate
rlabel metal3 s 27520 27208 28000 27328 6 chanx_right_out[8]
port 33 nsew default tristate
rlabel metal2 s 386 0 442 480 6 chany_bottom_in[0]
port 34 nsew default input
rlabel metal2 s 1122 0 1178 480 6 chany_bottom_in[1]
port 35 nsew default input
rlabel metal2 s 1858 0 1914 480 6 chany_bottom_in[2]
port 36 nsew default input
rlabel metal2 s 2686 0 2742 480 6 chany_bottom_in[3]
port 37 nsew default input
rlabel metal2 s 3422 0 3478 480 6 chany_bottom_in[4]
port 38 nsew default input
rlabel metal2 s 4250 0 4306 480 6 chany_bottom_in[5]
port 39 nsew default input
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_in[6]
port 40 nsew default input
rlabel metal2 s 5814 0 5870 480 6 chany_bottom_in[7]
port 41 nsew default input
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_in[8]
port 42 nsew default input
rlabel metal2 s 14370 0 14426 480 6 chany_bottom_out[0]
port 43 nsew default tristate
rlabel metal2 s 15106 0 15162 480 6 chany_bottom_out[1]
port 44 nsew default tristate
rlabel metal2 s 15842 0 15898 480 6 chany_bottom_out[2]
port 45 nsew default tristate
rlabel metal2 s 16670 0 16726 480 6 chany_bottom_out[3]
port 46 nsew default tristate
rlabel metal2 s 17406 0 17462 480 6 chany_bottom_out[4]
port 47 nsew default tristate
rlabel metal2 s 18234 0 18290 480 6 chany_bottom_out[5]
port 48 nsew default tristate
rlabel metal2 s 18970 0 19026 480 6 chany_bottom_out[6]
port 49 nsew default tristate
rlabel metal2 s 19798 0 19854 480 6 chany_bottom_out[7]
port 50 nsew default tristate
rlabel metal2 s 20534 0 20590 480 6 chany_bottom_out[8]
port 51 nsew default tristate
rlabel metal2 s 754 27520 810 28000 6 chany_top_in[0]
port 52 nsew default input
rlabel metal2 s 2226 27520 2282 28000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 3790 27520 3846 28000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 5354 27520 5410 28000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 6918 27520 6974 28000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 8482 27520 8538 28000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 10046 27520 10102 28000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 11610 27520 11666 28000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 13174 27520 13230 28000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 14738 27520 14794 28000 6 chany_top_out[0]
port 61 nsew default tristate
rlabel metal2 s 16210 27520 16266 28000 6 chany_top_out[1]
port 62 nsew default tristate
rlabel metal2 s 17774 27520 17830 28000 6 chany_top_out[2]
port 63 nsew default tristate
rlabel metal2 s 19338 27520 19394 28000 6 chany_top_out[3]
port 64 nsew default tristate
rlabel metal2 s 20902 27520 20958 28000 6 chany_top_out[4]
port 65 nsew default tristate
rlabel metal2 s 22466 27520 22522 28000 6 chany_top_out[5]
port 66 nsew default tristate
rlabel metal2 s 24030 27520 24086 28000 6 chany_top_out[6]
port 67 nsew default tristate
rlabel metal2 s 25594 27520 25650 28000 6 chany_top_out[7]
port 68 nsew default tristate
rlabel metal2 s 27158 27520 27214 28000 6 chany_top_out[8]
port 69 nsew default tristate
rlabel metal2 s 13542 0 13598 480 6 data_in
port 70 nsew default input
rlabel metal2 s 7378 0 7434 480 6 enable
port 71 nsew default input
rlabel metal3 s 27520 15104 28000 15224 6 right_bottom_grid_pin_12_
port 72 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 right_top_grid_pin_10_
port 73 nsew default input
rlabel metal3 s 0 19048 480 19168 6 top_left_grid_pin_11_
port 74 nsew default input
rlabel metal3 s 0 22584 480 22704 6 top_left_grid_pin_13_
port 75 nsew default input
rlabel metal3 s 0 26120 480 26240 6 top_left_grid_pin_15_
port 76 nsew default input
rlabel metal3 s 0 1640 480 1760 6 top_left_grid_pin_1_
port 77 nsew default input
rlabel metal3 s 0 5040 480 5160 6 top_left_grid_pin_3_
port 78 nsew default input
rlabel metal3 s 0 8576 480 8696 6 top_left_grid_pin_5_
port 79 nsew default input
rlabel metal3 s 0 12112 480 12232 6 top_left_grid_pin_7_
port 80 nsew default input
rlabel metal3 s 0 15648 480 15768 6 top_left_grid_pin_9_
port 81 nsew default input
rlabel metal3 s 27520 552 28000 672 6 top_right_grid_pin_11_
port 82 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 83 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 84 nsew default input
<< end >>
