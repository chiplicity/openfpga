magic
tech sky130A
magscale 1 2
timestamp 1604671380
<< locali >>
rect 33977 30039 34011 30277
rect 29009 26299 29043 26469
rect 32965 19159 32999 19465
rect 30021 16983 30055 17221
rect 31677 16439 31711 16745
rect 17693 15895 17727 16201
rect 31309 14399 31343 14569
rect 28917 11543 28951 11645
rect 7941 7191 7975 7293
<< viali >>
rect 35633 36329 35667 36363
rect 35449 36193 35483 36227
rect 35633 35785 35667 35819
rect 35449 35581 35483 35615
rect 33057 35445 33091 35479
rect 33425 35445 33459 35479
rect 35265 35445 35299 35479
rect 36001 35445 36035 35479
rect 33517 35241 33551 35275
rect 32404 35173 32438 35207
rect 34877 35105 34911 35139
rect 32137 35037 32171 35071
rect 34621 35037 34655 35071
rect 34529 34901 34563 34935
rect 36001 34901 36035 34935
rect 36277 34697 36311 34731
rect 37565 34697 37599 34731
rect 34253 34629 34287 34663
rect 34621 34629 34655 34663
rect 33517 34561 33551 34595
rect 34897 34561 34931 34595
rect 30481 34493 30515 34527
rect 32413 34493 32447 34527
rect 32873 34493 32907 34527
rect 37381 34493 37415 34527
rect 37933 34493 37967 34527
rect 30726 34425 30760 34459
rect 33333 34425 33367 34459
rect 35142 34425 35176 34459
rect 30297 34357 30331 34391
rect 31861 34357 31895 34391
rect 32965 34357 32999 34391
rect 33425 34357 33459 34391
rect 30573 34153 30607 34187
rect 33517 34153 33551 34187
rect 32382 34085 32416 34119
rect 34437 34085 34471 34119
rect 34888 34085 34922 34119
rect 32137 33949 32171 33983
rect 34621 33949 34655 33983
rect 30113 33813 30147 33847
rect 34069 33813 34103 33847
rect 36001 33813 36035 33847
rect 31401 33609 31435 33643
rect 34345 33609 34379 33643
rect 32137 33541 32171 33575
rect 32965 33473 32999 33507
rect 33149 33473 33183 33507
rect 30021 33405 30055 33439
rect 30277 33405 30311 33439
rect 32873 33405 32907 33439
rect 33517 33405 33551 33439
rect 35265 33405 35299 33439
rect 35521 33405 35555 33439
rect 29837 33269 29871 33303
rect 32505 33269 32539 33303
rect 34621 33269 34655 33303
rect 35081 33269 35115 33303
rect 36645 33269 36679 33303
rect 30849 33065 30883 33099
rect 32505 33065 32539 33099
rect 32873 33065 32907 33099
rect 33885 33065 33919 33099
rect 35081 33065 35115 33099
rect 29736 32929 29770 32963
rect 35440 32929 35474 32963
rect 29469 32861 29503 32895
rect 33977 32861 34011 32895
rect 34069 32861 34103 32895
rect 35173 32861 35207 32895
rect 33241 32725 33275 32759
rect 33517 32725 33551 32759
rect 36553 32725 36587 32759
rect 29837 32521 29871 32555
rect 30205 32521 30239 32555
rect 33241 32521 33275 32555
rect 34621 32521 34655 32555
rect 36553 32521 36587 32555
rect 36829 32521 36863 32555
rect 30389 32453 30423 32487
rect 31769 32453 31803 32487
rect 33609 32453 33643 32487
rect 36093 32453 36127 32487
rect 30941 32385 30975 32419
rect 32413 32385 32447 32419
rect 32597 32385 32631 32419
rect 35541 32385 35575 32419
rect 35633 32385 35667 32419
rect 30757 32317 30791 32351
rect 31493 32317 31527 32351
rect 32321 32317 32355 32351
rect 33701 32317 33735 32351
rect 36645 32317 36679 32351
rect 30849 32249 30883 32283
rect 29469 32181 29503 32215
rect 31953 32181 31987 32215
rect 33885 32181 33919 32215
rect 34345 32181 34379 32215
rect 35081 32181 35115 32215
rect 35449 32181 35483 32215
rect 37197 32181 37231 32215
rect 29653 31977 29687 32011
rect 30481 31977 30515 32011
rect 30849 31977 30883 32011
rect 31125 31977 31159 32011
rect 32689 31977 32723 32011
rect 33149 31977 33183 32011
rect 33701 31977 33735 32011
rect 34621 31977 34655 32011
rect 35081 31977 35115 32011
rect 36553 31977 36587 32011
rect 33057 31909 33091 31943
rect 28540 31841 28574 31875
rect 30941 31841 30975 31875
rect 35173 31841 35207 31875
rect 35440 31841 35474 31875
rect 28273 31773 28307 31807
rect 33241 31773 33275 31807
rect 31861 31637 31895 31671
rect 32505 31637 32539 31671
rect 34069 31637 34103 31671
rect 31033 31433 31067 31467
rect 31953 31433 31987 31467
rect 32229 31365 32263 31399
rect 32965 31365 32999 31399
rect 32597 31297 32631 31331
rect 33609 31297 33643 31331
rect 33793 31297 33827 31331
rect 35725 31297 35759 31331
rect 31585 31229 31619 31263
rect 32045 31229 32079 31263
rect 33517 31229 33551 31263
rect 34345 31229 34379 31263
rect 34713 31229 34747 31263
rect 35541 31229 35575 31263
rect 24869 31093 24903 31127
rect 27537 31093 27571 31127
rect 28365 31093 28399 31127
rect 28641 31093 28675 31127
rect 33149 31093 33183 31127
rect 35081 31093 35115 31127
rect 35449 31093 35483 31127
rect 36093 31093 36127 31127
rect 24777 30889 24811 30923
rect 25237 30889 25271 30923
rect 32781 30889 32815 30923
rect 33149 30889 33183 30923
rect 35909 30889 35943 30923
rect 27160 30753 27194 30787
rect 32137 30753 32171 30787
rect 33497 30753 33531 30787
rect 35541 30753 35575 30787
rect 35725 30753 35759 30787
rect 25329 30685 25363 30719
rect 25421 30685 25455 30719
rect 26893 30685 26927 30719
rect 33241 30685 33275 30719
rect 24409 30617 24443 30651
rect 35173 30617 35207 30651
rect 24869 30549 24903 30583
rect 28273 30549 28307 30583
rect 29285 30549 29319 30583
rect 29653 30549 29687 30583
rect 32321 30549 32355 30583
rect 34621 30549 34655 30583
rect 36369 30549 36403 30583
rect 33057 30345 33091 30379
rect 24041 30277 24075 30311
rect 24501 30277 24535 30311
rect 26985 30277 27019 30311
rect 32321 30277 32355 30311
rect 33977 30277 34011 30311
rect 34713 30277 34747 30311
rect 36645 30277 36679 30311
rect 28089 30209 28123 30243
rect 29745 30209 29779 30243
rect 29837 30209 29871 30243
rect 32689 30209 32723 30243
rect 33701 30209 33735 30243
rect 24961 30141 24995 30175
rect 25228 30141 25262 30175
rect 27813 30141 27847 30175
rect 28457 30141 28491 30175
rect 28825 30141 28859 30175
rect 29653 30141 29687 30175
rect 31953 30141 31987 30175
rect 27261 30073 27295 30107
rect 27905 30073 27939 30107
rect 33517 30073 33551 30107
rect 35541 30209 35575 30243
rect 35265 30141 35299 30175
rect 36277 30141 36311 30175
rect 36461 30141 36495 30175
rect 35357 30073 35391 30107
rect 37013 30073 37047 30107
rect 24777 30005 24811 30039
rect 26341 30005 26375 30039
rect 27445 30005 27479 30039
rect 29285 30005 29319 30039
rect 30297 30005 30331 30039
rect 33149 30005 33183 30039
rect 33609 30005 33643 30039
rect 33977 30005 34011 30039
rect 34253 30005 34287 30039
rect 34897 30005 34931 30039
rect 35909 30005 35943 30039
rect 25329 29801 25363 29835
rect 27905 29801 27939 29835
rect 28917 29801 28951 29835
rect 30389 29801 30423 29835
rect 35817 29801 35851 29835
rect 24216 29733 24250 29767
rect 26770 29733 26804 29767
rect 29276 29733 29310 29767
rect 33140 29733 33174 29767
rect 26525 29665 26559 29699
rect 29009 29665 29043 29699
rect 35725 29665 35759 29699
rect 23949 29597 23983 29631
rect 32873 29597 32907 29631
rect 35909 29597 35943 29631
rect 23857 29461 23891 29495
rect 26341 29461 26375 29495
rect 32781 29461 32815 29495
rect 34253 29461 34287 29495
rect 34989 29461 35023 29495
rect 35357 29461 35391 29495
rect 25329 29257 25363 29291
rect 25973 29257 26007 29291
rect 26433 29257 26467 29291
rect 32321 29257 32355 29291
rect 32965 29257 32999 29291
rect 36829 29257 36863 29291
rect 37565 29257 37599 29291
rect 27445 29189 27479 29223
rect 28181 29189 28215 29223
rect 30665 29189 30699 29223
rect 36277 29189 36311 29223
rect 26893 29121 26927 29155
rect 27077 29121 27111 29155
rect 33793 29121 33827 29155
rect 34621 29121 34655 29155
rect 34897 29121 34931 29155
rect 23949 29053 23983 29087
rect 24216 29053 24250 29087
rect 26801 29053 26835 29087
rect 27997 29053 28031 29087
rect 29285 29053 29319 29087
rect 32137 29053 32171 29087
rect 33609 29053 33643 29087
rect 37381 29053 37415 29087
rect 26249 28985 26283 29019
rect 29552 28985 29586 29019
rect 32045 28985 32079 29019
rect 33701 28985 33735 29019
rect 34345 28985 34379 29019
rect 35164 28985 35198 29019
rect 38025 28985 38059 29019
rect 23121 28917 23155 28951
rect 23489 28917 23523 28951
rect 27813 28917 27847 28951
rect 28733 28917 28767 28951
rect 29101 28917 29135 28951
rect 33241 28917 33275 28951
rect 24777 28713 24811 28747
rect 26341 28713 26375 28747
rect 29101 28713 29135 28747
rect 32965 28713 32999 28747
rect 34621 28713 34655 28747
rect 35357 28713 35391 28747
rect 35909 28713 35943 28747
rect 36277 28713 36311 28747
rect 26893 28645 26927 28679
rect 29460 28645 29494 28679
rect 23653 28577 23687 28611
rect 28089 28577 28123 28611
rect 33241 28577 33275 28611
rect 33508 28577 33542 28611
rect 35725 28577 35759 28611
rect 23397 28509 23431 28543
rect 26985 28509 27019 28543
rect 27169 28509 27203 28543
rect 29193 28509 29227 28543
rect 26525 28373 26559 28407
rect 27629 28373 27663 28407
rect 28273 28373 28307 28407
rect 30573 28373 30607 28407
rect 32597 28373 32631 28407
rect 22753 28169 22787 28203
rect 25053 28169 25087 28203
rect 26709 28169 26743 28203
rect 27077 28169 27111 28203
rect 27629 28169 27663 28203
rect 32597 28169 32631 28203
rect 33241 28169 33275 28203
rect 34253 28169 34287 28203
rect 35633 28169 35667 28203
rect 36737 28169 36771 28203
rect 25605 28101 25639 28135
rect 34621 28101 34655 28135
rect 28181 28033 28215 28067
rect 33149 28033 33183 28067
rect 33701 28033 33735 28067
rect 33885 28033 33919 28067
rect 23673 27965 23707 27999
rect 26157 27965 26191 27999
rect 27537 27965 27571 27999
rect 28089 27965 28123 27999
rect 29469 27965 29503 27999
rect 31953 27965 31987 27999
rect 33609 27965 33643 27999
rect 35449 27965 35483 27999
rect 36553 27965 36587 27999
rect 23121 27897 23155 27931
rect 23918 27897 23952 27931
rect 28733 27897 28767 27931
rect 29714 27897 29748 27931
rect 31861 27897 31895 27931
rect 23397 27829 23431 27863
rect 26065 27829 26099 27863
rect 26341 27829 26375 27863
rect 27997 27829 28031 27863
rect 29101 27829 29135 27863
rect 30849 27829 30883 27863
rect 32137 27829 32171 27863
rect 35265 27829 35299 27863
rect 36001 27829 36035 27863
rect 37197 27829 37231 27863
rect 24225 27625 24259 27659
rect 27721 27625 27755 27659
rect 28917 27625 28951 27659
rect 29377 27625 29411 27659
rect 28089 27557 28123 27591
rect 28825 27557 28859 27591
rect 32873 27557 32907 27591
rect 35418 27557 35452 27591
rect 26893 27489 26927 27523
rect 29285 27489 29319 27523
rect 30297 27489 30331 27523
rect 30481 27489 30515 27523
rect 30665 27489 30699 27523
rect 30849 27489 30883 27523
rect 32137 27489 32171 27523
rect 33701 27489 33735 27523
rect 33793 27489 33827 27523
rect 35173 27489 35207 27523
rect 24317 27421 24351 27455
rect 24501 27421 24535 27455
rect 26985 27421 27019 27455
rect 27169 27421 27203 27455
rect 29469 27421 29503 27455
rect 30021 27421 30055 27455
rect 33977 27421 34011 27455
rect 23397 27353 23431 27387
rect 26341 27353 26375 27387
rect 33241 27353 33275 27387
rect 23673 27285 23707 27319
rect 23857 27285 23891 27319
rect 26525 27285 26559 27319
rect 32321 27285 32355 27319
rect 33333 27285 33367 27319
rect 34437 27285 34471 27319
rect 36553 27285 36587 27319
rect 22385 27081 22419 27115
rect 25053 27081 25087 27115
rect 26341 27081 26375 27115
rect 26985 27081 27019 27115
rect 28365 27081 28399 27115
rect 31493 27081 31527 27115
rect 32321 27081 32355 27115
rect 33149 27081 33183 27115
rect 34253 27081 34287 27115
rect 28733 27013 28767 27047
rect 32781 27013 32815 27047
rect 33241 27013 33275 27047
rect 36829 27013 36863 27047
rect 27629 26945 27663 26979
rect 27813 26945 27847 26979
rect 33885 26945 33919 26979
rect 22477 26877 22511 26911
rect 23673 26877 23707 26911
rect 29561 26877 29595 26911
rect 29828 26877 29862 26911
rect 32045 26877 32079 26911
rect 32137 26877 32171 26911
rect 33701 26877 33735 26911
rect 35357 26877 35391 26911
rect 35449 26877 35483 26911
rect 35716 26877 35750 26911
rect 23121 26809 23155 26843
rect 23918 26809 23952 26843
rect 25605 26809 25639 26843
rect 27537 26809 27571 26843
rect 33609 26809 33643 26843
rect 34713 26809 34747 26843
rect 22661 26741 22695 26775
rect 23489 26741 23523 26775
rect 26617 26741 26651 26775
rect 27169 26741 27203 26775
rect 29101 26741 29135 26775
rect 30941 26741 30975 26775
rect 23489 26537 23523 26571
rect 24961 26537 24995 26571
rect 26525 26537 26559 26571
rect 28089 26537 28123 26571
rect 28549 26537 28583 26571
rect 29653 26537 29687 26571
rect 30665 26537 30699 26571
rect 31953 26537 31987 26571
rect 32505 26537 32539 26571
rect 35265 26537 35299 26571
rect 23826 26469 23860 26503
rect 26341 26469 26375 26503
rect 28457 26469 28491 26503
rect 29009 26469 29043 26503
rect 29193 26469 29227 26503
rect 32873 26469 32907 26503
rect 33232 26469 33266 26503
rect 35633 26469 35667 26503
rect 26893 26401 26927 26435
rect 26985 26401 27019 26435
rect 23581 26333 23615 26367
rect 25973 26333 26007 26367
rect 27169 26333 27203 26367
rect 27629 26333 27663 26367
rect 28733 26333 28767 26367
rect 30021 26401 30055 26435
rect 32965 26401 32999 26435
rect 35449 26401 35483 26435
rect 30113 26333 30147 26367
rect 30297 26333 30331 26367
rect 29009 26265 29043 26299
rect 29561 26265 29595 26299
rect 35817 26265 35851 26299
rect 34345 26197 34379 26231
rect 26525 25993 26559 26027
rect 28641 25993 28675 26027
rect 32781 25993 32815 26027
rect 33977 25993 34011 26027
rect 34621 25993 34655 26027
rect 35081 25993 35115 26027
rect 35909 25993 35943 26027
rect 36185 25993 36219 26027
rect 25421 25925 25455 25959
rect 26433 25925 26467 25959
rect 27997 25925 28031 25959
rect 32873 25925 32907 25959
rect 26985 25857 27019 25891
rect 27077 25857 27111 25891
rect 32413 25857 32447 25891
rect 33517 25857 33551 25891
rect 23489 25789 23523 25823
rect 24041 25789 24075 25823
rect 28089 25789 28123 25823
rect 29009 25789 29043 25823
rect 29929 25789 29963 25823
rect 32045 25789 32079 25823
rect 33333 25789 33367 25823
rect 34897 25789 34931 25823
rect 36001 25789 36035 25823
rect 36553 25789 36587 25823
rect 23121 25721 23155 25755
rect 24308 25721 24342 25755
rect 30196 25721 30230 25755
rect 23949 25653 23983 25687
rect 26065 25653 26099 25687
rect 26893 25653 26927 25687
rect 27629 25653 27663 25687
rect 28273 25653 28307 25687
rect 29745 25653 29779 25687
rect 31309 25653 31343 25687
rect 33241 25653 33275 25687
rect 35541 25653 35575 25687
rect 26341 25449 26375 25483
rect 27905 25449 27939 25483
rect 29745 25449 29779 25483
rect 30481 25449 30515 25483
rect 30849 25449 30883 25483
rect 31125 25449 31159 25483
rect 32137 25449 32171 25483
rect 32965 25449 32999 25483
rect 26792 25381 26826 25415
rect 28457 25381 28491 25415
rect 28825 25381 28859 25415
rect 33416 25381 33450 25415
rect 24216 25313 24250 25347
rect 25973 25313 26007 25347
rect 30941 25313 30975 25347
rect 33149 25313 33183 25347
rect 23949 25245 23983 25279
rect 26525 25245 26559 25279
rect 29837 25245 29871 25279
rect 30021 25245 30055 25279
rect 29377 25177 29411 25211
rect 23857 25109 23891 25143
rect 25329 25109 25363 25143
rect 29193 25109 29227 25143
rect 31769 25109 31803 25143
rect 34529 25109 34563 25143
rect 35173 25109 35207 25143
rect 26525 24905 26559 24939
rect 26893 24905 26927 24939
rect 31217 24905 31251 24939
rect 33149 24905 33183 24939
rect 33517 24905 33551 24939
rect 27997 24769 28031 24803
rect 29101 24769 29135 24803
rect 29285 24769 29319 24803
rect 32229 24769 32263 24803
rect 32321 24769 32355 24803
rect 34253 24769 34287 24803
rect 35449 24769 35483 24803
rect 24501 24701 24535 24735
rect 28089 24701 28123 24735
rect 28733 24701 28767 24735
rect 33701 24701 33735 24735
rect 35357 24701 35391 24735
rect 35909 24701 35943 24735
rect 24746 24633 24780 24667
rect 29552 24633 29586 24667
rect 31585 24633 31619 24667
rect 32137 24633 32171 24667
rect 35265 24633 35299 24667
rect 23949 24565 23983 24599
rect 24317 24565 24351 24599
rect 25881 24565 25915 24599
rect 28273 24565 28307 24599
rect 30665 24565 30699 24599
rect 31769 24565 31803 24599
rect 33885 24565 33919 24599
rect 34621 24565 34655 24599
rect 34897 24565 34931 24599
rect 24041 24361 24075 24395
rect 25053 24361 25087 24395
rect 30113 24361 30147 24395
rect 30573 24361 30607 24395
rect 31769 24361 31803 24395
rect 35357 24361 35391 24395
rect 24501 24293 24535 24327
rect 24961 24225 24995 24259
rect 28448 24225 28482 24259
rect 30665 24225 30699 24259
rect 34233 24225 34267 24259
rect 25237 24157 25271 24191
rect 28181 24157 28215 24191
rect 33977 24157 34011 24191
rect 36461 24157 36495 24191
rect 24593 24089 24627 24123
rect 30849 24089 30883 24123
rect 29561 24021 29595 24055
rect 35909 24021 35943 24055
rect 24685 23817 24719 23851
rect 25329 23817 25363 23851
rect 28089 23817 28123 23851
rect 28641 23817 28675 23851
rect 30573 23817 30607 23851
rect 34253 23817 34287 23851
rect 35265 23817 35299 23851
rect 36829 23817 36863 23851
rect 24961 23749 24995 23783
rect 30849 23749 30883 23783
rect 29929 23681 29963 23715
rect 31033 23681 31067 23715
rect 33793 23681 33827 23715
rect 35449 23681 35483 23715
rect 29101 23613 29135 23647
rect 29653 23613 29687 23647
rect 31300 23613 31334 23647
rect 35716 23613 35750 23647
rect 29745 23545 29779 23579
rect 34621 23545 34655 23579
rect 28181 23477 28215 23511
rect 29285 23477 29319 23511
rect 32413 23477 32447 23511
rect 28917 23273 28951 23307
rect 29009 23273 29043 23307
rect 29653 23273 29687 23307
rect 29929 23273 29963 23307
rect 30205 23273 30239 23307
rect 31125 23273 31159 23307
rect 33333 23273 33367 23307
rect 34529 23273 34563 23307
rect 36369 23273 36403 23307
rect 33701 23205 33735 23239
rect 34897 23205 34931 23239
rect 35256 23205 35290 23239
rect 34989 23137 35023 23171
rect 29101 23069 29135 23103
rect 33793 23069 33827 23103
rect 33885 23069 33919 23103
rect 28549 23001 28583 23035
rect 24041 22933 24075 22967
rect 26801 22933 26835 22967
rect 36921 22933 36955 22967
rect 28181 22729 28215 22763
rect 28549 22729 28583 22763
rect 33057 22729 33091 22763
rect 34621 22729 34655 22763
rect 36461 22729 36495 22763
rect 36553 22729 36587 22763
rect 25973 22661 26007 22695
rect 33701 22661 33735 22695
rect 34989 22661 35023 22695
rect 26893 22593 26927 22627
rect 26985 22593 27019 22627
rect 29745 22593 29779 22627
rect 35633 22593 35667 22627
rect 37013 22593 37047 22627
rect 37105 22593 37139 22627
rect 23949 22525 23983 22559
rect 24205 22525 24239 22559
rect 29285 22525 29319 22559
rect 30021 22525 30055 22559
rect 36921 22525 36955 22559
rect 26801 22457 26835 22491
rect 34253 22457 34287 22491
rect 35357 22457 35391 22491
rect 36001 22457 36035 22491
rect 25329 22389 25363 22423
rect 26249 22389 26283 22423
rect 26433 22389 26467 22423
rect 29101 22389 29135 22423
rect 29747 22389 29781 22423
rect 31125 22389 31159 22423
rect 33333 22389 33367 22423
rect 35449 22389 35483 22423
rect 28641 22185 28675 22219
rect 29745 22185 29779 22219
rect 32505 22185 32539 22219
rect 34161 22185 34195 22219
rect 36829 22185 36863 22219
rect 21465 22049 21499 22083
rect 22089 22049 22123 22083
rect 23949 22049 23983 22083
rect 24685 22049 24719 22083
rect 25697 22049 25731 22083
rect 26792 22049 26826 22083
rect 29285 22049 29319 22083
rect 30021 22049 30055 22083
rect 35081 22049 35115 22083
rect 21833 21981 21867 22015
rect 24777 21981 24811 22015
rect 24869 21981 24903 22015
rect 26525 21981 26559 22015
rect 32597 21981 32631 22015
rect 32689 21981 32723 22015
rect 34345 21981 34379 22015
rect 34668 21981 34702 22015
rect 34805 21981 34839 22015
rect 36185 21981 36219 22015
rect 29009 21913 29043 21947
rect 31953 21913 31987 21947
rect 23213 21845 23247 21879
rect 24317 21845 24351 21879
rect 25421 21845 25455 21879
rect 26157 21845 26191 21879
rect 27905 21845 27939 21879
rect 30205 21845 30239 21879
rect 30665 21845 30699 21879
rect 31033 21845 31067 21879
rect 32137 21845 32171 21879
rect 22385 21641 22419 21675
rect 23489 21641 23523 21675
rect 24409 21641 24443 21675
rect 26709 21641 26743 21675
rect 30113 21641 30147 21675
rect 30389 21641 30423 21675
rect 35909 21641 35943 21675
rect 21925 21505 21959 21539
rect 22753 21505 22787 21539
rect 23673 21505 23707 21539
rect 25329 21505 25363 21539
rect 30573 21505 30607 21539
rect 31033 21505 31067 21539
rect 35357 21505 35391 21539
rect 35541 21505 35575 21539
rect 36277 21505 36311 21539
rect 20913 21437 20947 21471
rect 21833 21437 21867 21471
rect 24869 21437 24903 21471
rect 25605 21437 25639 21471
rect 27629 21437 27663 21471
rect 31309 21437 31343 21471
rect 34345 21437 34379 21471
rect 36645 21437 36679 21471
rect 20361 21369 20395 21403
rect 21189 21369 21223 21403
rect 21741 21369 21775 21403
rect 27261 21369 27295 21403
rect 33517 21369 33551 21403
rect 34069 21369 34103 21403
rect 35265 21369 35299 21403
rect 21373 21301 21407 21335
rect 24777 21301 24811 21335
rect 25331 21301 25365 21335
rect 27813 21301 27847 21335
rect 31035 21301 31069 21335
rect 32413 21301 32447 21335
rect 32965 21301 32999 21335
rect 33333 21301 33367 21335
rect 34897 21301 34931 21335
rect 22293 21097 22327 21131
rect 24777 21097 24811 21131
rect 25697 21097 25731 21131
rect 26249 21097 26283 21131
rect 28457 21097 28491 21131
rect 29929 21097 29963 21131
rect 30941 21097 30975 21131
rect 32505 21097 32539 21131
rect 33885 21097 33919 21131
rect 23642 21029 23676 21063
rect 31953 21029 31987 21063
rect 34244 21029 34278 21063
rect 20913 20961 20947 20995
rect 21180 20961 21214 20995
rect 23397 20961 23431 20995
rect 26617 20961 26651 20995
rect 26940 20961 26974 20995
rect 30297 20961 30331 20995
rect 27077 20893 27111 20927
rect 27353 20893 27387 20927
rect 30389 20893 30423 20927
rect 30573 20893 30607 20927
rect 32597 20893 32631 20927
rect 32781 20893 32815 20927
rect 33977 20893 34011 20927
rect 32137 20825 32171 20859
rect 20085 20757 20119 20791
rect 25329 20757 25363 20791
rect 31493 20757 31527 20791
rect 35357 20757 35391 20791
rect 36001 20757 36035 20791
rect 19901 20553 19935 20587
rect 22293 20553 22327 20587
rect 23489 20553 23523 20587
rect 24869 20553 24903 20587
rect 26433 20553 26467 20587
rect 30757 20553 30791 20587
rect 31309 20553 31343 20587
rect 31677 20553 31711 20587
rect 34621 20553 34655 20587
rect 21925 20485 21959 20519
rect 29009 20485 29043 20519
rect 36645 20485 36679 20519
rect 19993 20417 20027 20451
rect 25053 20417 25087 20451
rect 28089 20417 28123 20451
rect 29377 20417 29411 20451
rect 32321 20417 32355 20451
rect 32597 20417 32631 20451
rect 20249 20349 20283 20383
rect 22477 20349 22511 20383
rect 23029 20349 23063 20383
rect 23673 20349 23707 20383
rect 24225 20349 24259 20383
rect 25320 20349 25354 20383
rect 27077 20349 27111 20383
rect 31861 20349 31895 20383
rect 32184 20349 32218 20383
rect 35265 20349 35299 20383
rect 27445 20281 27479 20315
rect 27905 20281 27939 20315
rect 29622 20281 29656 20315
rect 35532 20281 35566 20315
rect 21373 20213 21407 20247
rect 22661 20213 22695 20247
rect 23857 20213 23891 20247
rect 27537 20213 27571 20247
rect 27997 20213 28031 20247
rect 28549 20213 28583 20247
rect 33701 20213 33735 20247
rect 34345 20213 34379 20247
rect 35081 20213 35115 20247
rect 19717 20009 19751 20043
rect 20913 20009 20947 20043
rect 21281 20009 21315 20043
rect 23489 20009 23523 20043
rect 23765 20009 23799 20043
rect 24133 20009 24167 20043
rect 24225 20009 24259 20043
rect 25145 20009 25179 20043
rect 25421 20009 25455 20043
rect 26341 20009 26375 20043
rect 28457 20009 28491 20043
rect 29469 20009 29503 20043
rect 29837 20009 29871 20043
rect 29929 20009 29963 20043
rect 30389 20009 30423 20043
rect 30757 20009 30791 20043
rect 31585 20009 31619 20043
rect 31861 20009 31895 20043
rect 33701 20009 33735 20043
rect 27344 19941 27378 19975
rect 35072 19941 35106 19975
rect 18593 19873 18627 19907
rect 22477 19873 22511 19907
rect 26801 19873 26835 19907
rect 32588 19873 32622 19907
rect 18337 19805 18371 19839
rect 21373 19805 21407 19839
rect 21557 19805 21591 19839
rect 24317 19805 24351 19839
rect 27077 19805 27111 19839
rect 32321 19805 32355 19839
rect 34805 19805 34839 19839
rect 16497 19669 16531 19703
rect 16865 19669 16899 19703
rect 18153 19669 18187 19703
rect 20637 19669 20671 19703
rect 22661 19669 22695 19703
rect 36185 19669 36219 19703
rect 20453 19465 20487 19499
rect 21557 19465 21591 19499
rect 21925 19465 21959 19499
rect 24225 19465 24259 19499
rect 25053 19465 25087 19499
rect 26709 19465 26743 19499
rect 27721 19465 27755 19499
rect 28089 19465 28123 19499
rect 31861 19465 31895 19499
rect 32689 19465 32723 19499
rect 32965 19465 32999 19499
rect 34621 19465 34655 19499
rect 36093 19465 36127 19499
rect 16957 19329 16991 19363
rect 17877 19329 17911 19363
rect 18061 19329 18095 19363
rect 21189 19329 21223 19363
rect 23949 19329 23983 19363
rect 25605 19329 25639 19363
rect 26249 19329 26283 19363
rect 27353 19329 27387 19363
rect 16773 19261 16807 19295
rect 20085 19261 20119 19295
rect 20913 19261 20947 19295
rect 22201 19261 22235 19295
rect 22753 19261 22787 19295
rect 25421 19261 25455 19295
rect 25513 19261 25547 19295
rect 27169 19261 27203 19295
rect 16313 19193 16347 19227
rect 16865 19193 16899 19227
rect 18328 19193 18362 19227
rect 21005 19193 21039 19227
rect 26617 19193 26651 19227
rect 27077 19193 27111 19227
rect 33885 19329 33919 19363
rect 35633 19329 35667 19363
rect 33149 19261 33183 19295
rect 33701 19261 33735 19295
rect 34345 19261 34379 19295
rect 35541 19193 35575 19227
rect 15853 19125 15887 19159
rect 16405 19125 16439 19159
rect 19441 19125 19475 19159
rect 20545 19125 20579 19159
rect 22385 19125 22419 19159
rect 23121 19125 23155 19159
rect 24961 19125 24995 19159
rect 32321 19125 32355 19159
rect 32965 19125 32999 19159
rect 33241 19125 33275 19159
rect 33609 19125 33643 19159
rect 35081 19125 35115 19159
rect 35449 19125 35483 19159
rect 15669 18921 15703 18955
rect 18705 18921 18739 18955
rect 20637 18921 20671 18955
rect 21281 18921 21315 18955
rect 23765 18921 23799 18955
rect 25053 18921 25087 18955
rect 27537 18921 27571 18955
rect 33241 18921 33275 18955
rect 33701 18921 33735 18955
rect 35173 18921 35207 18955
rect 35265 18921 35299 18955
rect 35725 18921 35759 18955
rect 9956 18853 9990 18887
rect 18337 18853 18371 18887
rect 20913 18853 20947 18887
rect 27169 18853 27203 18887
rect 16385 18785 16419 18819
rect 19625 18785 19659 18819
rect 21097 18785 21131 18819
rect 22109 18785 22143 18819
rect 9689 18717 9723 18751
rect 16129 18717 16163 18751
rect 19717 18717 19751 18751
rect 19901 18717 19935 18751
rect 32137 18717 32171 18751
rect 19257 18649 19291 18683
rect 21649 18649 21683 18683
rect 22293 18649 22327 18683
rect 11069 18581 11103 18615
rect 14933 18581 14967 18615
rect 15945 18581 15979 18615
rect 17509 18581 17543 18615
rect 22017 18581 22051 18615
rect 26801 18581 26835 18615
rect 30665 18581 30699 18615
rect 32689 18581 32723 18615
rect 7389 18377 7423 18411
rect 10057 18377 10091 18411
rect 14841 18377 14875 18411
rect 17877 18377 17911 18411
rect 19441 18377 19475 18411
rect 20545 18377 20579 18411
rect 20913 18377 20947 18411
rect 21373 18377 21407 18411
rect 26525 18377 26559 18411
rect 32045 18377 32079 18411
rect 26709 18309 26743 18343
rect 30573 18309 30607 18343
rect 15485 18241 15519 18275
rect 16957 18241 16991 18275
rect 18061 18241 18095 18275
rect 21833 18241 21867 18275
rect 22017 18241 22051 18275
rect 26249 18241 26283 18275
rect 27261 18241 27295 18275
rect 31125 18241 31159 18275
rect 32781 18241 32815 18275
rect 7573 18173 7607 18207
rect 7829 18173 7863 18207
rect 14749 18173 14783 18207
rect 15301 18173 15335 18207
rect 16773 18173 16807 18207
rect 16865 18173 16899 18207
rect 27169 18173 27203 18207
rect 32505 18173 32539 18207
rect 17417 18105 17451 18139
rect 18306 18105 18340 18139
rect 19993 18105 20027 18139
rect 27077 18105 27111 18139
rect 30481 18105 30515 18139
rect 30941 18105 30975 18139
rect 8953 18037 8987 18071
rect 9689 18037 9723 18071
rect 15209 18037 15243 18071
rect 16221 18037 16255 18071
rect 16405 18037 16439 18071
rect 21741 18037 21775 18071
rect 22477 18037 22511 18071
rect 22845 18037 22879 18071
rect 24409 18037 24443 18071
rect 30021 18037 30055 18071
rect 31033 18037 31067 18071
rect 31585 18037 31619 18071
rect 32137 18037 32171 18071
rect 32597 18037 32631 18071
rect 14933 17833 14967 17867
rect 15577 17833 15611 17867
rect 17877 17833 17911 17867
rect 18797 17833 18831 17867
rect 19165 17833 19199 17867
rect 19533 17833 19567 17867
rect 23029 17833 23063 17867
rect 30941 17833 30975 17867
rect 33517 17833 33551 17867
rect 20637 17765 20671 17799
rect 32382 17765 32416 17799
rect 16764 17697 16798 17731
rect 18981 17697 19015 17731
rect 21649 17697 21683 17731
rect 22845 17697 22879 17731
rect 24685 17697 24719 17731
rect 28320 17697 28354 17731
rect 28733 17697 28767 17731
rect 35449 17697 35483 17731
rect 16497 17629 16531 17663
rect 19993 17629 20027 17663
rect 21741 17629 21775 17663
rect 21925 17629 21959 17663
rect 24777 17629 24811 17663
rect 24869 17629 24903 17663
rect 26617 17629 26651 17663
rect 27997 17629 28031 17663
rect 28457 17629 28491 17663
rect 32137 17629 32171 17663
rect 7665 17561 7699 17595
rect 23765 17561 23799 17595
rect 24317 17561 24351 17595
rect 30757 17561 30791 17595
rect 35633 17561 35667 17595
rect 8401 17493 8435 17527
rect 16221 17493 16255 17527
rect 18429 17493 18463 17527
rect 21189 17493 21223 17527
rect 21281 17493 21315 17527
rect 24133 17493 24167 17527
rect 29837 17493 29871 17527
rect 30389 17493 30423 17527
rect 16865 17289 16899 17323
rect 19809 17289 19843 17323
rect 22017 17289 22051 17323
rect 23673 17289 23707 17323
rect 24961 17289 24995 17323
rect 26985 17289 27019 17323
rect 28457 17289 28491 17323
rect 32137 17289 32171 17323
rect 33057 17289 33091 17323
rect 33241 17289 33275 17323
rect 35449 17289 35483 17323
rect 18061 17221 18095 17255
rect 19073 17221 19107 17255
rect 23397 17221 23431 17255
rect 25421 17221 25455 17255
rect 30021 17221 30055 17255
rect 30113 17221 30147 17255
rect 18705 17153 18739 17187
rect 21465 17153 21499 17187
rect 21557 17153 21591 17187
rect 24133 17153 24167 17187
rect 24225 17153 24259 17187
rect 25605 17153 25639 17187
rect 29837 17153 29871 17187
rect 8217 17085 8251 17119
rect 8401 17085 8435 17119
rect 15393 17085 15427 17119
rect 15485 17085 15519 17119
rect 15752 17085 15786 17119
rect 19625 17085 19659 17119
rect 20177 17085 20211 17119
rect 8646 17017 8680 17051
rect 17785 17017 17819 17051
rect 18521 17017 18555 17051
rect 23121 17017 23155 17051
rect 24041 17017 24075 17051
rect 25850 17017 25884 17051
rect 28733 17017 28767 17051
rect 30757 17153 30791 17187
rect 33701 17153 33735 17187
rect 33885 17153 33919 17187
rect 30297 17085 30331 17119
rect 31033 17085 31067 17119
rect 33609 17085 33643 17119
rect 34253 17085 34287 17119
rect 9781 16949 9815 16983
rect 17417 16949 17451 16983
rect 18429 16949 18463 16983
rect 20821 16949 20855 16983
rect 21005 16949 21039 16983
rect 21373 16949 21407 16983
rect 22385 16949 22419 16983
rect 27721 16949 27755 16983
rect 27997 16949 28031 16983
rect 30021 16949 30055 16983
rect 30759 16949 30793 16983
rect 32781 16949 32815 16983
rect 5457 16745 5491 16779
rect 8033 16745 8067 16779
rect 8401 16745 8435 16779
rect 11069 16745 11103 16779
rect 15301 16745 15335 16779
rect 15669 16745 15703 16779
rect 16497 16745 16531 16779
rect 18245 16745 18279 16779
rect 23029 16745 23063 16779
rect 23489 16745 23523 16779
rect 25697 16745 25731 16779
rect 27905 16745 27939 16779
rect 29377 16745 29411 16779
rect 30941 16745 30975 16779
rect 31493 16745 31527 16779
rect 31677 16745 31711 16779
rect 31953 16745 31987 16779
rect 34069 16745 34103 16779
rect 5917 16677 5951 16711
rect 7941 16677 7975 16711
rect 8493 16677 8527 16711
rect 21342 16677 21376 16711
rect 29828 16677 29862 16711
rect 5825 16609 5859 16643
rect 9956 16609 9990 16643
rect 17121 16609 17155 16643
rect 20637 16609 20671 16643
rect 23581 16609 23615 16643
rect 23848 16609 23882 16643
rect 26781 16609 26815 16643
rect 29561 16609 29595 16643
rect 4997 16541 5031 16575
rect 6009 16541 6043 16575
rect 8585 16541 8619 16575
rect 9689 16541 9723 16575
rect 15761 16541 15795 16575
rect 15945 16541 15979 16575
rect 16865 16541 16899 16575
rect 21097 16541 21131 16575
rect 26525 16541 26559 16575
rect 32137 16609 32171 16643
rect 32404 16609 32438 16643
rect 5365 16405 5399 16439
rect 7205 16405 7239 16439
rect 7481 16405 7515 16439
rect 18797 16405 18831 16439
rect 22477 16405 22511 16439
rect 24961 16405 24995 16439
rect 31677 16405 31711 16439
rect 33517 16405 33551 16439
rect 4905 16201 4939 16235
rect 8493 16201 8527 16235
rect 10057 16201 10091 16235
rect 10701 16201 10735 16235
rect 15393 16201 15427 16235
rect 15761 16201 15795 16235
rect 16405 16201 16439 16235
rect 17693 16201 17727 16235
rect 20637 16201 20671 16235
rect 20913 16201 20947 16235
rect 22477 16201 22511 16235
rect 23949 16201 23983 16235
rect 24409 16201 24443 16235
rect 24685 16201 24719 16235
rect 26249 16201 26283 16235
rect 27169 16201 27203 16235
rect 29377 16201 29411 16235
rect 30389 16201 30423 16235
rect 30757 16201 30791 16235
rect 32321 16201 32355 16235
rect 33241 16201 33275 16235
rect 15025 16133 15059 16167
rect 4445 16065 4479 16099
rect 5549 16065 5583 16099
rect 7573 16065 7607 16099
rect 7665 16065 7699 16099
rect 8217 16065 8251 16099
rect 17049 16065 17083 16099
rect 7481 15997 7515 16031
rect 8677 15997 8711 16031
rect 8944 15997 8978 16031
rect 5365 15929 5399 15963
rect 16313 15929 16347 15963
rect 16865 15929 16899 15963
rect 26801 16133 26835 16167
rect 27353 16133 27387 16167
rect 18061 16065 18095 16099
rect 21097 16065 21131 16099
rect 24869 16065 24903 16099
rect 27905 16065 27939 16099
rect 28365 16065 28399 16099
rect 29101 16065 29135 16099
rect 29837 16065 29871 16099
rect 30021 16065 30055 16099
rect 30941 16065 30975 16099
rect 18328 15997 18362 16031
rect 23489 15997 23523 16031
rect 23765 15997 23799 16031
rect 25136 15997 25170 16031
rect 27721 15997 27755 16031
rect 29745 15997 29779 16031
rect 20269 15929 20303 15963
rect 21342 15929 21376 15963
rect 27813 15929 27847 15963
rect 31186 15929 31220 15963
rect 4813 15861 4847 15895
rect 5273 15861 5307 15895
rect 6009 15861 6043 15895
rect 6285 15861 6319 15895
rect 7113 15861 7147 15895
rect 16773 15861 16807 15895
rect 17417 15861 17451 15895
rect 17693 15861 17727 15895
rect 17785 15861 17819 15895
rect 19441 15861 19475 15895
rect 32965 15861 32999 15895
rect 8493 15657 8527 15691
rect 9873 15657 9907 15691
rect 16129 15657 16163 15691
rect 16497 15657 16531 15691
rect 16957 15657 16991 15691
rect 18613 15657 18647 15691
rect 20729 15657 20763 15691
rect 22477 15657 22511 15691
rect 26341 15657 26375 15691
rect 27905 15657 27939 15691
rect 30021 15657 30055 15691
rect 33425 15657 33459 15691
rect 36553 15657 36587 15691
rect 7205 15589 7239 15623
rect 7941 15589 7975 15623
rect 17500 15589 17534 15623
rect 26792 15589 26826 15623
rect 5264 15521 5298 15555
rect 8401 15521 8435 15555
rect 21353 15521 21387 15555
rect 23949 15521 23983 15555
rect 24205 15521 24239 15555
rect 26525 15521 26559 15555
rect 30573 15521 30607 15555
rect 31309 15521 31343 15555
rect 31677 15521 31711 15555
rect 32137 15521 32171 15555
rect 32689 15521 32723 15555
rect 33241 15521 33275 15555
rect 35081 15521 35115 15555
rect 35440 15521 35474 15555
rect 4997 15453 5031 15487
rect 8677 15453 8711 15487
rect 17233 15453 17267 15487
rect 21097 15453 21131 15487
rect 30665 15453 30699 15487
rect 30849 15453 30883 15487
rect 35173 15453 35207 15487
rect 29653 15385 29687 15419
rect 4353 15317 4387 15351
rect 6377 15317 6411 15351
rect 7481 15317 7515 15351
rect 8033 15317 8067 15351
rect 14013 15317 14047 15351
rect 23673 15317 23707 15351
rect 25329 15317 25363 15351
rect 30205 15317 30239 15351
rect 32321 15317 32355 15351
rect 33793 15317 33827 15351
rect 7297 15113 7331 15147
rect 17601 15113 17635 15147
rect 20637 15113 20671 15147
rect 21005 15113 21039 15147
rect 23673 15113 23707 15147
rect 24777 15113 24811 15147
rect 26065 15113 26099 15147
rect 26525 15113 26559 15147
rect 26985 15113 27019 15147
rect 27445 15113 27479 15147
rect 29929 15113 29963 15147
rect 30573 15113 30607 15147
rect 30941 15113 30975 15147
rect 32413 15113 32447 15147
rect 25605 15045 25639 15079
rect 14565 14977 14599 15011
rect 21097 14977 21131 15011
rect 23489 14977 23523 15011
rect 24133 14977 24167 15011
rect 24225 14977 24259 15011
rect 30021 14977 30055 15011
rect 31033 14977 31067 15011
rect 4169 14909 4203 14943
rect 4261 14909 4295 14943
rect 6285 14909 6319 14943
rect 7665 14909 7699 14943
rect 7757 14909 7791 14943
rect 13461 14909 13495 14943
rect 23121 14909 23155 14943
rect 24041 14909 24075 14943
rect 25421 14909 25455 14943
rect 31300 14909 31334 14943
rect 33701 14909 33735 14943
rect 35173 14909 35207 14943
rect 4528 14841 4562 14875
rect 6653 14841 6687 14875
rect 8002 14841 8036 14875
rect 13829 14841 13863 14875
rect 14289 14841 14323 14875
rect 20269 14841 20303 14875
rect 21342 14841 21376 14875
rect 29561 14841 29595 14875
rect 35418 14841 35452 14875
rect 5641 14773 5675 14807
rect 9137 14773 9171 14807
rect 13921 14773 13955 14807
rect 14381 14773 14415 14807
rect 17233 14773 17267 14807
rect 22477 14773 22511 14807
rect 33241 14773 33275 14807
rect 33885 14773 33919 14807
rect 34253 14773 34287 14807
rect 34621 14773 34655 14807
rect 36553 14773 36587 14807
rect 7205 14569 7239 14603
rect 7849 14569 7883 14603
rect 8125 14569 8159 14603
rect 8861 14569 8895 14603
rect 14473 14569 14507 14603
rect 21097 14569 21131 14603
rect 21281 14569 21315 14603
rect 21741 14569 21775 14603
rect 24041 14569 24075 14603
rect 24317 14569 24351 14603
rect 30389 14569 30423 14603
rect 31309 14569 31343 14603
rect 32137 14569 32171 14603
rect 32505 14569 32539 14603
rect 35909 14569 35943 14603
rect 36829 14569 36863 14603
rect 21649 14501 21683 14535
rect 4517 14433 4551 14467
rect 7113 14433 7147 14467
rect 8309 14433 8343 14467
rect 9873 14433 9907 14467
rect 12541 14433 12575 14467
rect 12797 14433 12831 14467
rect 29377 14433 29411 14467
rect 30849 14433 30883 14467
rect 31953 14501 31987 14535
rect 36461 14501 36495 14535
rect 32597 14433 32631 14467
rect 33701 14433 33735 14467
rect 35265 14433 35299 14467
rect 36645 14433 36679 14467
rect 4261 14365 4295 14399
rect 7389 14365 7423 14399
rect 11529 14365 11563 14399
rect 21925 14365 21959 14399
rect 30941 14365 30975 14399
rect 31125 14365 31159 14399
rect 31309 14365 31343 14399
rect 31585 14365 31619 14399
rect 32781 14365 32815 14399
rect 34805 14365 34839 14399
rect 35357 14365 35391 14399
rect 35449 14365 35483 14399
rect 34897 14297 34931 14331
rect 5641 14229 5675 14263
rect 6745 14229 6779 14263
rect 8493 14229 8527 14263
rect 10057 14229 10091 14263
rect 10793 14229 10827 14263
rect 13921 14229 13955 14263
rect 19257 14229 19291 14263
rect 26985 14229 27019 14263
rect 29561 14229 29595 14263
rect 30481 14229 30515 14263
rect 33333 14229 33367 14263
rect 33885 14229 33919 14263
rect 34345 14229 34379 14263
rect 3525 14025 3559 14059
rect 3893 14025 3927 14059
rect 6561 14025 6595 14059
rect 7389 14025 7423 14059
rect 8309 14025 8343 14059
rect 10701 14025 10735 14059
rect 12633 14025 12667 14059
rect 16221 14025 16255 14059
rect 21373 14025 21407 14059
rect 22109 14025 22143 14059
rect 26709 14025 26743 14059
rect 29101 14025 29135 14059
rect 29469 14025 29503 14059
rect 30573 14025 30607 14059
rect 31217 14025 31251 14059
rect 32321 14025 32355 14059
rect 36461 14025 36495 14059
rect 37105 14025 37139 14059
rect 6285 13957 6319 13991
rect 7021 13957 7055 13991
rect 7849 13957 7883 13991
rect 8401 13957 8435 13991
rect 10793 13957 10827 13991
rect 21649 13957 21683 13991
rect 25605 13957 25639 13991
rect 31033 13957 31067 13991
rect 33885 13957 33919 13991
rect 3157 13889 3191 13923
rect 8861 13889 8895 13923
rect 8953 13889 8987 13923
rect 11345 13889 11379 13923
rect 11805 13889 11839 13923
rect 12265 13889 12299 13923
rect 13277 13889 13311 13923
rect 13461 13889 13495 13923
rect 13921 13889 13955 13923
rect 14887 13889 14921 13923
rect 19717 13889 19751 13923
rect 26433 13889 26467 13923
rect 27445 13889 27479 13923
rect 31677 13889 31711 13923
rect 31769 13889 31803 13923
rect 33425 13889 33459 13923
rect 34345 13889 34379 13923
rect 3985 13821 4019 13855
rect 4241 13821 4275 13855
rect 6837 13821 6871 13855
rect 9413 13821 9447 13855
rect 9873 13821 9907 13855
rect 11161 13821 11195 13855
rect 14381 13821 14415 13855
rect 15117 13821 15151 13855
rect 18613 13821 18647 13855
rect 19073 13821 19107 13855
rect 19625 13821 19659 13855
rect 25789 13821 25823 13855
rect 27261 13821 27295 13855
rect 28733 13821 28767 13855
rect 29285 13821 29319 13855
rect 30205 13821 30239 13855
rect 31585 13821 31619 13855
rect 35081 13821 35115 13855
rect 35348 13821 35382 13855
rect 8769 13753 8803 13787
rect 19533 13753 19567 13787
rect 25513 13753 25547 13787
rect 27353 13753 27387 13787
rect 32689 13753 32723 13787
rect 33241 13753 33275 13787
rect 5365 13685 5399 13719
rect 11253 13685 11287 13719
rect 12817 13685 12851 13719
rect 13185 13685 13219 13719
rect 14197 13685 14231 13719
rect 14843 13685 14877 13719
rect 19165 13685 19199 13719
rect 26893 13685 26927 13719
rect 32781 13685 32815 13719
rect 33149 13685 33183 13719
rect 34713 13685 34747 13719
rect 4261 13481 4295 13515
rect 5089 13481 5123 13515
rect 6929 13481 6963 13515
rect 8309 13481 8343 13515
rect 9689 13481 9723 13515
rect 10057 13481 10091 13515
rect 10885 13481 10919 13515
rect 12633 13481 12667 13515
rect 13553 13481 13587 13515
rect 14105 13481 14139 13515
rect 16681 13481 16715 13515
rect 18521 13481 18555 13515
rect 18981 13481 19015 13515
rect 27905 13481 27939 13515
rect 29009 13481 29043 13515
rect 29469 13481 29503 13515
rect 30757 13481 30791 13515
rect 31309 13481 31343 13515
rect 31953 13481 31987 13515
rect 32413 13481 32447 13515
rect 32873 13481 32907 13515
rect 33793 13481 33827 13515
rect 34897 13481 34931 13515
rect 36553 13481 36587 13515
rect 26770 13413 26804 13447
rect 33241 13413 33275 13447
rect 33701 13413 33735 13447
rect 4997 13345 5031 13379
rect 8493 13345 8527 13379
rect 9505 13345 9539 13379
rect 11509 13345 11543 13379
rect 15557 13345 15591 13379
rect 18153 13345 18187 13379
rect 21925 13345 21959 13379
rect 22192 13345 22226 13379
rect 26525 13345 26559 13379
rect 29377 13345 29411 13379
rect 30573 13345 30607 13379
rect 32229 13345 32263 13379
rect 34345 13345 34379 13379
rect 34805 13345 34839 13379
rect 35265 13345 35299 13379
rect 5273 13277 5307 13311
rect 10149 13277 10183 13311
rect 10333 13277 10367 13311
rect 11260 13277 11294 13311
rect 15301 13277 15335 13311
rect 19073 13277 19107 13311
rect 19165 13277 19199 13311
rect 29561 13277 29595 13311
rect 33977 13277 34011 13311
rect 35357 13277 35391 13311
rect 35449 13277 35483 13311
rect 8677 13209 8711 13243
rect 28917 13209 28951 13243
rect 33333 13209 33367 13243
rect 4629 13141 4663 13175
rect 7389 13141 7423 13175
rect 13277 13141 13311 13175
rect 14657 13141 14691 13175
rect 18613 13141 18647 13175
rect 21833 13141 21867 13175
rect 23305 13141 23339 13175
rect 30481 13141 30515 13175
rect 36001 13141 36035 13175
rect 3801 12937 3835 12971
rect 5273 12937 5307 12971
rect 6561 12937 6595 12971
rect 9045 12937 9079 12971
rect 11253 12937 11287 12971
rect 12173 12937 12207 12971
rect 15761 12937 15795 12971
rect 19441 12937 19475 12971
rect 25697 12937 25731 12971
rect 26525 12937 26559 12971
rect 30849 12937 30883 12971
rect 32229 12937 32263 12971
rect 32597 12937 32631 12971
rect 36553 12937 36587 12971
rect 9781 12869 9815 12903
rect 19993 12869 20027 12903
rect 29285 12869 29319 12903
rect 30297 12869 30331 12903
rect 3433 12801 3467 12835
rect 7849 12801 7883 12835
rect 9873 12801 9907 12835
rect 16313 12801 16347 12835
rect 16773 12801 16807 12835
rect 18061 12801 18095 12835
rect 26617 12801 26651 12835
rect 29837 12801 29871 12835
rect 31401 12801 31435 12835
rect 33241 12801 33275 12835
rect 3893 12733 3927 12767
rect 4160 12733 4194 12767
rect 7665 12733 7699 12767
rect 8585 12733 8619 12767
rect 11805 12733 11839 12767
rect 13093 12733 13127 12767
rect 13277 12733 13311 12767
rect 15301 12733 15335 12767
rect 16129 12733 16163 12767
rect 20453 12733 20487 12767
rect 20545 12733 20579 12767
rect 22477 12733 22511 12767
rect 35173 12733 35207 12767
rect 35440 12733 35474 12767
rect 7205 12665 7239 12699
rect 7757 12665 7791 12699
rect 9413 12665 9447 12699
rect 10118 12665 10152 12699
rect 12817 12665 12851 12699
rect 13522 12665 13556 12699
rect 18306 12665 18340 12699
rect 20790 12665 20824 12699
rect 22845 12665 22879 12699
rect 24317 12665 24351 12699
rect 24409 12665 24443 12699
rect 26884 12665 26918 12699
rect 28733 12665 28767 12699
rect 29653 12665 29687 12699
rect 30757 12665 30791 12699
rect 31309 12665 31343 12699
rect 32965 12665 32999 12699
rect 33609 12665 33643 12699
rect 5825 12597 5859 12631
rect 7297 12597 7331 12631
rect 14657 12597 14691 12631
rect 16221 12597 16255 12631
rect 17785 12597 17819 12631
rect 21925 12597 21959 12631
rect 27997 12597 28031 12631
rect 29009 12597 29043 12631
rect 29745 12597 29779 12631
rect 31217 12597 31251 12631
rect 31953 12597 31987 12631
rect 33057 12597 33091 12631
rect 34345 12597 34379 12631
rect 34713 12597 34747 12631
rect 4721 12393 4755 12427
rect 5641 12393 5675 12427
rect 9413 12393 9447 12427
rect 9689 12393 9723 12427
rect 12725 12393 12759 12427
rect 13645 12393 13679 12427
rect 16221 12393 16255 12427
rect 16681 12393 16715 12427
rect 20637 12393 20671 12427
rect 26801 12393 26835 12427
rect 27445 12393 27479 12427
rect 29561 12393 29595 12427
rect 29929 12393 29963 12427
rect 30113 12393 30147 12427
rect 31585 12393 31619 12427
rect 31861 12393 31895 12427
rect 32597 12393 32631 12427
rect 33057 12393 33091 12427
rect 33425 12393 33459 12427
rect 33517 12393 33551 12427
rect 34621 12393 34655 12427
rect 36553 12393 36587 12427
rect 4997 12325 5031 12359
rect 11437 12325 11471 12359
rect 15853 12325 15887 12359
rect 17049 12325 17083 12359
rect 18512 12325 18546 12359
rect 21465 12325 21499 12359
rect 22928 12325 22962 12359
rect 27077 12325 27111 12359
rect 27896 12325 27930 12359
rect 4353 12257 4387 12291
rect 5549 12257 5583 12291
rect 6745 12257 6779 12291
rect 8401 12257 8435 12291
rect 10057 12257 10091 12291
rect 11253 12257 11287 12291
rect 13553 12257 13587 12291
rect 15301 12257 15335 12291
rect 30481 12257 30515 12291
rect 32413 12257 32447 12291
rect 33885 12257 33919 12291
rect 35440 12257 35474 12291
rect 5825 12189 5859 12223
rect 8493 12189 8527 12223
rect 8677 12189 8711 12223
rect 10149 12189 10183 12223
rect 10333 12189 10367 12223
rect 13093 12189 13127 12223
rect 13737 12189 13771 12223
rect 17141 12189 17175 12223
rect 17325 12189 17359 12223
rect 18245 12189 18279 12223
rect 21557 12189 21591 12223
rect 21741 12189 21775 12223
rect 22661 12189 22695 12223
rect 27629 12189 27663 12223
rect 30573 12189 30607 12223
rect 30665 12189 30699 12223
rect 33977 12189 34011 12223
rect 34161 12189 34195 12223
rect 35173 12189 35207 12223
rect 5181 12121 5215 12155
rect 7297 12121 7331 12155
rect 29009 12121 29043 12155
rect 6929 12053 6963 12087
rect 7665 12053 7699 12087
rect 8033 12053 8067 12087
rect 9045 12053 9079 12087
rect 10793 12053 10827 12087
rect 11621 12053 11655 12087
rect 13185 12053 13219 12087
rect 15025 12053 15059 12087
rect 18153 12053 18187 12087
rect 19625 12053 19659 12087
rect 21097 12053 21131 12087
rect 22201 12053 22235 12087
rect 22569 12053 22603 12087
rect 24041 12053 24075 12087
rect 31125 12053 31159 12087
rect 34989 12053 35023 12087
rect 3893 11849 3927 11883
rect 6837 11849 6871 11883
rect 8033 11849 8067 11883
rect 8953 11849 8987 11883
rect 10425 11849 10459 11883
rect 11621 11849 11655 11883
rect 12725 11849 12759 11883
rect 16773 11849 16807 11883
rect 17141 11849 17175 11883
rect 20637 11849 20671 11883
rect 21281 11849 21315 11883
rect 21741 11849 21775 11883
rect 23029 11849 23063 11883
rect 23397 11849 23431 11883
rect 26617 11849 26651 11883
rect 28089 11849 28123 11883
rect 31401 11849 31435 11883
rect 32321 11849 32355 11883
rect 33609 11849 33643 11883
rect 36277 11849 36311 11883
rect 36829 11849 36863 11883
rect 3525 11713 3559 11747
rect 7481 11713 7515 11747
rect 12265 11713 12299 11747
rect 22569 11713 22603 11747
rect 23673 11713 23707 11747
rect 26709 11713 26743 11747
rect 32965 11713 32999 11747
rect 33977 11713 34011 11747
rect 34345 11713 34379 11747
rect 3985 11645 4019 11679
rect 4252 11645 4286 11679
rect 9045 11645 9079 11679
rect 13185 11645 13219 11679
rect 13452 11645 13486 11679
rect 19257 11645 19291 11679
rect 21925 11645 21959 11679
rect 23940 11645 23974 11679
rect 28917 11645 28951 11679
rect 29285 11645 29319 11679
rect 34897 11645 34931 11679
rect 6653 11577 6687 11611
rect 7297 11577 7331 11611
rect 9312 11577 9346 11611
rect 13001 11577 13035 11611
rect 19073 11577 19107 11611
rect 19502 11577 19536 11611
rect 21649 11577 21683 11611
rect 22477 11577 22511 11611
rect 26954 11577 26988 11611
rect 28733 11577 28767 11611
rect 29552 11577 29586 11611
rect 32229 11577 32263 11611
rect 32781 11577 32815 11611
rect 35164 11577 35198 11611
rect 5365 11509 5399 11543
rect 6285 11509 6319 11543
rect 7205 11509 7239 11543
rect 8401 11509 8435 11543
rect 11345 11509 11379 11543
rect 14565 11509 14599 11543
rect 17509 11509 17543 11543
rect 18245 11509 18279 11543
rect 18705 11509 18739 11543
rect 22017 11509 22051 11543
rect 22385 11509 22419 11543
rect 25053 11509 25087 11543
rect 28917 11509 28951 11543
rect 29009 11509 29043 11543
rect 30665 11509 30699 11543
rect 31861 11509 31895 11543
rect 32689 11509 32723 11543
rect 34621 11509 34655 11543
rect 4721 11305 4755 11339
rect 5181 11305 5215 11339
rect 5733 11305 5767 11339
rect 6193 11305 6227 11339
rect 9505 11305 9539 11339
rect 11069 11305 11103 11339
rect 14105 11305 14139 11339
rect 19257 11305 19291 11339
rect 19809 11305 19843 11339
rect 21741 11305 21775 11339
rect 22661 11305 22695 11339
rect 23397 11305 23431 11339
rect 26801 11305 26835 11339
rect 27629 11305 27663 11339
rect 28089 11305 28123 11339
rect 29561 11305 29595 11339
rect 30481 11305 30515 11339
rect 30849 11305 30883 11339
rect 33517 11305 33551 11339
rect 36001 11305 36035 11339
rect 6552 11237 6586 11271
rect 8309 11237 8343 11271
rect 21649 11237 21683 11271
rect 23756 11237 23790 11271
rect 28448 11237 28482 11271
rect 30205 11237 30239 11271
rect 32404 11237 32438 11271
rect 34866 11237 34900 11271
rect 4629 11169 4663 11203
rect 5089 11169 5123 11203
rect 9956 11169 9990 11203
rect 12981 11169 13015 11203
rect 17877 11169 17911 11203
rect 18144 11169 18178 11203
rect 21189 11169 21223 11203
rect 28181 11169 28215 11203
rect 5273 11101 5307 11135
rect 6285 11101 6319 11135
rect 9689 11101 9723 11135
rect 12725 11101 12759 11135
rect 21833 11101 21867 11135
rect 23489 11101 23523 11135
rect 32137 11101 32171 11135
rect 34621 11101 34655 11135
rect 7665 11033 7699 11067
rect 8677 11033 8711 11067
rect 20637 11033 20671 11067
rect 24869 11033 24903 11067
rect 34161 11033 34195 11067
rect 9045 10965 9079 10999
rect 21281 10965 21315 10999
rect 23029 10965 23063 10999
rect 3801 10761 3835 10795
rect 4077 10761 4111 10795
rect 5641 10761 5675 10795
rect 7297 10761 7331 10795
rect 9597 10761 9631 10795
rect 10149 10761 10183 10795
rect 10517 10761 10551 10795
rect 17141 10761 17175 10795
rect 19441 10761 19475 10795
rect 21005 10761 21039 10795
rect 21281 10761 21315 10795
rect 23029 10761 23063 10795
rect 23397 10761 23431 10795
rect 28181 10761 28215 10795
rect 28641 10761 28675 10795
rect 31585 10761 31619 10795
rect 33517 10761 33551 10795
rect 34621 10761 34655 10795
rect 35081 10761 35115 10795
rect 6377 10693 6411 10727
rect 8125 10693 8159 10727
rect 11345 10693 11379 10727
rect 13185 10693 13219 10727
rect 29469 10693 29503 10727
rect 35633 10693 35667 10727
rect 4261 10625 4295 10659
rect 8217 10625 8251 10659
rect 12725 10625 12759 10659
rect 14197 10625 14231 10659
rect 22569 10625 22603 10659
rect 29653 10625 29687 10659
rect 7113 10557 7147 10591
rect 7665 10557 7699 10591
rect 8484 10557 8518 10591
rect 11161 10557 11195 10591
rect 11713 10557 11747 10591
rect 13737 10557 13771 10591
rect 14473 10557 14507 10591
rect 17785 10557 17819 10591
rect 18061 10557 18095 10591
rect 21925 10557 21959 10591
rect 22477 10557 22511 10591
rect 23673 10557 23707 10591
rect 23940 10557 23974 10591
rect 29920 10557 29954 10591
rect 32137 10557 32171 10591
rect 35449 10557 35483 10591
rect 36001 10557 36035 10591
rect 4528 10489 4562 10523
rect 17417 10489 17451 10523
rect 18306 10489 18340 10523
rect 29101 10489 29135 10523
rect 32404 10489 32438 10523
rect 12265 10421 12299 10455
rect 13645 10421 13679 10455
rect 14199 10421 14233 10455
rect 15577 10421 15611 10455
rect 20637 10421 20671 10455
rect 22017 10421 22051 10455
rect 22385 10421 22419 10455
rect 25053 10421 25087 10455
rect 31033 10421 31067 10455
rect 32045 10421 32079 10455
rect 4353 10217 4387 10251
rect 4813 10217 4847 10251
rect 6469 10217 6503 10251
rect 7021 10217 7055 10251
rect 7941 10217 7975 10251
rect 8401 10217 8435 10251
rect 9873 10217 9907 10251
rect 10977 10217 11011 10251
rect 23213 10217 23247 10251
rect 29653 10217 29687 10251
rect 30113 10217 30147 10251
rect 32413 10217 32447 10251
rect 32689 10217 32723 10251
rect 34345 10217 34379 10251
rect 5356 10149 5390 10183
rect 12992 10149 13026 10183
rect 22109 10149 22143 10183
rect 23572 10149 23606 10183
rect 33232 10149 33266 10183
rect 5089 10081 5123 10115
rect 8309 10081 8343 10115
rect 9689 10081 9723 10115
rect 10793 10081 10827 10115
rect 12725 10081 12759 10115
rect 17121 10081 17155 10115
rect 19349 10081 19383 10115
rect 20913 10081 20947 10115
rect 30021 10081 30055 10115
rect 35449 10081 35483 10115
rect 8585 10013 8619 10047
rect 16865 10013 16899 10047
rect 23305 10013 23339 10047
rect 30205 10013 30239 10047
rect 32965 10013 32999 10047
rect 35633 9945 35667 9979
rect 14105 9877 14139 9911
rect 14657 9877 14691 9911
rect 16497 9877 16531 9911
rect 18245 9877 18279 9911
rect 18797 9877 18831 9911
rect 19533 9877 19567 9911
rect 21097 9877 21131 9911
rect 21557 9877 21591 9911
rect 22477 9877 22511 9911
rect 24685 9877 24719 9911
rect 5089 9673 5123 9707
rect 5457 9673 5491 9707
rect 9229 9673 9263 9707
rect 10885 9673 10919 9707
rect 12725 9673 12759 9707
rect 14013 9673 14047 9707
rect 17417 9673 17451 9707
rect 19441 9673 19475 9707
rect 21005 9673 21039 9707
rect 23029 9673 23063 9707
rect 24685 9673 24719 9707
rect 30021 9673 30055 9707
rect 32965 9673 32999 9707
rect 33425 9673 33459 9707
rect 35449 9673 35483 9707
rect 7113 9605 7147 9639
rect 8217 9605 8251 9639
rect 12173 9605 12207 9639
rect 16313 9605 16347 9639
rect 23673 9605 23707 9639
rect 29745 9605 29779 9639
rect 30481 9605 30515 9639
rect 13461 9537 13495 9571
rect 15577 9537 15611 9571
rect 17049 9537 17083 9571
rect 17877 9537 17911 9571
rect 18521 9537 18555 9571
rect 18705 9537 18739 9571
rect 21373 9537 21407 9571
rect 21925 9537 21959 9571
rect 22017 9537 22051 9571
rect 24133 9537 24167 9571
rect 24317 9537 24351 9571
rect 25421 9537 25455 9571
rect 7205 9469 7239 9503
rect 8309 9469 8343 9503
rect 13277 9469 13311 9503
rect 14473 9469 14507 9503
rect 18429 9469 18463 9503
rect 20637 9469 20671 9503
rect 21833 9469 21867 9503
rect 11897 9401 11931 9435
rect 13369 9401 13403 9435
rect 14289 9401 14323 9435
rect 15945 9401 15979 9435
rect 16865 9401 16899 9435
rect 7389 9333 7423 9367
rect 7849 9333 7883 9367
rect 8493 9333 8527 9367
rect 8953 9333 8987 9367
rect 9781 9333 9815 9367
rect 12909 9333 12943 9367
rect 16405 9333 16439 9367
rect 16773 9333 16807 9367
rect 18061 9333 18095 9367
rect 21465 9333 21499 9367
rect 23305 9333 23339 9367
rect 24041 9333 24075 9367
rect 25053 9333 25087 9367
rect 13093 9129 13127 9163
rect 13461 9129 13495 9163
rect 13553 9129 13587 9163
rect 17601 9129 17635 9163
rect 18245 9129 18279 9163
rect 18613 9129 18647 9163
rect 19257 9129 19291 9163
rect 21373 9129 21407 9163
rect 24041 9129 24075 9163
rect 13001 9061 13035 9095
rect 16488 9061 16522 9095
rect 22928 9061 22962 9095
rect 7288 8993 7322 9027
rect 10517 8993 10551 9027
rect 10876 8993 10910 9027
rect 16221 8993 16255 9027
rect 21281 8993 21315 9027
rect 27997 8993 28031 9027
rect 28253 8993 28287 9027
rect 7021 8925 7055 8959
rect 10609 8925 10643 8959
rect 13645 8925 13679 8959
rect 19349 8925 19383 8959
rect 19533 8925 19567 8959
rect 21465 8925 21499 8959
rect 22661 8925 22695 8959
rect 6929 8789 6963 8823
rect 8401 8789 8435 8823
rect 11989 8789 12023 8823
rect 18889 8789 18923 8823
rect 19993 8789 20027 8823
rect 20913 8789 20947 8823
rect 25237 8789 25271 8823
rect 29377 8789 29411 8823
rect 11437 8585 11471 8619
rect 12173 8585 12207 8619
rect 14381 8585 14415 8619
rect 16405 8585 16439 8619
rect 17417 8585 17451 8619
rect 18245 8585 18279 8619
rect 18981 8585 19015 8619
rect 19349 8585 19383 8619
rect 20637 8585 20671 8619
rect 21281 8585 21315 8619
rect 23121 8585 23155 8619
rect 26617 8585 26651 8619
rect 28089 8585 28123 8619
rect 28641 8585 28675 8619
rect 8217 8517 8251 8551
rect 10425 8517 10459 8551
rect 13829 8517 13863 8551
rect 19625 8517 19659 8551
rect 20913 8517 20947 8551
rect 21649 8517 21683 8551
rect 10241 8449 10275 8483
rect 10885 8449 10919 8483
rect 10977 8449 11011 8483
rect 12449 8449 12483 8483
rect 17049 8449 17083 8483
rect 24685 8449 24719 8483
rect 25697 8449 25731 8483
rect 26709 8449 26743 8483
rect 6837 8381 6871 8415
rect 9965 8381 9999 8415
rect 10793 8381 10827 8415
rect 17785 8381 17819 8415
rect 18061 8381 18095 8415
rect 19441 8381 19475 8415
rect 20729 8381 20763 8415
rect 25513 8381 25547 8415
rect 7104 8313 7138 8347
rect 12694 8313 12728 8347
rect 14933 8313 14967 8347
rect 15577 8313 15611 8347
rect 15853 8313 15887 8347
rect 16865 8313 16899 8347
rect 20085 8313 20119 8347
rect 25053 8313 25087 8347
rect 25605 8313 25639 8347
rect 26954 8313 26988 8347
rect 6193 8245 6227 8279
rect 6561 8245 6595 8279
rect 9505 8245 9539 8279
rect 16313 8245 16347 8279
rect 16773 8245 16807 8279
rect 22753 8245 22787 8279
rect 25145 8245 25179 8279
rect 8309 8041 8343 8075
rect 12541 8041 12575 8075
rect 13553 8041 13587 8075
rect 16681 8041 16715 8075
rect 17325 8041 17359 8075
rect 17969 8041 18003 8075
rect 19625 8041 19659 8075
rect 21189 8041 21223 8075
rect 26893 8041 26927 8075
rect 27261 8041 27295 8075
rect 28089 8041 28123 8075
rect 5273 7973 5307 8007
rect 5724 7973 5758 8007
rect 12725 7973 12759 8007
rect 21732 7973 21766 8007
rect 23857 7973 23891 8007
rect 24194 7973 24228 8007
rect 26801 7973 26835 8007
rect 27353 7973 27387 8007
rect 29000 7973 29034 8007
rect 5457 7905 5491 7939
rect 10232 7905 10266 7939
rect 13277 7905 13311 7939
rect 15301 7905 15335 7939
rect 15557 7905 15591 7939
rect 17785 7905 17819 7939
rect 28733 7905 28767 7939
rect 7481 7837 7515 7871
rect 8401 7837 8435 7871
rect 8585 7837 8619 7871
rect 9965 7837 9999 7871
rect 13737 7837 13771 7871
rect 19717 7837 19751 7871
rect 19901 7837 19935 7871
rect 21465 7837 21499 7871
rect 23949 7837 23983 7871
rect 27445 7837 27479 7871
rect 18981 7769 19015 7803
rect 6837 7701 6871 7735
rect 7941 7701 7975 7735
rect 11345 7701 11379 7735
rect 19257 7701 19291 7735
rect 22845 7701 22879 7735
rect 25329 7701 25363 7735
rect 30113 7701 30147 7735
rect 7389 7497 7423 7531
rect 9597 7497 9631 7531
rect 10149 7497 10183 7531
rect 10517 7497 10551 7531
rect 17509 7497 17543 7531
rect 20821 7497 20855 7531
rect 21833 7497 21867 7531
rect 25329 7497 25363 7531
rect 25973 7497 26007 7531
rect 26341 7497 26375 7531
rect 27813 7497 27847 7531
rect 28457 7497 28491 7531
rect 28733 7497 28767 7531
rect 5089 7361 5123 7395
rect 5825 7361 5859 7395
rect 11161 7361 11195 7395
rect 11253 7361 11287 7395
rect 29285 7361 29319 7395
rect 4721 7293 4755 7327
rect 5549 7293 5583 7327
rect 5641 7293 5675 7327
rect 7941 7293 7975 7327
rect 8217 7293 8251 7327
rect 11713 7293 11747 7327
rect 12449 7293 12483 7327
rect 13001 7293 13035 7327
rect 13829 7293 13863 7327
rect 13921 7293 13955 7327
rect 16865 7293 16899 7327
rect 18705 7293 18739 7327
rect 18889 7293 18923 7327
rect 19156 7293 19190 7327
rect 21557 7293 21591 7327
rect 23121 7293 23155 7327
rect 23489 7293 23523 7327
rect 23949 7293 23983 7327
rect 26433 7293 26467 7327
rect 26689 7293 26723 7327
rect 29552 7293 29586 7327
rect 4353 7225 4387 7259
rect 7757 7225 7791 7259
rect 8462 7225 8496 7259
rect 11069 7225 11103 7259
rect 12081 7225 12115 7259
rect 13461 7225 13495 7259
rect 14166 7225 14200 7259
rect 15945 7225 15979 7259
rect 18337 7225 18371 7259
rect 24216 7225 24250 7259
rect 5181 7157 5215 7191
rect 6193 7157 6227 7191
rect 7941 7157 7975 7191
rect 8033 7157 8067 7191
rect 10701 7157 10735 7191
rect 12633 7157 12667 7191
rect 15301 7157 15335 7191
rect 17049 7157 17083 7191
rect 17877 7157 17911 7191
rect 20269 7157 20303 7191
rect 30665 7157 30699 7191
rect 7757 6953 7791 6987
rect 7849 6953 7883 6987
rect 8493 6953 8527 6987
rect 11713 6953 11747 6987
rect 14013 6953 14047 6987
rect 19993 6953 20027 6987
rect 27261 6953 27295 6987
rect 29193 6953 29227 6987
rect 24041 6885 24075 6919
rect 27629 6885 27663 6919
rect 5172 6817 5206 6851
rect 10333 6817 10367 6851
rect 10600 6817 10634 6851
rect 16957 6817 16991 6851
rect 17969 6817 18003 6851
rect 18317 6817 18351 6851
rect 20913 6817 20947 6851
rect 21097 6817 21131 6851
rect 23213 6817 23247 6851
rect 24133 6817 24167 6851
rect 25329 6817 25363 6851
rect 26617 6817 26651 6851
rect 28089 6817 28123 6851
rect 28825 6817 28859 6851
rect 29285 6817 29319 6851
rect 29552 6817 29586 6851
rect 4905 6749 4939 6783
rect 8033 6749 8067 6783
rect 13553 6749 13587 6783
rect 14105 6749 14139 6783
rect 14197 6749 14231 6783
rect 15485 6749 15519 6783
rect 15945 6749 15979 6783
rect 18061 6749 18095 6783
rect 21281 6749 21315 6783
rect 23581 6749 23615 6783
rect 24317 6749 24351 6783
rect 28181 6749 28215 6783
rect 28273 6749 28307 6783
rect 22845 6681 22879 6715
rect 25973 6681 26007 6715
rect 26341 6681 26375 6715
rect 6285 6613 6319 6647
rect 7389 6613 7423 6647
rect 8769 6613 8803 6647
rect 10149 6613 10183 6647
rect 13645 6613 13679 6647
rect 14749 6613 14783 6647
rect 17141 6613 17175 6647
rect 17601 6613 17635 6647
rect 19441 6613 19475 6647
rect 23673 6613 23707 6647
rect 24777 6613 24811 6647
rect 25513 6613 25547 6647
rect 26801 6613 26835 6647
rect 27721 6613 27755 6647
rect 30665 6613 30699 6647
rect 4905 6409 4939 6443
rect 5365 6409 5399 6443
rect 8217 6409 8251 6443
rect 10885 6409 10919 6443
rect 13461 6409 13495 6443
rect 16865 6409 16899 6443
rect 17417 6409 17451 6443
rect 19165 6409 19199 6443
rect 19441 6409 19475 6443
rect 21741 6409 21775 6443
rect 25053 6409 25087 6443
rect 25605 6409 25639 6443
rect 26157 6409 26191 6443
rect 27629 6409 27663 6443
rect 28365 6409 28399 6443
rect 28733 6409 28767 6443
rect 30389 6409 30423 6443
rect 30665 6409 30699 6443
rect 6561 6341 6595 6375
rect 13093 6341 13127 6375
rect 19625 6341 19659 6375
rect 25973 6341 26007 6375
rect 29101 6341 29135 6375
rect 6837 6273 6871 6307
rect 9781 6273 9815 6307
rect 10333 6273 10367 6307
rect 10517 6273 10551 6307
rect 14381 6273 14415 6307
rect 18521 6273 18555 6307
rect 18705 6273 18739 6307
rect 20085 6273 20119 6307
rect 20269 6273 20303 6307
rect 26617 6273 26651 6307
rect 26801 6273 26835 6307
rect 29745 6273 29779 6307
rect 29929 6273 29963 6307
rect 7104 6205 7138 6239
rect 10241 6205 10275 6239
rect 12449 6205 12483 6239
rect 13921 6205 13955 6239
rect 14657 6205 14691 6239
rect 18429 6205 18463 6239
rect 19993 6205 20027 6239
rect 21189 6205 21223 6239
rect 22385 6205 22419 6239
rect 22477 6205 22511 6239
rect 23673 6205 23707 6239
rect 26525 6205 26559 6239
rect 27721 6205 27755 6239
rect 29653 6205 29687 6239
rect 8861 6137 8895 6171
rect 9413 6137 9447 6171
rect 21005 6137 21039 6171
rect 23121 6137 23155 6171
rect 23940 6137 23974 6171
rect 9873 6069 9907 6103
rect 12173 6069 12207 6103
rect 12633 6069 12667 6103
rect 13829 6069 13863 6103
rect 14383 6069 14417 6103
rect 15761 6069 15795 6103
rect 16957 6069 16991 6103
rect 17877 6069 17911 6103
rect 18061 6069 18095 6103
rect 21373 6069 21407 6103
rect 22661 6069 22695 6103
rect 23397 6069 23431 6103
rect 27261 6069 27295 6103
rect 27905 6069 27939 6103
rect 29285 6069 29319 6103
rect 31125 6069 31159 6103
rect 33333 6069 33367 6103
rect 4353 5865 4387 5899
rect 6009 5865 6043 5899
rect 6929 5865 6963 5899
rect 7757 5865 7791 5899
rect 9965 5865 9999 5899
rect 10425 5865 10459 5899
rect 11805 5865 11839 5899
rect 13645 5865 13679 5899
rect 14657 5865 14691 5899
rect 15761 5865 15795 5899
rect 17877 5865 17911 5899
rect 19993 5865 20027 5899
rect 20269 5865 20303 5899
rect 21373 5865 21407 5899
rect 21833 5865 21867 5899
rect 22109 5865 22143 5899
rect 24409 5865 24443 5899
rect 26249 5865 26283 5899
rect 27261 5865 27295 5899
rect 27813 5865 27847 5899
rect 28365 5865 28399 5899
rect 28825 5865 28859 5899
rect 6101 5797 6135 5831
rect 13553 5797 13587 5831
rect 18236 5797 18270 5831
rect 23274 5797 23308 5831
rect 29460 5797 29494 5831
rect 8217 5729 8251 5763
rect 10517 5729 10551 5763
rect 11621 5729 11655 5763
rect 14013 5729 14047 5763
rect 15669 5729 15703 5763
rect 17969 5729 18003 5763
rect 21925 5729 21959 5763
rect 26893 5729 26927 5763
rect 27721 5729 27755 5763
rect 34345 5729 34379 5763
rect 6193 5661 6227 5695
rect 7205 5661 7239 5695
rect 8033 5661 8067 5695
rect 14105 5661 14139 5695
rect 14289 5661 14323 5695
rect 15853 5661 15887 5695
rect 16957 5661 16991 5695
rect 20913 5661 20947 5695
rect 23029 5661 23063 5695
rect 27905 5661 27939 5695
rect 29193 5661 29227 5695
rect 32689 5661 32723 5695
rect 34437 5661 34471 5695
rect 34529 5661 34563 5695
rect 9505 5593 9539 5627
rect 12817 5593 12851 5627
rect 16313 5593 16347 5627
rect 16865 5593 16899 5627
rect 27353 5593 27387 5627
rect 31953 5593 31987 5627
rect 5641 5525 5675 5559
rect 8401 5525 8435 5559
rect 10701 5525 10735 5559
rect 11069 5525 11103 5559
rect 13185 5525 13219 5559
rect 15025 5525 15059 5559
rect 15301 5525 15335 5559
rect 17509 5525 17543 5559
rect 19349 5525 19383 5559
rect 22477 5525 22511 5559
rect 22937 5525 22971 5559
rect 24961 5525 24995 5559
rect 30573 5525 30607 5559
rect 31217 5525 31251 5559
rect 32321 5525 32355 5559
rect 33149 5525 33183 5559
rect 33977 5525 34011 5559
rect 4169 5321 4203 5355
rect 6193 5321 6227 5355
rect 7849 5321 7883 5355
rect 8861 5321 8895 5355
rect 10609 5321 10643 5355
rect 12633 5321 12667 5355
rect 13461 5321 13495 5355
rect 15301 5321 15335 5355
rect 16221 5321 16255 5355
rect 18061 5321 18095 5355
rect 19073 5321 19107 5355
rect 19441 5321 19475 5355
rect 19809 5321 19843 5355
rect 20637 5321 20671 5355
rect 20913 5321 20947 5355
rect 23029 5321 23063 5355
rect 23397 5321 23431 5355
rect 25605 5321 25639 5355
rect 25973 5321 26007 5355
rect 29101 5321 29135 5355
rect 30389 5321 30423 5355
rect 32505 5321 32539 5355
rect 33977 5321 34011 5355
rect 34345 5321 34379 5355
rect 4261 5185 4295 5219
rect 9321 5185 9355 5219
rect 9873 5185 9907 5219
rect 10057 5185 10091 5219
rect 18705 5185 18739 5219
rect 22477 5185 22511 5219
rect 22569 5185 22603 5219
rect 23673 5185 23707 5219
rect 28273 5185 28307 5219
rect 29929 5185 29963 5219
rect 31401 5185 31435 5219
rect 32137 5185 32171 5219
rect 33149 5185 33183 5219
rect 6837 5117 6871 5151
rect 7941 5117 7975 5151
rect 8493 5117 8527 5151
rect 10977 5117 11011 5151
rect 12449 5117 12483 5151
rect 13921 5117 13955 5151
rect 14177 5117 14211 5151
rect 16405 5117 16439 5151
rect 16957 5117 16991 5151
rect 19625 5117 19659 5151
rect 20269 5117 20303 5151
rect 20729 5117 20763 5151
rect 21281 5117 21315 5151
rect 22385 5117 22419 5151
rect 26157 5117 26191 5151
rect 26709 5117 26743 5151
rect 27169 5117 27203 5151
rect 32965 5117 32999 5151
rect 4528 5049 4562 5083
rect 7481 5049 7515 5083
rect 9781 5049 9815 5083
rect 13737 5049 13771 5083
rect 17877 5049 17911 5083
rect 21925 5049 21959 5083
rect 23940 5049 23974 5083
rect 28089 5049 28123 5083
rect 28733 5049 28767 5083
rect 29653 5049 29687 5083
rect 31309 5049 31343 5083
rect 33057 5049 33091 5083
rect 33701 5049 33735 5083
rect 5641 4981 5675 5015
rect 6561 4981 6595 5015
rect 7021 4981 7055 5015
rect 8125 4981 8159 5015
rect 9413 4981 9447 5015
rect 11161 4981 11195 5015
rect 11713 4981 11747 5015
rect 12265 4981 12299 5015
rect 13093 4981 13127 5015
rect 15853 4981 15887 5015
rect 16589 4981 16623 5015
rect 17509 4981 17543 5015
rect 18429 4981 18463 5015
rect 18521 4981 18555 5015
rect 22017 4981 22051 5015
rect 25053 4981 25087 5015
rect 26341 4981 26375 5015
rect 27445 4981 27479 5015
rect 27629 4981 27663 5015
rect 27997 4981 28031 5015
rect 29285 4981 29319 5015
rect 29745 4981 29779 5015
rect 30665 4981 30699 5015
rect 30849 4981 30883 5015
rect 31217 4981 31251 5015
rect 32597 4981 32631 5015
rect 34897 4981 34931 5015
rect 4537 4777 4571 4811
rect 4997 4777 5031 4811
rect 6561 4777 6595 4811
rect 8401 4777 8435 4811
rect 9413 4777 9447 4811
rect 10149 4777 10183 4811
rect 13829 4777 13863 4811
rect 13921 4777 13955 4811
rect 15761 4777 15795 4811
rect 18153 4777 18187 4811
rect 19625 4777 19659 4811
rect 22293 4777 22327 4811
rect 23949 4777 23983 4811
rect 24317 4777 24351 4811
rect 24777 4777 24811 4811
rect 25237 4777 25271 4811
rect 25881 4777 25915 4811
rect 26249 4777 26283 4811
rect 28457 4777 28491 4811
rect 29193 4777 29227 4811
rect 29653 4777 29687 4811
rect 29929 4777 29963 4811
rect 31401 4777 31435 4811
rect 31769 4777 31803 4811
rect 33057 4777 33091 4811
rect 33517 4777 33551 4811
rect 34529 4777 34563 4811
rect 35173 4777 35207 4811
rect 6469 4709 6503 4743
rect 8769 4709 8803 4743
rect 10517 4709 10551 4743
rect 10793 4709 10827 4743
rect 16773 4709 16807 4743
rect 23121 4709 23155 4743
rect 26792 4709 26826 4743
rect 30757 4709 30791 4743
rect 4905 4641 4939 4675
rect 5733 4641 5767 4675
rect 7757 4641 7791 4675
rect 9781 4641 9815 4675
rect 9965 4641 9999 4675
rect 10977 4641 11011 4675
rect 11244 4641 11278 4675
rect 15669 4641 15703 4675
rect 18061 4641 18095 4675
rect 20637 4641 20671 4675
rect 20913 4641 20947 4675
rect 21180 4641 21214 4675
rect 23397 4641 23431 4675
rect 29009 4641 29043 4675
rect 30665 4641 30699 4675
rect 32137 4641 32171 4675
rect 35081 4641 35115 4675
rect 4353 4573 4387 4607
rect 5089 4573 5123 4607
rect 6745 4573 6779 4607
rect 13369 4573 13403 4607
rect 14013 4573 14047 4607
rect 15853 4573 15887 4607
rect 17601 4573 17635 4607
rect 18337 4573 18371 4607
rect 18705 4573 18739 4607
rect 19717 4573 19751 4607
rect 19809 4573 19843 4607
rect 25329 4573 25363 4607
rect 25421 4573 25455 4607
rect 26525 4573 26559 4607
rect 30849 4573 30883 4607
rect 33609 4573 33643 4607
rect 33793 4573 33827 4607
rect 35357 4573 35391 4607
rect 15025 4505 15059 4539
rect 16313 4505 16347 4539
rect 17233 4505 17267 4539
rect 17693 4505 17727 4539
rect 19165 4505 19199 4539
rect 27905 4505 27939 4539
rect 32689 4505 32723 4539
rect 33149 4505 33183 4539
rect 34713 4505 34747 4539
rect 6101 4437 6135 4471
rect 7205 4437 7239 4471
rect 7481 4437 7515 4471
rect 7941 4437 7975 4471
rect 12357 4437 12391 4471
rect 12909 4437 12943 4471
rect 13461 4437 13495 4471
rect 14473 4437 14507 4471
rect 15301 4437 15335 4471
rect 19257 4437 19291 4471
rect 20361 4437 20395 4471
rect 23581 4437 23615 4471
rect 24869 4437 24903 4471
rect 30297 4437 30331 4471
rect 34253 4437 34287 4471
rect 35725 4437 35759 4471
rect 4077 4233 4111 4267
rect 6193 4233 6227 4267
rect 6561 4233 6595 4267
rect 6837 4233 6871 4267
rect 11069 4233 11103 4267
rect 11345 4233 11379 4267
rect 14105 4233 14139 4267
rect 16221 4233 16255 4267
rect 19993 4233 20027 4267
rect 22109 4233 22143 4267
rect 27537 4233 27571 4267
rect 28273 4233 28307 4267
rect 28641 4233 28675 4267
rect 29469 4233 29503 4267
rect 30389 4233 30423 4267
rect 34713 4233 34747 4267
rect 3065 4097 3099 4131
rect 3801 4097 3835 4131
rect 7389 4097 7423 4131
rect 7941 4097 7975 4131
rect 9045 4097 9079 4131
rect 10425 4097 10459 4131
rect 10609 4097 10643 4131
rect 13001 4097 13035 4131
rect 13553 4097 13587 4131
rect 14289 4097 14323 4131
rect 17785 4097 17819 4131
rect 21649 4097 21683 4131
rect 22845 4097 22879 4131
rect 24225 4097 24259 4131
rect 24685 4097 24719 4131
rect 25145 4097 25179 4131
rect 27905 4097 27939 4131
rect 29009 4097 29043 4131
rect 30021 4097 30055 4131
rect 31401 4097 31435 4131
rect 3157 4029 3191 4063
rect 4261 4029 4295 4063
rect 4528 4029 4562 4063
rect 7205 4029 7239 4063
rect 8769 4029 8803 4063
rect 10333 4029 10367 4063
rect 12173 4029 12207 4063
rect 12817 4029 12851 4063
rect 14556 4029 14590 4063
rect 16773 4029 16807 4063
rect 17325 4029 17359 4063
rect 18613 4029 18647 4063
rect 18880 4029 18914 4063
rect 21005 4029 21039 4063
rect 21465 4029 21499 4063
rect 22477 4029 22511 4063
rect 24041 4029 24075 4063
rect 24133 4029 24167 4063
rect 25421 4029 25455 4063
rect 25605 4029 25639 4063
rect 25872 4029 25906 4063
rect 28089 4029 28123 4063
rect 29285 4029 29319 4063
rect 31125 4029 31159 4063
rect 32321 4029 32355 4063
rect 32577 4029 32611 4063
rect 35357 4029 35391 4063
rect 35449 4029 35483 4063
rect 35716 4029 35750 4063
rect 8309 3961 8343 3995
rect 8861 3961 8895 3995
rect 9505 3961 9539 3995
rect 20637 3961 20671 3995
rect 23489 3961 23523 3995
rect 3341 3893 3375 3927
rect 5641 3893 5675 3927
rect 7297 3893 7331 3927
rect 8401 3893 8435 3927
rect 9781 3893 9815 3927
rect 9965 3893 9999 3927
rect 11897 3893 11931 3927
rect 12449 3893 12483 3927
rect 12909 3893 12943 3927
rect 15669 3893 15703 3927
rect 16681 3893 16715 3927
rect 16957 3893 16991 3927
rect 18429 3893 18463 3927
rect 21097 3893 21131 3927
rect 21557 3893 21591 3927
rect 23673 3893 23707 3927
rect 26985 3893 27019 3927
rect 30757 3893 30791 3927
rect 31217 3893 31251 3927
rect 31861 3893 31895 3927
rect 32137 3893 32171 3927
rect 33701 3893 33735 3927
rect 34345 3893 34379 3927
rect 36829 3893 36863 3927
rect 4813 3689 4847 3723
rect 5181 3689 5215 3723
rect 7849 3689 7883 3723
rect 9229 3689 9263 3723
rect 10517 3689 10551 3723
rect 10885 3689 10919 3723
rect 14933 3689 14967 3723
rect 15853 3689 15887 3723
rect 16221 3689 16255 3723
rect 16865 3689 16899 3723
rect 17879 3689 17913 3723
rect 19901 3689 19935 3723
rect 23305 3689 23339 3723
rect 23673 3689 23707 3723
rect 23949 3689 23983 3723
rect 24869 3689 24903 3723
rect 25329 3689 25363 3723
rect 25973 3689 26007 3723
rect 26893 3689 26927 3723
rect 26985 3689 27019 3723
rect 29837 3689 29871 3723
rect 30389 3689 30423 3723
rect 31493 3689 31527 3723
rect 35449 3689 35483 3723
rect 5610 3621 5644 3655
rect 10425 3621 10459 3655
rect 12602 3621 12636 3655
rect 14565 3621 14599 3655
rect 27629 3621 27663 3655
rect 35357 3621 35391 3655
rect 35909 3621 35943 3655
rect 4261 3553 4295 3587
rect 5365 3553 5399 3587
rect 7757 3553 7791 3587
rect 8217 3553 8251 3587
rect 10977 3553 11011 3587
rect 16313 3553 16347 3587
rect 17233 3553 17267 3587
rect 21261 3553 21295 3587
rect 23765 3553 23799 3587
rect 25237 3553 25271 3587
rect 26341 3553 26375 3587
rect 28713 3553 28747 3587
rect 30941 3553 30975 3587
rect 33241 3553 33275 3587
rect 35817 3553 35851 3587
rect 8309 3485 8343 3519
rect 8401 3485 8435 3519
rect 8861 3485 8895 3519
rect 11161 3485 11195 3519
rect 11529 3485 11563 3519
rect 11897 3485 11931 3519
rect 12357 3485 12391 3519
rect 16405 3485 16439 3519
rect 17417 3485 17451 3519
rect 17877 3485 17911 3519
rect 18153 3485 18187 3519
rect 19257 3485 19291 3519
rect 21005 3485 21039 3519
rect 25513 3485 25547 3519
rect 27169 3485 27203 3519
rect 27905 3485 27939 3519
rect 28457 3485 28491 3519
rect 32505 3485 32539 3519
rect 32828 3485 32862 3519
rect 32965 3485 32999 3519
rect 36001 3485 36035 3519
rect 36829 3485 36863 3519
rect 4445 3417 4479 3451
rect 20177 3417 20211 3451
rect 20729 3417 20763 3451
rect 30849 3417 30883 3451
rect 31953 3417 31987 3451
rect 34989 3417 35023 3451
rect 3801 3349 3835 3383
rect 6745 3349 6779 3383
rect 7297 3349 7331 3383
rect 9965 3349 9999 3383
rect 13737 3349 13771 3383
rect 15577 3349 15611 3383
rect 22385 3349 22419 3383
rect 24409 3349 24443 3383
rect 24777 3349 24811 3383
rect 26525 3349 26559 3383
rect 28273 3349 28307 3383
rect 31125 3349 31159 3383
rect 32321 3349 32355 3383
rect 34345 3349 34379 3383
rect 36553 3349 36587 3383
rect 2053 3145 2087 3179
rect 3801 3145 3835 3179
rect 6193 3145 6227 3179
rect 6561 3145 6595 3179
rect 8217 3145 8251 3179
rect 8769 3145 8803 3179
rect 9413 3145 9447 3179
rect 11253 3145 11287 3179
rect 11897 3145 11931 3179
rect 16405 3145 16439 3179
rect 17049 3145 17083 3179
rect 17509 3145 17543 3179
rect 19993 3145 20027 3179
rect 23305 3145 23339 3179
rect 24225 3145 24259 3179
rect 25605 3145 25639 3179
rect 27169 3145 27203 3179
rect 27721 3145 27755 3179
rect 28549 3145 28583 3179
rect 29101 3145 29135 3179
rect 30757 3145 30791 3179
rect 31309 3145 31343 3179
rect 34621 3145 34655 3179
rect 35265 3145 35299 3179
rect 36829 3145 36863 3179
rect 37381 3145 37415 3179
rect 3341 3077 3375 3111
rect 4169 3077 4203 3111
rect 33701 3077 33735 3111
rect 4261 3009 4295 3043
rect 6837 3009 6871 3043
rect 12633 3009 12667 3043
rect 13461 3009 13495 3043
rect 13645 3009 13679 3043
rect 14105 3009 14139 3043
rect 15025 3009 15059 3043
rect 21005 3009 21039 3043
rect 24685 3009 24719 3043
rect 24777 3009 24811 3043
rect 25789 3009 25823 3043
rect 29377 3009 29411 3043
rect 31861 3009 31895 3043
rect 32321 3009 32355 3043
rect 32597 3009 32631 3043
rect 35449 3009 35483 3043
rect 1409 2941 1443 2975
rect 3157 2941 3191 2975
rect 4528 2941 4562 2975
rect 9781 2941 9815 2975
rect 9873 2941 9907 2975
rect 12265 2941 12299 2975
rect 13369 2941 13403 2975
rect 14565 2941 14599 2975
rect 15301 2941 15335 2975
rect 17877 2941 17911 2975
rect 18061 2941 18095 2975
rect 20545 2941 20579 2975
rect 21281 2941 21315 2975
rect 25237 2941 25271 2975
rect 29644 2941 29678 2975
rect 35716 2941 35750 2975
rect 7082 2873 7116 2907
rect 10140 2873 10174 2907
rect 18306 2873 18340 2907
rect 23949 2873 23983 2907
rect 24593 2873 24627 2907
rect 26034 2873 26068 2907
rect 1593 2805 1627 2839
rect 5641 2805 5675 2839
rect 13001 2805 13035 2839
rect 14473 2805 14507 2839
rect 15027 2805 15061 2839
rect 19441 2805 19475 2839
rect 20453 2805 20487 2839
rect 21007 2805 21041 2839
rect 22385 2805 22419 2839
rect 23029 2805 23063 2839
rect 28181 2805 28215 2839
rect 31769 2805 31803 2839
rect 32323 2805 32357 2839
rect 34253 2805 34287 2839
rect 2421 2601 2455 2635
rect 3157 2601 3191 2635
rect 5089 2601 5123 2635
rect 5273 2601 5307 2635
rect 6653 2601 6687 2635
rect 8585 2601 8619 2635
rect 9137 2601 9171 2635
rect 11161 2601 11195 2635
rect 12357 2601 12391 2635
rect 14289 2601 14323 2635
rect 14841 2601 14875 2635
rect 16865 2601 16899 2635
rect 17417 2601 17451 2635
rect 19993 2601 20027 2635
rect 22661 2601 22695 2635
rect 23857 2601 23891 2635
rect 24501 2601 24535 2635
rect 25053 2601 25087 2635
rect 25973 2601 26007 2635
rect 26617 2601 26651 2635
rect 28273 2601 28307 2635
rect 29469 2601 29503 2635
rect 31953 2601 31987 2635
rect 32321 2601 32355 2635
rect 34253 2601 34287 2635
rect 36829 2601 36863 2635
rect 3893 2533 3927 2567
rect 5733 2533 5767 2567
rect 6285 2533 6319 2567
rect 7472 2533 7506 2567
rect 10048 2533 10082 2567
rect 11713 2533 11747 2567
rect 13176 2533 13210 2567
rect 15730 2533 15764 2567
rect 18880 2533 18914 2567
rect 21548 2533 21582 2567
rect 24409 2533 24443 2567
rect 25605 2533 25639 2567
rect 27160 2533 27194 2567
rect 30082 2533 30116 2567
rect 33140 2533 33174 2567
rect 34805 2533 34839 2567
rect 35716 2533 35750 2567
rect 37381 2533 37415 2567
rect 1409 2465 1443 2499
rect 2053 2465 2087 2499
rect 2513 2465 2547 2499
rect 4169 2465 4203 2499
rect 5641 2465 5675 2499
rect 7205 2465 7239 2499
rect 9505 2465 9539 2499
rect 9781 2465 9815 2499
rect 12909 2465 12943 2499
rect 15209 2465 15243 2499
rect 15485 2465 15519 2499
rect 18153 2465 18187 2499
rect 18613 2465 18647 2499
rect 20637 2465 20671 2499
rect 21005 2465 21039 2499
rect 21281 2465 21315 2499
rect 25789 2465 25823 2499
rect 26893 2465 26927 2499
rect 29837 2465 29871 2499
rect 32873 2465 32907 2499
rect 35173 2465 35207 2499
rect 35449 2465 35483 2499
rect 3525 2397 3559 2431
rect 5825 2397 5859 2431
rect 23489 2397 23523 2431
rect 24593 2397 24627 2431
rect 25513 2397 25547 2431
rect 4353 2329 4387 2363
rect 29193 2329 29227 2363
rect 1593 2261 1627 2295
rect 2697 2261 2731 2295
rect 4813 2261 4847 2295
rect 24041 2261 24075 2295
rect 26249 2261 26283 2295
rect 31217 2261 31251 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 38824 37562
rect 1104 37488 38824 37510
rect 1104 37018 38824 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 38824 37018
rect 1104 36944 38824 36966
rect 1104 36474 38824 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 38824 36474
rect 1104 36400 38824 36422
rect 35618 36360 35624 36372
rect 35579 36332 35624 36360
rect 35618 36320 35624 36332
rect 35676 36320 35682 36372
rect 35437 36227 35495 36233
rect 35437 36193 35449 36227
rect 35483 36224 35495 36227
rect 35802 36224 35808 36236
rect 35483 36196 35808 36224
rect 35483 36193 35495 36196
rect 35437 36187 35495 36193
rect 35802 36184 35808 36196
rect 35860 36184 35866 36236
rect 1104 35930 38824 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 38824 35930
rect 1104 35856 38824 35878
rect 35621 35819 35679 35825
rect 35621 35785 35633 35819
rect 35667 35816 35679 35819
rect 35710 35816 35716 35828
rect 35667 35788 35716 35816
rect 35667 35785 35679 35788
rect 35621 35779 35679 35785
rect 35710 35776 35716 35788
rect 35768 35776 35774 35828
rect 35437 35615 35495 35621
rect 35437 35612 35449 35615
rect 35268 35584 35449 35612
rect 33042 35476 33048 35488
rect 33003 35448 33048 35476
rect 33042 35436 33048 35448
rect 33100 35436 33106 35488
rect 33410 35476 33416 35488
rect 33371 35448 33416 35476
rect 33410 35436 33416 35448
rect 33468 35436 33474 35488
rect 34790 35436 34796 35488
rect 34848 35476 34854 35488
rect 35268 35485 35296 35584
rect 35437 35581 35449 35584
rect 35483 35581 35495 35615
rect 35437 35575 35495 35581
rect 35253 35479 35311 35485
rect 35253 35476 35265 35479
rect 34848 35448 35265 35476
rect 34848 35436 34854 35448
rect 35253 35445 35265 35448
rect 35299 35445 35311 35479
rect 35253 35439 35311 35445
rect 35894 35436 35900 35488
rect 35952 35476 35958 35488
rect 35989 35479 36047 35485
rect 35989 35476 36001 35479
rect 35952 35448 36001 35476
rect 35952 35436 35958 35448
rect 35989 35445 36001 35448
rect 36035 35445 36047 35479
rect 35989 35439 36047 35445
rect 1104 35386 38824 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 38824 35386
rect 1104 35312 38824 35334
rect 33410 35232 33416 35284
rect 33468 35272 33474 35284
rect 33505 35275 33563 35281
rect 33505 35272 33517 35275
rect 33468 35244 33517 35272
rect 33468 35232 33474 35244
rect 33505 35241 33517 35244
rect 33551 35241 33563 35275
rect 33505 35235 33563 35241
rect 32392 35207 32450 35213
rect 32392 35173 32404 35207
rect 32438 35204 32450 35207
rect 33042 35204 33048 35216
rect 32438 35176 33048 35204
rect 32438 35173 32450 35176
rect 32392 35167 32450 35173
rect 33042 35164 33048 35176
rect 33100 35164 33106 35216
rect 34514 35096 34520 35148
rect 34572 35136 34578 35148
rect 34865 35139 34923 35145
rect 34865 35136 34877 35139
rect 34572 35108 34877 35136
rect 34572 35096 34578 35108
rect 34865 35105 34877 35108
rect 34911 35105 34923 35139
rect 34865 35099 34923 35105
rect 32122 35068 32128 35080
rect 32083 35040 32128 35068
rect 32122 35028 32128 35040
rect 32180 35028 32186 35080
rect 34606 35068 34612 35080
rect 34567 35040 34612 35068
rect 34606 35028 34612 35040
rect 34664 35028 34670 35080
rect 34514 34932 34520 34944
rect 34475 34904 34520 34932
rect 34514 34892 34520 34904
rect 34572 34892 34578 34944
rect 35894 34892 35900 34944
rect 35952 34932 35958 34944
rect 35989 34935 36047 34941
rect 35989 34932 36001 34935
rect 35952 34904 36001 34932
rect 35952 34892 35958 34904
rect 35989 34901 36001 34904
rect 36035 34901 36047 34935
rect 35989 34895 36047 34901
rect 1104 34842 38824 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 38824 34842
rect 1104 34768 38824 34790
rect 34514 34688 34520 34740
rect 34572 34728 34578 34740
rect 36265 34731 36323 34737
rect 36265 34728 36277 34731
rect 34572 34700 36277 34728
rect 34572 34688 34578 34700
rect 36265 34697 36277 34700
rect 36311 34697 36323 34731
rect 37550 34728 37556 34740
rect 37511 34700 37556 34728
rect 36265 34691 36323 34697
rect 37550 34688 37556 34700
rect 37608 34688 37614 34740
rect 34241 34663 34299 34669
rect 34241 34660 34253 34663
rect 32416 34632 34253 34660
rect 30469 34527 30527 34533
rect 30469 34524 30481 34527
rect 30300 34496 30481 34524
rect 30006 34348 30012 34400
rect 30064 34388 30070 34400
rect 30300 34397 30328 34496
rect 30469 34493 30481 34496
rect 30515 34524 30527 34527
rect 32122 34524 32128 34536
rect 30515 34496 32128 34524
rect 30515 34493 30527 34496
rect 30469 34487 30527 34493
rect 32122 34484 32128 34496
rect 32180 34524 32186 34536
rect 32416 34533 32444 34632
rect 34241 34629 34253 34632
rect 34287 34660 34299 34663
rect 34606 34660 34612 34672
rect 34287 34632 34612 34660
rect 34287 34629 34299 34632
rect 34241 34623 34299 34629
rect 34606 34620 34612 34632
rect 34664 34660 34670 34672
rect 34664 34632 34928 34660
rect 34664 34620 34670 34632
rect 33226 34552 33232 34604
rect 33284 34592 33290 34604
rect 34900 34601 34928 34632
rect 33505 34595 33563 34601
rect 33505 34592 33517 34595
rect 33284 34564 33517 34592
rect 33284 34552 33290 34564
rect 33505 34561 33517 34564
rect 33551 34561 33563 34595
rect 33505 34555 33563 34561
rect 34885 34595 34943 34601
rect 34885 34561 34897 34595
rect 34931 34561 34943 34595
rect 34885 34555 34943 34561
rect 32401 34527 32459 34533
rect 32401 34524 32413 34527
rect 32180 34496 32413 34524
rect 32180 34484 32186 34496
rect 32401 34493 32413 34496
rect 32447 34493 32459 34527
rect 32401 34487 32459 34493
rect 32861 34527 32919 34533
rect 32861 34493 32873 34527
rect 32907 34524 32919 34527
rect 33042 34524 33048 34536
rect 32907 34496 33048 34524
rect 32907 34493 32919 34496
rect 32861 34487 32919 34493
rect 33042 34484 33048 34496
rect 33100 34524 33106 34536
rect 37369 34527 37427 34533
rect 33100 34496 33456 34524
rect 33100 34484 33106 34496
rect 30558 34416 30564 34468
rect 30616 34456 30622 34468
rect 30714 34459 30772 34465
rect 30714 34456 30726 34459
rect 30616 34428 30726 34456
rect 30616 34416 30622 34428
rect 30714 34425 30726 34428
rect 30760 34425 30772 34459
rect 33318 34456 33324 34468
rect 33279 34428 33324 34456
rect 30714 34419 30772 34425
rect 33318 34416 33324 34428
rect 33376 34416 33382 34468
rect 30285 34391 30343 34397
rect 30285 34388 30297 34391
rect 30064 34360 30297 34388
rect 30064 34348 30070 34360
rect 30285 34357 30297 34360
rect 30331 34357 30343 34391
rect 31846 34388 31852 34400
rect 31807 34360 31852 34388
rect 30285 34351 30343 34357
rect 31846 34348 31852 34360
rect 31904 34348 31910 34400
rect 32950 34388 32956 34400
rect 32911 34360 32956 34388
rect 32950 34348 32956 34360
rect 33008 34348 33014 34400
rect 33428 34397 33456 34496
rect 37369 34493 37381 34527
rect 37415 34524 37427 34527
rect 37826 34524 37832 34536
rect 37415 34496 37832 34524
rect 37415 34493 37427 34496
rect 37369 34487 37427 34493
rect 37826 34484 37832 34496
rect 37884 34524 37890 34536
rect 37921 34527 37979 34533
rect 37921 34524 37933 34527
rect 37884 34496 37933 34524
rect 37884 34484 37890 34496
rect 37921 34493 37933 34496
rect 37967 34493 37979 34527
rect 37921 34487 37979 34493
rect 34422 34416 34428 34468
rect 34480 34456 34486 34468
rect 35130 34459 35188 34465
rect 35130 34456 35142 34459
rect 34480 34428 35142 34456
rect 34480 34416 34486 34428
rect 35130 34425 35142 34428
rect 35176 34425 35188 34459
rect 35130 34419 35188 34425
rect 33413 34391 33471 34397
rect 33413 34357 33425 34391
rect 33459 34388 33471 34391
rect 33502 34388 33508 34400
rect 33459 34360 33508 34388
rect 33459 34357 33471 34360
rect 33413 34351 33471 34357
rect 33502 34348 33508 34360
rect 33560 34348 33566 34400
rect 1104 34298 38824 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 38824 34298
rect 1104 34224 38824 34246
rect 30558 34184 30564 34196
rect 30519 34156 30564 34184
rect 30558 34144 30564 34156
rect 30616 34144 30622 34196
rect 33502 34184 33508 34196
rect 33463 34156 33508 34184
rect 33502 34144 33508 34156
rect 33560 34144 33566 34196
rect 31846 34076 31852 34128
rect 31904 34116 31910 34128
rect 32370 34119 32428 34125
rect 32370 34116 32382 34119
rect 31904 34088 32382 34116
rect 31904 34076 31910 34088
rect 32370 34085 32382 34088
rect 32416 34116 32428 34119
rect 32858 34116 32864 34128
rect 32416 34088 32864 34116
rect 32416 34085 32428 34088
rect 32370 34079 32428 34085
rect 32858 34076 32864 34088
rect 32916 34076 32922 34128
rect 33318 34076 33324 34128
rect 33376 34116 33382 34128
rect 34422 34116 34428 34128
rect 33376 34088 34428 34116
rect 33376 34076 33382 34088
rect 34422 34076 34428 34088
rect 34480 34076 34486 34128
rect 34514 34076 34520 34128
rect 34572 34116 34578 34128
rect 34876 34119 34934 34125
rect 34876 34116 34888 34119
rect 34572 34088 34888 34116
rect 34572 34076 34578 34088
rect 34876 34085 34888 34088
rect 34922 34116 34934 34119
rect 35802 34116 35808 34128
rect 34922 34088 35808 34116
rect 34922 34085 34934 34088
rect 34876 34079 34934 34085
rect 35802 34076 35808 34088
rect 35860 34076 35866 34128
rect 32122 33980 32128 33992
rect 32083 33952 32128 33980
rect 32122 33940 32128 33952
rect 32180 33940 32186 33992
rect 34606 33980 34612 33992
rect 34567 33952 34612 33980
rect 34606 33940 34612 33952
rect 34664 33940 34670 33992
rect 30098 33844 30104 33856
rect 30059 33816 30104 33844
rect 30098 33804 30104 33816
rect 30156 33804 30162 33856
rect 33226 33804 33232 33856
rect 33284 33844 33290 33856
rect 34057 33847 34115 33853
rect 34057 33844 34069 33847
rect 33284 33816 34069 33844
rect 33284 33804 33290 33816
rect 34057 33813 34069 33816
rect 34103 33813 34115 33847
rect 35986 33844 35992 33856
rect 35947 33816 35992 33844
rect 34057 33807 34115 33813
rect 35986 33804 35992 33816
rect 36044 33804 36050 33856
rect 1104 33754 38824 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 38824 33754
rect 1104 33680 38824 33702
rect 30650 33600 30656 33652
rect 30708 33640 30714 33652
rect 31389 33643 31447 33649
rect 31389 33640 31401 33643
rect 30708 33612 31401 33640
rect 30708 33600 30714 33612
rect 31389 33609 31401 33612
rect 31435 33640 31447 33643
rect 32490 33640 32496 33652
rect 31435 33612 32496 33640
rect 31435 33609 31447 33612
rect 31389 33603 31447 33609
rect 32490 33600 32496 33612
rect 32548 33600 32554 33652
rect 33870 33600 33876 33652
rect 33928 33640 33934 33652
rect 34333 33643 34391 33649
rect 34333 33640 34345 33643
rect 33928 33612 34345 33640
rect 33928 33600 33934 33612
rect 34333 33609 34345 33612
rect 34379 33640 34391 33643
rect 34514 33640 34520 33652
rect 34379 33612 34520 33640
rect 34379 33609 34391 33612
rect 34333 33603 34391 33609
rect 34514 33600 34520 33612
rect 34572 33600 34578 33652
rect 32122 33572 32128 33584
rect 32083 33544 32128 33572
rect 32122 33532 32128 33544
rect 32180 33532 32186 33584
rect 32490 33464 32496 33516
rect 32548 33504 32554 33516
rect 32953 33507 33011 33513
rect 32953 33504 32965 33507
rect 32548 33476 32965 33504
rect 32548 33464 32554 33476
rect 32953 33473 32965 33476
rect 32999 33473 33011 33507
rect 32953 33467 33011 33473
rect 33137 33507 33195 33513
rect 33137 33473 33149 33507
rect 33183 33504 33195 33507
rect 33226 33504 33232 33516
rect 33183 33476 33232 33504
rect 33183 33473 33195 33476
rect 33137 33467 33195 33473
rect 33226 33464 33232 33476
rect 33284 33464 33290 33516
rect 30006 33436 30012 33448
rect 29840 33408 30012 33436
rect 29454 33260 29460 33312
rect 29512 33300 29518 33312
rect 29840 33309 29868 33408
rect 30006 33396 30012 33408
rect 30064 33396 30070 33448
rect 30098 33396 30104 33448
rect 30156 33436 30162 33448
rect 30282 33445 30288 33448
rect 30265 33439 30288 33445
rect 30265 33436 30277 33439
rect 30156 33408 30277 33436
rect 30156 33396 30162 33408
rect 30265 33405 30277 33408
rect 30340 33436 30346 33448
rect 32858 33436 32864 33448
rect 30340 33408 30413 33436
rect 32819 33408 32864 33436
rect 30265 33399 30288 33405
rect 30282 33396 30288 33399
rect 30340 33396 30346 33408
rect 32858 33396 32864 33408
rect 32916 33436 32922 33448
rect 33505 33439 33563 33445
rect 33505 33436 33517 33439
rect 32916 33408 33517 33436
rect 32916 33396 32922 33408
rect 33505 33405 33517 33408
rect 33551 33405 33563 33439
rect 35253 33439 35311 33445
rect 35253 33436 35265 33439
rect 33505 33399 33563 33405
rect 35084 33408 35265 33436
rect 29825 33303 29883 33309
rect 29825 33300 29837 33303
rect 29512 33272 29837 33300
rect 29512 33260 29518 33272
rect 29825 33269 29837 33272
rect 29871 33269 29883 33303
rect 29825 33263 29883 33269
rect 32306 33260 32312 33312
rect 32364 33300 32370 33312
rect 32493 33303 32551 33309
rect 32493 33300 32505 33303
rect 32364 33272 32505 33300
rect 32364 33260 32370 33272
rect 32493 33269 32505 33272
rect 32539 33269 32551 33303
rect 34606 33300 34612 33312
rect 34567 33272 34612 33300
rect 32493 33263 32551 33269
rect 34606 33260 34612 33272
rect 34664 33300 34670 33312
rect 35084 33309 35112 33408
rect 35253 33405 35265 33408
rect 35299 33405 35311 33439
rect 35253 33399 35311 33405
rect 35342 33396 35348 33448
rect 35400 33436 35406 33448
rect 35509 33439 35567 33445
rect 35509 33436 35521 33439
rect 35400 33408 35521 33436
rect 35400 33396 35406 33408
rect 35509 33405 35521 33408
rect 35555 33436 35567 33439
rect 35986 33436 35992 33448
rect 35555 33408 35992 33436
rect 35555 33405 35567 33408
rect 35509 33399 35567 33405
rect 35986 33396 35992 33408
rect 36044 33396 36050 33448
rect 35069 33303 35127 33309
rect 35069 33300 35081 33303
rect 34664 33272 35081 33300
rect 34664 33260 34670 33272
rect 35069 33269 35081 33272
rect 35115 33269 35127 33303
rect 36630 33300 36636 33312
rect 36591 33272 36636 33300
rect 35069 33263 35127 33269
rect 36630 33260 36636 33272
rect 36688 33260 36694 33312
rect 1104 33210 38824 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 38824 33210
rect 1104 33136 38824 33158
rect 30374 33056 30380 33108
rect 30432 33096 30438 33108
rect 30742 33096 30748 33108
rect 30432 33068 30748 33096
rect 30432 33056 30438 33068
rect 30742 33056 30748 33068
rect 30800 33096 30806 33108
rect 30837 33099 30895 33105
rect 30837 33096 30849 33099
rect 30800 33068 30849 33096
rect 30800 33056 30806 33068
rect 30837 33065 30849 33068
rect 30883 33065 30895 33099
rect 32490 33096 32496 33108
rect 32451 33068 32496 33096
rect 30837 33059 30895 33065
rect 32490 33056 32496 33068
rect 32548 33056 32554 33108
rect 32858 33096 32864 33108
rect 32819 33068 32864 33096
rect 32858 33056 32864 33068
rect 32916 33056 32922 33108
rect 33870 33096 33876 33108
rect 33831 33068 33876 33096
rect 33870 33056 33876 33068
rect 33928 33056 33934 33108
rect 35069 33099 35127 33105
rect 35069 33065 35081 33099
rect 35115 33096 35127 33099
rect 35342 33096 35348 33108
rect 35115 33068 35348 33096
rect 35115 33065 35127 33068
rect 35069 33059 35127 33065
rect 35342 33056 35348 33068
rect 35400 33056 35406 33108
rect 29730 32969 29736 32972
rect 29724 32923 29736 32969
rect 29788 32960 29794 32972
rect 34330 32960 34336 32972
rect 29788 32932 29824 32960
rect 33980 32932 34336 32960
rect 29730 32920 29736 32923
rect 29788 32920 29794 32932
rect 29454 32892 29460 32904
rect 29415 32864 29460 32892
rect 29454 32852 29460 32864
rect 29512 32852 29518 32904
rect 33594 32852 33600 32904
rect 33652 32892 33658 32904
rect 33980 32901 34008 32932
rect 34330 32920 34336 32932
rect 34388 32920 34394 32972
rect 35434 32969 35440 32972
rect 35428 32960 35440 32969
rect 35395 32932 35440 32960
rect 35428 32923 35440 32932
rect 35492 32960 35498 32972
rect 36630 32960 36636 32972
rect 35492 32932 36636 32960
rect 35434 32920 35440 32923
rect 35492 32920 35498 32932
rect 36630 32920 36636 32932
rect 36688 32920 36694 32972
rect 33965 32895 34023 32901
rect 33965 32892 33977 32895
rect 33652 32864 33977 32892
rect 33652 32852 33658 32864
rect 33965 32861 33977 32864
rect 34011 32861 34023 32895
rect 33965 32855 34023 32861
rect 34057 32895 34115 32901
rect 34057 32861 34069 32895
rect 34103 32861 34115 32895
rect 34057 32855 34115 32861
rect 34072 32824 34100 32855
rect 34606 32852 34612 32904
rect 34664 32892 34670 32904
rect 35161 32895 35219 32901
rect 35161 32892 35173 32895
rect 34664 32864 35173 32892
rect 34664 32852 34670 32864
rect 35161 32861 35173 32864
rect 35207 32861 35219 32895
rect 35161 32855 35219 32861
rect 33244 32796 34100 32824
rect 33244 32768 33272 32796
rect 30926 32716 30932 32768
rect 30984 32756 30990 32768
rect 33226 32756 33232 32768
rect 30984 32728 33232 32756
rect 30984 32716 30990 32728
rect 33226 32716 33232 32728
rect 33284 32716 33290 32768
rect 33502 32756 33508 32768
rect 33463 32728 33508 32756
rect 33502 32716 33508 32728
rect 33560 32716 33566 32768
rect 35802 32716 35808 32768
rect 35860 32756 35866 32768
rect 36541 32759 36599 32765
rect 36541 32756 36553 32759
rect 35860 32728 36553 32756
rect 35860 32716 35866 32728
rect 36541 32725 36553 32728
rect 36587 32725 36599 32759
rect 36541 32719 36599 32725
rect 1104 32666 38824 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 38824 32666
rect 1104 32592 38824 32614
rect 29730 32512 29736 32564
rect 29788 32552 29794 32564
rect 29825 32555 29883 32561
rect 29825 32552 29837 32555
rect 29788 32524 29837 32552
rect 29788 32512 29794 32524
rect 29825 32521 29837 32524
rect 29871 32552 29883 32555
rect 30193 32555 30251 32561
rect 30193 32552 30205 32555
rect 29871 32524 30205 32552
rect 29871 32521 29883 32524
rect 29825 32515 29883 32521
rect 30193 32521 30205 32524
rect 30239 32521 30251 32555
rect 30193 32515 30251 32521
rect 33229 32555 33287 32561
rect 33229 32521 33241 32555
rect 33275 32552 33287 32555
rect 33870 32552 33876 32564
rect 33275 32524 33876 32552
rect 33275 32521 33287 32524
rect 33229 32515 33287 32521
rect 30208 32280 30236 32515
rect 33870 32512 33876 32524
rect 33928 32512 33934 32564
rect 34606 32552 34612 32564
rect 34567 32524 34612 32552
rect 34606 32512 34612 32524
rect 34664 32512 34670 32564
rect 36541 32555 36599 32561
rect 36541 32521 36553 32555
rect 36587 32552 36599 32555
rect 36630 32552 36636 32564
rect 36587 32524 36636 32552
rect 36587 32521 36599 32524
rect 36541 32515 36599 32521
rect 36630 32512 36636 32524
rect 36688 32512 36694 32564
rect 36814 32552 36820 32564
rect 36775 32524 36820 32552
rect 36814 32512 36820 32524
rect 36872 32512 36878 32564
rect 30377 32487 30435 32493
rect 30377 32453 30389 32487
rect 30423 32484 30435 32487
rect 31757 32487 31815 32493
rect 31757 32484 31769 32487
rect 30423 32456 31769 32484
rect 30423 32453 30435 32456
rect 30377 32447 30435 32453
rect 31757 32453 31769 32456
rect 31803 32484 31815 32487
rect 33594 32484 33600 32496
rect 31803 32456 32444 32484
rect 33555 32456 33600 32484
rect 31803 32453 31815 32456
rect 31757 32447 31815 32453
rect 30926 32416 30932 32428
rect 30887 32388 30932 32416
rect 30926 32376 30932 32388
rect 30984 32376 30990 32428
rect 32416 32425 32444 32456
rect 33594 32444 33600 32456
rect 33652 32444 33658 32496
rect 35986 32484 35992 32496
rect 35544 32456 35992 32484
rect 32401 32419 32459 32425
rect 32401 32385 32413 32419
rect 32447 32385 32459 32419
rect 32582 32416 32588 32428
rect 32543 32388 32588 32416
rect 32401 32379 32459 32385
rect 32582 32376 32588 32388
rect 32640 32376 32646 32428
rect 35544 32425 35572 32456
rect 35986 32444 35992 32456
rect 36044 32484 36050 32496
rect 36081 32487 36139 32493
rect 36081 32484 36093 32487
rect 36044 32456 36093 32484
rect 36044 32444 36050 32456
rect 36081 32453 36093 32456
rect 36127 32453 36139 32487
rect 36081 32447 36139 32453
rect 35529 32419 35587 32425
rect 35529 32385 35541 32419
rect 35575 32385 35587 32419
rect 35529 32379 35587 32385
rect 35618 32376 35624 32428
rect 35676 32416 35682 32428
rect 35676 32388 35721 32416
rect 35676 32376 35682 32388
rect 30742 32348 30748 32360
rect 30703 32320 30748 32348
rect 30742 32308 30748 32320
rect 30800 32308 30806 32360
rect 31481 32351 31539 32357
rect 31481 32317 31493 32351
rect 31527 32348 31539 32351
rect 32306 32348 32312 32360
rect 31527 32320 32312 32348
rect 31527 32317 31539 32320
rect 31481 32311 31539 32317
rect 32306 32308 32312 32320
rect 32364 32308 32370 32360
rect 33689 32351 33747 32357
rect 33689 32317 33701 32351
rect 33735 32348 33747 32351
rect 36633 32351 36691 32357
rect 33735 32320 34376 32348
rect 33735 32317 33747 32320
rect 33689 32311 33747 32317
rect 30837 32283 30895 32289
rect 30837 32280 30849 32283
rect 30208 32252 30849 32280
rect 30837 32249 30849 32252
rect 30883 32249 30895 32283
rect 30837 32243 30895 32249
rect 34348 32224 34376 32320
rect 36633 32317 36645 32351
rect 36679 32348 36691 32351
rect 36679 32320 37136 32348
rect 36679 32317 36691 32320
rect 36633 32311 36691 32317
rect 37108 32224 37136 32320
rect 28442 32172 28448 32224
rect 28500 32212 28506 32224
rect 29454 32212 29460 32224
rect 28500 32184 29460 32212
rect 28500 32172 28506 32184
rect 29454 32172 29460 32184
rect 29512 32172 29518 32224
rect 31938 32212 31944 32224
rect 31899 32184 31944 32212
rect 31938 32172 31944 32184
rect 31996 32172 32002 32224
rect 33873 32215 33931 32221
rect 33873 32181 33885 32215
rect 33919 32212 33931 32215
rect 33962 32212 33968 32224
rect 33919 32184 33968 32212
rect 33919 32181 33931 32184
rect 33873 32175 33931 32181
rect 33962 32172 33968 32184
rect 34020 32172 34026 32224
rect 34330 32212 34336 32224
rect 34291 32184 34336 32212
rect 34330 32172 34336 32184
rect 34388 32172 34394 32224
rect 34698 32172 34704 32224
rect 34756 32212 34762 32224
rect 35069 32215 35127 32221
rect 35069 32212 35081 32215
rect 34756 32184 35081 32212
rect 34756 32172 34762 32184
rect 35069 32181 35081 32184
rect 35115 32181 35127 32215
rect 35434 32212 35440 32224
rect 35395 32184 35440 32212
rect 35069 32175 35127 32181
rect 35434 32172 35440 32184
rect 35492 32172 35498 32224
rect 37090 32172 37096 32224
rect 37148 32212 37154 32224
rect 37185 32215 37243 32221
rect 37185 32212 37197 32215
rect 37148 32184 37197 32212
rect 37148 32172 37154 32184
rect 37185 32181 37197 32184
rect 37231 32181 37243 32215
rect 37185 32175 37243 32181
rect 1104 32122 38824 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 38824 32122
rect 1104 32048 38824 32070
rect 29641 32011 29699 32017
rect 29641 31977 29653 32011
rect 29687 32008 29699 32011
rect 29730 32008 29736 32020
rect 29687 31980 29736 32008
rect 29687 31977 29699 31980
rect 29641 31971 29699 31977
rect 29730 31968 29736 31980
rect 29788 31968 29794 32020
rect 30469 32011 30527 32017
rect 30469 31977 30481 32011
rect 30515 32008 30527 32011
rect 30742 32008 30748 32020
rect 30515 31980 30748 32008
rect 30515 31977 30527 31980
rect 30469 31971 30527 31977
rect 30742 31968 30748 31980
rect 30800 31968 30806 32020
rect 30837 32011 30895 32017
rect 30837 31977 30849 32011
rect 30883 32008 30895 32011
rect 30926 32008 30932 32020
rect 30883 31980 30932 32008
rect 30883 31977 30895 31980
rect 30837 31971 30895 31977
rect 30926 31968 30932 31980
rect 30984 31968 30990 32020
rect 31113 32011 31171 32017
rect 31113 31977 31125 32011
rect 31159 32008 31171 32011
rect 31662 32008 31668 32020
rect 31159 31980 31668 32008
rect 31159 31977 31171 31980
rect 31113 31971 31171 31977
rect 31662 31968 31668 31980
rect 31720 31968 31726 32020
rect 32677 32011 32735 32017
rect 32677 31977 32689 32011
rect 32723 31977 32735 32011
rect 32677 31971 32735 31977
rect 28534 31881 28540 31884
rect 28528 31872 28540 31881
rect 28495 31844 28540 31872
rect 28528 31835 28540 31844
rect 28534 31832 28540 31835
rect 28592 31832 28598 31884
rect 30929 31875 30987 31881
rect 30929 31841 30941 31875
rect 30975 31872 30987 31875
rect 31018 31872 31024 31884
rect 30975 31844 31024 31872
rect 30975 31841 30987 31844
rect 30929 31835 30987 31841
rect 31018 31832 31024 31844
rect 31076 31872 31082 31884
rect 32692 31872 32720 31971
rect 32950 31968 32956 32020
rect 33008 32008 33014 32020
rect 33137 32011 33195 32017
rect 33137 32008 33149 32011
rect 33008 31980 33149 32008
rect 33008 31968 33014 31980
rect 33137 31977 33149 31980
rect 33183 31977 33195 32011
rect 33137 31971 33195 31977
rect 33226 31968 33232 32020
rect 33284 32008 33290 32020
rect 33689 32011 33747 32017
rect 33689 32008 33701 32011
rect 33284 31980 33701 32008
rect 33284 31968 33290 31980
rect 33689 31977 33701 31980
rect 33735 32008 33747 32011
rect 34606 32008 34612 32020
rect 33735 31980 34612 32008
rect 33735 31977 33747 31980
rect 33689 31971 33747 31977
rect 34606 31968 34612 31980
rect 34664 31968 34670 32020
rect 35069 32011 35127 32017
rect 35069 31977 35081 32011
rect 35115 32008 35127 32011
rect 35434 32008 35440 32020
rect 35115 31980 35440 32008
rect 35115 31977 35127 31980
rect 35069 31971 35127 31977
rect 35434 31968 35440 31980
rect 35492 31968 35498 32020
rect 35894 31968 35900 32020
rect 35952 32008 35958 32020
rect 36541 32011 36599 32017
rect 36541 32008 36553 32011
rect 35952 31980 36553 32008
rect 35952 31968 35958 31980
rect 36541 31977 36553 31980
rect 36587 31977 36599 32011
rect 36541 31971 36599 31977
rect 32766 31900 32772 31952
rect 32824 31940 32830 31952
rect 33045 31943 33103 31949
rect 33045 31940 33057 31943
rect 32824 31912 33057 31940
rect 32824 31900 32830 31912
rect 33045 31909 33057 31912
rect 33091 31940 33103 31943
rect 33502 31940 33508 31952
rect 33091 31912 33508 31940
rect 33091 31909 33103 31912
rect 33045 31903 33103 31909
rect 33502 31900 33508 31912
rect 33560 31900 33566 31952
rect 31076 31844 32720 31872
rect 31076 31832 31082 31844
rect 34514 31832 34520 31884
rect 34572 31872 34578 31884
rect 35161 31875 35219 31881
rect 35161 31872 35173 31875
rect 34572 31844 35173 31872
rect 34572 31832 34578 31844
rect 35161 31841 35173 31844
rect 35207 31841 35219 31875
rect 35161 31835 35219 31841
rect 35428 31875 35486 31881
rect 35428 31841 35440 31875
rect 35474 31872 35486 31875
rect 35802 31872 35808 31884
rect 35474 31844 35808 31872
rect 35474 31841 35486 31844
rect 35428 31835 35486 31841
rect 35802 31832 35808 31844
rect 35860 31832 35866 31884
rect 28261 31807 28319 31813
rect 28261 31773 28273 31807
rect 28307 31773 28319 31807
rect 32582 31804 32588 31816
rect 32495 31776 32588 31804
rect 28261 31767 28319 31773
rect 28276 31668 28304 31767
rect 28442 31668 28448 31680
rect 28276 31640 28448 31668
rect 28442 31628 28448 31640
rect 28500 31628 28506 31680
rect 31846 31668 31852 31680
rect 31807 31640 31852 31668
rect 31846 31628 31852 31640
rect 31904 31668 31910 31680
rect 32508 31677 32536 31776
rect 32582 31764 32588 31776
rect 32640 31804 32646 31816
rect 33229 31807 33287 31813
rect 33229 31804 33241 31807
rect 32640 31776 33241 31804
rect 32640 31764 32646 31776
rect 33229 31773 33241 31776
rect 33275 31773 33287 31807
rect 33229 31767 33287 31773
rect 32493 31671 32551 31677
rect 32493 31668 32505 31671
rect 31904 31640 32505 31668
rect 31904 31628 31910 31640
rect 32493 31637 32505 31640
rect 32539 31637 32551 31671
rect 34054 31668 34060 31680
rect 34015 31640 34060 31668
rect 32493 31631 32551 31637
rect 34054 31628 34060 31640
rect 34112 31628 34118 31680
rect 1104 31578 38824 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 38824 31578
rect 1104 31504 38824 31526
rect 31018 31464 31024 31476
rect 30979 31436 31024 31464
rect 31018 31424 31024 31436
rect 31076 31424 31082 31476
rect 31941 31467 31999 31473
rect 31941 31433 31953 31467
rect 31987 31464 31999 31467
rect 32766 31464 32772 31476
rect 31987 31436 32772 31464
rect 31987 31433 31999 31436
rect 31941 31427 31999 31433
rect 32766 31424 32772 31436
rect 32824 31424 32830 31476
rect 32217 31399 32275 31405
rect 32217 31365 32229 31399
rect 32263 31396 32275 31399
rect 32953 31399 33011 31405
rect 32953 31396 32965 31399
rect 32263 31368 32965 31396
rect 32263 31365 32275 31368
rect 32217 31359 32275 31365
rect 32953 31365 32965 31368
rect 32999 31396 33011 31399
rect 32999 31368 33640 31396
rect 32999 31365 33011 31368
rect 32953 31359 33011 31365
rect 31754 31288 31760 31340
rect 31812 31328 31818 31340
rect 33612 31337 33640 31368
rect 35342 31356 35348 31408
rect 35400 31396 35406 31408
rect 35618 31396 35624 31408
rect 35400 31368 35624 31396
rect 35400 31356 35406 31368
rect 35618 31356 35624 31368
rect 35676 31356 35682 31408
rect 32585 31331 32643 31337
rect 32585 31328 32597 31331
rect 31812 31300 32597 31328
rect 31812 31288 31818 31300
rect 32585 31297 32597 31300
rect 32631 31328 32643 31331
rect 33597 31331 33655 31337
rect 32631 31300 33548 31328
rect 32631 31297 32643 31300
rect 32585 31291 32643 31297
rect 31573 31263 31631 31269
rect 31573 31229 31585 31263
rect 31619 31260 31631 31263
rect 31938 31260 31944 31272
rect 31619 31232 31944 31260
rect 31619 31229 31631 31232
rect 31573 31223 31631 31229
rect 31938 31220 31944 31232
rect 31996 31260 32002 31272
rect 33520 31269 33548 31300
rect 33597 31297 33609 31331
rect 33643 31297 33655 31331
rect 33597 31291 33655 31297
rect 33781 31331 33839 31337
rect 33781 31297 33793 31331
rect 33827 31328 33839 31331
rect 34054 31328 34060 31340
rect 33827 31300 34060 31328
rect 33827 31297 33839 31300
rect 33781 31291 33839 31297
rect 34054 31288 34060 31300
rect 34112 31328 34118 31340
rect 34422 31328 34428 31340
rect 34112 31300 34428 31328
rect 34112 31288 34118 31300
rect 34422 31288 34428 31300
rect 34480 31288 34486 31340
rect 34606 31288 34612 31340
rect 34664 31328 34670 31340
rect 35710 31328 35716 31340
rect 34664 31300 35716 31328
rect 34664 31288 34670 31300
rect 35710 31288 35716 31300
rect 35768 31328 35774 31340
rect 36078 31328 36084 31340
rect 35768 31300 36084 31328
rect 35768 31288 35774 31300
rect 36078 31288 36084 31300
rect 36136 31288 36142 31340
rect 32033 31263 32091 31269
rect 32033 31260 32045 31263
rect 31996 31232 32045 31260
rect 31996 31220 32002 31232
rect 32033 31229 32045 31232
rect 32079 31229 32091 31263
rect 32033 31223 32091 31229
rect 33505 31263 33563 31269
rect 33505 31229 33517 31263
rect 33551 31229 33563 31263
rect 33505 31223 33563 31229
rect 34333 31263 34391 31269
rect 34333 31229 34345 31263
rect 34379 31260 34391 31263
rect 34701 31263 34759 31269
rect 34701 31260 34713 31263
rect 34379 31232 34713 31260
rect 34379 31229 34391 31232
rect 34333 31223 34391 31229
rect 34701 31229 34713 31232
rect 34747 31260 34759 31263
rect 35529 31263 35587 31269
rect 35529 31260 35541 31263
rect 34747 31232 35541 31260
rect 34747 31229 34759 31232
rect 34701 31223 34759 31229
rect 35529 31229 35541 31232
rect 35575 31260 35587 31263
rect 35802 31260 35808 31272
rect 35575 31232 35808 31260
rect 35575 31229 35587 31232
rect 35529 31223 35587 31229
rect 35802 31220 35808 31232
rect 35860 31220 35866 31272
rect 24854 31124 24860 31136
rect 24815 31096 24860 31124
rect 24854 31084 24860 31096
rect 24912 31084 24918 31136
rect 27522 31124 27528 31136
rect 27483 31096 27528 31124
rect 27522 31084 27528 31096
rect 27580 31084 27586 31136
rect 28353 31127 28411 31133
rect 28353 31093 28365 31127
rect 28399 31124 28411 31127
rect 28442 31124 28448 31136
rect 28399 31096 28448 31124
rect 28399 31093 28411 31096
rect 28353 31087 28411 31093
rect 28442 31084 28448 31096
rect 28500 31084 28506 31136
rect 28534 31084 28540 31136
rect 28592 31124 28598 31136
rect 28629 31127 28687 31133
rect 28629 31124 28641 31127
rect 28592 31096 28641 31124
rect 28592 31084 28598 31096
rect 28629 31093 28641 31096
rect 28675 31093 28687 31127
rect 28629 31087 28687 31093
rect 33137 31127 33195 31133
rect 33137 31093 33149 31127
rect 33183 31124 33195 31127
rect 33318 31124 33324 31136
rect 33183 31096 33324 31124
rect 33183 31093 33195 31096
rect 33137 31087 33195 31093
rect 33318 31084 33324 31096
rect 33376 31084 33382 31136
rect 35069 31127 35127 31133
rect 35069 31093 35081 31127
rect 35115 31124 35127 31127
rect 35250 31124 35256 31136
rect 35115 31096 35256 31124
rect 35115 31093 35127 31096
rect 35069 31087 35127 31093
rect 35250 31084 35256 31096
rect 35308 31084 35314 31136
rect 35434 31124 35440 31136
rect 35395 31096 35440 31124
rect 35434 31084 35440 31096
rect 35492 31124 35498 31136
rect 35894 31124 35900 31136
rect 35492 31096 35900 31124
rect 35492 31084 35498 31096
rect 35894 31084 35900 31096
rect 35952 31084 35958 31136
rect 36078 31124 36084 31136
rect 36039 31096 36084 31124
rect 36078 31084 36084 31096
rect 36136 31084 36142 31136
rect 1104 31034 38824 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 38824 31034
rect 1104 30960 38824 30982
rect 24765 30923 24823 30929
rect 24765 30889 24777 30923
rect 24811 30920 24823 30923
rect 24854 30920 24860 30932
rect 24811 30892 24860 30920
rect 24811 30889 24823 30892
rect 24765 30883 24823 30889
rect 24854 30880 24860 30892
rect 24912 30920 24918 30932
rect 25222 30920 25228 30932
rect 24912 30892 25228 30920
rect 24912 30880 24918 30892
rect 25222 30880 25228 30892
rect 25280 30880 25286 30932
rect 32769 30923 32827 30929
rect 32769 30889 32781 30923
rect 32815 30920 32827 30923
rect 32950 30920 32956 30932
rect 32815 30892 32956 30920
rect 32815 30889 32827 30892
rect 32769 30883 32827 30889
rect 32950 30880 32956 30892
rect 33008 30880 33014 30932
rect 33137 30923 33195 30929
rect 33137 30889 33149 30923
rect 33183 30920 33195 30923
rect 33226 30920 33232 30932
rect 33183 30892 33232 30920
rect 33183 30889 33195 30892
rect 33137 30883 33195 30889
rect 33226 30880 33232 30892
rect 33284 30880 33290 30932
rect 35897 30923 35955 30929
rect 35897 30889 35909 30923
rect 35943 30920 35955 30923
rect 35986 30920 35992 30932
rect 35943 30892 35992 30920
rect 35943 30889 35955 30892
rect 35897 30883 35955 30889
rect 35986 30880 35992 30892
rect 36044 30880 36050 30932
rect 27148 30787 27206 30793
rect 27148 30753 27160 30787
rect 27194 30784 27206 30787
rect 27614 30784 27620 30796
rect 27194 30756 27620 30784
rect 27194 30753 27206 30756
rect 27148 30747 27206 30753
rect 27614 30744 27620 30756
rect 27672 30744 27678 30796
rect 32122 30784 32128 30796
rect 32083 30756 32128 30784
rect 32122 30744 32128 30756
rect 32180 30744 32186 30796
rect 33134 30744 33140 30796
rect 33192 30784 33198 30796
rect 33485 30787 33543 30793
rect 33485 30784 33497 30787
rect 33192 30756 33497 30784
rect 33192 30744 33198 30756
rect 33485 30753 33497 30756
rect 33531 30784 33543 30787
rect 35434 30784 35440 30796
rect 33531 30756 35440 30784
rect 33531 30753 33543 30756
rect 33485 30747 33543 30753
rect 35434 30744 35440 30756
rect 35492 30784 35498 30796
rect 35529 30787 35587 30793
rect 35529 30784 35541 30787
rect 35492 30756 35541 30784
rect 35492 30744 35498 30756
rect 35529 30753 35541 30756
rect 35575 30753 35587 30787
rect 35529 30747 35587 30753
rect 35713 30787 35771 30793
rect 35713 30753 35725 30787
rect 35759 30784 35771 30787
rect 35802 30784 35808 30796
rect 35759 30756 35808 30784
rect 35759 30753 35771 30756
rect 35713 30747 35771 30753
rect 35802 30744 35808 30756
rect 35860 30744 35866 30796
rect 24854 30676 24860 30728
rect 24912 30716 24918 30728
rect 25317 30719 25375 30725
rect 25317 30716 25329 30719
rect 24912 30688 25329 30716
rect 24912 30676 24918 30688
rect 25317 30685 25329 30688
rect 25363 30685 25375 30719
rect 25317 30679 25375 30685
rect 25409 30719 25467 30725
rect 25409 30685 25421 30719
rect 25455 30685 25467 30719
rect 26878 30716 26884 30728
rect 26839 30688 26884 30716
rect 25409 30679 25467 30685
rect 24397 30651 24455 30657
rect 24397 30617 24409 30651
rect 24443 30648 24455 30651
rect 24946 30648 24952 30660
rect 24443 30620 24952 30648
rect 24443 30617 24455 30620
rect 24397 30611 24455 30617
rect 24946 30608 24952 30620
rect 25004 30648 25010 30660
rect 25424 30648 25452 30679
rect 26878 30676 26884 30688
rect 26936 30676 26942 30728
rect 33229 30719 33287 30725
rect 33229 30685 33241 30719
rect 33275 30685 33287 30719
rect 33229 30679 33287 30685
rect 25004 30620 25452 30648
rect 25004 30608 25010 30620
rect 24857 30583 24915 30589
rect 24857 30549 24869 30583
rect 24903 30580 24915 30583
rect 26234 30580 26240 30592
rect 24903 30552 26240 30580
rect 24903 30549 24915 30552
rect 24857 30543 24915 30549
rect 26234 30540 26240 30552
rect 26292 30540 26298 30592
rect 28261 30583 28319 30589
rect 28261 30549 28273 30583
rect 28307 30580 28319 30583
rect 29270 30580 29276 30592
rect 28307 30552 29276 30580
rect 28307 30549 28319 30552
rect 28261 30543 28319 30549
rect 29270 30540 29276 30552
rect 29328 30540 29334 30592
rect 29638 30580 29644 30592
rect 29599 30552 29644 30580
rect 29638 30540 29644 30552
rect 29696 30540 29702 30592
rect 32306 30580 32312 30592
rect 32267 30552 32312 30580
rect 32306 30540 32312 30552
rect 32364 30540 32370 30592
rect 33134 30540 33140 30592
rect 33192 30580 33198 30592
rect 33244 30580 33272 30679
rect 35161 30651 35219 30657
rect 35161 30648 35173 30651
rect 34256 30620 35173 30648
rect 34146 30580 34152 30592
rect 33192 30552 34152 30580
rect 33192 30540 33198 30552
rect 34146 30540 34152 30552
rect 34204 30580 34210 30592
rect 34256 30580 34284 30620
rect 35161 30617 35173 30620
rect 35207 30617 35219 30651
rect 35161 30611 35219 30617
rect 34606 30580 34612 30592
rect 34204 30552 34284 30580
rect 34567 30552 34612 30580
rect 34204 30540 34210 30552
rect 34606 30540 34612 30552
rect 34664 30540 34670 30592
rect 35986 30540 35992 30592
rect 36044 30580 36050 30592
rect 36357 30583 36415 30589
rect 36357 30580 36369 30583
rect 36044 30552 36369 30580
rect 36044 30540 36050 30552
rect 36357 30549 36369 30552
rect 36403 30580 36415 30583
rect 37182 30580 37188 30592
rect 36403 30552 37188 30580
rect 36403 30549 36415 30552
rect 36357 30543 36415 30549
rect 37182 30540 37188 30552
rect 37240 30540 37246 30592
rect 1104 30490 38824 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 38824 30490
rect 1104 30416 38824 30438
rect 27890 30336 27896 30388
rect 27948 30376 27954 30388
rect 28534 30376 28540 30388
rect 27948 30348 28540 30376
rect 27948 30336 27954 30348
rect 28534 30336 28540 30348
rect 28592 30336 28598 30388
rect 33045 30379 33103 30385
rect 33045 30345 33057 30379
rect 33091 30376 33103 30379
rect 33134 30376 33140 30388
rect 33091 30348 33140 30376
rect 33091 30345 33103 30348
rect 33045 30339 33103 30345
rect 33134 30336 33140 30348
rect 33192 30336 33198 30388
rect 34606 30376 34612 30388
rect 34440 30348 34612 30376
rect 24029 30311 24087 30317
rect 24029 30277 24041 30311
rect 24075 30308 24087 30311
rect 24210 30308 24216 30320
rect 24075 30280 24216 30308
rect 24075 30277 24087 30280
rect 24029 30271 24087 30277
rect 24210 30268 24216 30280
rect 24268 30308 24274 30320
rect 24489 30311 24547 30317
rect 24489 30308 24501 30311
rect 24268 30280 24501 30308
rect 24268 30268 24274 30280
rect 24489 30277 24501 30280
rect 24535 30308 24547 30311
rect 24854 30308 24860 30320
rect 24535 30280 24860 30308
rect 24535 30277 24547 30280
rect 24489 30271 24547 30277
rect 24854 30268 24860 30280
rect 24912 30268 24918 30320
rect 26878 30268 26884 30320
rect 26936 30308 26942 30320
rect 26973 30311 27031 30317
rect 26973 30308 26985 30311
rect 26936 30280 26985 30308
rect 26936 30268 26942 30280
rect 26973 30277 26985 30280
rect 27019 30308 27031 30311
rect 28442 30308 28448 30320
rect 27019 30280 28448 30308
rect 27019 30277 27031 30280
rect 26973 30271 27031 30277
rect 28442 30268 28448 30280
rect 28500 30268 28506 30320
rect 32309 30311 32367 30317
rect 32309 30277 32321 30311
rect 32355 30308 32367 30311
rect 33965 30311 34023 30317
rect 33965 30308 33977 30311
rect 32355 30280 33977 30308
rect 32355 30277 32367 30280
rect 32309 30271 32367 30277
rect 33965 30277 33977 30280
rect 34011 30308 34023 30311
rect 34440 30308 34468 30348
rect 34606 30336 34612 30348
rect 34664 30336 34670 30388
rect 35986 30376 35992 30388
rect 35912 30348 35992 30376
rect 34698 30308 34704 30320
rect 34011 30280 34468 30308
rect 34659 30280 34704 30308
rect 34011 30277 34023 30280
rect 33965 30271 34023 30277
rect 34698 30268 34704 30280
rect 34756 30308 34762 30320
rect 35158 30308 35164 30320
rect 34756 30280 35164 30308
rect 34756 30268 34762 30280
rect 35158 30268 35164 30280
rect 35216 30268 35222 30320
rect 35912 30308 35940 30348
rect 35986 30336 35992 30348
rect 36044 30336 36050 30388
rect 35544 30280 35940 30308
rect 36633 30311 36691 30317
rect 27522 30200 27528 30252
rect 27580 30240 27586 30252
rect 28077 30243 28135 30249
rect 28077 30240 28089 30243
rect 27580 30212 28089 30240
rect 27580 30200 27586 30212
rect 28077 30209 28089 30212
rect 28123 30240 28135 30243
rect 28123 30212 28948 30240
rect 28123 30209 28135 30212
rect 28077 30203 28135 30209
rect 25222 30181 25228 30184
rect 24949 30175 25007 30181
rect 24949 30172 24961 30175
rect 24780 30144 24961 30172
rect 23934 29996 23940 30048
rect 23992 30036 23998 30048
rect 24780 30045 24808 30144
rect 24949 30141 24961 30144
rect 24995 30141 25007 30175
rect 25216 30172 25228 30181
rect 25183 30144 25228 30172
rect 24949 30135 25007 30141
rect 25216 30135 25228 30144
rect 25222 30132 25228 30135
rect 25280 30132 25286 30184
rect 27614 30132 27620 30184
rect 27672 30172 27678 30184
rect 27801 30175 27859 30181
rect 27801 30172 27813 30175
rect 27672 30144 27813 30172
rect 27672 30132 27678 30144
rect 27801 30141 27813 30144
rect 27847 30172 27859 30175
rect 28445 30175 28503 30181
rect 28445 30172 28457 30175
rect 27847 30144 28457 30172
rect 27847 30141 27859 30144
rect 27801 30135 27859 30141
rect 28445 30141 28457 30144
rect 28491 30172 28503 30175
rect 28813 30175 28871 30181
rect 28813 30172 28825 30175
rect 28491 30144 28825 30172
rect 28491 30141 28503 30144
rect 28445 30135 28503 30141
rect 28813 30141 28825 30144
rect 28859 30141 28871 30175
rect 28813 30135 28871 30141
rect 27249 30107 27307 30113
rect 27249 30104 27261 30107
rect 26344 30076 27261 30104
rect 26344 30048 26372 30076
rect 27249 30073 27261 30076
rect 27295 30104 27307 30107
rect 27893 30107 27951 30113
rect 27893 30104 27905 30107
rect 27295 30076 27905 30104
rect 27295 30073 27307 30076
rect 27249 30067 27307 30073
rect 27893 30073 27905 30076
rect 27939 30073 27951 30107
rect 28920 30104 28948 30212
rect 29270 30200 29276 30252
rect 29328 30240 29334 30252
rect 29733 30243 29791 30249
rect 29733 30240 29745 30243
rect 29328 30212 29745 30240
rect 29328 30200 29334 30212
rect 29733 30209 29745 30212
rect 29779 30209 29791 30243
rect 29733 30203 29791 30209
rect 29825 30243 29883 30249
rect 29825 30209 29837 30243
rect 29871 30209 29883 30243
rect 29825 30203 29883 30209
rect 32677 30243 32735 30249
rect 32677 30209 32689 30243
rect 32723 30240 32735 30243
rect 33042 30240 33048 30252
rect 32723 30212 33048 30240
rect 32723 30209 32735 30212
rect 32677 30203 32735 30209
rect 29638 30172 29644 30184
rect 29599 30144 29644 30172
rect 29638 30132 29644 30144
rect 29696 30132 29702 30184
rect 28920 30076 29500 30104
rect 27893 30067 27951 30073
rect 29472 30048 29500 30076
rect 24765 30039 24823 30045
rect 24765 30036 24777 30039
rect 23992 30008 24777 30036
rect 23992 29996 23998 30008
rect 24765 30005 24777 30008
rect 24811 30005 24823 30039
rect 26326 30036 26332 30048
rect 26287 30008 26332 30036
rect 24765 29999 24823 30005
rect 26326 29996 26332 30008
rect 26384 29996 26390 30048
rect 27430 30036 27436 30048
rect 27391 30008 27436 30036
rect 27430 29996 27436 30008
rect 27488 29996 27494 30048
rect 28994 29996 29000 30048
rect 29052 30036 29058 30048
rect 29273 30039 29331 30045
rect 29273 30036 29285 30039
rect 29052 30008 29285 30036
rect 29052 29996 29058 30008
rect 29273 30005 29285 30008
rect 29319 30005 29331 30039
rect 29273 29999 29331 30005
rect 29454 29996 29460 30048
rect 29512 30036 29518 30048
rect 29840 30036 29868 30203
rect 33042 30200 33048 30212
rect 33100 30200 33106 30252
rect 33226 30200 33232 30252
rect 33284 30240 33290 30252
rect 33689 30243 33747 30249
rect 33689 30240 33701 30243
rect 33284 30212 33701 30240
rect 33284 30200 33290 30212
rect 33689 30209 33701 30212
rect 33735 30240 33747 30243
rect 33778 30240 33784 30252
rect 33735 30212 33784 30240
rect 33735 30209 33747 30212
rect 33689 30203 33747 30209
rect 33778 30200 33784 30212
rect 33836 30200 33842 30252
rect 34330 30200 34336 30252
rect 34388 30240 34394 30252
rect 35544 30249 35572 30280
rect 36633 30277 36645 30311
rect 36679 30308 36691 30311
rect 36722 30308 36728 30320
rect 36679 30280 36728 30308
rect 36679 30277 36691 30280
rect 36633 30271 36691 30277
rect 36722 30268 36728 30280
rect 36780 30268 36786 30320
rect 35529 30243 35587 30249
rect 35529 30240 35541 30243
rect 34388 30212 35541 30240
rect 34388 30200 34394 30212
rect 35529 30209 35541 30212
rect 35575 30209 35587 30243
rect 35529 30203 35587 30209
rect 31941 30175 31999 30181
rect 31941 30141 31953 30175
rect 31987 30172 31999 30175
rect 32122 30172 32128 30184
rect 31987 30144 32128 30172
rect 31987 30141 31999 30144
rect 31941 30135 31999 30141
rect 32122 30132 32128 30144
rect 32180 30172 32186 30184
rect 35250 30172 35256 30184
rect 32180 30144 34928 30172
rect 35211 30144 35256 30172
rect 32180 30132 32186 30144
rect 33505 30107 33563 30113
rect 33505 30073 33517 30107
rect 33551 30104 33563 30107
rect 33551 30076 34284 30104
rect 33551 30073 33563 30076
rect 33505 30067 33563 30073
rect 34256 30048 34284 30076
rect 30285 30039 30343 30045
rect 30285 30036 30297 30039
rect 29512 30008 30297 30036
rect 29512 29996 29518 30008
rect 30285 30005 30297 30008
rect 30331 30005 30343 30039
rect 30285 29999 30343 30005
rect 33137 30039 33195 30045
rect 33137 30005 33149 30039
rect 33183 30036 33195 30039
rect 33410 30036 33416 30048
rect 33183 30008 33416 30036
rect 33183 30005 33195 30008
rect 33137 29999 33195 30005
rect 33410 29996 33416 30008
rect 33468 29996 33474 30048
rect 33594 29996 33600 30048
rect 33652 30036 33658 30048
rect 33965 30039 34023 30045
rect 33965 30036 33977 30039
rect 33652 30008 33977 30036
rect 33652 29996 33658 30008
rect 33965 30005 33977 30008
rect 34011 30005 34023 30039
rect 34238 30036 34244 30048
rect 34199 30008 34244 30036
rect 33965 29999 34023 30005
rect 34238 29996 34244 30008
rect 34296 29996 34302 30048
rect 34900 30045 34928 30144
rect 35250 30132 35256 30144
rect 35308 30172 35314 30184
rect 36265 30175 36323 30181
rect 36265 30172 36277 30175
rect 35308 30144 36277 30172
rect 35308 30132 35314 30144
rect 36265 30141 36277 30144
rect 36311 30141 36323 30175
rect 36265 30135 36323 30141
rect 36449 30175 36507 30181
rect 36449 30141 36461 30175
rect 36495 30141 36507 30175
rect 36449 30135 36507 30141
rect 35158 30064 35164 30116
rect 35216 30104 35222 30116
rect 35345 30107 35403 30113
rect 35345 30104 35357 30107
rect 35216 30076 35357 30104
rect 35216 30064 35222 30076
rect 35345 30073 35357 30076
rect 35391 30073 35403 30107
rect 35345 30067 35403 30073
rect 36170 30064 36176 30116
rect 36228 30104 36234 30116
rect 36464 30104 36492 30135
rect 37001 30107 37059 30113
rect 37001 30104 37013 30107
rect 36228 30076 37013 30104
rect 36228 30064 36234 30076
rect 37001 30073 37013 30076
rect 37047 30073 37059 30107
rect 37001 30067 37059 30073
rect 34885 30039 34943 30045
rect 34885 30005 34897 30039
rect 34931 30005 34943 30039
rect 35894 30036 35900 30048
rect 35855 30008 35900 30036
rect 34885 29999 34943 30005
rect 35894 29996 35900 30008
rect 35952 29996 35958 30048
rect 1104 29946 38824 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 38824 29946
rect 1104 29872 38824 29894
rect 25222 29792 25228 29844
rect 25280 29832 25286 29844
rect 25317 29835 25375 29841
rect 25317 29832 25329 29835
rect 25280 29804 25329 29832
rect 25280 29792 25286 29804
rect 25317 29801 25329 29804
rect 25363 29801 25375 29835
rect 25317 29795 25375 29801
rect 27614 29792 27620 29844
rect 27672 29832 27678 29844
rect 27893 29835 27951 29841
rect 27893 29832 27905 29835
rect 27672 29804 27905 29832
rect 27672 29792 27678 29804
rect 27893 29801 27905 29804
rect 27939 29801 27951 29835
rect 27893 29795 27951 29801
rect 28905 29835 28963 29841
rect 28905 29801 28917 29835
rect 28951 29832 28963 29835
rect 29638 29832 29644 29844
rect 28951 29804 29644 29832
rect 28951 29801 28963 29804
rect 28905 29795 28963 29801
rect 29638 29792 29644 29804
rect 29696 29832 29702 29844
rect 30377 29835 30435 29841
rect 30377 29832 30389 29835
rect 29696 29804 30389 29832
rect 29696 29792 29702 29804
rect 30377 29801 30389 29804
rect 30423 29801 30435 29835
rect 30377 29795 30435 29801
rect 34514 29792 34520 29844
rect 34572 29832 34578 29844
rect 35342 29832 35348 29844
rect 34572 29804 35348 29832
rect 34572 29792 34578 29804
rect 35342 29792 35348 29804
rect 35400 29832 35406 29844
rect 35805 29835 35863 29841
rect 35805 29832 35817 29835
rect 35400 29804 35817 29832
rect 35400 29792 35406 29804
rect 35805 29801 35817 29804
rect 35851 29801 35863 29835
rect 35805 29795 35863 29801
rect 24210 29773 24216 29776
rect 24204 29764 24216 29773
rect 24171 29736 24216 29764
rect 24204 29727 24216 29736
rect 24210 29724 24216 29727
rect 24268 29724 24274 29776
rect 26326 29724 26332 29776
rect 26384 29764 26390 29776
rect 26758 29767 26816 29773
rect 26758 29764 26770 29767
rect 26384 29736 26770 29764
rect 26384 29724 26390 29736
rect 26758 29733 26770 29736
rect 26804 29733 26816 29767
rect 26758 29727 26816 29733
rect 26878 29724 26884 29776
rect 26936 29724 26942 29776
rect 29270 29773 29276 29776
rect 29264 29764 29276 29773
rect 29231 29736 29276 29764
rect 29264 29727 29276 29736
rect 29270 29724 29276 29727
rect 29328 29724 29334 29776
rect 32950 29724 32956 29776
rect 33008 29764 33014 29776
rect 33128 29767 33186 29773
rect 33128 29764 33140 29767
rect 33008 29736 33140 29764
rect 33008 29724 33014 29736
rect 33128 29733 33140 29736
rect 33174 29764 33186 29767
rect 33594 29764 33600 29776
rect 33174 29736 33600 29764
rect 33174 29733 33186 29736
rect 33128 29727 33186 29733
rect 33594 29724 33600 29736
rect 33652 29724 33658 29776
rect 26510 29696 26516 29708
rect 26423 29668 26516 29696
rect 26510 29656 26516 29668
rect 26568 29696 26574 29708
rect 26896 29696 26924 29724
rect 26568 29668 26924 29696
rect 26568 29656 26574 29668
rect 28442 29656 28448 29708
rect 28500 29696 28506 29708
rect 28997 29699 29055 29705
rect 28997 29696 29009 29699
rect 28500 29668 29009 29696
rect 28500 29656 28506 29668
rect 28997 29665 29009 29668
rect 29043 29696 29055 29699
rect 29086 29696 29092 29708
rect 29043 29668 29092 29696
rect 29043 29665 29055 29668
rect 28997 29659 29055 29665
rect 29086 29656 29092 29668
rect 29144 29656 29150 29708
rect 34514 29656 34520 29708
rect 34572 29696 34578 29708
rect 35710 29696 35716 29708
rect 34572 29668 35471 29696
rect 35671 29668 35716 29696
rect 34572 29656 34578 29668
rect 23934 29628 23940 29640
rect 23895 29600 23940 29628
rect 23934 29588 23940 29600
rect 23992 29588 23998 29640
rect 32858 29628 32864 29640
rect 32819 29600 32864 29628
rect 32858 29588 32864 29600
rect 32916 29588 32922 29640
rect 34606 29588 34612 29640
rect 34664 29628 34670 29640
rect 35443 29628 35471 29668
rect 35710 29656 35716 29668
rect 35768 29656 35774 29708
rect 35897 29631 35955 29637
rect 35897 29628 35909 29631
rect 34664 29600 35388 29628
rect 35443 29600 35909 29628
rect 34664 29588 34670 29600
rect 23845 29495 23903 29501
rect 23845 29461 23857 29495
rect 23891 29492 23903 29495
rect 24210 29492 24216 29504
rect 23891 29464 24216 29492
rect 23891 29461 23903 29464
rect 23845 29455 23903 29461
rect 24210 29452 24216 29464
rect 24268 29452 24274 29504
rect 26329 29495 26387 29501
rect 26329 29461 26341 29495
rect 26375 29492 26387 29495
rect 27522 29492 27528 29504
rect 26375 29464 27528 29492
rect 26375 29461 26387 29464
rect 26329 29455 26387 29461
rect 27522 29452 27528 29464
rect 27580 29452 27586 29504
rect 32769 29495 32827 29501
rect 32769 29461 32781 29495
rect 32815 29492 32827 29495
rect 33594 29492 33600 29504
rect 32815 29464 33600 29492
rect 32815 29461 32827 29464
rect 32769 29455 32827 29461
rect 33594 29452 33600 29464
rect 33652 29452 33658 29504
rect 34238 29492 34244 29504
rect 34199 29464 34244 29492
rect 34238 29452 34244 29464
rect 34296 29452 34302 29504
rect 34977 29495 35035 29501
rect 34977 29461 34989 29495
rect 35023 29492 35035 29495
rect 35250 29492 35256 29504
rect 35023 29464 35256 29492
rect 35023 29461 35035 29464
rect 34977 29455 35035 29461
rect 35250 29452 35256 29464
rect 35308 29452 35314 29504
rect 35360 29501 35388 29600
rect 35897 29597 35909 29600
rect 35943 29628 35955 29631
rect 35986 29628 35992 29640
rect 35943 29600 35992 29628
rect 35943 29597 35955 29600
rect 35897 29591 35955 29597
rect 35986 29588 35992 29600
rect 36044 29588 36050 29640
rect 35345 29495 35403 29501
rect 35345 29461 35357 29495
rect 35391 29461 35403 29495
rect 35345 29455 35403 29461
rect 1104 29402 38824 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 38824 29402
rect 1104 29328 38824 29350
rect 24854 29248 24860 29300
rect 24912 29288 24918 29300
rect 25317 29291 25375 29297
rect 25317 29288 25329 29291
rect 24912 29260 25329 29288
rect 24912 29248 24918 29260
rect 25317 29257 25329 29260
rect 25363 29257 25375 29291
rect 25317 29251 25375 29257
rect 25961 29291 26019 29297
rect 25961 29257 25973 29291
rect 26007 29288 26019 29291
rect 26326 29288 26332 29300
rect 26007 29260 26332 29288
rect 26007 29257 26019 29260
rect 25961 29251 26019 29257
rect 26326 29248 26332 29260
rect 26384 29248 26390 29300
rect 26421 29291 26479 29297
rect 26421 29257 26433 29291
rect 26467 29288 26479 29291
rect 27614 29288 27620 29300
rect 26467 29260 27620 29288
rect 26467 29257 26479 29260
rect 26421 29251 26479 29257
rect 27614 29248 27620 29260
rect 27672 29248 27678 29300
rect 32306 29288 32312 29300
rect 32267 29260 32312 29288
rect 32306 29248 32312 29260
rect 32364 29248 32370 29300
rect 32858 29248 32864 29300
rect 32916 29288 32922 29300
rect 32953 29291 33011 29297
rect 32953 29288 32965 29291
rect 32916 29260 32965 29288
rect 32916 29248 32922 29260
rect 32953 29257 32965 29260
rect 32999 29288 33011 29291
rect 33042 29288 33048 29300
rect 32999 29260 33048 29288
rect 32999 29257 33011 29260
rect 32953 29251 33011 29257
rect 33042 29248 33048 29260
rect 33100 29248 33106 29300
rect 35802 29248 35808 29300
rect 35860 29288 35866 29300
rect 36817 29291 36875 29297
rect 36817 29288 36829 29291
rect 35860 29260 36829 29288
rect 35860 29248 35866 29260
rect 36817 29257 36829 29260
rect 36863 29257 36875 29291
rect 36817 29251 36875 29257
rect 37182 29248 37188 29300
rect 37240 29288 37246 29300
rect 37553 29291 37611 29297
rect 37553 29288 37565 29291
rect 37240 29260 37565 29288
rect 37240 29248 37246 29260
rect 37553 29257 37565 29260
rect 37599 29257 37611 29291
rect 37553 29251 37611 29257
rect 27433 29223 27491 29229
rect 27433 29220 27445 29223
rect 26896 29192 27445 29220
rect 26234 29112 26240 29164
rect 26292 29152 26298 29164
rect 26896 29161 26924 29192
rect 27433 29189 27445 29192
rect 27479 29189 27491 29223
rect 27433 29183 27491 29189
rect 28169 29223 28227 29229
rect 28169 29189 28181 29223
rect 28215 29220 28227 29223
rect 28442 29220 28448 29232
rect 28215 29192 28448 29220
rect 28215 29189 28227 29192
rect 28169 29183 28227 29189
rect 28442 29180 28448 29192
rect 28500 29180 28506 29232
rect 30282 29180 30288 29232
rect 30340 29220 30346 29232
rect 30653 29223 30711 29229
rect 30653 29220 30665 29223
rect 30340 29192 30665 29220
rect 30340 29180 30346 29192
rect 30653 29189 30665 29192
rect 30699 29189 30711 29223
rect 36262 29220 36268 29232
rect 36223 29192 36268 29220
rect 30653 29183 30711 29189
rect 36262 29180 36268 29192
rect 36320 29180 36326 29232
rect 26881 29155 26939 29161
rect 26881 29152 26893 29155
rect 26292 29124 26893 29152
rect 26292 29112 26298 29124
rect 26881 29121 26893 29124
rect 26927 29121 26939 29155
rect 26881 29115 26939 29121
rect 27065 29155 27123 29161
rect 27065 29121 27077 29155
rect 27111 29152 27123 29155
rect 27522 29152 27528 29164
rect 27111 29124 27528 29152
rect 27111 29121 27123 29124
rect 27065 29115 27123 29121
rect 27522 29112 27528 29124
rect 27580 29112 27586 29164
rect 32858 29152 32864 29164
rect 30300 29124 32864 29152
rect 23934 29084 23940 29096
rect 23584 29056 23940 29084
rect 23584 28960 23612 29056
rect 23934 29044 23940 29056
rect 23992 29044 23998 29096
rect 24210 29093 24216 29096
rect 24204 29084 24216 29093
rect 24171 29056 24216 29084
rect 24204 29047 24216 29056
rect 24210 29044 24216 29047
rect 24268 29044 24274 29096
rect 26326 29044 26332 29096
rect 26384 29084 26390 29096
rect 26789 29087 26847 29093
rect 26789 29084 26801 29087
rect 26384 29056 26801 29084
rect 26384 29044 26390 29056
rect 26789 29053 26801 29056
rect 26835 29084 26847 29087
rect 27430 29084 27436 29096
rect 26835 29056 27436 29084
rect 26835 29053 26847 29056
rect 26789 29047 26847 29053
rect 27430 29044 27436 29056
rect 27488 29044 27494 29096
rect 27985 29087 28043 29093
rect 27985 29084 27997 29087
rect 27816 29056 27997 29084
rect 26237 29019 26295 29025
rect 26237 28985 26249 29019
rect 26283 29016 26295 29019
rect 26510 29016 26516 29028
rect 26283 28988 26516 29016
rect 26283 28985 26295 28988
rect 26237 28979 26295 28985
rect 26510 28976 26516 28988
rect 26568 28976 26574 29028
rect 27816 28960 27844 29056
rect 27985 29053 27997 29056
rect 28031 29053 28043 29087
rect 29273 29087 29331 29093
rect 29273 29084 29285 29087
rect 27985 29047 28043 29053
rect 29196 29056 29285 29084
rect 29196 29016 29224 29056
rect 29273 29053 29285 29056
rect 29319 29084 29331 29087
rect 30300 29084 30328 29124
rect 32858 29112 32864 29124
rect 32916 29112 32922 29164
rect 33778 29152 33784 29164
rect 33739 29124 33784 29152
rect 33778 29112 33784 29124
rect 33836 29112 33842 29164
rect 34146 29112 34152 29164
rect 34204 29152 34210 29164
rect 34609 29155 34667 29161
rect 34609 29152 34621 29155
rect 34204 29124 34621 29152
rect 34204 29112 34210 29124
rect 34609 29121 34621 29124
rect 34655 29152 34667 29155
rect 34885 29155 34943 29161
rect 34885 29152 34897 29155
rect 34655 29124 34897 29152
rect 34655 29121 34667 29124
rect 34609 29115 34667 29121
rect 34885 29121 34897 29124
rect 34931 29121 34943 29155
rect 34885 29115 34943 29121
rect 29319 29056 30328 29084
rect 32125 29087 32183 29093
rect 29319 29053 29331 29056
rect 29273 29047 29331 29053
rect 32125 29053 32137 29087
rect 32171 29084 32183 29087
rect 33594 29084 33600 29096
rect 32171 29056 32205 29084
rect 33555 29056 33600 29084
rect 32171 29053 32183 29056
rect 32125 29047 32183 29053
rect 29104 28988 29224 29016
rect 29540 29019 29598 29025
rect 29104 28960 29132 28988
rect 29540 28985 29552 29019
rect 29586 29016 29598 29019
rect 29638 29016 29644 29028
rect 29586 28988 29644 29016
rect 29586 28985 29598 28988
rect 29540 28979 29598 28985
rect 29638 28976 29644 28988
rect 29696 28976 29702 29028
rect 32033 29019 32091 29025
rect 32033 28985 32045 29019
rect 32079 29016 32091 29019
rect 32140 29016 32168 29047
rect 33594 29044 33600 29056
rect 33652 29044 33658 29096
rect 34900 29084 34928 29115
rect 34974 29084 34980 29096
rect 34900 29056 34980 29084
rect 34974 29044 34980 29056
rect 35032 29044 35038 29096
rect 37369 29087 37427 29093
rect 37369 29053 37381 29087
rect 37415 29053 37427 29087
rect 37369 29047 37427 29053
rect 33042 29016 33048 29028
rect 32079 28988 33048 29016
rect 32079 28985 32091 28988
rect 32033 28979 32091 28985
rect 33042 28976 33048 28988
rect 33100 28976 33106 29028
rect 33689 29019 33747 29025
rect 33689 28985 33701 29019
rect 33735 29016 33747 29019
rect 34333 29019 34391 29025
rect 34333 29016 34345 29019
rect 33735 28988 34345 29016
rect 33735 28985 33747 28988
rect 33689 28979 33747 28985
rect 34333 28985 34345 28988
rect 34379 29016 34391 29019
rect 34514 29016 34520 29028
rect 34379 28988 34520 29016
rect 34379 28985 34391 28988
rect 34333 28979 34391 28985
rect 34514 28976 34520 28988
rect 34572 29016 34578 29028
rect 35152 29019 35210 29025
rect 35152 29016 35164 29019
rect 34572 28988 35164 29016
rect 34572 28976 34578 28988
rect 35152 28985 35164 28988
rect 35198 29016 35210 29019
rect 35250 29016 35256 29028
rect 35198 28988 35256 29016
rect 35198 28985 35210 28988
rect 35152 28979 35210 28985
rect 35250 28976 35256 28988
rect 35308 28976 35314 29028
rect 37384 29016 37412 29047
rect 38010 29016 38016 29028
rect 37384 28988 38016 29016
rect 38010 28976 38016 28988
rect 38068 28976 38074 29028
rect 23109 28951 23167 28957
rect 23109 28917 23121 28951
rect 23155 28948 23167 28951
rect 23477 28951 23535 28957
rect 23477 28948 23489 28951
rect 23155 28920 23489 28948
rect 23155 28917 23167 28920
rect 23109 28911 23167 28917
rect 23477 28917 23489 28920
rect 23523 28948 23535 28951
rect 23566 28948 23572 28960
rect 23523 28920 23572 28948
rect 23523 28917 23535 28920
rect 23477 28911 23535 28917
rect 23566 28908 23572 28920
rect 23624 28908 23630 28960
rect 27798 28948 27804 28960
rect 27759 28920 27804 28948
rect 27798 28908 27804 28920
rect 27856 28908 27862 28960
rect 28442 28908 28448 28960
rect 28500 28948 28506 28960
rect 28534 28948 28540 28960
rect 28500 28920 28540 28948
rect 28500 28908 28506 28920
rect 28534 28908 28540 28920
rect 28592 28908 28598 28960
rect 28721 28951 28779 28957
rect 28721 28917 28733 28951
rect 28767 28948 28779 28951
rect 29086 28948 29092 28960
rect 28767 28920 29092 28948
rect 28767 28917 28779 28920
rect 28721 28911 28779 28917
rect 29086 28908 29092 28920
rect 29144 28908 29150 28960
rect 33226 28948 33232 28960
rect 33187 28920 33232 28948
rect 33226 28908 33232 28920
rect 33284 28908 33290 28960
rect 1104 28858 38824 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 38824 28858
rect 1104 28784 38824 28806
rect 24210 28704 24216 28756
rect 24268 28744 24274 28756
rect 24765 28747 24823 28753
rect 24765 28744 24777 28747
rect 24268 28716 24777 28744
rect 24268 28704 24274 28716
rect 24765 28713 24777 28716
rect 24811 28713 24823 28747
rect 26326 28744 26332 28756
rect 26287 28716 26332 28744
rect 24765 28707 24823 28713
rect 24780 28676 24808 28707
rect 26326 28704 26332 28716
rect 26384 28704 26390 28756
rect 29089 28747 29147 28753
rect 29089 28713 29101 28747
rect 29135 28744 29147 28747
rect 29270 28744 29276 28756
rect 29135 28716 29276 28744
rect 29135 28713 29147 28716
rect 29089 28707 29147 28713
rect 29270 28704 29276 28716
rect 29328 28704 29334 28756
rect 32950 28744 32956 28756
rect 32911 28716 32956 28744
rect 32950 28704 32956 28716
rect 33008 28704 33014 28756
rect 34514 28704 34520 28756
rect 34572 28744 34578 28756
rect 34609 28747 34667 28753
rect 34609 28744 34621 28747
rect 34572 28716 34621 28744
rect 34572 28704 34578 28716
rect 34609 28713 34621 28716
rect 34655 28713 34667 28747
rect 35342 28744 35348 28756
rect 35303 28716 35348 28744
rect 34609 28707 34667 28713
rect 35342 28704 35348 28716
rect 35400 28704 35406 28756
rect 35897 28747 35955 28753
rect 35897 28713 35909 28747
rect 35943 28744 35955 28747
rect 35986 28744 35992 28756
rect 35943 28716 35992 28744
rect 35943 28713 35955 28716
rect 35897 28707 35955 28713
rect 35986 28704 35992 28716
rect 36044 28744 36050 28756
rect 36265 28747 36323 28753
rect 36265 28744 36277 28747
rect 36044 28716 36277 28744
rect 36044 28704 36050 28716
rect 36265 28713 36277 28716
rect 36311 28713 36323 28747
rect 36265 28707 36323 28713
rect 26881 28679 26939 28685
rect 26881 28676 26893 28679
rect 24780 28648 26893 28676
rect 26881 28645 26893 28648
rect 26927 28676 26939 28679
rect 27062 28676 27068 28688
rect 26927 28648 27068 28676
rect 26927 28645 26939 28648
rect 26881 28639 26939 28645
rect 27062 28636 27068 28648
rect 27120 28636 27126 28688
rect 29448 28679 29506 28685
rect 29448 28645 29460 28679
rect 29494 28676 29506 28679
rect 29546 28676 29552 28688
rect 29494 28648 29552 28676
rect 29494 28645 29506 28648
rect 29448 28639 29506 28645
rect 29546 28636 29552 28648
rect 29604 28676 29610 28688
rect 30282 28676 30288 28688
rect 29604 28648 30288 28676
rect 29604 28636 29610 28648
rect 30282 28636 30288 28648
rect 30340 28636 30346 28688
rect 23474 28568 23480 28620
rect 23532 28608 23538 28620
rect 23641 28611 23699 28617
rect 23641 28608 23653 28611
rect 23532 28580 23653 28608
rect 23532 28568 23538 28580
rect 23641 28577 23653 28580
rect 23687 28577 23699 28611
rect 23641 28571 23699 28577
rect 27614 28568 27620 28620
rect 27672 28608 27678 28620
rect 28074 28608 28080 28620
rect 27672 28580 28080 28608
rect 27672 28568 27678 28580
rect 28074 28568 28080 28580
rect 28132 28568 28138 28620
rect 32858 28568 32864 28620
rect 32916 28608 32922 28620
rect 33042 28608 33048 28620
rect 32916 28580 33048 28608
rect 32916 28568 32922 28580
rect 33042 28568 33048 28580
rect 33100 28608 33106 28620
rect 33229 28611 33287 28617
rect 33229 28608 33241 28611
rect 33100 28580 33241 28608
rect 33100 28568 33106 28580
rect 33229 28577 33241 28580
rect 33275 28577 33287 28611
rect 33229 28571 33287 28577
rect 33496 28611 33554 28617
rect 33496 28577 33508 28611
rect 33542 28608 33554 28611
rect 34238 28608 34244 28620
rect 33542 28580 34244 28608
rect 33542 28577 33554 28580
rect 33496 28571 33554 28577
rect 34238 28568 34244 28580
rect 34296 28568 34302 28620
rect 35713 28611 35771 28617
rect 35713 28577 35725 28611
rect 35759 28608 35771 28611
rect 35986 28608 35992 28620
rect 35759 28580 35992 28608
rect 35759 28577 35771 28580
rect 35713 28571 35771 28577
rect 35986 28568 35992 28580
rect 36044 28568 36050 28620
rect 23385 28543 23443 28549
rect 23385 28509 23397 28543
rect 23431 28509 23443 28543
rect 26970 28540 26976 28552
rect 26931 28512 26976 28540
rect 23385 28503 23443 28509
rect 23400 28404 23428 28503
rect 26970 28500 26976 28512
rect 27028 28500 27034 28552
rect 27154 28540 27160 28552
rect 27115 28512 27160 28540
rect 27154 28500 27160 28512
rect 27212 28500 27218 28552
rect 29086 28500 29092 28552
rect 29144 28540 29150 28552
rect 29181 28543 29239 28549
rect 29181 28540 29193 28543
rect 29144 28512 29193 28540
rect 29144 28500 29150 28512
rect 29181 28509 29193 28512
rect 29227 28509 29239 28543
rect 29181 28503 29239 28509
rect 23566 28404 23572 28416
rect 23400 28376 23572 28404
rect 23566 28364 23572 28376
rect 23624 28364 23630 28416
rect 26326 28364 26332 28416
rect 26384 28404 26390 28416
rect 26513 28407 26571 28413
rect 26513 28404 26525 28407
rect 26384 28376 26525 28404
rect 26384 28364 26390 28376
rect 26513 28373 26525 28376
rect 26559 28373 26571 28407
rect 27614 28404 27620 28416
rect 27575 28376 27620 28404
rect 26513 28367 26571 28373
rect 27614 28364 27620 28376
rect 27672 28364 27678 28416
rect 28258 28404 28264 28416
rect 28219 28376 28264 28404
rect 28258 28364 28264 28376
rect 28316 28364 28322 28416
rect 30282 28364 30288 28416
rect 30340 28404 30346 28416
rect 30561 28407 30619 28413
rect 30561 28404 30573 28407
rect 30340 28376 30573 28404
rect 30340 28364 30346 28376
rect 30561 28373 30573 28376
rect 30607 28373 30619 28407
rect 30561 28367 30619 28373
rect 32585 28407 32643 28413
rect 32585 28373 32597 28407
rect 32631 28404 32643 28407
rect 36078 28404 36084 28416
rect 32631 28376 36084 28404
rect 32631 28373 32643 28376
rect 32585 28367 32643 28373
rect 36078 28364 36084 28376
rect 36136 28404 36142 28416
rect 36722 28404 36728 28416
rect 36136 28376 36728 28404
rect 36136 28364 36142 28376
rect 36722 28364 36728 28376
rect 36780 28364 36786 28416
rect 1104 28314 38824 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 38824 28314
rect 1104 28240 38824 28262
rect 22741 28203 22799 28209
rect 22741 28169 22753 28203
rect 22787 28200 22799 28203
rect 23474 28200 23480 28212
rect 22787 28172 23480 28200
rect 22787 28169 22799 28172
rect 22741 28163 22799 28169
rect 23474 28160 23480 28172
rect 23532 28200 23538 28212
rect 25041 28203 25099 28209
rect 25041 28200 25053 28203
rect 23532 28172 25053 28200
rect 23532 28160 23538 28172
rect 25041 28169 25053 28172
rect 25087 28200 25099 28203
rect 26697 28203 26755 28209
rect 26697 28200 26709 28203
rect 25087 28172 26709 28200
rect 25087 28169 25099 28172
rect 25041 28163 25099 28169
rect 26697 28169 26709 28172
rect 26743 28200 26755 28203
rect 26970 28200 26976 28212
rect 26743 28172 26976 28200
rect 26743 28169 26755 28172
rect 26697 28163 26755 28169
rect 26970 28160 26976 28172
rect 27028 28160 27034 28212
rect 27062 28160 27068 28212
rect 27120 28200 27126 28212
rect 27617 28203 27675 28209
rect 27120 28172 27165 28200
rect 27120 28160 27126 28172
rect 27617 28169 27629 28203
rect 27663 28200 27675 28203
rect 27798 28200 27804 28212
rect 27663 28172 27804 28200
rect 27663 28169 27675 28172
rect 27617 28163 27675 28169
rect 27798 28160 27804 28172
rect 27856 28160 27862 28212
rect 32582 28200 32588 28212
rect 32543 28172 32588 28200
rect 32582 28160 32588 28172
rect 32640 28160 32646 28212
rect 33134 28160 33140 28212
rect 33192 28200 33198 28212
rect 33229 28203 33287 28209
rect 33229 28200 33241 28203
rect 33192 28172 33241 28200
rect 33192 28160 33198 28172
rect 33229 28169 33241 28172
rect 33275 28169 33287 28203
rect 34238 28200 34244 28212
rect 34199 28172 34244 28200
rect 33229 28163 33287 28169
rect 34238 28160 34244 28172
rect 34296 28160 34302 28212
rect 35526 28160 35532 28212
rect 35584 28200 35590 28212
rect 35621 28203 35679 28209
rect 35621 28200 35633 28203
rect 35584 28172 35633 28200
rect 35584 28160 35590 28172
rect 35621 28169 35633 28172
rect 35667 28169 35679 28203
rect 36722 28200 36728 28212
rect 36683 28172 36728 28200
rect 35621 28163 35679 28169
rect 36722 28160 36728 28172
rect 36780 28160 36786 28212
rect 24854 28092 24860 28144
rect 24912 28132 24918 28144
rect 25593 28135 25651 28141
rect 25593 28132 25605 28135
rect 24912 28104 25605 28132
rect 24912 28092 24918 28104
rect 25593 28101 25605 28104
rect 25639 28132 25651 28135
rect 27154 28132 27160 28144
rect 25639 28104 27160 28132
rect 25639 28101 25651 28104
rect 25593 28095 25651 28101
rect 27154 28092 27160 28104
rect 27212 28092 27218 28144
rect 34609 28135 34667 28141
rect 34609 28132 34621 28135
rect 33704 28104 34621 28132
rect 27614 28024 27620 28076
rect 27672 28064 27678 28076
rect 28169 28067 28227 28073
rect 28169 28064 28181 28067
rect 27672 28036 28181 28064
rect 27672 28024 27678 28036
rect 28169 28033 28181 28036
rect 28215 28033 28227 28067
rect 33134 28064 33140 28076
rect 33095 28036 33140 28064
rect 28169 28027 28227 28033
rect 33134 28024 33140 28036
rect 33192 28024 33198 28076
rect 33410 28024 33416 28076
rect 33468 28064 33474 28076
rect 33704 28073 33732 28104
rect 34609 28101 34621 28104
rect 34655 28101 34667 28135
rect 34609 28095 34667 28101
rect 33689 28067 33747 28073
rect 33689 28064 33701 28067
rect 33468 28036 33701 28064
rect 33468 28024 33474 28036
rect 33689 28033 33701 28036
rect 33735 28033 33747 28067
rect 33689 28027 33747 28033
rect 33873 28067 33931 28073
rect 33873 28033 33885 28067
rect 33919 28064 33931 28067
rect 34330 28064 34336 28076
rect 33919 28036 34336 28064
rect 33919 28033 33931 28036
rect 33873 28027 33931 28033
rect 23566 27956 23572 28008
rect 23624 27996 23630 28008
rect 23661 27999 23719 28005
rect 23661 27996 23673 27999
rect 23624 27968 23673 27996
rect 23624 27956 23630 27968
rect 23661 27965 23673 27968
rect 23707 27965 23719 27999
rect 23661 27959 23719 27965
rect 26145 27999 26203 28005
rect 26145 27965 26157 27999
rect 26191 27965 26203 27999
rect 26145 27959 26203 27965
rect 27525 27999 27583 28005
rect 27525 27965 27537 27999
rect 27571 27996 27583 27999
rect 28077 27999 28135 28005
rect 28077 27996 28089 27999
rect 27571 27968 28089 27996
rect 27571 27965 27583 27968
rect 27525 27959 27583 27965
rect 28077 27965 28089 27968
rect 28123 27996 28135 27999
rect 28902 27996 28908 28008
rect 28123 27968 28908 27996
rect 28123 27965 28135 27968
rect 28077 27959 28135 27965
rect 23109 27931 23167 27937
rect 23109 27897 23121 27931
rect 23155 27928 23167 27931
rect 23474 27928 23480 27940
rect 23155 27900 23480 27928
rect 23155 27897 23167 27900
rect 23109 27891 23167 27897
rect 23474 27888 23480 27900
rect 23532 27928 23538 27940
rect 23906 27931 23964 27937
rect 23906 27928 23918 27931
rect 23532 27900 23918 27928
rect 23532 27888 23538 27900
rect 23906 27897 23918 27900
rect 23952 27928 23964 27931
rect 24210 27928 24216 27940
rect 23952 27900 24216 27928
rect 23952 27897 23964 27900
rect 23906 27891 23964 27897
rect 24210 27888 24216 27900
rect 24268 27888 24274 27940
rect 26160 27872 26188 27959
rect 28902 27956 28908 27968
rect 28960 27956 28966 28008
rect 29457 27999 29515 28005
rect 29457 27996 29469 27999
rect 29104 27968 29469 27996
rect 28721 27931 28779 27937
rect 28721 27897 28733 27931
rect 28767 27928 28779 27931
rect 29104 27928 29132 27968
rect 29457 27965 29469 27968
rect 29503 27965 29515 27999
rect 29457 27959 29515 27965
rect 31941 27999 31999 28005
rect 31941 27965 31953 27999
rect 31987 27996 31999 27999
rect 32582 27996 32588 28008
rect 31987 27968 32588 27996
rect 31987 27965 31999 27968
rect 31941 27959 31999 27965
rect 32582 27956 32588 27968
rect 32640 27956 32646 28008
rect 33226 27956 33232 28008
rect 33284 27996 33290 28008
rect 33597 27999 33655 28005
rect 33597 27996 33609 27999
rect 33284 27968 33609 27996
rect 33284 27956 33290 27968
rect 33597 27965 33609 27968
rect 33643 27965 33655 27999
rect 33597 27959 33655 27965
rect 28767 27900 29132 27928
rect 28767 27897 28779 27900
rect 28721 27891 28779 27897
rect 29104 27872 29132 27900
rect 29270 27888 29276 27940
rect 29328 27928 29334 27940
rect 29702 27931 29760 27937
rect 29702 27928 29714 27931
rect 29328 27900 29714 27928
rect 29328 27888 29334 27900
rect 29702 27897 29714 27900
rect 29748 27897 29760 27931
rect 31846 27928 31852 27940
rect 31759 27900 31852 27928
rect 29702 27891 29760 27897
rect 31846 27888 31852 27900
rect 31904 27928 31910 27940
rect 33888 27928 33916 28027
rect 34330 28024 34336 28036
rect 34388 28024 34394 28076
rect 35437 27999 35495 28005
rect 35437 27996 35449 27999
rect 31904 27900 33916 27928
rect 35268 27968 35449 27996
rect 31904 27888 31910 27900
rect 23385 27863 23443 27869
rect 23385 27829 23397 27863
rect 23431 27860 23443 27863
rect 23566 27860 23572 27872
rect 23431 27832 23572 27860
rect 23431 27829 23443 27832
rect 23385 27823 23443 27829
rect 23566 27820 23572 27832
rect 23624 27820 23630 27872
rect 26053 27863 26111 27869
rect 26053 27829 26065 27863
rect 26099 27860 26111 27863
rect 26142 27860 26148 27872
rect 26099 27832 26148 27860
rect 26099 27829 26111 27832
rect 26053 27823 26111 27829
rect 26142 27820 26148 27832
rect 26200 27820 26206 27872
rect 26329 27863 26387 27869
rect 26329 27829 26341 27863
rect 26375 27860 26387 27863
rect 26602 27860 26608 27872
rect 26375 27832 26608 27860
rect 26375 27829 26387 27832
rect 26329 27823 26387 27829
rect 26602 27820 26608 27832
rect 26660 27820 26666 27872
rect 27982 27860 27988 27872
rect 27943 27832 27988 27860
rect 27982 27820 27988 27832
rect 28040 27820 28046 27872
rect 29086 27860 29092 27872
rect 29047 27832 29092 27860
rect 29086 27820 29092 27832
rect 29144 27820 29150 27872
rect 30650 27820 30656 27872
rect 30708 27860 30714 27872
rect 30837 27863 30895 27869
rect 30837 27860 30849 27863
rect 30708 27832 30849 27860
rect 30708 27820 30714 27832
rect 30837 27829 30849 27832
rect 30883 27829 30895 27863
rect 32122 27860 32128 27872
rect 32083 27832 32128 27860
rect 30837 27823 30895 27829
rect 32122 27820 32128 27832
rect 32180 27820 32186 27872
rect 34606 27820 34612 27872
rect 34664 27860 34670 27872
rect 35268 27869 35296 27968
rect 35437 27965 35449 27968
rect 35483 27965 35495 27999
rect 35437 27959 35495 27965
rect 36541 27999 36599 28005
rect 36541 27965 36553 27999
rect 36587 27996 36599 27999
rect 36587 27968 37228 27996
rect 36587 27965 36599 27968
rect 36541 27959 36599 27965
rect 37200 27872 37228 27968
rect 35253 27863 35311 27869
rect 35253 27860 35265 27863
rect 34664 27832 35265 27860
rect 34664 27820 34670 27832
rect 35253 27829 35265 27832
rect 35299 27829 35311 27863
rect 35986 27860 35992 27872
rect 35947 27832 35992 27860
rect 35253 27823 35311 27829
rect 35986 27820 35992 27832
rect 36044 27820 36050 27872
rect 37182 27860 37188 27872
rect 37143 27832 37188 27860
rect 37182 27820 37188 27832
rect 37240 27820 37246 27872
rect 1104 27770 38824 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 38824 27770
rect 1104 27696 38824 27718
rect 24210 27656 24216 27668
rect 24171 27628 24216 27656
rect 24210 27616 24216 27628
rect 24268 27616 24274 27668
rect 27709 27659 27767 27665
rect 27709 27625 27721 27659
rect 27755 27656 27767 27659
rect 27982 27656 27988 27668
rect 27755 27628 27988 27656
rect 27755 27625 27767 27628
rect 27709 27619 27767 27625
rect 27982 27616 27988 27628
rect 28040 27656 28046 27668
rect 28905 27659 28963 27665
rect 28905 27656 28917 27659
rect 28040 27628 28917 27656
rect 28040 27616 28046 27628
rect 28905 27625 28917 27628
rect 28951 27625 28963 27659
rect 28905 27619 28963 27625
rect 29365 27659 29423 27665
rect 29365 27625 29377 27659
rect 29411 27656 29423 27659
rect 29546 27656 29552 27668
rect 29411 27628 29552 27656
rect 29411 27625 29423 27628
rect 29365 27619 29423 27625
rect 24854 27548 24860 27600
rect 24912 27548 24918 27600
rect 28074 27588 28080 27600
rect 28035 27560 28080 27588
rect 28074 27548 28080 27560
rect 28132 27548 28138 27600
rect 28718 27548 28724 27600
rect 28776 27588 28782 27600
rect 28813 27591 28871 27597
rect 28813 27588 28825 27591
rect 28776 27560 28825 27588
rect 28776 27548 28782 27560
rect 28813 27557 28825 27560
rect 28859 27588 28871 27591
rect 29380 27588 29408 27619
rect 29546 27616 29552 27628
rect 29604 27616 29610 27668
rect 33226 27656 33232 27668
rect 33060 27628 33232 27656
rect 28859 27560 29408 27588
rect 32861 27591 32919 27597
rect 28859 27557 28871 27560
rect 28813 27551 28871 27557
rect 32861 27557 32873 27591
rect 32907 27588 32919 27591
rect 33060 27588 33088 27628
rect 33226 27616 33232 27628
rect 33284 27616 33290 27668
rect 32907 27560 33088 27588
rect 32907 27557 32919 27560
rect 32861 27551 32919 27557
rect 33594 27548 33600 27600
rect 33652 27588 33658 27600
rect 35406 27591 35464 27597
rect 35406 27588 35418 27591
rect 33652 27560 35418 27588
rect 33652 27548 33658 27560
rect 35406 27557 35418 27560
rect 35452 27557 35464 27591
rect 35406 27551 35464 27557
rect 35526 27548 35532 27600
rect 35584 27548 35590 27600
rect 24302 27452 24308 27464
rect 24263 27424 24308 27452
rect 24302 27412 24308 27424
rect 24360 27412 24366 27464
rect 24489 27455 24547 27461
rect 24489 27421 24501 27455
rect 24535 27452 24547 27455
rect 24872 27452 24900 27548
rect 26326 27480 26332 27532
rect 26384 27520 26390 27532
rect 26881 27523 26939 27529
rect 26881 27520 26893 27523
rect 26384 27492 26893 27520
rect 26384 27480 26390 27492
rect 26881 27489 26893 27492
rect 26927 27489 26939 27523
rect 29270 27520 29276 27532
rect 29231 27492 29276 27520
rect 26881 27483 26939 27489
rect 29270 27480 29276 27492
rect 29328 27520 29334 27532
rect 30282 27520 30288 27532
rect 29328 27492 30288 27520
rect 29328 27480 29334 27492
rect 30282 27480 30288 27492
rect 30340 27480 30346 27532
rect 30466 27520 30472 27532
rect 30427 27492 30472 27520
rect 30466 27480 30472 27492
rect 30524 27480 30530 27532
rect 30650 27520 30656 27532
rect 30611 27492 30656 27520
rect 30650 27480 30656 27492
rect 30708 27480 30714 27532
rect 30837 27523 30895 27529
rect 30837 27489 30849 27523
rect 30883 27520 30895 27523
rect 31938 27520 31944 27532
rect 30883 27492 31944 27520
rect 30883 27489 30895 27492
rect 30837 27483 30895 27489
rect 31938 27480 31944 27492
rect 31996 27520 32002 27532
rect 32125 27523 32183 27529
rect 32125 27520 32137 27523
rect 31996 27492 32137 27520
rect 31996 27480 32002 27492
rect 32125 27489 32137 27492
rect 32171 27489 32183 27523
rect 32125 27483 32183 27489
rect 33134 27480 33140 27532
rect 33192 27520 33198 27532
rect 33689 27523 33747 27529
rect 33689 27520 33701 27523
rect 33192 27492 33701 27520
rect 33192 27480 33198 27492
rect 33689 27489 33701 27492
rect 33735 27489 33747 27523
rect 33689 27483 33747 27489
rect 33781 27523 33839 27529
rect 33781 27489 33793 27523
rect 33827 27520 33839 27523
rect 35161 27523 35219 27529
rect 33827 27492 34744 27520
rect 33827 27489 33839 27492
rect 33781 27483 33839 27489
rect 24535 27424 24900 27452
rect 24535 27421 24547 27424
rect 24489 27415 24547 27421
rect 23385 27387 23443 27393
rect 23385 27353 23397 27387
rect 23431 27384 23443 27387
rect 24504 27384 24532 27415
rect 26418 27412 26424 27464
rect 26476 27452 26482 27464
rect 26973 27455 27031 27461
rect 26973 27452 26985 27455
rect 26476 27424 26985 27452
rect 26476 27412 26482 27424
rect 26973 27421 26985 27424
rect 27019 27421 27031 27455
rect 27154 27452 27160 27464
rect 27115 27424 27160 27452
rect 26973 27415 27031 27421
rect 27154 27412 27160 27424
rect 27212 27452 27218 27464
rect 27522 27452 27528 27464
rect 27212 27424 27528 27452
rect 27212 27412 27218 27424
rect 27522 27412 27528 27424
rect 27580 27412 27586 27464
rect 29454 27452 29460 27464
rect 29415 27424 29460 27452
rect 29454 27412 29460 27424
rect 29512 27412 29518 27464
rect 30009 27455 30067 27461
rect 30009 27421 30021 27455
rect 30055 27452 30067 27455
rect 30668 27452 30696 27480
rect 30055 27424 30696 27452
rect 30055 27421 30067 27424
rect 30009 27415 30067 27421
rect 32766 27412 32772 27464
rect 32824 27452 32830 27464
rect 33796 27452 33824 27483
rect 34716 27464 34744 27492
rect 35161 27489 35173 27523
rect 35207 27520 35219 27523
rect 35250 27520 35256 27532
rect 35207 27492 35256 27520
rect 35207 27489 35219 27492
rect 35161 27483 35219 27489
rect 35250 27480 35256 27492
rect 35308 27520 35314 27532
rect 35544 27520 35572 27548
rect 35308 27492 35572 27520
rect 35308 27480 35314 27492
rect 32824 27424 33824 27452
rect 33965 27455 34023 27461
rect 32824 27412 32830 27424
rect 33965 27421 33977 27455
rect 34011 27452 34023 27455
rect 34011 27424 34468 27452
rect 34011 27421 34023 27424
rect 33965 27415 34023 27421
rect 23431 27356 24532 27384
rect 26329 27387 26387 27393
rect 23431 27353 23443 27356
rect 23385 27347 23443 27353
rect 26329 27353 26341 27387
rect 26375 27384 26387 27387
rect 27172 27384 27200 27412
rect 33226 27384 33232 27396
rect 26375 27356 27200 27384
rect 33187 27356 33232 27384
rect 26375 27353 26387 27356
rect 26329 27347 26387 27353
rect 33226 27344 33232 27356
rect 33284 27344 33290 27396
rect 34440 27328 34468 27424
rect 34698 27412 34704 27464
rect 34756 27412 34762 27464
rect 23566 27276 23572 27328
rect 23624 27316 23630 27328
rect 23661 27319 23719 27325
rect 23661 27316 23673 27319
rect 23624 27288 23673 27316
rect 23624 27276 23630 27288
rect 23661 27285 23673 27288
rect 23707 27285 23719 27319
rect 23842 27316 23848 27328
rect 23803 27288 23848 27316
rect 23661 27279 23719 27285
rect 23842 27276 23848 27288
rect 23900 27276 23906 27328
rect 26510 27316 26516 27328
rect 26471 27288 26516 27316
rect 26510 27276 26516 27288
rect 26568 27276 26574 27328
rect 32306 27316 32312 27328
rect 32267 27288 32312 27316
rect 32306 27276 32312 27288
rect 32364 27276 32370 27328
rect 33318 27316 33324 27328
rect 33279 27288 33324 27316
rect 33318 27276 33324 27288
rect 33376 27276 33382 27328
rect 34422 27316 34428 27328
rect 34383 27288 34428 27316
rect 34422 27276 34428 27288
rect 34480 27276 34486 27328
rect 36538 27316 36544 27328
rect 36499 27288 36544 27316
rect 36538 27276 36544 27288
rect 36596 27276 36602 27328
rect 1104 27226 38824 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 38824 27226
rect 1104 27152 38824 27174
rect 22370 27112 22376 27124
rect 22331 27084 22376 27112
rect 22370 27072 22376 27084
rect 22428 27072 22434 27124
rect 23474 27072 23480 27124
rect 23532 27112 23538 27124
rect 25041 27115 25099 27121
rect 25041 27112 25053 27115
rect 23532 27084 25053 27112
rect 23532 27072 23538 27084
rect 25041 27081 25053 27084
rect 25087 27081 25099 27115
rect 25041 27075 25099 27081
rect 26329 27115 26387 27121
rect 26329 27081 26341 27115
rect 26375 27112 26387 27115
rect 26418 27112 26424 27124
rect 26375 27084 26424 27112
rect 26375 27081 26387 27084
rect 26329 27075 26387 27081
rect 26418 27072 26424 27084
rect 26476 27072 26482 27124
rect 26602 27072 26608 27124
rect 26660 27112 26666 27124
rect 26973 27115 27031 27121
rect 26973 27112 26985 27115
rect 26660 27084 26985 27112
rect 26660 27072 26666 27084
rect 26973 27081 26985 27084
rect 27019 27081 27031 27115
rect 26973 27075 27031 27081
rect 28353 27115 28411 27121
rect 28353 27081 28365 27115
rect 28399 27112 28411 27115
rect 29270 27112 29276 27124
rect 28399 27084 29276 27112
rect 28399 27081 28411 27084
rect 28353 27075 28411 27081
rect 26988 26976 27016 27075
rect 29270 27072 29276 27084
rect 29328 27072 29334 27124
rect 30650 27072 30656 27124
rect 30708 27112 30714 27124
rect 31481 27115 31539 27121
rect 31481 27112 31493 27115
rect 30708 27084 31493 27112
rect 30708 27072 30714 27084
rect 31481 27081 31493 27084
rect 31527 27081 31539 27115
rect 31481 27075 31539 27081
rect 32309 27115 32367 27121
rect 32309 27081 32321 27115
rect 32355 27112 32367 27115
rect 33134 27112 33140 27124
rect 32355 27084 33140 27112
rect 32355 27081 32367 27084
rect 32309 27075 32367 27081
rect 33134 27072 33140 27084
rect 33192 27072 33198 27124
rect 33594 27072 33600 27124
rect 33652 27112 33658 27124
rect 34241 27115 34299 27121
rect 34241 27112 34253 27115
rect 33652 27084 34253 27112
rect 33652 27072 33658 27084
rect 34241 27081 34253 27084
rect 34287 27081 34299 27115
rect 34241 27075 34299 27081
rect 35710 27072 35716 27124
rect 35768 27112 35774 27124
rect 36446 27112 36452 27124
rect 35768 27084 36452 27112
rect 35768 27072 35774 27084
rect 36446 27072 36452 27084
rect 36504 27072 36510 27124
rect 28718 27044 28724 27056
rect 28679 27016 28724 27044
rect 28718 27004 28724 27016
rect 28776 27004 28782 27056
rect 32766 27044 32772 27056
rect 32727 27016 32772 27044
rect 32766 27004 32772 27016
rect 32824 27004 32830 27056
rect 33229 27047 33287 27053
rect 33229 27013 33241 27047
rect 33275 27044 33287 27047
rect 34514 27044 34520 27056
rect 33275 27016 34520 27044
rect 33275 27013 33287 27016
rect 33229 27007 33287 27013
rect 34514 27004 34520 27016
rect 34572 27004 34578 27056
rect 36814 27044 36820 27056
rect 36775 27016 36820 27044
rect 36814 27004 36820 27016
rect 36872 27004 36878 27056
rect 27617 26979 27675 26985
rect 27617 26976 27629 26979
rect 26988 26948 27629 26976
rect 27617 26945 27629 26948
rect 27663 26945 27675 26979
rect 27798 26976 27804 26988
rect 27759 26948 27804 26976
rect 27617 26939 27675 26945
rect 27798 26936 27804 26948
rect 27856 26936 27862 26988
rect 33870 26976 33876 26988
rect 33831 26948 33876 26976
rect 33870 26936 33876 26948
rect 33928 26936 33934 26988
rect 22370 26868 22376 26920
rect 22428 26908 22434 26920
rect 22465 26911 22523 26917
rect 22465 26908 22477 26911
rect 22428 26880 22477 26908
rect 22428 26868 22434 26880
rect 22465 26877 22477 26880
rect 22511 26877 22523 26911
rect 22465 26871 22523 26877
rect 23566 26868 23572 26920
rect 23624 26908 23630 26920
rect 23661 26911 23719 26917
rect 23661 26908 23673 26911
rect 23624 26880 23673 26908
rect 23624 26868 23630 26880
rect 23661 26877 23673 26880
rect 23707 26877 23719 26911
rect 29549 26911 29607 26917
rect 29549 26908 29561 26911
rect 23661 26871 23719 26877
rect 29288 26880 29561 26908
rect 23109 26843 23167 26849
rect 23109 26809 23121 26843
rect 23155 26840 23167 26843
rect 23906 26843 23964 26849
rect 23906 26840 23918 26843
rect 23155 26812 23918 26840
rect 23155 26809 23167 26812
rect 23109 26803 23167 26809
rect 23906 26809 23918 26812
rect 23952 26840 23964 26843
rect 24302 26840 24308 26852
rect 23952 26812 24308 26840
rect 23952 26809 23964 26812
rect 23906 26803 23964 26809
rect 24302 26800 24308 26812
rect 24360 26840 24366 26852
rect 25593 26843 25651 26849
rect 25593 26840 25605 26843
rect 24360 26812 25605 26840
rect 24360 26800 24366 26812
rect 25593 26809 25605 26812
rect 25639 26809 25651 26843
rect 27525 26843 27583 26849
rect 27525 26840 27537 26843
rect 25593 26803 25651 26809
rect 26620 26812 27537 26840
rect 26620 26784 26648 26812
rect 27525 26809 27537 26812
rect 27571 26809 27583 26843
rect 27525 26803 27583 26809
rect 29288 26784 29316 26880
rect 29549 26877 29561 26880
rect 29595 26877 29607 26911
rect 29549 26871 29607 26877
rect 29816 26911 29874 26917
rect 29816 26877 29828 26911
rect 29862 26908 29874 26911
rect 30650 26908 30656 26920
rect 29862 26880 30656 26908
rect 29862 26877 29874 26880
rect 29816 26871 29874 26877
rect 30650 26868 30656 26880
rect 30708 26868 30714 26920
rect 32033 26911 32091 26917
rect 32033 26877 32045 26911
rect 32079 26908 32091 26911
rect 32125 26911 32183 26917
rect 32125 26908 32137 26911
rect 32079 26880 32137 26908
rect 32079 26877 32091 26880
rect 32033 26871 32091 26877
rect 32125 26877 32137 26880
rect 32171 26908 32183 26911
rect 33226 26908 33232 26920
rect 32171 26880 33232 26908
rect 32171 26877 32183 26880
rect 32125 26871 32183 26877
rect 33226 26868 33232 26880
rect 33284 26908 33290 26920
rect 33689 26911 33747 26917
rect 33689 26908 33701 26911
rect 33284 26880 33701 26908
rect 33284 26868 33290 26880
rect 33689 26877 33701 26880
rect 33735 26877 33747 26911
rect 33689 26871 33747 26877
rect 35345 26911 35403 26917
rect 35345 26877 35357 26911
rect 35391 26908 35403 26911
rect 35437 26911 35495 26917
rect 35437 26908 35449 26911
rect 35391 26880 35449 26908
rect 35391 26877 35403 26880
rect 35345 26871 35403 26877
rect 35437 26877 35449 26880
rect 35483 26908 35495 26911
rect 35526 26908 35532 26920
rect 35483 26880 35532 26908
rect 35483 26877 35495 26880
rect 35437 26871 35495 26877
rect 35526 26868 35532 26880
rect 35584 26868 35590 26920
rect 35710 26917 35716 26920
rect 35704 26908 35716 26917
rect 35623 26880 35716 26908
rect 32858 26800 32864 26852
rect 32916 26840 32922 26852
rect 33597 26843 33655 26849
rect 33597 26840 33609 26843
rect 32916 26812 33609 26840
rect 32916 26800 32922 26812
rect 33597 26809 33609 26812
rect 33643 26840 33655 26843
rect 34330 26840 34336 26852
rect 33643 26812 34336 26840
rect 33643 26809 33655 26812
rect 33597 26803 33655 26809
rect 34330 26800 34336 26812
rect 34388 26800 34394 26852
rect 34701 26843 34759 26849
rect 34701 26809 34713 26843
rect 34747 26840 34759 26843
rect 35636 26840 35664 26880
rect 35704 26871 35716 26880
rect 35768 26908 35774 26920
rect 36538 26908 36544 26920
rect 35768 26880 36544 26908
rect 35710 26868 35716 26871
rect 35768 26868 35774 26880
rect 36538 26868 36544 26880
rect 36596 26868 36602 26920
rect 34747 26812 35664 26840
rect 34747 26809 34759 26812
rect 34701 26803 34759 26809
rect 22646 26772 22652 26784
rect 22607 26744 22652 26772
rect 22646 26732 22652 26744
rect 22704 26732 22710 26784
rect 23477 26775 23535 26781
rect 23477 26741 23489 26775
rect 23523 26772 23535 26775
rect 23566 26772 23572 26784
rect 23523 26744 23572 26772
rect 23523 26741 23535 26744
rect 23477 26735 23535 26741
rect 23566 26732 23572 26744
rect 23624 26732 23630 26784
rect 26602 26772 26608 26784
rect 26563 26744 26608 26772
rect 26602 26732 26608 26744
rect 26660 26732 26666 26784
rect 27157 26775 27215 26781
rect 27157 26741 27169 26775
rect 27203 26772 27215 26775
rect 27706 26772 27712 26784
rect 27203 26744 27712 26772
rect 27203 26741 27215 26744
rect 27157 26735 27215 26741
rect 27706 26732 27712 26744
rect 27764 26732 27770 26784
rect 29086 26772 29092 26784
rect 28999 26744 29092 26772
rect 29086 26732 29092 26744
rect 29144 26772 29150 26784
rect 29270 26772 29276 26784
rect 29144 26744 29276 26772
rect 29144 26732 29150 26744
rect 29270 26732 29276 26744
rect 29328 26732 29334 26784
rect 30834 26732 30840 26784
rect 30892 26772 30898 26784
rect 30929 26775 30987 26781
rect 30929 26772 30941 26775
rect 30892 26744 30941 26772
rect 30892 26732 30898 26744
rect 30929 26741 30941 26744
rect 30975 26741 30987 26775
rect 30929 26735 30987 26741
rect 1104 26682 38824 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 38824 26682
rect 1104 26608 38824 26630
rect 23474 26568 23480 26580
rect 23435 26540 23480 26568
rect 23474 26528 23480 26540
rect 23532 26528 23538 26580
rect 24302 26528 24308 26580
rect 24360 26568 24366 26580
rect 24949 26571 25007 26577
rect 24949 26568 24961 26571
rect 24360 26540 24961 26568
rect 24360 26528 24366 26540
rect 24949 26537 24961 26540
rect 24995 26537 25007 26571
rect 24949 26531 25007 26537
rect 26234 26528 26240 26580
rect 26292 26568 26298 26580
rect 26513 26571 26571 26577
rect 26513 26568 26525 26571
rect 26292 26540 26525 26568
rect 26292 26528 26298 26540
rect 26513 26537 26525 26540
rect 26559 26537 26571 26571
rect 26513 26531 26571 26537
rect 28077 26571 28135 26577
rect 28077 26537 28089 26571
rect 28123 26537 28135 26571
rect 28077 26531 28135 26537
rect 23750 26460 23756 26512
rect 23808 26509 23814 26512
rect 23808 26503 23872 26509
rect 23808 26469 23826 26503
rect 23860 26469 23872 26503
rect 26326 26500 26332 26512
rect 26287 26472 26332 26500
rect 23808 26463 23872 26469
rect 23808 26460 23814 26463
rect 26326 26460 26332 26472
rect 26384 26460 26390 26512
rect 26878 26432 26884 26444
rect 26839 26404 26884 26432
rect 26878 26392 26884 26404
rect 26936 26392 26942 26444
rect 26973 26435 27031 26441
rect 26973 26401 26985 26435
rect 27019 26432 27031 26435
rect 27522 26432 27528 26444
rect 27019 26404 27528 26432
rect 27019 26401 27031 26404
rect 26973 26395 27031 26401
rect 27522 26392 27528 26404
rect 27580 26392 27586 26444
rect 28092 26432 28120 26531
rect 28258 26528 28264 26580
rect 28316 26568 28322 26580
rect 28537 26571 28595 26577
rect 28537 26568 28549 26571
rect 28316 26540 28549 26568
rect 28316 26528 28322 26540
rect 28537 26537 28549 26540
rect 28583 26537 28595 26571
rect 28537 26531 28595 26537
rect 28810 26528 28816 26580
rect 28868 26568 28874 26580
rect 29641 26571 29699 26577
rect 29641 26568 29653 26571
rect 28868 26540 29653 26568
rect 28868 26528 28874 26540
rect 29641 26537 29653 26540
rect 29687 26537 29699 26571
rect 29641 26531 29699 26537
rect 30466 26528 30472 26580
rect 30524 26568 30530 26580
rect 30653 26571 30711 26577
rect 30653 26568 30665 26571
rect 30524 26540 30665 26568
rect 30524 26528 30530 26540
rect 30653 26537 30665 26540
rect 30699 26537 30711 26571
rect 31938 26568 31944 26580
rect 31899 26540 31944 26568
rect 30653 26531 30711 26537
rect 31938 26528 31944 26540
rect 31996 26528 32002 26580
rect 32493 26571 32551 26577
rect 32493 26537 32505 26571
rect 32539 26568 32551 26571
rect 33870 26568 33876 26580
rect 32539 26540 33876 26568
rect 32539 26537 32551 26540
rect 32493 26531 32551 26537
rect 33870 26528 33876 26540
rect 33928 26528 33934 26580
rect 35253 26571 35311 26577
rect 35253 26537 35265 26571
rect 35299 26568 35311 26571
rect 35526 26568 35532 26580
rect 35299 26540 35532 26568
rect 35299 26537 35311 26540
rect 35253 26531 35311 26537
rect 35526 26528 35532 26540
rect 35584 26528 35590 26580
rect 28442 26500 28448 26512
rect 28403 26472 28448 26500
rect 28442 26460 28448 26472
rect 28500 26460 28506 26512
rect 28997 26503 29055 26509
rect 28997 26469 29009 26503
rect 29043 26500 29055 26503
rect 29181 26503 29239 26509
rect 29181 26500 29193 26503
rect 29043 26472 29193 26500
rect 29043 26469 29055 26472
rect 28997 26463 29055 26469
rect 29181 26469 29193 26472
rect 29227 26500 29239 26503
rect 29454 26500 29460 26512
rect 29227 26472 29460 26500
rect 29227 26469 29239 26472
rect 29181 26463 29239 26469
rect 29454 26460 29460 26472
rect 29512 26500 29518 26512
rect 30374 26500 30380 26512
rect 29512 26472 30380 26500
rect 29512 26460 29518 26472
rect 30374 26460 30380 26472
rect 30432 26460 30438 26512
rect 32858 26500 32864 26512
rect 32819 26472 32864 26500
rect 32858 26460 32864 26472
rect 32916 26460 32922 26512
rect 33220 26503 33278 26509
rect 33220 26469 33232 26503
rect 33266 26500 33278 26503
rect 34422 26500 34428 26512
rect 33266 26472 34428 26500
rect 33266 26469 33278 26472
rect 33220 26463 33278 26469
rect 34422 26460 34428 26472
rect 34480 26460 34486 26512
rect 35621 26503 35679 26509
rect 35621 26469 35633 26503
rect 35667 26500 35679 26503
rect 35710 26500 35716 26512
rect 35667 26472 35716 26500
rect 35667 26469 35679 26472
rect 35621 26463 35679 26469
rect 35710 26460 35716 26472
rect 35768 26500 35774 26512
rect 35986 26500 35992 26512
rect 35768 26472 35992 26500
rect 35768 26460 35774 26472
rect 35986 26460 35992 26472
rect 36044 26460 36050 26512
rect 30009 26435 30067 26441
rect 30009 26432 30021 26435
rect 28092 26404 30021 26432
rect 30009 26401 30021 26404
rect 30055 26432 30067 26435
rect 30190 26432 30196 26444
rect 30055 26404 30196 26432
rect 30055 26401 30067 26404
rect 30009 26395 30067 26401
rect 30190 26392 30196 26404
rect 30248 26392 30254 26444
rect 32953 26435 33011 26441
rect 32953 26401 32965 26435
rect 32999 26432 33011 26435
rect 33042 26432 33048 26444
rect 32999 26404 33048 26432
rect 32999 26401 33011 26404
rect 32953 26395 33011 26401
rect 33042 26392 33048 26404
rect 33100 26392 33106 26444
rect 35437 26435 35495 26441
rect 35437 26401 35449 26435
rect 35483 26432 35495 26435
rect 35526 26432 35532 26444
rect 35483 26404 35532 26432
rect 35483 26401 35495 26404
rect 35437 26395 35495 26401
rect 35526 26392 35532 26404
rect 35584 26392 35590 26444
rect 23566 26364 23572 26376
rect 23527 26336 23572 26364
rect 23566 26324 23572 26336
rect 23624 26324 23630 26376
rect 25961 26367 26019 26373
rect 25961 26333 25973 26367
rect 26007 26364 26019 26367
rect 27154 26364 27160 26376
rect 26007 26336 27160 26364
rect 26007 26333 26019 26336
rect 25961 26327 26019 26333
rect 27154 26324 27160 26336
rect 27212 26324 27218 26376
rect 27617 26367 27675 26373
rect 27617 26333 27629 26367
rect 27663 26364 27675 26367
rect 27798 26364 27804 26376
rect 27663 26336 27804 26364
rect 27663 26333 27675 26336
rect 27617 26327 27675 26333
rect 27798 26324 27804 26336
rect 27856 26364 27862 26376
rect 28718 26364 28724 26376
rect 27856 26336 28724 26364
rect 27856 26324 27862 26336
rect 28718 26324 28724 26336
rect 28776 26324 28782 26376
rect 29822 26324 29828 26376
rect 29880 26364 29886 26376
rect 30101 26367 30159 26373
rect 30101 26364 30113 26367
rect 29880 26336 30113 26364
rect 29880 26324 29886 26336
rect 30101 26333 30113 26336
rect 30147 26333 30159 26367
rect 30282 26364 30288 26376
rect 30243 26336 30288 26364
rect 30101 26327 30159 26333
rect 30282 26324 30288 26336
rect 30340 26324 30346 26376
rect 27062 26256 27068 26308
rect 27120 26296 27126 26308
rect 28997 26299 29055 26305
rect 28997 26296 29009 26299
rect 27120 26268 29009 26296
rect 27120 26256 27126 26268
rect 28997 26265 29009 26268
rect 29043 26265 29055 26299
rect 28997 26259 29055 26265
rect 29549 26299 29607 26305
rect 29549 26265 29561 26299
rect 29595 26296 29607 26299
rect 30300 26296 30328 26324
rect 29595 26268 30328 26296
rect 35805 26299 35863 26305
rect 29595 26265 29607 26268
rect 29549 26259 29607 26265
rect 35805 26265 35817 26299
rect 35851 26296 35863 26299
rect 35894 26296 35900 26308
rect 35851 26268 35900 26296
rect 35851 26265 35863 26268
rect 35805 26259 35863 26265
rect 35894 26256 35900 26268
rect 35952 26256 35958 26308
rect 34330 26228 34336 26240
rect 34291 26200 34336 26228
rect 34330 26188 34336 26200
rect 34388 26188 34394 26240
rect 1104 26138 38824 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 38824 26138
rect 1104 26064 38824 26086
rect 26326 25984 26332 26036
rect 26384 26024 26390 26036
rect 26513 26027 26571 26033
rect 26513 26024 26525 26027
rect 26384 25996 26525 26024
rect 26384 25984 26390 25996
rect 26513 25993 26525 25996
rect 26559 26024 26571 26027
rect 26878 26024 26884 26036
rect 26559 25996 26884 26024
rect 26559 25993 26571 25996
rect 26513 25987 26571 25993
rect 26878 25984 26884 25996
rect 26936 25984 26942 26036
rect 28258 25984 28264 26036
rect 28316 26024 28322 26036
rect 28629 26027 28687 26033
rect 28629 26024 28641 26027
rect 28316 25996 28641 26024
rect 28316 25984 28322 25996
rect 28629 25993 28641 25996
rect 28675 25993 28687 26027
rect 28629 25987 28687 25993
rect 32769 26027 32827 26033
rect 32769 25993 32781 26027
rect 32815 26024 32827 26027
rect 32950 26024 32956 26036
rect 32815 25996 32956 26024
rect 32815 25993 32827 25996
rect 32769 25987 32827 25993
rect 32950 25984 32956 25996
rect 33008 25984 33014 26036
rect 33965 26027 34023 26033
rect 33965 25993 33977 26027
rect 34011 26024 34023 26027
rect 34422 26024 34428 26036
rect 34011 25996 34428 26024
rect 34011 25993 34023 25996
rect 33965 25987 34023 25993
rect 34422 25984 34428 25996
rect 34480 25984 34486 26036
rect 34514 25984 34520 26036
rect 34572 26024 34578 26036
rect 34609 26027 34667 26033
rect 34609 26024 34621 26027
rect 34572 25996 34621 26024
rect 34572 25984 34578 25996
rect 34609 25993 34621 25996
rect 34655 25993 34667 26027
rect 34609 25987 34667 25993
rect 25409 25959 25467 25965
rect 25409 25925 25421 25959
rect 25455 25956 25467 25959
rect 26421 25959 26479 25965
rect 26421 25956 26433 25959
rect 25455 25928 26433 25956
rect 25455 25925 25467 25928
rect 25409 25919 25467 25925
rect 26421 25925 26433 25928
rect 26467 25956 26479 25959
rect 26786 25956 26792 25968
rect 26467 25928 26792 25956
rect 26467 25925 26479 25928
rect 26421 25919 26479 25925
rect 26786 25916 26792 25928
rect 26844 25956 26850 25968
rect 27985 25959 28043 25965
rect 26844 25928 27016 25956
rect 26844 25916 26850 25928
rect 26988 25897 27016 25928
rect 27985 25925 27997 25959
rect 28031 25956 28043 25959
rect 28442 25956 28448 25968
rect 28031 25928 28448 25956
rect 28031 25925 28043 25928
rect 27985 25919 28043 25925
rect 28442 25916 28448 25928
rect 28500 25916 28506 25968
rect 32861 25959 32919 25965
rect 32861 25925 32873 25959
rect 32907 25956 32919 25959
rect 33042 25956 33048 25968
rect 32907 25928 33048 25956
rect 32907 25925 32919 25928
rect 32861 25919 32919 25925
rect 33042 25916 33048 25928
rect 33100 25916 33106 25968
rect 26973 25891 27031 25897
rect 26973 25857 26985 25891
rect 27019 25857 27031 25891
rect 26973 25851 27031 25857
rect 27062 25848 27068 25900
rect 27120 25888 27126 25900
rect 32401 25891 32459 25897
rect 27120 25860 27165 25888
rect 27120 25848 27126 25860
rect 32401 25857 32413 25891
rect 32447 25888 32459 25891
rect 33502 25888 33508 25900
rect 32447 25860 33508 25888
rect 32447 25857 32459 25860
rect 32401 25851 32459 25857
rect 33502 25848 33508 25860
rect 33560 25888 33566 25900
rect 34330 25888 34336 25900
rect 33560 25860 34336 25888
rect 33560 25848 33566 25860
rect 34330 25848 34336 25860
rect 34388 25848 34394 25900
rect 23477 25823 23535 25829
rect 23477 25789 23489 25823
rect 23523 25820 23535 25823
rect 23566 25820 23572 25832
rect 23523 25792 23572 25820
rect 23523 25789 23535 25792
rect 23477 25783 23535 25789
rect 23566 25780 23572 25792
rect 23624 25820 23630 25832
rect 23934 25820 23940 25832
rect 23624 25792 23940 25820
rect 23624 25780 23630 25792
rect 23934 25780 23940 25792
rect 23992 25820 23998 25832
rect 24029 25823 24087 25829
rect 24029 25820 24041 25823
rect 23992 25792 24041 25820
rect 23992 25780 23998 25792
rect 24029 25789 24041 25792
rect 24075 25789 24087 25823
rect 24029 25783 24087 25789
rect 27706 25780 27712 25832
rect 27764 25820 27770 25832
rect 28077 25823 28135 25829
rect 28077 25820 28089 25823
rect 27764 25792 28089 25820
rect 27764 25780 27770 25792
rect 28077 25789 28089 25792
rect 28123 25820 28135 25823
rect 28442 25820 28448 25832
rect 28123 25792 28448 25820
rect 28123 25789 28135 25792
rect 28077 25783 28135 25789
rect 28442 25780 28448 25792
rect 28500 25820 28506 25832
rect 28997 25823 29055 25829
rect 28997 25820 29009 25823
rect 28500 25792 29009 25820
rect 28500 25780 28506 25792
rect 28997 25789 29009 25792
rect 29043 25820 29055 25823
rect 29822 25820 29828 25832
rect 29043 25792 29828 25820
rect 29043 25789 29055 25792
rect 28997 25783 29055 25789
rect 29822 25780 29828 25792
rect 29880 25780 29886 25832
rect 29917 25823 29975 25829
rect 29917 25789 29929 25823
rect 29963 25789 29975 25823
rect 29917 25783 29975 25789
rect 32033 25823 32091 25829
rect 32033 25789 32045 25823
rect 32079 25820 32091 25823
rect 33318 25820 33324 25832
rect 32079 25792 33324 25820
rect 32079 25789 32091 25792
rect 32033 25783 32091 25789
rect 23109 25755 23167 25761
rect 23109 25721 23121 25755
rect 23155 25752 23167 25755
rect 23750 25752 23756 25764
rect 23155 25724 23756 25752
rect 23155 25721 23167 25724
rect 23109 25715 23167 25721
rect 23750 25712 23756 25724
rect 23808 25752 23814 25764
rect 24302 25761 24308 25764
rect 24296 25752 24308 25761
rect 23808 25724 24072 25752
rect 24263 25724 24308 25752
rect 23808 25712 23814 25724
rect 23934 25684 23940 25696
rect 23895 25656 23940 25684
rect 23934 25644 23940 25656
rect 23992 25644 23998 25696
rect 24044 25684 24072 25724
rect 24296 25715 24308 25724
rect 24302 25712 24308 25715
rect 24360 25712 24366 25764
rect 29932 25752 29960 25783
rect 33318 25780 33324 25792
rect 33376 25780 33382 25832
rect 34624 25820 34652 25987
rect 34698 25984 34704 26036
rect 34756 26024 34762 26036
rect 35069 26027 35127 26033
rect 35069 26024 35081 26027
rect 34756 25996 35081 26024
rect 34756 25984 34762 25996
rect 35069 25993 35081 25996
rect 35115 25993 35127 26027
rect 35069 25987 35127 25993
rect 35897 26027 35955 26033
rect 35897 25993 35909 26027
rect 35943 26024 35955 26027
rect 35986 26024 35992 26036
rect 35943 25996 35992 26024
rect 35943 25993 35955 25996
rect 35897 25987 35955 25993
rect 35986 25984 35992 25996
rect 36044 25984 36050 26036
rect 36170 26024 36176 26036
rect 36131 25996 36176 26024
rect 36170 25984 36176 25996
rect 36228 25984 36234 26036
rect 34885 25823 34943 25829
rect 34885 25820 34897 25823
rect 34624 25792 34897 25820
rect 34885 25789 34897 25792
rect 34931 25789 34943 25823
rect 34885 25783 34943 25789
rect 35894 25780 35900 25832
rect 35952 25820 35958 25832
rect 35989 25823 36047 25829
rect 35989 25820 36001 25823
rect 35952 25792 36001 25820
rect 35952 25780 35958 25792
rect 35989 25789 36001 25792
rect 36035 25820 36047 25823
rect 36541 25823 36599 25829
rect 36541 25820 36553 25823
rect 36035 25792 36553 25820
rect 36035 25789 36047 25792
rect 35989 25783 36047 25789
rect 36541 25789 36553 25792
rect 36587 25789 36599 25823
rect 36541 25783 36599 25789
rect 29748 25724 29960 25752
rect 26053 25687 26111 25693
rect 26053 25684 26065 25687
rect 24044 25656 26065 25684
rect 26053 25653 26065 25656
rect 26099 25684 26111 25687
rect 26878 25684 26884 25696
rect 26099 25656 26884 25684
rect 26099 25653 26111 25656
rect 26053 25647 26111 25653
rect 26878 25644 26884 25656
rect 26936 25644 26942 25696
rect 27614 25684 27620 25696
rect 27575 25656 27620 25684
rect 27614 25644 27620 25656
rect 27672 25644 27678 25696
rect 28258 25684 28264 25696
rect 28219 25656 28264 25684
rect 28258 25644 28264 25656
rect 28316 25644 28322 25696
rect 29270 25644 29276 25696
rect 29328 25684 29334 25696
rect 29748 25693 29776 25724
rect 30006 25712 30012 25764
rect 30064 25752 30070 25764
rect 30184 25755 30242 25761
rect 30184 25752 30196 25755
rect 30064 25724 30196 25752
rect 30064 25712 30070 25724
rect 30184 25721 30196 25724
rect 30230 25752 30242 25755
rect 30834 25752 30840 25764
rect 30230 25724 30840 25752
rect 30230 25721 30242 25724
rect 30184 25715 30242 25721
rect 30834 25712 30840 25724
rect 30892 25712 30898 25764
rect 29733 25687 29791 25693
rect 29733 25684 29745 25687
rect 29328 25656 29745 25684
rect 29328 25644 29334 25656
rect 29733 25653 29745 25656
rect 29779 25653 29791 25687
rect 31294 25684 31300 25696
rect 31255 25656 31300 25684
rect 29733 25647 29791 25653
rect 31294 25644 31300 25656
rect 31352 25644 31358 25696
rect 32950 25644 32956 25696
rect 33008 25684 33014 25696
rect 33229 25687 33287 25693
rect 33229 25684 33241 25687
rect 33008 25656 33241 25684
rect 33008 25644 33014 25656
rect 33229 25653 33241 25656
rect 33275 25653 33287 25687
rect 35526 25684 35532 25696
rect 35487 25656 35532 25684
rect 33229 25647 33287 25653
rect 35526 25644 35532 25656
rect 35584 25644 35590 25696
rect 1104 25594 38824 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 38824 25594
rect 1104 25520 38824 25542
rect 26326 25480 26332 25492
rect 26287 25452 26332 25480
rect 26326 25440 26332 25452
rect 26384 25440 26390 25492
rect 26878 25440 26884 25492
rect 26936 25480 26942 25492
rect 27893 25483 27951 25489
rect 27893 25480 27905 25483
rect 26936 25452 27905 25480
rect 26936 25440 26942 25452
rect 27893 25449 27905 25452
rect 27939 25449 27951 25483
rect 27893 25443 27951 25449
rect 28258 25440 28264 25492
rect 28316 25480 28322 25492
rect 29733 25483 29791 25489
rect 29733 25480 29745 25483
rect 28316 25452 29745 25480
rect 28316 25440 28322 25452
rect 29733 25449 29745 25452
rect 29779 25480 29791 25483
rect 30098 25480 30104 25492
rect 29779 25452 30104 25480
rect 29779 25449 29791 25452
rect 29733 25443 29791 25449
rect 30098 25440 30104 25452
rect 30156 25440 30162 25492
rect 30190 25440 30196 25492
rect 30248 25480 30254 25492
rect 30469 25483 30527 25489
rect 30469 25480 30481 25483
rect 30248 25452 30481 25480
rect 30248 25440 30254 25452
rect 30469 25449 30481 25452
rect 30515 25449 30527 25483
rect 30834 25480 30840 25492
rect 30795 25452 30840 25480
rect 30469 25443 30527 25449
rect 30834 25440 30840 25452
rect 30892 25440 30898 25492
rect 31113 25483 31171 25489
rect 31113 25449 31125 25483
rect 31159 25449 31171 25483
rect 31113 25443 31171 25449
rect 32125 25483 32183 25489
rect 32125 25449 32137 25483
rect 32171 25480 32183 25483
rect 32950 25480 32956 25492
rect 32171 25452 32956 25480
rect 32171 25449 32183 25452
rect 32125 25443 32183 25449
rect 26786 25421 26792 25424
rect 26780 25412 26792 25421
rect 26747 25384 26792 25412
rect 26780 25375 26792 25384
rect 26786 25372 26792 25375
rect 26844 25372 26850 25424
rect 28442 25412 28448 25424
rect 28403 25384 28448 25412
rect 28442 25372 28448 25384
rect 28500 25372 28506 25424
rect 28718 25372 28724 25424
rect 28776 25412 28782 25424
rect 28813 25415 28871 25421
rect 28813 25412 28825 25415
rect 28776 25384 28825 25412
rect 28776 25372 28782 25384
rect 28813 25381 28825 25384
rect 28859 25381 28871 25415
rect 28813 25375 28871 25381
rect 30374 25372 30380 25424
rect 30432 25412 30438 25424
rect 31128 25412 31156 25443
rect 32950 25440 32956 25452
rect 33008 25440 33014 25492
rect 30432 25384 31156 25412
rect 33404 25415 33462 25421
rect 30432 25372 30438 25384
rect 33404 25381 33416 25415
rect 33450 25412 33462 25415
rect 33502 25412 33508 25424
rect 33450 25384 33508 25412
rect 33450 25381 33462 25384
rect 33404 25375 33462 25381
rect 33502 25372 33508 25384
rect 33560 25372 33566 25424
rect 24210 25353 24216 25356
rect 24204 25344 24216 25353
rect 24171 25316 24216 25344
rect 24204 25307 24216 25316
rect 24210 25304 24216 25307
rect 24268 25304 24274 25356
rect 25222 25304 25228 25356
rect 25280 25344 25286 25356
rect 25961 25347 26019 25353
rect 25961 25344 25973 25347
rect 25280 25316 25973 25344
rect 25280 25304 25286 25316
rect 25961 25313 25973 25316
rect 26007 25344 26019 25347
rect 27062 25344 27068 25356
rect 26007 25316 27068 25344
rect 26007 25313 26019 25316
rect 25961 25307 26019 25313
rect 27062 25304 27068 25316
rect 27120 25304 27126 25356
rect 30926 25344 30932 25356
rect 30887 25316 30932 25344
rect 30926 25304 30932 25316
rect 30984 25304 30990 25356
rect 33134 25344 33140 25356
rect 33095 25316 33140 25344
rect 33134 25304 33140 25316
rect 33192 25304 33198 25356
rect 23934 25276 23940 25288
rect 23895 25248 23940 25276
rect 23934 25236 23940 25248
rect 23992 25236 23998 25288
rect 26510 25276 26516 25288
rect 26471 25248 26516 25276
rect 26510 25236 26516 25248
rect 26568 25236 26574 25288
rect 29825 25279 29883 25285
rect 29825 25276 29837 25279
rect 29196 25248 29837 25276
rect 23845 25143 23903 25149
rect 23845 25109 23857 25143
rect 23891 25140 23903 25143
rect 24302 25140 24308 25152
rect 23891 25112 24308 25140
rect 23891 25109 23903 25112
rect 23845 25103 23903 25109
rect 24302 25100 24308 25112
rect 24360 25140 24366 25152
rect 24946 25140 24952 25152
rect 24360 25112 24952 25140
rect 24360 25100 24366 25112
rect 24946 25100 24952 25112
rect 25004 25140 25010 25152
rect 25317 25143 25375 25149
rect 25317 25140 25329 25143
rect 25004 25112 25329 25140
rect 25004 25100 25010 25112
rect 25317 25109 25329 25112
rect 25363 25109 25375 25143
rect 25317 25103 25375 25109
rect 28994 25100 29000 25152
rect 29052 25140 29058 25152
rect 29196 25149 29224 25248
rect 29825 25245 29837 25248
rect 29871 25245 29883 25279
rect 30006 25276 30012 25288
rect 29967 25248 30012 25276
rect 29825 25239 29883 25245
rect 30006 25236 30012 25248
rect 30064 25236 30070 25288
rect 29365 25211 29423 25217
rect 29365 25177 29377 25211
rect 29411 25208 29423 25211
rect 29411 25180 31800 25208
rect 29411 25177 29423 25180
rect 29365 25171 29423 25177
rect 31772 25152 31800 25180
rect 29181 25143 29239 25149
rect 29181 25140 29193 25143
rect 29052 25112 29193 25140
rect 29052 25100 29058 25112
rect 29181 25109 29193 25112
rect 29227 25109 29239 25143
rect 29181 25103 29239 25109
rect 31754 25100 31760 25152
rect 31812 25140 31818 25152
rect 34514 25140 34520 25152
rect 31812 25112 31857 25140
rect 34475 25112 34520 25140
rect 31812 25100 31818 25112
rect 34514 25100 34520 25112
rect 34572 25100 34578 25152
rect 35161 25143 35219 25149
rect 35161 25109 35173 25143
rect 35207 25140 35219 25143
rect 35434 25140 35440 25152
rect 35207 25112 35440 25140
rect 35207 25109 35219 25112
rect 35161 25103 35219 25109
rect 35434 25100 35440 25112
rect 35492 25100 35498 25152
rect 1104 25050 38824 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 38824 25050
rect 1104 24976 38824 24998
rect 26510 24936 26516 24948
rect 26471 24908 26516 24936
rect 26510 24896 26516 24908
rect 26568 24896 26574 24948
rect 26786 24896 26792 24948
rect 26844 24936 26850 24948
rect 26881 24939 26939 24945
rect 26881 24936 26893 24939
rect 26844 24908 26893 24936
rect 26844 24896 26850 24908
rect 26881 24905 26893 24908
rect 26927 24905 26939 24939
rect 26881 24899 26939 24905
rect 30926 24896 30932 24948
rect 30984 24936 30990 24948
rect 31205 24939 31263 24945
rect 31205 24936 31217 24939
rect 30984 24908 31217 24936
rect 30984 24896 30990 24908
rect 31205 24905 31217 24908
rect 31251 24905 31263 24939
rect 33134 24936 33140 24948
rect 33095 24908 33140 24936
rect 31205 24899 31263 24905
rect 33134 24896 33140 24908
rect 33192 24896 33198 24948
rect 33502 24936 33508 24948
rect 33463 24908 33508 24936
rect 33502 24896 33508 24908
rect 33560 24896 33566 24948
rect 31294 24828 31300 24880
rect 31352 24868 31358 24880
rect 31352 24840 32352 24868
rect 31352 24828 31358 24840
rect 27985 24803 28043 24809
rect 27985 24769 27997 24803
rect 28031 24800 28043 24803
rect 28810 24800 28816 24812
rect 28031 24772 28816 24800
rect 28031 24769 28043 24772
rect 27985 24763 28043 24769
rect 28092 24741 28120 24772
rect 28810 24760 28816 24772
rect 28868 24760 28874 24812
rect 29089 24803 29147 24809
rect 29089 24769 29101 24803
rect 29135 24800 29147 24803
rect 29270 24800 29276 24812
rect 29135 24772 29276 24800
rect 29135 24769 29147 24772
rect 29089 24763 29147 24769
rect 29270 24760 29276 24772
rect 29328 24760 29334 24812
rect 31754 24760 31760 24812
rect 31812 24800 31818 24812
rect 32324 24809 32352 24840
rect 32217 24803 32275 24809
rect 32217 24800 32229 24803
rect 31812 24772 32229 24800
rect 31812 24760 31818 24772
rect 32217 24769 32229 24772
rect 32263 24769 32275 24803
rect 32217 24763 32275 24769
rect 32309 24803 32367 24809
rect 32309 24769 32321 24803
rect 32355 24769 32367 24803
rect 34238 24800 34244 24812
rect 32309 24763 32367 24769
rect 33704 24772 34244 24800
rect 33704 24741 33732 24772
rect 34238 24760 34244 24772
rect 34296 24760 34302 24812
rect 35434 24800 35440 24812
rect 35395 24772 35440 24800
rect 35434 24760 35440 24772
rect 35492 24760 35498 24812
rect 24489 24735 24547 24741
rect 24489 24732 24501 24735
rect 24320 24704 24501 24732
rect 23934 24596 23940 24608
rect 23895 24568 23940 24596
rect 23934 24556 23940 24568
rect 23992 24596 23998 24608
rect 24320 24605 24348 24704
rect 24489 24701 24501 24704
rect 24535 24701 24547 24735
rect 24489 24695 24547 24701
rect 28077 24735 28135 24741
rect 28077 24701 28089 24735
rect 28123 24732 28135 24735
rect 28721 24735 28779 24741
rect 28123 24704 28157 24732
rect 28123 24701 28135 24704
rect 28077 24695 28135 24701
rect 28721 24701 28733 24735
rect 28767 24732 28779 24735
rect 33689 24735 33747 24741
rect 28767 24704 29224 24732
rect 28767 24701 28779 24704
rect 28721 24695 28779 24701
rect 24670 24624 24676 24676
rect 24728 24673 24734 24676
rect 24728 24667 24792 24673
rect 24728 24633 24746 24667
rect 24780 24633 24792 24667
rect 28902 24664 28908 24676
rect 24728 24627 24792 24633
rect 28276 24636 28908 24664
rect 24728 24624 24734 24627
rect 24305 24599 24363 24605
rect 24305 24596 24317 24599
rect 23992 24568 24317 24596
rect 23992 24556 23998 24568
rect 24305 24565 24317 24568
rect 24351 24565 24363 24599
rect 24305 24559 24363 24565
rect 25038 24556 25044 24608
rect 25096 24596 25102 24608
rect 28276 24605 28304 24636
rect 28902 24624 28908 24636
rect 28960 24624 28966 24676
rect 29196 24664 29224 24704
rect 33689 24701 33701 24735
rect 33735 24701 33747 24735
rect 33689 24695 33747 24701
rect 34422 24692 34428 24744
rect 34480 24732 34486 24744
rect 35345 24735 35403 24741
rect 35345 24732 35357 24735
rect 34480 24704 35357 24732
rect 34480 24692 34486 24704
rect 35345 24701 35357 24704
rect 35391 24732 35403 24735
rect 35897 24735 35955 24741
rect 35897 24732 35909 24735
rect 35391 24704 35909 24732
rect 35391 24701 35403 24704
rect 35345 24695 35403 24701
rect 35897 24701 35909 24704
rect 35943 24701 35955 24735
rect 35897 24695 35955 24701
rect 29546 24673 29552 24676
rect 29540 24664 29552 24673
rect 29196 24636 29552 24664
rect 29540 24627 29552 24636
rect 29546 24624 29552 24627
rect 29604 24624 29610 24676
rect 30374 24624 30380 24676
rect 30432 24664 30438 24676
rect 31573 24667 31631 24673
rect 31573 24664 31585 24667
rect 30432 24636 31585 24664
rect 30432 24624 30438 24636
rect 31573 24633 31585 24636
rect 31619 24664 31631 24667
rect 32125 24667 32183 24673
rect 32125 24664 32137 24667
rect 31619 24636 32137 24664
rect 31619 24633 31631 24636
rect 31573 24627 31631 24633
rect 32125 24633 32137 24636
rect 32171 24633 32183 24667
rect 34330 24664 34336 24676
rect 32125 24627 32183 24633
rect 33888 24636 34336 24664
rect 25869 24599 25927 24605
rect 25869 24596 25881 24599
rect 25096 24568 25881 24596
rect 25096 24556 25102 24568
rect 25869 24565 25881 24568
rect 25915 24565 25927 24599
rect 25869 24559 25927 24565
rect 28261 24599 28319 24605
rect 28261 24565 28273 24599
rect 28307 24565 28319 24599
rect 28261 24559 28319 24565
rect 29914 24556 29920 24608
rect 29972 24596 29978 24608
rect 30653 24599 30711 24605
rect 30653 24596 30665 24599
rect 29972 24568 30665 24596
rect 29972 24556 29978 24568
rect 30653 24565 30665 24568
rect 30699 24565 30711 24599
rect 30653 24559 30711 24565
rect 31754 24556 31760 24608
rect 31812 24596 31818 24608
rect 33888 24605 33916 24636
rect 34330 24624 34336 24636
rect 34388 24624 34394 24676
rect 35253 24667 35311 24673
rect 35253 24664 35265 24667
rect 34624 24636 35265 24664
rect 34624 24608 34652 24636
rect 35253 24633 35265 24636
rect 35299 24633 35311 24667
rect 35253 24627 35311 24633
rect 33873 24599 33931 24605
rect 31812 24568 31857 24596
rect 31812 24556 31818 24568
rect 33873 24565 33885 24599
rect 33919 24565 33931 24599
rect 34606 24596 34612 24608
rect 34567 24568 34612 24596
rect 33873 24559 33931 24565
rect 34606 24556 34612 24568
rect 34664 24556 34670 24608
rect 34882 24596 34888 24608
rect 34843 24568 34888 24596
rect 34882 24556 34888 24568
rect 34940 24556 34946 24608
rect 1104 24506 38824 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 38824 24506
rect 1104 24432 38824 24454
rect 24029 24395 24087 24401
rect 24029 24361 24041 24395
rect 24075 24392 24087 24395
rect 24210 24392 24216 24404
rect 24075 24364 24216 24392
rect 24075 24361 24087 24364
rect 24029 24355 24087 24361
rect 24210 24352 24216 24364
rect 24268 24392 24274 24404
rect 25038 24392 25044 24404
rect 24268 24364 25044 24392
rect 24268 24352 24274 24364
rect 25038 24352 25044 24364
rect 25096 24352 25102 24404
rect 30098 24392 30104 24404
rect 30059 24364 30104 24392
rect 30098 24352 30104 24364
rect 30156 24352 30162 24404
rect 30561 24395 30619 24401
rect 30561 24361 30573 24395
rect 30607 24392 30619 24395
rect 30834 24392 30840 24404
rect 30607 24364 30840 24392
rect 30607 24361 30619 24364
rect 30561 24355 30619 24361
rect 30834 24352 30840 24364
rect 30892 24352 30898 24404
rect 31294 24352 31300 24404
rect 31352 24392 31358 24404
rect 31757 24395 31815 24401
rect 31757 24392 31769 24395
rect 31352 24364 31769 24392
rect 31352 24352 31358 24364
rect 31757 24361 31769 24364
rect 31803 24361 31815 24395
rect 31757 24355 31815 24361
rect 35345 24395 35403 24401
rect 35345 24361 35357 24395
rect 35391 24392 35403 24395
rect 35434 24392 35440 24404
rect 35391 24364 35440 24392
rect 35391 24361 35403 24364
rect 35345 24355 35403 24361
rect 35434 24352 35440 24364
rect 35492 24352 35498 24404
rect 24489 24327 24547 24333
rect 24489 24293 24501 24327
rect 24535 24324 24547 24327
rect 24670 24324 24676 24336
rect 24535 24296 24676 24324
rect 24535 24293 24547 24296
rect 24489 24287 24547 24293
rect 24670 24284 24676 24296
rect 24728 24284 24734 24336
rect 24946 24256 24952 24268
rect 24907 24228 24952 24256
rect 24946 24216 24952 24228
rect 25004 24216 25010 24268
rect 28074 24216 28080 24268
rect 28132 24256 28138 24268
rect 28436 24259 28494 24265
rect 28436 24256 28448 24259
rect 28132 24228 28448 24256
rect 28132 24216 28138 24228
rect 28436 24225 28448 24228
rect 28482 24256 28494 24259
rect 29914 24256 29920 24268
rect 28482 24228 29920 24256
rect 28482 24225 28494 24228
rect 28436 24219 28494 24225
rect 29914 24216 29920 24228
rect 29972 24216 29978 24268
rect 30650 24256 30656 24268
rect 30611 24228 30656 24256
rect 30650 24216 30656 24228
rect 30708 24216 30714 24268
rect 33870 24216 33876 24268
rect 33928 24256 33934 24268
rect 34221 24259 34279 24265
rect 34221 24256 34233 24259
rect 33928 24228 34233 24256
rect 33928 24216 33934 24228
rect 34221 24225 34233 24228
rect 34267 24256 34279 24259
rect 34514 24256 34520 24268
rect 34267 24228 34520 24256
rect 34267 24225 34279 24228
rect 34221 24219 34279 24225
rect 34514 24216 34520 24228
rect 34572 24216 34578 24268
rect 25222 24188 25228 24200
rect 25183 24160 25228 24188
rect 25222 24148 25228 24160
rect 25280 24148 25286 24200
rect 26510 24148 26516 24200
rect 26568 24188 26574 24200
rect 27246 24188 27252 24200
rect 26568 24160 27252 24188
rect 26568 24148 26574 24160
rect 27246 24148 27252 24160
rect 27304 24188 27310 24200
rect 28166 24188 28172 24200
rect 27304 24160 28172 24188
rect 27304 24148 27310 24160
rect 28166 24148 28172 24160
rect 28224 24148 28230 24200
rect 33134 24148 33140 24200
rect 33192 24188 33198 24200
rect 33962 24188 33968 24200
rect 33192 24160 33968 24188
rect 33192 24148 33198 24160
rect 33962 24148 33968 24160
rect 34020 24148 34026 24200
rect 36446 24188 36452 24200
rect 36407 24160 36452 24188
rect 36446 24148 36452 24160
rect 36504 24148 36510 24200
rect 24578 24120 24584 24132
rect 24539 24092 24584 24120
rect 24578 24080 24584 24092
rect 24636 24080 24642 24132
rect 30466 24080 30472 24132
rect 30524 24120 30530 24132
rect 30837 24123 30895 24129
rect 30837 24120 30849 24123
rect 30524 24092 30849 24120
rect 30524 24080 30530 24092
rect 30837 24089 30849 24092
rect 30883 24089 30895 24123
rect 30837 24083 30895 24089
rect 28902 24012 28908 24064
rect 28960 24052 28966 24064
rect 29549 24055 29607 24061
rect 29549 24052 29561 24055
rect 28960 24024 29561 24052
rect 28960 24012 28966 24024
rect 29549 24021 29561 24024
rect 29595 24021 29607 24055
rect 29549 24015 29607 24021
rect 35710 24012 35716 24064
rect 35768 24052 35774 24064
rect 35897 24055 35955 24061
rect 35897 24052 35909 24055
rect 35768 24024 35909 24052
rect 35768 24012 35774 24024
rect 35897 24021 35909 24024
rect 35943 24021 35955 24055
rect 35897 24015 35955 24021
rect 1104 23962 38824 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 38824 23962
rect 1104 23888 38824 23910
rect 24673 23851 24731 23857
rect 24673 23817 24685 23851
rect 24719 23848 24731 23851
rect 25038 23848 25044 23860
rect 24719 23820 25044 23848
rect 24719 23817 24731 23820
rect 24673 23811 24731 23817
rect 25038 23808 25044 23820
rect 25096 23808 25102 23860
rect 25222 23808 25228 23860
rect 25280 23848 25286 23860
rect 25317 23851 25375 23857
rect 25317 23848 25329 23851
rect 25280 23820 25329 23848
rect 25280 23808 25286 23820
rect 25317 23817 25329 23820
rect 25363 23817 25375 23851
rect 28074 23848 28080 23860
rect 28035 23820 28080 23848
rect 25317 23811 25375 23817
rect 28074 23808 28080 23820
rect 28132 23808 28138 23860
rect 28166 23808 28172 23860
rect 28224 23848 28230 23860
rect 28629 23851 28687 23857
rect 28629 23848 28641 23851
rect 28224 23820 28641 23848
rect 28224 23808 28230 23820
rect 28629 23817 28641 23820
rect 28675 23817 28687 23851
rect 28629 23811 28687 23817
rect 30561 23851 30619 23857
rect 30561 23817 30573 23851
rect 30607 23848 30619 23851
rect 30650 23848 30656 23860
rect 30607 23820 30656 23848
rect 30607 23817 30619 23820
rect 30561 23811 30619 23817
rect 24946 23780 24952 23792
rect 24907 23752 24952 23780
rect 24946 23740 24952 23752
rect 25004 23740 25010 23792
rect 28644 23780 28672 23811
rect 30650 23808 30656 23820
rect 30708 23808 30714 23860
rect 33962 23808 33968 23860
rect 34020 23848 34026 23860
rect 34241 23851 34299 23857
rect 34241 23848 34253 23851
rect 34020 23820 34253 23848
rect 34020 23808 34026 23820
rect 34241 23817 34253 23820
rect 34287 23848 34299 23851
rect 35253 23851 35311 23857
rect 35253 23848 35265 23851
rect 34287 23820 35265 23848
rect 34287 23817 34299 23820
rect 34241 23811 34299 23817
rect 34992 23792 35020 23820
rect 35253 23817 35265 23820
rect 35299 23817 35311 23851
rect 36814 23848 36820 23860
rect 36775 23820 36820 23848
rect 35253 23811 35311 23817
rect 30837 23783 30895 23789
rect 30837 23780 30849 23783
rect 28644 23752 30849 23780
rect 30837 23749 30849 23752
rect 30883 23780 30895 23783
rect 30883 23752 31064 23780
rect 30883 23749 30895 23752
rect 30837 23743 30895 23749
rect 29914 23712 29920 23724
rect 29875 23684 29920 23712
rect 29914 23672 29920 23684
rect 29972 23672 29978 23724
rect 31036 23721 31064 23752
rect 34974 23740 34980 23792
rect 35032 23740 35038 23792
rect 31021 23715 31079 23721
rect 31021 23681 31033 23715
rect 31067 23681 31079 23715
rect 31021 23675 31079 23681
rect 33781 23715 33839 23721
rect 33781 23681 33793 23715
rect 33827 23712 33839 23715
rect 34606 23712 34612 23724
rect 33827 23684 34612 23712
rect 33827 23681 33839 23684
rect 33781 23675 33839 23681
rect 29089 23647 29147 23653
rect 29089 23613 29101 23647
rect 29135 23644 29147 23647
rect 29270 23644 29276 23656
rect 29135 23616 29276 23644
rect 29135 23613 29147 23616
rect 29089 23607 29147 23613
rect 29270 23604 29276 23616
rect 29328 23644 29334 23656
rect 29641 23647 29699 23653
rect 29641 23644 29653 23647
rect 29328 23616 29653 23644
rect 29328 23604 29334 23616
rect 29641 23613 29653 23616
rect 29687 23644 29699 23647
rect 30006 23644 30012 23656
rect 29687 23616 30012 23644
rect 29687 23613 29699 23616
rect 29641 23607 29699 23613
rect 30006 23604 30012 23616
rect 30064 23604 30070 23656
rect 29730 23576 29736 23588
rect 29691 23548 29736 23576
rect 29730 23536 29736 23548
rect 29788 23536 29794 23588
rect 31036 23576 31064 23675
rect 34606 23672 34612 23684
rect 34664 23672 34670 23724
rect 35268 23712 35296 23811
rect 36814 23808 36820 23820
rect 36872 23808 36878 23860
rect 35437 23715 35495 23721
rect 35437 23712 35449 23715
rect 35268 23684 35449 23712
rect 35437 23681 35449 23684
rect 35483 23681 35495 23715
rect 35437 23675 35495 23681
rect 31294 23653 31300 23656
rect 31288 23644 31300 23653
rect 31255 23616 31300 23644
rect 31288 23607 31300 23616
rect 31294 23604 31300 23607
rect 31352 23604 31358 23656
rect 35710 23653 35716 23656
rect 35704 23644 35716 23653
rect 35671 23616 35716 23644
rect 35704 23607 35716 23616
rect 35710 23604 35716 23607
rect 35768 23604 35774 23656
rect 33134 23576 33140 23588
rect 31036 23548 33140 23576
rect 33134 23536 33140 23548
rect 33192 23536 33198 23588
rect 33870 23536 33876 23588
rect 33928 23576 33934 23588
rect 34609 23579 34667 23585
rect 34609 23576 34621 23579
rect 33928 23548 34621 23576
rect 33928 23536 33934 23548
rect 34609 23545 34621 23548
rect 34655 23545 34667 23579
rect 34609 23539 34667 23545
rect 28166 23508 28172 23520
rect 28127 23480 28172 23508
rect 28166 23468 28172 23480
rect 28224 23468 28230 23520
rect 29086 23468 29092 23520
rect 29144 23508 29150 23520
rect 29273 23511 29331 23517
rect 29273 23508 29285 23511
rect 29144 23480 29285 23508
rect 29144 23468 29150 23480
rect 29273 23477 29285 23480
rect 29319 23477 29331 23511
rect 29273 23471 29331 23477
rect 31938 23468 31944 23520
rect 31996 23508 32002 23520
rect 32401 23511 32459 23517
rect 32401 23508 32413 23511
rect 31996 23480 32413 23508
rect 31996 23468 32002 23480
rect 32401 23477 32413 23480
rect 32447 23477 32459 23511
rect 32401 23471 32459 23477
rect 1104 23418 38824 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 38824 23418
rect 1104 23344 38824 23366
rect 28166 23264 28172 23316
rect 28224 23304 28230 23316
rect 28534 23304 28540 23316
rect 28224 23276 28540 23304
rect 28224 23264 28230 23276
rect 28534 23264 28540 23276
rect 28592 23304 28598 23316
rect 28905 23307 28963 23313
rect 28905 23304 28917 23307
rect 28592 23276 28917 23304
rect 28592 23264 28598 23276
rect 28905 23273 28917 23276
rect 28951 23273 28963 23307
rect 28905 23267 28963 23273
rect 28997 23307 29055 23313
rect 28997 23273 29009 23307
rect 29043 23304 29055 23307
rect 29086 23304 29092 23316
rect 29043 23276 29092 23304
rect 29043 23273 29055 23276
rect 28997 23267 29055 23273
rect 29086 23264 29092 23276
rect 29144 23264 29150 23316
rect 29641 23307 29699 23313
rect 29641 23273 29653 23307
rect 29687 23304 29699 23307
rect 29730 23304 29736 23316
rect 29687 23276 29736 23304
rect 29687 23273 29699 23276
rect 29641 23267 29699 23273
rect 29730 23264 29736 23276
rect 29788 23264 29794 23316
rect 29914 23304 29920 23316
rect 29875 23276 29920 23304
rect 29914 23264 29920 23276
rect 29972 23264 29978 23316
rect 30193 23307 30251 23313
rect 30193 23273 30205 23307
rect 30239 23304 30251 23307
rect 30282 23304 30288 23316
rect 30239 23276 30288 23304
rect 30239 23273 30251 23276
rect 30193 23267 30251 23273
rect 30282 23264 30288 23276
rect 30340 23264 30346 23316
rect 31113 23307 31171 23313
rect 31113 23273 31125 23307
rect 31159 23304 31171 23307
rect 31294 23304 31300 23316
rect 31159 23276 31300 23304
rect 31159 23273 31171 23276
rect 31113 23267 31171 23273
rect 31294 23264 31300 23276
rect 31352 23264 31358 23316
rect 33321 23307 33379 23313
rect 33321 23273 33333 23307
rect 33367 23304 33379 23307
rect 34422 23304 34428 23316
rect 33367 23276 34428 23304
rect 33367 23273 33379 23276
rect 33321 23267 33379 23273
rect 34422 23264 34428 23276
rect 34480 23264 34486 23316
rect 34517 23307 34575 23313
rect 34517 23273 34529 23307
rect 34563 23304 34575 23307
rect 35710 23304 35716 23316
rect 34563 23276 35716 23304
rect 34563 23273 34575 23276
rect 34517 23267 34575 23273
rect 35710 23264 35716 23276
rect 35768 23304 35774 23316
rect 36357 23307 36415 23313
rect 36357 23304 36369 23307
rect 35768 23276 36369 23304
rect 35768 23264 35774 23276
rect 36357 23273 36369 23276
rect 36403 23273 36415 23307
rect 36357 23267 36415 23273
rect 33134 23196 33140 23248
rect 33192 23236 33198 23248
rect 33686 23236 33692 23248
rect 33192 23208 33692 23236
rect 33192 23196 33198 23208
rect 33686 23196 33692 23208
rect 33744 23196 33750 23248
rect 34885 23239 34943 23245
rect 34885 23205 34897 23239
rect 34931 23236 34943 23239
rect 35244 23239 35302 23245
rect 35244 23236 35256 23239
rect 34931 23208 35256 23236
rect 34931 23205 34943 23208
rect 34885 23199 34943 23205
rect 35244 23205 35256 23208
rect 35290 23236 35302 23239
rect 35434 23236 35440 23248
rect 35290 23208 35440 23236
rect 35290 23205 35302 23208
rect 35244 23199 35302 23205
rect 35434 23196 35440 23208
rect 35492 23196 35498 23248
rect 34514 23128 34520 23180
rect 34572 23168 34578 23180
rect 34974 23168 34980 23180
rect 34572 23140 34980 23168
rect 34572 23128 34578 23140
rect 34974 23128 34980 23140
rect 35032 23128 35038 23180
rect 28074 23060 28080 23112
rect 28132 23100 28138 23112
rect 28902 23100 28908 23112
rect 28132 23072 28908 23100
rect 28132 23060 28138 23072
rect 28902 23060 28908 23072
rect 28960 23100 28966 23112
rect 29089 23103 29147 23109
rect 29089 23100 29101 23103
rect 28960 23072 29101 23100
rect 28960 23060 28966 23072
rect 29089 23069 29101 23072
rect 29135 23069 29147 23103
rect 33778 23100 33784 23112
rect 33739 23072 33784 23100
rect 29089 23063 29147 23069
rect 33778 23060 33784 23072
rect 33836 23060 33842 23112
rect 33870 23060 33876 23112
rect 33928 23100 33934 23112
rect 33928 23072 33973 23100
rect 33928 23060 33934 23072
rect 28537 23035 28595 23041
rect 28537 23001 28549 23035
rect 28583 23032 28595 23035
rect 29730 23032 29736 23044
rect 28583 23004 29736 23032
rect 28583 23001 28595 23004
rect 28537 22995 28595 23001
rect 29730 22992 29736 23004
rect 29788 22992 29794 23044
rect 24026 22964 24032 22976
rect 23987 22936 24032 22964
rect 24026 22924 24032 22936
rect 24084 22924 24090 22976
rect 26786 22964 26792 22976
rect 26747 22936 26792 22964
rect 26786 22924 26792 22936
rect 26844 22924 26850 22976
rect 34698 22924 34704 22976
rect 34756 22964 34762 22976
rect 35342 22964 35348 22976
rect 34756 22936 35348 22964
rect 34756 22924 34762 22936
rect 35342 22924 35348 22936
rect 35400 22924 35406 22976
rect 36906 22964 36912 22976
rect 36867 22936 36912 22964
rect 36906 22924 36912 22936
rect 36964 22924 36970 22976
rect 1104 22874 38824 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 38824 22874
rect 1104 22800 38824 22822
rect 28074 22720 28080 22772
rect 28132 22760 28138 22772
rect 28169 22763 28227 22769
rect 28169 22760 28181 22763
rect 28132 22732 28181 22760
rect 28132 22720 28138 22732
rect 28169 22729 28181 22732
rect 28215 22729 28227 22763
rect 28534 22760 28540 22772
rect 28495 22732 28540 22760
rect 28169 22723 28227 22729
rect 28534 22720 28540 22732
rect 28592 22720 28598 22772
rect 33045 22763 33103 22769
rect 33045 22729 33057 22763
rect 33091 22760 33103 22763
rect 33870 22760 33876 22772
rect 33091 22732 33876 22760
rect 33091 22729 33103 22732
rect 33045 22723 33103 22729
rect 33870 22720 33876 22732
rect 33928 22720 33934 22772
rect 34514 22720 34520 22772
rect 34572 22760 34578 22772
rect 34609 22763 34667 22769
rect 34609 22760 34621 22763
rect 34572 22732 34621 22760
rect 34572 22720 34578 22732
rect 34609 22729 34621 22732
rect 34655 22729 34667 22763
rect 36446 22760 36452 22772
rect 36407 22732 36452 22760
rect 34609 22723 34667 22729
rect 36446 22720 36452 22732
rect 36504 22720 36510 22772
rect 36538 22720 36544 22772
rect 36596 22760 36602 22772
rect 36596 22732 36641 22760
rect 36596 22720 36602 22732
rect 36814 22720 36820 22772
rect 36872 22760 36878 22772
rect 36872 22732 37136 22760
rect 36872 22720 36878 22732
rect 25961 22695 26019 22701
rect 25961 22661 25973 22695
rect 26007 22692 26019 22695
rect 26694 22692 26700 22704
rect 26007 22664 26700 22692
rect 26007 22661 26019 22664
rect 25961 22655 26019 22661
rect 26694 22652 26700 22664
rect 26752 22692 26758 22704
rect 33686 22692 33692 22704
rect 26752 22664 27016 22692
rect 33647 22664 33692 22692
rect 26752 22652 26758 22664
rect 26326 22584 26332 22636
rect 26384 22624 26390 22636
rect 26786 22624 26792 22636
rect 26384 22596 26792 22624
rect 26384 22584 26390 22596
rect 26786 22584 26792 22596
rect 26844 22624 26850 22636
rect 26988 22633 27016 22664
rect 33686 22652 33692 22664
rect 33744 22652 33750 22704
rect 34977 22695 35035 22701
rect 34977 22661 34989 22695
rect 35023 22692 35035 22695
rect 36906 22692 36912 22704
rect 35023 22664 36912 22692
rect 35023 22661 35035 22664
rect 34977 22655 35035 22661
rect 36906 22652 36912 22664
rect 36964 22692 36970 22704
rect 36964 22664 37044 22692
rect 36964 22652 36970 22664
rect 26881 22627 26939 22633
rect 26881 22624 26893 22627
rect 26844 22596 26893 22624
rect 26844 22584 26850 22596
rect 26881 22593 26893 22596
rect 26927 22593 26939 22627
rect 26881 22587 26939 22593
rect 26973 22627 27031 22633
rect 26973 22593 26985 22627
rect 27019 22593 27031 22627
rect 26973 22587 27031 22593
rect 29730 22584 29736 22636
rect 29788 22624 29794 22636
rect 35621 22627 35679 22633
rect 29788 22596 29833 22624
rect 29788 22584 29794 22596
rect 35621 22593 35633 22627
rect 35667 22624 35679 22627
rect 35710 22624 35716 22636
rect 35667 22596 35716 22624
rect 35667 22593 35679 22596
rect 35621 22587 35679 22593
rect 35710 22584 35716 22596
rect 35768 22584 35774 22636
rect 37016 22633 37044 22664
rect 37108 22633 37136 22732
rect 37001 22627 37059 22633
rect 37001 22593 37013 22627
rect 37047 22593 37059 22627
rect 37001 22587 37059 22593
rect 37093 22627 37151 22633
rect 37093 22593 37105 22627
rect 37139 22593 37151 22627
rect 37093 22587 37151 22593
rect 23934 22556 23940 22568
rect 23895 22528 23940 22556
rect 23934 22516 23940 22528
rect 23992 22516 23998 22568
rect 24026 22516 24032 22568
rect 24084 22556 24090 22568
rect 24193 22559 24251 22565
rect 24193 22556 24205 22559
rect 24084 22528 24205 22556
rect 24084 22516 24090 22528
rect 24193 22525 24205 22528
rect 24239 22525 24251 22559
rect 24193 22519 24251 22525
rect 29178 22516 29184 22568
rect 29236 22556 29242 22568
rect 29273 22559 29331 22565
rect 29273 22556 29285 22559
rect 29236 22528 29285 22556
rect 29236 22516 29242 22528
rect 29273 22525 29285 22528
rect 29319 22525 29331 22559
rect 29273 22519 29331 22525
rect 30006 22516 30012 22568
rect 30064 22556 30070 22568
rect 30064 22528 30109 22556
rect 30064 22516 30070 22528
rect 36446 22516 36452 22568
rect 36504 22556 36510 22568
rect 36909 22559 36967 22565
rect 36909 22556 36921 22559
rect 36504 22528 36921 22556
rect 36504 22516 36510 22528
rect 36909 22525 36921 22528
rect 36955 22525 36967 22559
rect 36909 22519 36967 22525
rect 26789 22491 26847 22497
rect 26789 22488 26801 22491
rect 26252 22460 26801 22488
rect 26252 22432 26280 22460
rect 26789 22457 26801 22460
rect 26835 22457 26847 22491
rect 26789 22451 26847 22457
rect 33134 22448 33140 22500
rect 33192 22488 33198 22500
rect 34241 22491 34299 22497
rect 34241 22488 34253 22491
rect 33192 22460 34253 22488
rect 33192 22448 33198 22460
rect 34241 22457 34253 22460
rect 34287 22457 34299 22491
rect 34241 22451 34299 22457
rect 25314 22420 25320 22432
rect 25275 22392 25320 22420
rect 25314 22380 25320 22392
rect 25372 22380 25378 22432
rect 26234 22420 26240 22432
rect 26195 22392 26240 22420
rect 26234 22380 26240 22392
rect 26292 22380 26298 22432
rect 26418 22420 26424 22432
rect 26379 22392 26424 22420
rect 26418 22380 26424 22392
rect 26476 22380 26482 22432
rect 29089 22423 29147 22429
rect 29089 22389 29101 22423
rect 29135 22420 29147 22423
rect 29735 22423 29793 22429
rect 29735 22420 29747 22423
rect 29135 22392 29747 22420
rect 29135 22389 29147 22392
rect 29089 22383 29147 22389
rect 29735 22389 29747 22392
rect 29781 22420 29793 22423
rect 30374 22420 30380 22432
rect 29781 22392 30380 22420
rect 29781 22389 29793 22392
rect 29735 22383 29793 22389
rect 30374 22380 30380 22392
rect 30432 22380 30438 22432
rect 31113 22423 31171 22429
rect 31113 22389 31125 22423
rect 31159 22420 31171 22423
rect 33321 22423 33379 22429
rect 33321 22420 33333 22423
rect 31159 22392 33333 22420
rect 31159 22389 31171 22392
rect 31113 22383 31171 22389
rect 33321 22389 33333 22392
rect 33367 22420 33379 22423
rect 33778 22420 33784 22432
rect 33367 22392 33784 22420
rect 33367 22389 33379 22392
rect 33321 22383 33379 22389
rect 33778 22380 33784 22392
rect 33836 22420 33842 22432
rect 34146 22420 34152 22432
rect 33836 22392 34152 22420
rect 33836 22380 33842 22392
rect 34146 22380 34152 22392
rect 34204 22380 34210 22432
rect 34256 22420 34284 22451
rect 34514 22448 34520 22500
rect 34572 22488 34578 22500
rect 34882 22488 34888 22500
rect 34572 22460 34888 22488
rect 34572 22448 34578 22460
rect 34882 22448 34888 22460
rect 34940 22488 34946 22500
rect 35345 22491 35403 22497
rect 35345 22488 35357 22491
rect 34940 22460 35357 22488
rect 34940 22448 34946 22460
rect 35345 22457 35357 22460
rect 35391 22488 35403 22491
rect 35894 22488 35900 22500
rect 35391 22460 35900 22488
rect 35391 22457 35403 22460
rect 35345 22451 35403 22457
rect 35894 22448 35900 22460
rect 35952 22488 35958 22500
rect 35989 22491 36047 22497
rect 35989 22488 36001 22491
rect 35952 22460 36001 22488
rect 35952 22448 35958 22460
rect 35989 22457 36001 22460
rect 36035 22457 36047 22491
rect 35989 22451 36047 22457
rect 35434 22420 35440 22432
rect 34256 22392 35440 22420
rect 35434 22380 35440 22392
rect 35492 22380 35498 22432
rect 35526 22380 35532 22432
rect 35584 22420 35590 22432
rect 36538 22420 36544 22432
rect 35584 22392 36544 22420
rect 35584 22380 35590 22392
rect 36538 22380 36544 22392
rect 36596 22380 36602 22432
rect 1104 22330 38824 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 38824 22330
rect 1104 22256 38824 22278
rect 28629 22219 28687 22225
rect 28629 22185 28641 22219
rect 28675 22216 28687 22219
rect 28902 22216 28908 22228
rect 28675 22188 28908 22216
rect 28675 22185 28687 22188
rect 28629 22179 28687 22185
rect 28902 22176 28908 22188
rect 28960 22176 28966 22228
rect 29730 22216 29736 22228
rect 29691 22188 29736 22216
rect 29730 22176 29736 22188
rect 29788 22176 29794 22228
rect 31754 22176 31760 22228
rect 31812 22216 31818 22228
rect 32398 22216 32404 22228
rect 31812 22188 32404 22216
rect 31812 22176 31818 22188
rect 32398 22176 32404 22188
rect 32456 22216 32462 22228
rect 32493 22219 32551 22225
rect 32493 22216 32505 22219
rect 32456 22188 32505 22216
rect 32456 22176 32462 22188
rect 32493 22185 32505 22188
rect 32539 22185 32551 22219
rect 34146 22216 34152 22228
rect 34107 22188 34152 22216
rect 32493 22179 32551 22185
rect 34146 22176 34152 22188
rect 34204 22176 34210 22228
rect 35434 22176 35440 22228
rect 35492 22216 35498 22228
rect 36814 22216 36820 22228
rect 35492 22188 35848 22216
rect 36775 22188 36820 22216
rect 35492 22176 35498 22188
rect 21453 22083 21511 22089
rect 21453 22049 21465 22083
rect 21499 22080 21511 22083
rect 21910 22080 21916 22092
rect 21499 22052 21916 22080
rect 21499 22049 21511 22052
rect 21453 22043 21511 22049
rect 21910 22040 21916 22052
rect 21968 22080 21974 22092
rect 22077 22083 22135 22089
rect 22077 22080 22089 22083
rect 21968 22052 22089 22080
rect 21968 22040 21974 22052
rect 22077 22049 22089 22052
rect 22123 22049 22135 22083
rect 23934 22080 23940 22092
rect 23895 22052 23940 22080
rect 22077 22043 22135 22049
rect 23934 22040 23940 22052
rect 23992 22040 23998 22092
rect 24670 22080 24676 22092
rect 24631 22052 24676 22080
rect 24670 22040 24676 22052
rect 24728 22040 24734 22092
rect 26786 22089 26792 22092
rect 25685 22083 25743 22089
rect 25685 22080 25697 22083
rect 24780 22052 25697 22080
rect 21818 22012 21824 22024
rect 21779 21984 21824 22012
rect 21818 21972 21824 21984
rect 21876 21972 21882 22024
rect 23750 21972 23756 22024
rect 23808 22012 23814 22024
rect 24780 22021 24808 22052
rect 25685 22049 25697 22052
rect 25731 22049 25743 22083
rect 26780 22080 26792 22089
rect 26747 22052 26792 22080
rect 25685 22043 25743 22049
rect 26780 22043 26792 22052
rect 26786 22040 26792 22043
rect 26844 22040 26850 22092
rect 29270 22080 29276 22092
rect 29231 22052 29276 22080
rect 29270 22040 29276 22052
rect 29328 22040 29334 22092
rect 30009 22083 30067 22089
rect 30009 22049 30021 22083
rect 30055 22080 30067 22083
rect 30190 22080 30196 22092
rect 30055 22052 30196 22080
rect 30055 22049 30067 22052
rect 30009 22043 30067 22049
rect 30190 22040 30196 22052
rect 30248 22040 30254 22092
rect 34164 22080 34192 22176
rect 35820 22148 35848 22188
rect 36814 22176 36820 22188
rect 36872 22176 36878 22228
rect 35820 22120 35940 22148
rect 35069 22083 35127 22089
rect 35069 22080 35081 22083
rect 34164 22052 35081 22080
rect 35069 22049 35081 22052
rect 35115 22049 35127 22083
rect 35912 22080 35940 22120
rect 35912 22052 36216 22080
rect 35069 22043 35127 22049
rect 24765 22015 24823 22021
rect 24765 22012 24777 22015
rect 23808 21984 24777 22012
rect 23808 21972 23814 21984
rect 24765 21981 24777 21984
rect 24811 21981 24823 22015
rect 24765 21975 24823 21981
rect 24857 22015 24915 22021
rect 24857 21981 24869 22015
rect 24903 21981 24915 22015
rect 26510 22012 26516 22024
rect 26471 21984 26516 22012
rect 24857 21975 24915 21981
rect 24026 21904 24032 21956
rect 24084 21944 24090 21956
rect 24872 21944 24900 21975
rect 26510 21972 26516 21984
rect 26568 21972 26574 22024
rect 32582 22012 32588 22024
rect 32543 21984 32588 22012
rect 32582 21972 32588 21984
rect 32640 21972 32646 22024
rect 32674 21972 32680 22024
rect 32732 22012 32738 22024
rect 34330 22012 34336 22024
rect 32732 21984 32777 22012
rect 34291 21984 34336 22012
rect 32732 21972 32738 21984
rect 34330 21972 34336 21984
rect 34388 21972 34394 22024
rect 34514 21972 34520 22024
rect 34572 22012 34578 22024
rect 34656 22015 34714 22021
rect 34656 22012 34668 22015
rect 34572 21984 34668 22012
rect 34572 21972 34578 21984
rect 34656 21981 34668 21984
rect 34702 21981 34714 22015
rect 34656 21975 34714 21981
rect 34793 22015 34851 22021
rect 34793 21981 34805 22015
rect 34839 22012 34851 22015
rect 34882 22012 34888 22024
rect 34839 21984 34888 22012
rect 34839 21981 34851 21984
rect 34793 21975 34851 21981
rect 34882 21972 34888 21984
rect 34940 21972 34946 22024
rect 36188 22021 36216 22052
rect 36173 22015 36231 22021
rect 36173 21981 36185 22015
rect 36219 21981 36231 22015
rect 36173 21975 36231 21981
rect 28997 21947 29055 21953
rect 28997 21944 29009 21947
rect 24084 21916 24900 21944
rect 27540 21916 29009 21944
rect 24084 21904 24090 21916
rect 24780 21888 24808 21916
rect 23198 21876 23204 21888
rect 23159 21848 23204 21876
rect 23198 21836 23204 21848
rect 23256 21836 23262 21888
rect 24302 21876 24308 21888
rect 24263 21848 24308 21876
rect 24302 21836 24308 21848
rect 24360 21836 24366 21888
rect 24762 21836 24768 21888
rect 24820 21836 24826 21888
rect 25409 21879 25467 21885
rect 25409 21845 25421 21879
rect 25455 21876 25467 21879
rect 25590 21876 25596 21888
rect 25455 21848 25596 21876
rect 25455 21845 25467 21848
rect 25409 21839 25467 21845
rect 25590 21836 25596 21848
rect 25648 21836 25654 21888
rect 26145 21879 26203 21885
rect 26145 21845 26157 21879
rect 26191 21876 26203 21879
rect 26234 21876 26240 21888
rect 26191 21848 26240 21876
rect 26191 21845 26203 21848
rect 26145 21839 26203 21845
rect 26234 21836 26240 21848
rect 26292 21876 26298 21888
rect 27540 21876 27568 21916
rect 28997 21913 29009 21916
rect 29043 21944 29055 21947
rect 29178 21944 29184 21956
rect 29043 21916 29184 21944
rect 29043 21913 29055 21916
rect 28997 21907 29055 21913
rect 29178 21904 29184 21916
rect 29236 21944 29242 21956
rect 31938 21944 31944 21956
rect 29236 21916 30788 21944
rect 31851 21916 31944 21944
rect 29236 21904 29242 21916
rect 30760 21888 30788 21916
rect 31938 21904 31944 21916
rect 31996 21944 32002 21956
rect 32692 21944 32720 21972
rect 31996 21916 32720 21944
rect 31996 21904 32002 21916
rect 27890 21876 27896 21888
rect 26292 21848 27568 21876
rect 27851 21848 27896 21876
rect 26292 21836 26298 21848
rect 27890 21836 27896 21848
rect 27948 21836 27954 21888
rect 30190 21876 30196 21888
rect 30151 21848 30196 21876
rect 30190 21836 30196 21848
rect 30248 21836 30254 21888
rect 30650 21876 30656 21888
rect 30611 21848 30656 21876
rect 30650 21836 30656 21848
rect 30708 21836 30714 21888
rect 30742 21836 30748 21888
rect 30800 21876 30806 21888
rect 31021 21879 31079 21885
rect 31021 21876 31033 21879
rect 30800 21848 31033 21876
rect 30800 21836 30806 21848
rect 31021 21845 31033 21848
rect 31067 21876 31079 21879
rect 31662 21876 31668 21888
rect 31067 21848 31668 21876
rect 31067 21845 31079 21848
rect 31021 21839 31079 21845
rect 31662 21836 31668 21848
rect 31720 21836 31726 21888
rect 32122 21876 32128 21888
rect 32083 21848 32128 21876
rect 32122 21836 32128 21848
rect 32180 21836 32186 21888
rect 1104 21786 38824 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 38824 21786
rect 1104 21712 38824 21734
rect 21818 21632 21824 21684
rect 21876 21672 21882 21684
rect 22373 21675 22431 21681
rect 22373 21672 22385 21675
rect 21876 21644 22385 21672
rect 21876 21632 21882 21644
rect 22373 21641 22385 21644
rect 22419 21641 22431 21675
rect 22373 21635 22431 21641
rect 23477 21675 23535 21681
rect 23477 21641 23489 21675
rect 23523 21672 23535 21675
rect 24026 21672 24032 21684
rect 23523 21644 24032 21672
rect 23523 21641 23535 21644
rect 23477 21635 23535 21641
rect 24026 21632 24032 21644
rect 24084 21632 24090 21684
rect 24397 21675 24455 21681
rect 24397 21641 24409 21675
rect 24443 21672 24455 21675
rect 24670 21672 24676 21684
rect 24443 21644 24676 21672
rect 24443 21641 24455 21644
rect 24397 21635 24455 21641
rect 21910 21536 21916 21548
rect 21871 21508 21916 21536
rect 21910 21496 21916 21508
rect 21968 21536 21974 21548
rect 22741 21539 22799 21545
rect 22741 21536 22753 21539
rect 21968 21508 22753 21536
rect 21968 21496 21974 21508
rect 22741 21505 22753 21508
rect 22787 21505 22799 21539
rect 22741 21499 22799 21505
rect 23661 21539 23719 21545
rect 23661 21505 23673 21539
rect 23707 21536 23719 21539
rect 24412 21536 24440 21635
rect 24670 21632 24676 21644
rect 24728 21632 24734 21684
rect 26050 21632 26056 21684
rect 26108 21672 26114 21684
rect 26694 21672 26700 21684
rect 26108 21644 26700 21672
rect 26108 21632 26114 21644
rect 26694 21632 26700 21644
rect 26752 21632 26758 21684
rect 30098 21672 30104 21684
rect 30059 21644 30104 21672
rect 30098 21632 30104 21644
rect 30156 21632 30162 21684
rect 30374 21672 30380 21684
rect 30335 21644 30380 21672
rect 30374 21632 30380 21644
rect 30432 21632 30438 21684
rect 35894 21672 35900 21684
rect 35855 21644 35900 21672
rect 35894 21632 35900 21644
rect 35952 21632 35958 21684
rect 23707 21508 24440 21536
rect 23707 21505 23719 21508
rect 23661 21499 23719 21505
rect 25038 21496 25044 21548
rect 25096 21536 25102 21548
rect 25317 21539 25375 21545
rect 25317 21536 25329 21539
rect 25096 21508 25329 21536
rect 25096 21496 25102 21508
rect 25317 21505 25329 21508
rect 25363 21505 25375 21539
rect 26234 21536 26240 21548
rect 25317 21499 25375 21505
rect 25516 21508 26240 21536
rect 20898 21468 20904 21480
rect 20811 21440 20904 21468
rect 20898 21428 20904 21440
rect 20956 21468 20962 21480
rect 21821 21471 21879 21477
rect 21821 21468 21833 21471
rect 20956 21440 21833 21468
rect 20956 21428 20962 21440
rect 21821 21437 21833 21440
rect 21867 21437 21879 21471
rect 21821 21431 21879 21437
rect 24857 21471 24915 21477
rect 24857 21437 24869 21471
rect 24903 21468 24915 21471
rect 25516 21468 25544 21508
rect 26234 21496 26240 21508
rect 26292 21496 26298 21548
rect 30561 21539 30619 21545
rect 30561 21505 30573 21539
rect 30607 21536 30619 21539
rect 30742 21536 30748 21548
rect 30607 21508 30748 21536
rect 30607 21505 30619 21508
rect 30561 21499 30619 21505
rect 30742 21496 30748 21508
rect 30800 21496 30806 21548
rect 31018 21536 31024 21548
rect 30979 21508 31024 21536
rect 31018 21496 31024 21508
rect 31076 21496 31082 21548
rect 35342 21536 35348 21548
rect 35303 21508 35348 21536
rect 35342 21496 35348 21508
rect 35400 21496 35406 21548
rect 35434 21496 35440 21548
rect 35492 21536 35498 21548
rect 35529 21539 35587 21545
rect 35529 21536 35541 21539
rect 35492 21508 35541 21536
rect 35492 21496 35498 21508
rect 35529 21505 35541 21508
rect 35575 21536 35587 21539
rect 36265 21539 36323 21545
rect 36265 21536 36277 21539
rect 35575 21508 36277 21536
rect 35575 21505 35587 21508
rect 35529 21499 35587 21505
rect 36265 21505 36277 21508
rect 36311 21505 36323 21539
rect 36265 21499 36323 21505
rect 24903 21440 25544 21468
rect 24903 21437 24915 21440
rect 24857 21431 24915 21437
rect 25590 21428 25596 21480
rect 25648 21468 25654 21480
rect 25648 21440 25693 21468
rect 25648 21428 25654 21440
rect 26786 21428 26792 21480
rect 26844 21468 26850 21480
rect 27617 21471 27675 21477
rect 27617 21468 27629 21471
rect 26844 21440 27629 21468
rect 26844 21428 26850 21440
rect 27617 21437 27629 21440
rect 27663 21437 27675 21471
rect 27617 21431 27675 21437
rect 30650 21428 30656 21480
rect 30708 21468 30714 21480
rect 31294 21468 31300 21480
rect 30708 21440 31300 21468
rect 30708 21428 30714 21440
rect 31294 21428 31300 21440
rect 31352 21428 31358 21480
rect 34333 21471 34391 21477
rect 34333 21468 34345 21471
rect 31956 21440 34345 21468
rect 20349 21403 20407 21409
rect 20349 21369 20361 21403
rect 20395 21400 20407 21403
rect 21177 21403 21235 21409
rect 21177 21400 21189 21403
rect 20395 21372 21189 21400
rect 20395 21369 20407 21372
rect 20349 21363 20407 21369
rect 21177 21369 21189 21372
rect 21223 21400 21235 21403
rect 21729 21403 21787 21409
rect 21729 21400 21741 21403
rect 21223 21372 21741 21400
rect 21223 21369 21235 21372
rect 21177 21363 21235 21369
rect 21729 21369 21741 21372
rect 21775 21369 21787 21403
rect 21729 21363 21787 21369
rect 26510 21360 26516 21412
rect 26568 21400 26574 21412
rect 27246 21400 27252 21412
rect 26568 21372 27252 21400
rect 26568 21360 26574 21372
rect 27246 21360 27252 21372
rect 27304 21360 27310 21412
rect 21358 21332 21364 21344
rect 21319 21304 21364 21332
rect 21358 21292 21364 21304
rect 21416 21292 21422 21344
rect 24765 21335 24823 21341
rect 24765 21301 24777 21335
rect 24811 21332 24823 21335
rect 25319 21335 25377 21341
rect 25319 21332 25331 21335
rect 24811 21304 25331 21332
rect 24811 21301 24823 21304
rect 24765 21295 24823 21301
rect 25319 21301 25331 21304
rect 25365 21332 25377 21335
rect 26970 21332 26976 21344
rect 25365 21304 26976 21332
rect 25365 21301 25377 21304
rect 25319 21295 25377 21301
rect 26970 21292 26976 21304
rect 27028 21292 27034 21344
rect 27430 21292 27436 21344
rect 27488 21332 27494 21344
rect 27801 21335 27859 21341
rect 27801 21332 27813 21335
rect 27488 21304 27813 21332
rect 27488 21292 27494 21304
rect 27801 21301 27813 21304
rect 27847 21301 27859 21335
rect 27801 21295 27859 21301
rect 30374 21292 30380 21344
rect 30432 21332 30438 21344
rect 31023 21335 31081 21341
rect 31023 21332 31035 21335
rect 30432 21304 31035 21332
rect 30432 21292 30438 21304
rect 31023 21301 31035 21304
rect 31069 21332 31081 21335
rect 31570 21332 31576 21344
rect 31069 21304 31576 21332
rect 31069 21301 31081 21304
rect 31023 21295 31081 21301
rect 31570 21292 31576 21304
rect 31628 21332 31634 21344
rect 31956 21332 31984 21440
rect 34333 21437 34345 21440
rect 34379 21468 34391 21471
rect 34514 21468 34520 21480
rect 34379 21440 34520 21468
rect 34379 21437 34391 21440
rect 34333 21431 34391 21437
rect 34514 21428 34520 21440
rect 34572 21428 34578 21480
rect 35360 21468 35388 21496
rect 36633 21471 36691 21477
rect 36633 21468 36645 21471
rect 35360 21440 36645 21468
rect 36633 21437 36645 21440
rect 36679 21437 36691 21471
rect 36633 21431 36691 21437
rect 33505 21403 33563 21409
rect 33505 21369 33517 21403
rect 33551 21400 33563 21403
rect 34057 21403 34115 21409
rect 34057 21400 34069 21403
rect 33551 21372 34069 21400
rect 33551 21369 33563 21372
rect 33505 21363 33563 21369
rect 34057 21369 34069 21372
rect 34103 21400 34115 21403
rect 35253 21403 35311 21409
rect 35253 21400 35265 21403
rect 34103 21372 35265 21400
rect 34103 21369 34115 21372
rect 34057 21363 34115 21369
rect 35253 21369 35265 21372
rect 35299 21369 35311 21403
rect 35253 21363 35311 21369
rect 31628 21304 31984 21332
rect 32401 21335 32459 21341
rect 31628 21292 31634 21304
rect 32401 21301 32413 21335
rect 32447 21332 32459 21335
rect 32582 21332 32588 21344
rect 32447 21304 32588 21332
rect 32447 21301 32459 21304
rect 32401 21295 32459 21301
rect 32582 21292 32588 21304
rect 32640 21332 32646 21344
rect 32953 21335 33011 21341
rect 32953 21332 32965 21335
rect 32640 21304 32965 21332
rect 32640 21292 32646 21304
rect 32953 21301 32965 21304
rect 32999 21301 33011 21335
rect 33318 21332 33324 21344
rect 33279 21304 33324 21332
rect 32953 21295 33011 21301
rect 33318 21292 33324 21304
rect 33376 21292 33382 21344
rect 34790 21292 34796 21344
rect 34848 21332 34854 21344
rect 34885 21335 34943 21341
rect 34885 21332 34897 21335
rect 34848 21304 34897 21332
rect 34848 21292 34854 21304
rect 34885 21301 34897 21304
rect 34931 21301 34943 21335
rect 34885 21295 34943 21301
rect 1104 21242 38824 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 38824 21242
rect 1104 21168 38824 21190
rect 21910 21088 21916 21140
rect 21968 21128 21974 21140
rect 22281 21131 22339 21137
rect 22281 21128 22293 21131
rect 21968 21100 22293 21128
rect 21968 21088 21974 21100
rect 22281 21097 22293 21100
rect 22327 21097 22339 21131
rect 24762 21128 24768 21140
rect 24723 21100 24768 21128
rect 22281 21091 22339 21097
rect 24762 21088 24768 21100
rect 24820 21088 24826 21140
rect 25314 21088 25320 21140
rect 25372 21128 25378 21140
rect 25685 21131 25743 21137
rect 25685 21128 25697 21131
rect 25372 21100 25697 21128
rect 25372 21088 25378 21100
rect 25685 21097 25697 21100
rect 25731 21097 25743 21131
rect 26234 21128 26240 21140
rect 26195 21100 26240 21128
rect 25685 21091 25743 21097
rect 26234 21088 26240 21100
rect 26292 21088 26298 21140
rect 28442 21128 28448 21140
rect 28403 21100 28448 21128
rect 28442 21088 28448 21100
rect 28500 21088 28506 21140
rect 29917 21131 29975 21137
rect 29917 21097 29929 21131
rect 29963 21128 29975 21131
rect 30929 21131 30987 21137
rect 30929 21128 30941 21131
rect 29963 21100 30941 21128
rect 29963 21097 29975 21100
rect 29917 21091 29975 21097
rect 30929 21097 30941 21100
rect 30975 21128 30987 21131
rect 31018 21128 31024 21140
rect 30975 21100 31024 21128
rect 30975 21097 30987 21100
rect 30929 21091 30987 21097
rect 31018 21088 31024 21100
rect 31076 21088 31082 21140
rect 31294 21088 31300 21140
rect 31352 21128 31358 21140
rect 32493 21131 32551 21137
rect 32493 21128 32505 21131
rect 31352 21100 32505 21128
rect 31352 21088 31358 21100
rect 32493 21097 32505 21100
rect 32539 21128 32551 21131
rect 33042 21128 33048 21140
rect 32539 21100 33048 21128
rect 32539 21097 32551 21100
rect 32493 21091 32551 21097
rect 33042 21088 33048 21100
rect 33100 21088 33106 21140
rect 33873 21131 33931 21137
rect 33873 21097 33885 21131
rect 33919 21128 33931 21131
rect 34330 21128 34336 21140
rect 33919 21100 34336 21128
rect 33919 21097 33931 21100
rect 33873 21091 33931 21097
rect 34330 21088 34336 21100
rect 34388 21088 34394 21140
rect 21818 21060 21824 21072
rect 20916 21032 21824 21060
rect 20916 21001 20944 21032
rect 21818 21020 21824 21032
rect 21876 21020 21882 21072
rect 23198 21020 23204 21072
rect 23256 21060 23262 21072
rect 23474 21060 23480 21072
rect 23256 21032 23480 21060
rect 23256 21020 23262 21032
rect 23474 21020 23480 21032
rect 23532 21060 23538 21072
rect 23630 21063 23688 21069
rect 23630 21060 23642 21063
rect 23532 21032 23642 21060
rect 23532 21020 23538 21032
rect 23630 21029 23642 21032
rect 23676 21029 23688 21063
rect 23630 21023 23688 21029
rect 20901 20995 20959 21001
rect 20901 20961 20913 20995
rect 20947 20961 20959 20995
rect 20901 20955 20959 20961
rect 21168 20995 21226 21001
rect 21168 20961 21180 20995
rect 21214 20992 21226 20995
rect 21542 20992 21548 21004
rect 21214 20964 21548 20992
rect 21214 20961 21226 20964
rect 21168 20955 21226 20961
rect 21542 20952 21548 20964
rect 21600 20952 21606 21004
rect 23385 20995 23443 21001
rect 23385 20961 23397 20995
rect 23431 20992 23443 20995
rect 23934 20992 23940 21004
rect 23431 20964 23940 20992
rect 23431 20961 23443 20964
rect 23385 20955 23443 20961
rect 23934 20952 23940 20964
rect 23992 20952 23998 21004
rect 26252 20992 26280 21088
rect 31941 21063 31999 21069
rect 31941 21029 31953 21063
rect 31987 21060 31999 21063
rect 32582 21060 32588 21072
rect 31987 21032 32588 21060
rect 31987 21029 31999 21032
rect 31941 21023 31999 21029
rect 32582 21020 32588 21032
rect 32640 21020 32646 21072
rect 34232 21063 34290 21069
rect 34232 21029 34244 21063
rect 34278 21060 34290 21063
rect 34606 21060 34612 21072
rect 34278 21032 34612 21060
rect 34278 21029 34290 21032
rect 34232 21023 34290 21029
rect 34606 21020 34612 21032
rect 34664 21060 34670 21072
rect 35434 21060 35440 21072
rect 34664 21032 35440 21060
rect 34664 21020 34670 21032
rect 35434 21020 35440 21032
rect 35492 21020 35498 21072
rect 26970 21001 26976 21004
rect 26605 20995 26663 21001
rect 26605 20992 26617 20995
rect 26252 20964 26617 20992
rect 26605 20961 26617 20964
rect 26651 20961 26663 20995
rect 26605 20955 26663 20961
rect 26928 20995 26976 21001
rect 26928 20961 26940 20995
rect 26974 20961 26976 20995
rect 26928 20955 26976 20961
rect 26970 20952 26976 20955
rect 27028 20952 27034 21004
rect 30282 20992 30288 21004
rect 30243 20964 30288 20992
rect 30282 20952 30288 20964
rect 30340 20952 30346 21004
rect 32398 20952 32404 21004
rect 32456 20992 32462 21004
rect 33318 20992 33324 21004
rect 32456 20964 33324 20992
rect 32456 20952 32462 20964
rect 27062 20924 27068 20936
rect 27023 20896 27068 20924
rect 27062 20884 27068 20896
rect 27120 20884 27126 20936
rect 27338 20924 27344 20936
rect 27299 20896 27344 20924
rect 27338 20884 27344 20896
rect 27396 20884 27402 20936
rect 29822 20884 29828 20936
rect 29880 20924 29886 20936
rect 30377 20927 30435 20933
rect 30377 20924 30389 20927
rect 29880 20896 30389 20924
rect 29880 20884 29886 20896
rect 30377 20893 30389 20896
rect 30423 20893 30435 20927
rect 30377 20887 30435 20893
rect 30561 20927 30619 20933
rect 30561 20893 30573 20927
rect 30607 20924 30619 20927
rect 30742 20924 30748 20936
rect 30607 20896 30748 20924
rect 30607 20893 30619 20896
rect 30561 20887 30619 20893
rect 30392 20856 30420 20887
rect 30742 20884 30748 20896
rect 30800 20884 30806 20936
rect 31662 20884 31668 20936
rect 31720 20924 31726 20936
rect 32600 20933 32628 20964
rect 33318 20952 33324 20964
rect 33376 20952 33382 21004
rect 32585 20927 32643 20933
rect 32585 20924 32597 20927
rect 31720 20896 32597 20924
rect 31720 20884 31726 20896
rect 32585 20893 32597 20896
rect 32631 20893 32643 20927
rect 32766 20924 32772 20936
rect 32727 20896 32772 20924
rect 32585 20887 32643 20893
rect 32766 20884 32772 20896
rect 32824 20884 32830 20936
rect 33965 20927 34023 20933
rect 33965 20893 33977 20927
rect 34011 20893 34023 20927
rect 33965 20887 34023 20893
rect 32125 20859 32183 20865
rect 32125 20856 32137 20859
rect 30392 20828 32137 20856
rect 32125 20825 32137 20828
rect 32171 20825 32183 20859
rect 32125 20819 32183 20825
rect 20070 20788 20076 20800
rect 20031 20760 20076 20788
rect 20070 20748 20076 20760
rect 20128 20748 20134 20800
rect 25038 20748 25044 20800
rect 25096 20788 25102 20800
rect 25317 20791 25375 20797
rect 25317 20788 25329 20791
rect 25096 20760 25329 20788
rect 25096 20748 25102 20760
rect 25317 20757 25329 20760
rect 25363 20757 25375 20791
rect 25317 20751 25375 20757
rect 30374 20748 30380 20800
rect 30432 20788 30438 20800
rect 31481 20791 31539 20797
rect 31481 20788 31493 20791
rect 30432 20760 31493 20788
rect 30432 20748 30438 20760
rect 31481 20757 31493 20760
rect 31527 20788 31539 20791
rect 32766 20788 32772 20800
rect 31527 20760 32772 20788
rect 31527 20757 31539 20760
rect 31481 20751 31539 20757
rect 32766 20748 32772 20760
rect 32824 20748 32830 20800
rect 33980 20788 34008 20887
rect 34330 20788 34336 20800
rect 33980 20760 34336 20788
rect 34330 20748 34336 20760
rect 34388 20748 34394 20800
rect 35342 20788 35348 20800
rect 35303 20760 35348 20788
rect 35342 20748 35348 20760
rect 35400 20748 35406 20800
rect 35989 20791 36047 20797
rect 35989 20757 36001 20791
rect 36035 20788 36047 20791
rect 36170 20788 36176 20800
rect 36035 20760 36176 20788
rect 36035 20757 36047 20760
rect 35989 20751 36047 20757
rect 36170 20748 36176 20760
rect 36228 20748 36234 20800
rect 1104 20698 38824 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 38824 20698
rect 1104 20624 38824 20646
rect 19889 20587 19947 20593
rect 19889 20553 19901 20587
rect 19935 20584 19947 20587
rect 19935 20556 20944 20584
rect 19935 20553 19947 20556
rect 19889 20547 19947 20553
rect 18322 20408 18328 20460
rect 18380 20448 18386 20460
rect 19996 20457 20024 20556
rect 20916 20516 20944 20556
rect 21542 20544 21548 20596
rect 21600 20584 21606 20596
rect 22281 20587 22339 20593
rect 22281 20584 22293 20587
rect 21600 20556 22293 20584
rect 21600 20544 21606 20556
rect 22281 20553 22293 20556
rect 22327 20553 22339 20587
rect 22281 20547 22339 20553
rect 23477 20587 23535 20593
rect 23477 20553 23489 20587
rect 23523 20584 23535 20587
rect 23934 20584 23940 20596
rect 23523 20556 23940 20584
rect 23523 20553 23535 20556
rect 23477 20547 23535 20553
rect 23934 20544 23940 20556
rect 23992 20584 23998 20596
rect 24857 20587 24915 20593
rect 24857 20584 24869 20587
rect 23992 20556 24869 20584
rect 23992 20544 23998 20556
rect 24857 20553 24869 20556
rect 24903 20584 24915 20587
rect 25406 20584 25412 20596
rect 24903 20556 25412 20584
rect 24903 20553 24915 20556
rect 24857 20547 24915 20553
rect 20990 20516 20996 20528
rect 20903 20488 20996 20516
rect 20990 20476 20996 20488
rect 21048 20516 21054 20528
rect 21818 20516 21824 20528
rect 21048 20488 21824 20516
rect 21048 20476 21054 20488
rect 21818 20476 21824 20488
rect 21876 20516 21882 20528
rect 21913 20519 21971 20525
rect 21913 20516 21925 20519
rect 21876 20488 21925 20516
rect 21876 20476 21882 20488
rect 21913 20485 21925 20488
rect 21959 20485 21971 20519
rect 21913 20479 21971 20485
rect 19981 20451 20039 20457
rect 19981 20448 19993 20451
rect 18380 20420 19993 20448
rect 18380 20408 18386 20420
rect 19981 20417 19993 20420
rect 20027 20417 20039 20451
rect 24872 20448 24900 20547
rect 25406 20544 25412 20556
rect 25464 20584 25470 20596
rect 26421 20587 26479 20593
rect 25464 20556 26372 20584
rect 25464 20544 25470 20556
rect 26344 20516 26372 20556
rect 26421 20553 26433 20587
rect 26467 20584 26479 20587
rect 26786 20584 26792 20596
rect 26467 20556 26792 20584
rect 26467 20553 26479 20556
rect 26421 20547 26479 20553
rect 26786 20544 26792 20556
rect 26844 20544 26850 20596
rect 30742 20584 30748 20596
rect 30703 20556 30748 20584
rect 30742 20544 30748 20556
rect 30800 20544 30806 20596
rect 31294 20584 31300 20596
rect 31255 20556 31300 20584
rect 31294 20544 31300 20556
rect 31352 20544 31358 20596
rect 31570 20544 31576 20596
rect 31628 20584 31634 20596
rect 31665 20587 31723 20593
rect 31665 20584 31677 20587
rect 31628 20556 31677 20584
rect 31628 20544 31634 20556
rect 31665 20553 31677 20556
rect 31711 20553 31723 20587
rect 34606 20584 34612 20596
rect 34567 20556 34612 20584
rect 31665 20547 31723 20553
rect 34606 20544 34612 20556
rect 34664 20544 34670 20596
rect 26510 20516 26516 20528
rect 26344 20488 26516 20516
rect 26510 20476 26516 20488
rect 26568 20516 26574 20528
rect 28997 20519 29055 20525
rect 28997 20516 29009 20519
rect 26568 20488 29009 20516
rect 26568 20476 26574 20488
rect 28997 20485 29009 20488
rect 29043 20516 29055 20519
rect 29043 20488 29408 20516
rect 29043 20485 29055 20488
rect 28997 20479 29055 20485
rect 25041 20451 25099 20457
rect 25041 20448 25053 20451
rect 24872 20420 25053 20448
rect 19981 20411 20039 20417
rect 25041 20417 25053 20420
rect 25087 20417 25099 20451
rect 25041 20411 25099 20417
rect 27890 20408 27896 20460
rect 27948 20448 27954 20460
rect 29380 20457 29408 20488
rect 31846 20476 31852 20528
rect 31904 20476 31910 20528
rect 36630 20516 36636 20528
rect 36591 20488 36636 20516
rect 36630 20476 36636 20488
rect 36688 20476 36694 20528
rect 28077 20451 28135 20457
rect 28077 20448 28089 20451
rect 27948 20420 28089 20448
rect 27948 20408 27954 20420
rect 28077 20417 28089 20420
rect 28123 20417 28135 20451
rect 28077 20411 28135 20417
rect 29365 20451 29423 20457
rect 29365 20417 29377 20451
rect 29411 20417 29423 20451
rect 31864 20448 31892 20476
rect 32309 20451 32367 20457
rect 32309 20448 32321 20451
rect 31864 20420 32321 20448
rect 29365 20411 29423 20417
rect 32309 20417 32321 20420
rect 32355 20417 32367 20451
rect 32582 20448 32588 20460
rect 32543 20420 32588 20448
rect 32309 20411 32367 20417
rect 32582 20408 32588 20420
rect 32640 20408 32646 20460
rect 20070 20340 20076 20392
rect 20128 20380 20134 20392
rect 20237 20383 20295 20389
rect 20237 20380 20249 20383
rect 20128 20352 20249 20380
rect 20128 20340 20134 20352
rect 20237 20349 20249 20352
rect 20283 20349 20295 20383
rect 22462 20380 22468 20392
rect 22423 20352 22468 20380
rect 20237 20343 20295 20349
rect 22462 20340 22468 20352
rect 22520 20380 22526 20392
rect 23017 20383 23075 20389
rect 23017 20380 23029 20383
rect 22520 20352 23029 20380
rect 22520 20340 22526 20352
rect 23017 20349 23029 20352
rect 23063 20349 23075 20383
rect 23658 20380 23664 20392
rect 23619 20352 23664 20380
rect 23017 20343 23075 20349
rect 23658 20340 23664 20352
rect 23716 20380 23722 20392
rect 25314 20389 25320 20392
rect 24213 20383 24271 20389
rect 24213 20380 24225 20383
rect 23716 20352 24225 20380
rect 23716 20340 23722 20352
rect 24213 20349 24225 20352
rect 24259 20349 24271 20383
rect 25308 20380 25320 20389
rect 25275 20352 25320 20380
rect 24213 20343 24271 20349
rect 25308 20343 25320 20352
rect 25314 20340 25320 20343
rect 25372 20340 25378 20392
rect 26970 20340 26976 20392
rect 27028 20380 27034 20392
rect 27065 20383 27123 20389
rect 27065 20380 27077 20383
rect 27028 20352 27077 20380
rect 27028 20340 27034 20352
rect 27065 20349 27077 20352
rect 27111 20380 27123 20383
rect 27522 20380 27528 20392
rect 27111 20352 27528 20380
rect 27111 20349 27123 20352
rect 27065 20343 27123 20349
rect 27522 20340 27528 20352
rect 27580 20340 27586 20392
rect 31754 20340 31760 20392
rect 31812 20380 31818 20392
rect 31849 20383 31907 20389
rect 31849 20380 31861 20383
rect 31812 20352 31861 20380
rect 31812 20340 31818 20352
rect 31849 20349 31861 20352
rect 31895 20349 31907 20383
rect 32172 20383 32230 20389
rect 32172 20380 32184 20383
rect 31849 20343 31907 20349
rect 31956 20352 32184 20380
rect 27338 20272 27344 20324
rect 27396 20312 27402 20324
rect 27433 20315 27491 20321
rect 27433 20312 27445 20315
rect 27396 20284 27445 20312
rect 27396 20272 27402 20284
rect 27433 20281 27445 20284
rect 27479 20312 27491 20315
rect 27893 20315 27951 20321
rect 27893 20312 27905 20315
rect 27479 20284 27905 20312
rect 27479 20281 27491 20284
rect 27433 20275 27491 20281
rect 27893 20281 27905 20284
rect 27939 20312 27951 20315
rect 28074 20312 28080 20324
rect 27939 20284 28080 20312
rect 27939 20281 27951 20284
rect 27893 20275 27951 20281
rect 28074 20272 28080 20284
rect 28132 20272 28138 20324
rect 29454 20272 29460 20324
rect 29512 20312 29518 20324
rect 29610 20315 29668 20321
rect 29610 20312 29622 20315
rect 29512 20284 29622 20312
rect 29512 20272 29518 20284
rect 29610 20281 29622 20284
rect 29656 20312 29668 20315
rect 30374 20312 30380 20324
rect 29656 20284 30380 20312
rect 29656 20281 29668 20284
rect 29610 20275 29668 20281
rect 30374 20272 30380 20284
rect 30432 20272 30438 20324
rect 31570 20272 31576 20324
rect 31628 20312 31634 20324
rect 31956 20312 31984 20352
rect 32172 20349 32184 20352
rect 32218 20349 32230 20383
rect 35253 20383 35311 20389
rect 35253 20380 35265 20383
rect 32172 20343 32230 20349
rect 35084 20352 35265 20380
rect 31628 20284 31984 20312
rect 31628 20272 31634 20284
rect 21361 20247 21419 20253
rect 21361 20213 21373 20247
rect 21407 20244 21419 20247
rect 21542 20244 21548 20256
rect 21407 20216 21548 20244
rect 21407 20213 21419 20216
rect 21361 20207 21419 20213
rect 21542 20204 21548 20216
rect 21600 20204 21606 20256
rect 22646 20244 22652 20256
rect 22607 20216 22652 20244
rect 22646 20204 22652 20216
rect 22704 20204 22710 20256
rect 23842 20244 23848 20256
rect 23803 20216 23848 20244
rect 23842 20204 23848 20216
rect 23900 20204 23906 20256
rect 27522 20244 27528 20256
rect 27483 20216 27528 20244
rect 27522 20204 27528 20216
rect 27580 20204 27586 20256
rect 27982 20244 27988 20256
rect 27943 20216 27988 20244
rect 27982 20204 27988 20216
rect 28040 20244 28046 20256
rect 28537 20247 28595 20253
rect 28537 20244 28549 20247
rect 28040 20216 28549 20244
rect 28040 20204 28046 20216
rect 28537 20213 28549 20216
rect 28583 20213 28595 20247
rect 33686 20244 33692 20256
rect 33647 20216 33692 20244
rect 28537 20207 28595 20213
rect 33686 20204 33692 20216
rect 33744 20204 33750 20256
rect 34330 20244 34336 20256
rect 34291 20216 34336 20244
rect 34330 20204 34336 20216
rect 34388 20244 34394 20256
rect 35084 20253 35112 20352
rect 35253 20349 35265 20352
rect 35299 20349 35311 20383
rect 35253 20343 35311 20349
rect 35520 20315 35578 20321
rect 35520 20281 35532 20315
rect 35566 20312 35578 20315
rect 36170 20312 36176 20324
rect 35566 20284 36176 20312
rect 35566 20281 35578 20284
rect 35520 20275 35578 20281
rect 36170 20272 36176 20284
rect 36228 20272 36234 20324
rect 35069 20247 35127 20253
rect 35069 20244 35081 20247
rect 34388 20216 35081 20244
rect 34388 20204 34394 20216
rect 35069 20213 35081 20216
rect 35115 20213 35127 20247
rect 35069 20207 35127 20213
rect 1104 20154 38824 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 38824 20154
rect 1104 20080 38824 20102
rect 19705 20043 19763 20049
rect 19705 20009 19717 20043
rect 19751 20040 19763 20043
rect 20070 20040 20076 20052
rect 19751 20012 20076 20040
rect 19751 20009 19763 20012
rect 19705 20003 19763 20009
rect 20070 20000 20076 20012
rect 20128 20000 20134 20052
rect 20898 20040 20904 20052
rect 20859 20012 20904 20040
rect 20898 20000 20904 20012
rect 20956 20000 20962 20052
rect 21266 20040 21272 20052
rect 21227 20012 21272 20040
rect 21266 20000 21272 20012
rect 21324 20000 21330 20052
rect 22646 20040 22652 20052
rect 21376 20012 22652 20040
rect 17954 19864 17960 19916
rect 18012 19904 18018 19916
rect 18581 19907 18639 19913
rect 18581 19904 18593 19907
rect 18012 19876 18593 19904
rect 18012 19864 18018 19876
rect 18581 19873 18593 19876
rect 18627 19873 18639 19907
rect 18581 19867 18639 19873
rect 18046 19796 18052 19848
rect 18104 19836 18110 19848
rect 18322 19836 18328 19848
rect 18104 19808 18328 19836
rect 18104 19796 18110 19808
rect 18322 19796 18328 19808
rect 18380 19796 18386 19848
rect 21082 19796 21088 19848
rect 21140 19836 21146 19848
rect 21376 19845 21404 20012
rect 22646 20000 22652 20012
rect 22704 20000 22710 20052
rect 23474 20040 23480 20052
rect 23435 20012 23480 20040
rect 23474 20000 23480 20012
rect 23532 20000 23538 20052
rect 23750 20040 23756 20052
rect 23711 20012 23756 20040
rect 23750 20000 23756 20012
rect 23808 20000 23814 20052
rect 24118 20040 24124 20052
rect 24079 20012 24124 20040
rect 24118 20000 24124 20012
rect 24176 20000 24182 20052
rect 24210 20000 24216 20052
rect 24268 20040 24274 20052
rect 25133 20043 25191 20049
rect 24268 20012 24313 20040
rect 24268 20000 24274 20012
rect 25133 20009 25145 20043
rect 25179 20040 25191 20043
rect 25314 20040 25320 20052
rect 25179 20012 25320 20040
rect 25179 20009 25191 20012
rect 25133 20003 25191 20009
rect 25314 20000 25320 20012
rect 25372 20000 25378 20052
rect 25409 20043 25467 20049
rect 25409 20009 25421 20043
rect 25455 20040 25467 20043
rect 26142 20040 26148 20052
rect 25455 20012 26148 20040
rect 25455 20009 25467 20012
rect 25409 20003 25467 20009
rect 26142 20000 26148 20012
rect 26200 20000 26206 20052
rect 26329 20043 26387 20049
rect 26329 20009 26341 20043
rect 26375 20040 26387 20043
rect 26694 20040 26700 20052
rect 26375 20012 26700 20040
rect 26375 20009 26387 20012
rect 26329 20003 26387 20009
rect 26694 20000 26700 20012
rect 26752 20040 26758 20052
rect 27062 20040 27068 20052
rect 26752 20012 27068 20040
rect 26752 20000 26758 20012
rect 27062 20000 27068 20012
rect 27120 20000 27126 20052
rect 27798 20000 27804 20052
rect 27856 20040 27862 20052
rect 28445 20043 28503 20049
rect 28445 20040 28457 20043
rect 27856 20012 28457 20040
rect 27856 20000 27862 20012
rect 28445 20009 28457 20012
rect 28491 20009 28503 20043
rect 29454 20040 29460 20052
rect 29415 20012 29460 20040
rect 28445 20003 28503 20009
rect 29454 20000 29460 20012
rect 29512 20000 29518 20052
rect 29822 20040 29828 20052
rect 29783 20012 29828 20040
rect 29822 20000 29828 20012
rect 29880 20000 29886 20052
rect 29917 20043 29975 20049
rect 29917 20009 29929 20043
rect 29963 20040 29975 20043
rect 30282 20040 30288 20052
rect 29963 20012 30288 20040
rect 29963 20009 29975 20012
rect 29917 20003 29975 20009
rect 30282 20000 30288 20012
rect 30340 20040 30346 20052
rect 30377 20043 30435 20049
rect 30377 20040 30389 20043
rect 30340 20012 30389 20040
rect 30340 20000 30346 20012
rect 30377 20009 30389 20012
rect 30423 20009 30435 20043
rect 30742 20040 30748 20052
rect 30703 20012 30748 20040
rect 30377 20003 30435 20009
rect 30742 20000 30748 20012
rect 30800 20000 30806 20052
rect 31573 20043 31631 20049
rect 31573 20009 31585 20043
rect 31619 20040 31631 20043
rect 31662 20040 31668 20052
rect 31619 20012 31668 20040
rect 31619 20009 31631 20012
rect 31573 20003 31631 20009
rect 31662 20000 31668 20012
rect 31720 20000 31726 20052
rect 31846 20040 31852 20052
rect 31807 20012 31852 20040
rect 31846 20000 31852 20012
rect 31904 20040 31910 20052
rect 33226 20040 33232 20052
rect 31904 20012 33232 20040
rect 31904 20000 31910 20012
rect 33226 20000 33232 20012
rect 33284 20000 33290 20052
rect 33689 20043 33747 20049
rect 33689 20009 33701 20043
rect 33735 20040 33747 20043
rect 34606 20040 34612 20052
rect 33735 20012 34612 20040
rect 33735 20009 33747 20012
rect 33689 20003 33747 20009
rect 34606 20000 34612 20012
rect 34664 20000 34670 20052
rect 23492 19972 23520 20000
rect 27332 19975 27390 19981
rect 23492 19944 24256 19972
rect 22462 19904 22468 19916
rect 22423 19876 22468 19904
rect 22462 19864 22468 19876
rect 22520 19864 22526 19916
rect 24228 19904 24256 19944
rect 27332 19941 27344 19975
rect 27378 19972 27390 19975
rect 27890 19972 27896 19984
rect 27378 19944 27896 19972
rect 27378 19941 27390 19944
rect 27332 19935 27390 19941
rect 27890 19932 27896 19944
rect 27948 19932 27954 19984
rect 35060 19975 35118 19981
rect 35060 19941 35072 19975
rect 35106 19972 35118 19975
rect 35342 19972 35348 19984
rect 35106 19944 35348 19972
rect 35106 19941 35118 19944
rect 35060 19935 35118 19941
rect 35342 19932 35348 19944
rect 35400 19932 35406 19984
rect 26789 19907 26847 19913
rect 24228 19876 24348 19904
rect 21361 19839 21419 19845
rect 21361 19836 21373 19839
rect 21140 19808 21373 19836
rect 21140 19796 21146 19808
rect 21361 19805 21373 19808
rect 21407 19805 21419 19839
rect 21542 19836 21548 19848
rect 21455 19808 21548 19836
rect 21361 19799 21419 19805
rect 21542 19796 21548 19808
rect 21600 19836 21606 19848
rect 21910 19836 21916 19848
rect 21600 19808 21916 19836
rect 21600 19796 21606 19808
rect 21910 19796 21916 19808
rect 21968 19796 21974 19848
rect 24320 19845 24348 19876
rect 26789 19873 26801 19907
rect 26835 19904 26847 19907
rect 28074 19904 28080 19916
rect 26835 19876 28080 19904
rect 26835 19873 26847 19876
rect 26789 19867 26847 19873
rect 28074 19864 28080 19876
rect 28132 19864 28138 19916
rect 32582 19913 32588 19916
rect 32576 19904 32588 19913
rect 32543 19876 32588 19904
rect 32576 19867 32588 19876
rect 32582 19864 32588 19867
rect 32640 19864 32646 19916
rect 24305 19839 24363 19845
rect 24305 19805 24317 19839
rect 24351 19805 24363 19839
rect 24305 19799 24363 19805
rect 26510 19796 26516 19848
rect 26568 19836 26574 19848
rect 27062 19836 27068 19848
rect 26568 19808 27068 19836
rect 26568 19796 26574 19808
rect 27062 19796 27068 19808
rect 27120 19796 27126 19848
rect 32306 19836 32312 19848
rect 32267 19808 32312 19836
rect 32306 19796 32312 19808
rect 32364 19796 32370 19848
rect 34330 19796 34336 19848
rect 34388 19836 34394 19848
rect 34606 19836 34612 19848
rect 34388 19808 34612 19836
rect 34388 19796 34394 19808
rect 34606 19796 34612 19808
rect 34664 19836 34670 19848
rect 34793 19839 34851 19845
rect 34793 19836 34805 19839
rect 34664 19808 34805 19836
rect 34664 19796 34670 19808
rect 34793 19805 34805 19808
rect 34839 19805 34851 19839
rect 34793 19799 34851 19805
rect 16485 19703 16543 19709
rect 16485 19669 16497 19703
rect 16531 19700 16543 19703
rect 16574 19700 16580 19712
rect 16531 19672 16580 19700
rect 16531 19669 16543 19672
rect 16485 19663 16543 19669
rect 16574 19660 16580 19672
rect 16632 19660 16638 19712
rect 16853 19703 16911 19709
rect 16853 19669 16865 19703
rect 16899 19700 16911 19703
rect 16942 19700 16948 19712
rect 16899 19672 16948 19700
rect 16899 19669 16911 19672
rect 16853 19663 16911 19669
rect 16942 19660 16948 19672
rect 17000 19660 17006 19712
rect 18141 19703 18199 19709
rect 18141 19669 18153 19703
rect 18187 19700 18199 19703
rect 18322 19700 18328 19712
rect 18187 19672 18328 19700
rect 18187 19669 18199 19672
rect 18141 19663 18199 19669
rect 18322 19660 18328 19672
rect 18380 19660 18386 19712
rect 19334 19660 19340 19712
rect 19392 19700 19398 19712
rect 20622 19700 20628 19712
rect 19392 19672 20628 19700
rect 19392 19660 19398 19672
rect 20622 19660 20628 19672
rect 20680 19660 20686 19712
rect 21174 19660 21180 19712
rect 21232 19700 21238 19712
rect 22649 19703 22707 19709
rect 22649 19700 22661 19703
rect 21232 19672 22661 19700
rect 21232 19660 21238 19672
rect 22649 19669 22661 19672
rect 22695 19669 22707 19703
rect 36170 19700 36176 19712
rect 36131 19672 36176 19700
rect 22649 19663 22707 19669
rect 36170 19660 36176 19672
rect 36228 19660 36234 19712
rect 1104 19610 38824 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 38824 19610
rect 1104 19536 38824 19558
rect 20441 19499 20499 19505
rect 20441 19465 20453 19499
rect 20487 19496 20499 19499
rect 21082 19496 21088 19508
rect 20487 19468 21088 19496
rect 20487 19465 20499 19468
rect 20441 19459 20499 19465
rect 21082 19456 21088 19468
rect 21140 19456 21146 19508
rect 21266 19456 21272 19508
rect 21324 19496 21330 19508
rect 21545 19499 21603 19505
rect 21545 19496 21557 19499
rect 21324 19468 21557 19496
rect 21324 19456 21330 19468
rect 21545 19465 21557 19468
rect 21591 19465 21603 19499
rect 21910 19496 21916 19508
rect 21871 19468 21916 19496
rect 21545 19459 21603 19465
rect 21910 19456 21916 19468
rect 21968 19456 21974 19508
rect 24118 19456 24124 19508
rect 24176 19496 24182 19508
rect 24213 19499 24271 19505
rect 24213 19496 24225 19499
rect 24176 19468 24225 19496
rect 24176 19456 24182 19468
rect 24213 19465 24225 19468
rect 24259 19465 24271 19499
rect 24213 19459 24271 19465
rect 25041 19499 25099 19505
rect 25041 19465 25053 19499
rect 25087 19496 25099 19499
rect 26326 19496 26332 19508
rect 25087 19468 26332 19496
rect 25087 19465 25099 19468
rect 25041 19459 25099 19465
rect 26326 19456 26332 19468
rect 26384 19456 26390 19508
rect 26694 19496 26700 19508
rect 26655 19468 26700 19496
rect 26694 19456 26700 19468
rect 26752 19456 26758 19508
rect 27062 19456 27068 19508
rect 27120 19496 27126 19508
rect 27709 19499 27767 19505
rect 27709 19496 27721 19499
rect 27120 19468 27721 19496
rect 27120 19456 27126 19468
rect 27709 19465 27721 19468
rect 27755 19465 27767 19499
rect 27709 19459 27767 19465
rect 27890 19456 27896 19508
rect 27948 19496 27954 19508
rect 28077 19499 28135 19505
rect 28077 19496 28089 19499
rect 27948 19468 28089 19496
rect 27948 19456 27954 19468
rect 28077 19465 28089 19468
rect 28123 19465 28135 19499
rect 28077 19459 28135 19465
rect 31754 19456 31760 19508
rect 31812 19496 31818 19508
rect 31849 19499 31907 19505
rect 31849 19496 31861 19499
rect 31812 19468 31861 19496
rect 31812 19456 31818 19468
rect 31849 19465 31861 19468
rect 31895 19465 31907 19499
rect 31849 19459 31907 19465
rect 32582 19456 32588 19508
rect 32640 19496 32646 19508
rect 32677 19499 32735 19505
rect 32677 19496 32689 19499
rect 32640 19468 32689 19496
rect 32640 19456 32646 19468
rect 32677 19465 32689 19468
rect 32723 19465 32735 19499
rect 32677 19459 32735 19465
rect 32953 19499 33011 19505
rect 32953 19465 32965 19499
rect 32999 19496 33011 19499
rect 34606 19496 34612 19508
rect 32999 19468 34612 19496
rect 32999 19465 33011 19468
rect 32953 19459 33011 19465
rect 34606 19456 34612 19468
rect 34664 19456 34670 19508
rect 35342 19456 35348 19508
rect 35400 19496 35406 19508
rect 36081 19499 36139 19505
rect 36081 19496 36093 19499
rect 35400 19468 36093 19496
rect 35400 19456 35406 19468
rect 36081 19465 36093 19468
rect 36127 19465 36139 19499
rect 36081 19459 36139 19465
rect 35360 19428 35388 19456
rect 33888 19400 35388 19428
rect 33888 19372 33916 19400
rect 16666 19320 16672 19372
rect 16724 19360 16730 19372
rect 16945 19363 17003 19369
rect 16945 19360 16957 19363
rect 16724 19332 16957 19360
rect 16724 19320 16730 19332
rect 16945 19329 16957 19332
rect 16991 19329 17003 19363
rect 16945 19323 17003 19329
rect 17865 19363 17923 19369
rect 17865 19329 17877 19363
rect 17911 19360 17923 19363
rect 18046 19360 18052 19372
rect 17911 19332 18052 19360
rect 17911 19329 17923 19332
rect 17865 19323 17923 19329
rect 18046 19320 18052 19332
rect 18104 19320 18110 19372
rect 21174 19360 21180 19372
rect 20640 19332 21180 19360
rect 16574 19252 16580 19304
rect 16632 19292 16638 19304
rect 16761 19295 16819 19301
rect 16761 19292 16773 19295
rect 16632 19264 16773 19292
rect 16632 19252 16638 19264
rect 16761 19261 16773 19264
rect 16807 19292 16819 19295
rect 17954 19292 17960 19304
rect 16807 19264 17960 19292
rect 16807 19261 16819 19264
rect 16761 19255 16819 19261
rect 17954 19252 17960 19264
rect 18012 19252 18018 19304
rect 20073 19295 20131 19301
rect 20073 19261 20085 19295
rect 20119 19292 20131 19295
rect 20640 19292 20668 19332
rect 21174 19320 21180 19332
rect 21232 19320 21238 19372
rect 23937 19363 23995 19369
rect 23937 19329 23949 19363
rect 23983 19360 23995 19363
rect 24210 19360 24216 19372
rect 23983 19332 24216 19360
rect 23983 19329 23995 19332
rect 23937 19323 23995 19329
rect 24210 19320 24216 19332
rect 24268 19320 24274 19372
rect 25314 19320 25320 19372
rect 25372 19360 25378 19372
rect 25593 19363 25651 19369
rect 25593 19360 25605 19363
rect 25372 19332 25605 19360
rect 25372 19320 25378 19332
rect 25593 19329 25605 19332
rect 25639 19329 25651 19363
rect 25593 19323 25651 19329
rect 26237 19363 26295 19369
rect 26237 19329 26249 19363
rect 26283 19360 26295 19363
rect 27341 19363 27399 19369
rect 27341 19360 27353 19363
rect 26283 19332 27353 19360
rect 26283 19329 26295 19332
rect 26237 19323 26295 19329
rect 27341 19329 27353 19332
rect 27387 19360 27399 19363
rect 27798 19360 27804 19372
rect 27387 19332 27804 19360
rect 27387 19329 27399 19332
rect 27341 19323 27399 19329
rect 27798 19320 27804 19332
rect 27856 19320 27862 19372
rect 33870 19360 33876 19372
rect 33783 19332 33876 19360
rect 33870 19320 33876 19332
rect 33928 19320 33934 19372
rect 35621 19363 35679 19369
rect 35621 19360 35633 19363
rect 34440 19332 35633 19360
rect 20119 19264 20668 19292
rect 20119 19261 20131 19264
rect 20073 19255 20131 19261
rect 20714 19252 20720 19304
rect 20772 19292 20778 19304
rect 20901 19295 20959 19301
rect 20901 19292 20913 19295
rect 20772 19264 20913 19292
rect 20772 19252 20778 19264
rect 20901 19261 20913 19264
rect 20947 19292 20959 19295
rect 22189 19295 22247 19301
rect 22189 19292 22201 19295
rect 20947 19264 22201 19292
rect 20947 19261 20959 19264
rect 20901 19255 20959 19261
rect 22189 19261 22201 19264
rect 22235 19292 22247 19295
rect 22741 19295 22799 19301
rect 22741 19292 22753 19295
rect 22235 19264 22753 19292
rect 22235 19261 22247 19264
rect 22189 19255 22247 19261
rect 22741 19261 22753 19264
rect 22787 19261 22799 19295
rect 22741 19255 22799 19261
rect 25038 19252 25044 19304
rect 25096 19292 25102 19304
rect 25409 19295 25467 19301
rect 25409 19292 25421 19295
rect 25096 19264 25421 19292
rect 25096 19252 25102 19264
rect 25409 19261 25421 19264
rect 25455 19261 25467 19295
rect 25409 19255 25467 19261
rect 25498 19252 25504 19304
rect 25556 19292 25562 19304
rect 26050 19292 26056 19304
rect 25556 19264 26056 19292
rect 25556 19252 25562 19264
rect 26050 19252 26056 19264
rect 26108 19252 26114 19304
rect 27157 19295 27215 19301
rect 27157 19261 27169 19295
rect 27203 19292 27215 19295
rect 27522 19292 27528 19304
rect 27203 19264 27528 19292
rect 27203 19261 27215 19264
rect 27157 19255 27215 19261
rect 27522 19252 27528 19264
rect 27580 19252 27586 19304
rect 33134 19292 33140 19304
rect 33095 19264 33140 19292
rect 33134 19252 33140 19264
rect 33192 19292 33198 19304
rect 33686 19292 33692 19304
rect 33192 19264 33692 19292
rect 33192 19252 33198 19264
rect 33686 19252 33692 19264
rect 33744 19252 33750 19304
rect 34333 19295 34391 19301
rect 34333 19261 34345 19295
rect 34379 19292 34391 19295
rect 34440 19292 34468 19332
rect 35621 19329 35633 19332
rect 35667 19360 35679 19363
rect 36170 19360 36176 19372
rect 35667 19332 36176 19360
rect 35667 19329 35679 19332
rect 35621 19323 35679 19329
rect 36170 19320 36176 19332
rect 36228 19320 36234 19372
rect 34379 19264 34468 19292
rect 34379 19261 34391 19264
rect 34333 19255 34391 19261
rect 18322 19233 18328 19236
rect 16301 19227 16359 19233
rect 16301 19193 16313 19227
rect 16347 19224 16359 19227
rect 16853 19227 16911 19233
rect 16853 19224 16865 19227
rect 16347 19196 16865 19224
rect 16347 19193 16359 19196
rect 16301 19187 16359 19193
rect 16853 19193 16865 19196
rect 16899 19224 16911 19227
rect 18316 19224 18328 19233
rect 16899 19196 18328 19224
rect 16899 19193 16911 19196
rect 16853 19187 16911 19193
rect 18316 19187 18328 19196
rect 18322 19184 18328 19187
rect 18380 19184 18386 19236
rect 20990 19224 20996 19236
rect 20951 19196 20996 19224
rect 20990 19184 20996 19196
rect 21048 19184 21054 19236
rect 26605 19227 26663 19233
rect 26605 19193 26617 19227
rect 26651 19224 26663 19227
rect 27065 19227 27123 19233
rect 27065 19224 27077 19227
rect 26651 19196 27077 19224
rect 26651 19193 26663 19196
rect 26605 19187 26663 19193
rect 27065 19193 27077 19196
rect 27111 19224 27123 19227
rect 27430 19224 27436 19236
rect 27111 19196 27436 19224
rect 27111 19193 27123 19196
rect 27065 19187 27123 19193
rect 27430 19184 27436 19196
rect 27488 19184 27494 19236
rect 35529 19227 35587 19233
rect 35529 19224 35541 19227
rect 33244 19196 35541 19224
rect 15838 19156 15844 19168
rect 15799 19128 15844 19156
rect 15838 19116 15844 19128
rect 15896 19116 15902 19168
rect 16390 19156 16396 19168
rect 16351 19128 16396 19156
rect 16390 19116 16396 19128
rect 16448 19116 16454 19168
rect 19426 19156 19432 19168
rect 19387 19128 19432 19156
rect 19426 19116 19432 19128
rect 19484 19116 19490 19168
rect 20530 19156 20536 19168
rect 20491 19128 20536 19156
rect 20530 19116 20536 19128
rect 20588 19116 20594 19168
rect 22370 19156 22376 19168
rect 22331 19128 22376 19156
rect 22370 19116 22376 19128
rect 22428 19116 22434 19168
rect 23106 19156 23112 19168
rect 23067 19128 23112 19156
rect 23106 19116 23112 19128
rect 23164 19116 23170 19168
rect 24949 19159 25007 19165
rect 24949 19125 24961 19159
rect 24995 19156 25007 19159
rect 25498 19156 25504 19168
rect 24995 19128 25504 19156
rect 24995 19125 25007 19128
rect 24949 19119 25007 19125
rect 25498 19116 25504 19128
rect 25556 19116 25562 19168
rect 31938 19116 31944 19168
rect 31996 19156 32002 19168
rect 32306 19156 32312 19168
rect 31996 19128 32312 19156
rect 31996 19116 32002 19128
rect 32306 19116 32312 19128
rect 32364 19156 32370 19168
rect 33244 19165 33272 19196
rect 35529 19193 35541 19196
rect 35575 19224 35587 19227
rect 35710 19224 35716 19236
rect 35575 19196 35716 19224
rect 35575 19193 35587 19196
rect 35529 19187 35587 19193
rect 35710 19184 35716 19196
rect 35768 19184 35774 19236
rect 32953 19159 33011 19165
rect 32953 19156 32965 19159
rect 32364 19128 32965 19156
rect 32364 19116 32370 19128
rect 32953 19125 32965 19128
rect 32999 19125 33011 19159
rect 32953 19119 33011 19125
rect 33229 19159 33287 19165
rect 33229 19125 33241 19159
rect 33275 19125 33287 19159
rect 33229 19119 33287 19125
rect 33318 19116 33324 19168
rect 33376 19156 33382 19168
rect 33597 19159 33655 19165
rect 33597 19156 33609 19159
rect 33376 19128 33609 19156
rect 33376 19116 33382 19128
rect 33597 19125 33609 19128
rect 33643 19125 33655 19159
rect 33597 19119 33655 19125
rect 34698 19116 34704 19168
rect 34756 19156 34762 19168
rect 35069 19159 35127 19165
rect 35069 19156 35081 19159
rect 34756 19128 35081 19156
rect 34756 19116 34762 19128
rect 35069 19125 35081 19128
rect 35115 19125 35127 19159
rect 35069 19119 35127 19125
rect 35250 19116 35256 19168
rect 35308 19156 35314 19168
rect 35437 19159 35495 19165
rect 35437 19156 35449 19159
rect 35308 19128 35449 19156
rect 35308 19116 35314 19128
rect 35437 19125 35449 19128
rect 35483 19125 35495 19159
rect 35437 19119 35495 19125
rect 1104 19066 38824 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 38824 19066
rect 1104 18992 38824 19014
rect 15657 18955 15715 18961
rect 15657 18921 15669 18955
rect 15703 18952 15715 18955
rect 16390 18952 16396 18964
rect 15703 18924 16396 18952
rect 15703 18921 15715 18924
rect 15657 18915 15715 18921
rect 16390 18912 16396 18924
rect 16448 18912 16454 18964
rect 17954 18912 17960 18964
rect 18012 18952 18018 18964
rect 18693 18955 18751 18961
rect 18693 18952 18705 18955
rect 18012 18924 18705 18952
rect 18012 18912 18018 18924
rect 18693 18921 18705 18924
rect 18739 18952 18751 18955
rect 19426 18952 19432 18964
rect 18739 18924 19432 18952
rect 18739 18921 18751 18924
rect 18693 18915 18751 18921
rect 19426 18912 19432 18924
rect 19484 18912 19490 18964
rect 20625 18955 20683 18961
rect 20625 18921 20637 18955
rect 20671 18952 20683 18955
rect 20990 18952 20996 18964
rect 20671 18924 20996 18952
rect 20671 18921 20683 18924
rect 20625 18915 20683 18921
rect 20990 18912 20996 18924
rect 21048 18912 21054 18964
rect 21269 18955 21327 18961
rect 21269 18921 21281 18955
rect 21315 18952 21327 18955
rect 22462 18952 22468 18964
rect 21315 18924 22468 18952
rect 21315 18921 21327 18924
rect 21269 18915 21327 18921
rect 22462 18912 22468 18924
rect 22520 18952 22526 18964
rect 23106 18952 23112 18964
rect 22520 18924 23112 18952
rect 22520 18912 22526 18924
rect 23106 18912 23112 18924
rect 23164 18912 23170 18964
rect 23474 18912 23480 18964
rect 23532 18952 23538 18964
rect 23753 18955 23811 18961
rect 23753 18952 23765 18955
rect 23532 18924 23765 18952
rect 23532 18912 23538 18924
rect 23753 18921 23765 18924
rect 23799 18921 23811 18955
rect 25038 18952 25044 18964
rect 24999 18924 25044 18952
rect 23753 18915 23811 18921
rect 25038 18912 25044 18924
rect 25096 18912 25102 18964
rect 27522 18952 27528 18964
rect 27483 18924 27528 18952
rect 27522 18912 27528 18924
rect 27580 18912 27586 18964
rect 33226 18952 33232 18964
rect 33187 18924 33232 18952
rect 33226 18912 33232 18924
rect 33284 18912 33290 18964
rect 33689 18955 33747 18961
rect 33689 18921 33701 18955
rect 33735 18952 33747 18955
rect 33870 18952 33876 18964
rect 33735 18924 33876 18952
rect 33735 18921 33747 18924
rect 33689 18915 33747 18921
rect 33870 18912 33876 18924
rect 33928 18912 33934 18964
rect 35161 18955 35219 18961
rect 35161 18921 35173 18955
rect 35207 18952 35219 18955
rect 35250 18952 35256 18964
rect 35207 18924 35256 18952
rect 35207 18921 35219 18924
rect 35161 18915 35219 18921
rect 35250 18912 35256 18924
rect 35308 18912 35314 18964
rect 35710 18952 35716 18964
rect 35671 18924 35716 18952
rect 35710 18912 35716 18924
rect 35768 18912 35774 18964
rect 9950 18893 9956 18896
rect 9944 18884 9956 18893
rect 9911 18856 9956 18884
rect 9944 18847 9956 18856
rect 9950 18844 9956 18847
rect 10008 18844 10014 18896
rect 18046 18844 18052 18896
rect 18104 18884 18110 18896
rect 18325 18887 18383 18893
rect 18325 18884 18337 18887
rect 18104 18856 18337 18884
rect 18104 18844 18110 18856
rect 18325 18853 18337 18856
rect 18371 18853 18383 18887
rect 20898 18884 20904 18896
rect 20859 18856 20904 18884
rect 18325 18847 18383 18853
rect 20898 18844 20904 18856
rect 20956 18844 20962 18896
rect 27157 18887 27215 18893
rect 27157 18853 27169 18887
rect 27203 18884 27215 18887
rect 27890 18884 27896 18896
rect 27203 18856 27896 18884
rect 27203 18853 27215 18856
rect 27157 18847 27215 18853
rect 27890 18844 27896 18856
rect 27948 18844 27954 18896
rect 16206 18776 16212 18828
rect 16264 18816 16270 18828
rect 16373 18819 16431 18825
rect 16373 18816 16385 18819
rect 16264 18788 16385 18816
rect 16264 18776 16270 18788
rect 16373 18785 16385 18788
rect 16419 18785 16431 18819
rect 16373 18779 16431 18785
rect 19426 18776 19432 18828
rect 19484 18816 19490 18828
rect 19613 18819 19671 18825
rect 19613 18816 19625 18819
rect 19484 18788 19625 18816
rect 19484 18776 19490 18788
rect 19613 18785 19625 18788
rect 19659 18785 19671 18819
rect 19613 18779 19671 18785
rect 20070 18776 20076 18828
rect 20128 18816 20134 18828
rect 21085 18819 21143 18825
rect 21085 18816 21097 18819
rect 20128 18788 21097 18816
rect 20128 18776 20134 18788
rect 21085 18785 21097 18788
rect 21131 18785 21143 18819
rect 21085 18779 21143 18785
rect 22097 18819 22155 18825
rect 22097 18785 22109 18819
rect 22143 18816 22155 18819
rect 22830 18816 22836 18828
rect 22143 18788 22836 18816
rect 22143 18785 22155 18788
rect 22097 18779 22155 18785
rect 22830 18776 22836 18788
rect 22888 18776 22894 18828
rect 9674 18748 9680 18760
rect 9635 18720 9680 18748
rect 9674 18708 9680 18720
rect 9732 18708 9738 18760
rect 16117 18751 16175 18757
rect 16117 18717 16129 18751
rect 16163 18717 16175 18751
rect 19702 18748 19708 18760
rect 19663 18720 19708 18748
rect 16117 18711 16175 18717
rect 11054 18612 11060 18624
rect 11015 18584 11060 18612
rect 11054 18572 11060 18584
rect 11112 18572 11118 18624
rect 14918 18612 14924 18624
rect 14879 18584 14924 18612
rect 14918 18572 14924 18584
rect 14976 18572 14982 18624
rect 15930 18612 15936 18624
rect 15891 18584 15936 18612
rect 15930 18572 15936 18584
rect 15988 18572 15994 18624
rect 16132 18612 16160 18711
rect 19702 18708 19708 18720
rect 19760 18708 19766 18760
rect 19889 18751 19947 18757
rect 19889 18717 19901 18751
rect 19935 18748 19947 18751
rect 19978 18748 19984 18760
rect 19935 18720 19984 18748
rect 19935 18717 19947 18720
rect 19889 18711 19947 18717
rect 19978 18708 19984 18720
rect 20036 18708 20042 18760
rect 32030 18708 32036 18760
rect 32088 18748 32094 18760
rect 32125 18751 32183 18757
rect 32125 18748 32137 18751
rect 32088 18720 32137 18748
rect 32088 18708 32094 18720
rect 32125 18717 32137 18720
rect 32171 18717 32183 18751
rect 32125 18711 32183 18717
rect 19245 18683 19303 18689
rect 19245 18649 19257 18683
rect 19291 18680 19303 18683
rect 19334 18680 19340 18692
rect 19291 18652 19340 18680
rect 19291 18649 19303 18652
rect 19245 18643 19303 18649
rect 19334 18640 19340 18652
rect 19392 18640 19398 18692
rect 21637 18683 21695 18689
rect 21637 18649 21649 18683
rect 21683 18680 21695 18683
rect 21818 18680 21824 18692
rect 21683 18652 21824 18680
rect 21683 18649 21695 18652
rect 21637 18643 21695 18649
rect 21818 18640 21824 18652
rect 21876 18680 21882 18692
rect 22281 18683 22339 18689
rect 22281 18680 22293 18683
rect 21876 18652 22293 18680
rect 21876 18640 21882 18652
rect 22281 18649 22293 18652
rect 22327 18649 22339 18683
rect 22281 18643 22339 18649
rect 16298 18612 16304 18624
rect 16132 18584 16304 18612
rect 16298 18572 16304 18584
rect 16356 18572 16362 18624
rect 17494 18612 17500 18624
rect 17455 18584 17500 18612
rect 17494 18572 17500 18584
rect 17552 18572 17558 18624
rect 22002 18612 22008 18624
rect 21963 18584 22008 18612
rect 22002 18572 22008 18584
rect 22060 18572 22066 18624
rect 26789 18615 26847 18621
rect 26789 18581 26801 18615
rect 26835 18612 26847 18615
rect 27154 18612 27160 18624
rect 26835 18584 27160 18612
rect 26835 18581 26847 18584
rect 26789 18575 26847 18581
rect 27154 18572 27160 18584
rect 27212 18572 27218 18624
rect 30653 18615 30711 18621
rect 30653 18581 30665 18615
rect 30699 18612 30711 18615
rect 31110 18612 31116 18624
rect 30699 18584 31116 18612
rect 30699 18581 30711 18584
rect 30653 18575 30711 18581
rect 31110 18572 31116 18584
rect 31168 18572 31174 18624
rect 32674 18612 32680 18624
rect 32635 18584 32680 18612
rect 32674 18572 32680 18584
rect 32732 18572 32738 18624
rect 1104 18522 38824 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 38824 18522
rect 1104 18448 38824 18470
rect 7374 18408 7380 18420
rect 7335 18380 7380 18408
rect 7374 18368 7380 18380
rect 7432 18368 7438 18420
rect 9950 18368 9956 18420
rect 10008 18408 10014 18420
rect 10045 18411 10103 18417
rect 10045 18408 10057 18411
rect 10008 18380 10057 18408
rect 10008 18368 10014 18380
rect 10045 18377 10057 18380
rect 10091 18377 10103 18411
rect 10045 18371 10103 18377
rect 14829 18411 14887 18417
rect 14829 18377 14841 18411
rect 14875 18408 14887 18411
rect 15930 18408 15936 18420
rect 14875 18380 15936 18408
rect 14875 18377 14887 18380
rect 14829 18371 14887 18377
rect 15930 18368 15936 18380
rect 15988 18408 15994 18420
rect 16850 18408 16856 18420
rect 15988 18380 16856 18408
rect 15988 18368 15994 18380
rect 16850 18368 16856 18380
rect 16908 18368 16914 18420
rect 17865 18411 17923 18417
rect 17865 18377 17877 18411
rect 17911 18408 17923 18411
rect 18046 18408 18052 18420
rect 17911 18380 18052 18408
rect 17911 18377 17923 18380
rect 17865 18371 17923 18377
rect 18046 18368 18052 18380
rect 18104 18368 18110 18420
rect 18322 18368 18328 18420
rect 18380 18408 18386 18420
rect 19429 18411 19487 18417
rect 19429 18408 19441 18411
rect 18380 18380 19441 18408
rect 18380 18368 18386 18380
rect 19429 18377 19441 18380
rect 19475 18377 19487 18411
rect 19429 18371 19487 18377
rect 20070 18368 20076 18420
rect 20128 18408 20134 18420
rect 20533 18411 20591 18417
rect 20533 18408 20545 18411
rect 20128 18380 20545 18408
rect 20128 18368 20134 18380
rect 20533 18377 20545 18380
rect 20579 18377 20591 18411
rect 20898 18408 20904 18420
rect 20859 18380 20904 18408
rect 20533 18371 20591 18377
rect 20898 18368 20904 18380
rect 20956 18368 20962 18420
rect 20990 18368 20996 18420
rect 21048 18408 21054 18420
rect 21361 18411 21419 18417
rect 21361 18408 21373 18411
rect 21048 18380 21373 18408
rect 21048 18368 21054 18380
rect 21361 18377 21373 18380
rect 21407 18377 21419 18411
rect 26510 18408 26516 18420
rect 26471 18380 26516 18408
rect 21361 18371 21419 18377
rect 26510 18368 26516 18380
rect 26568 18368 26574 18420
rect 32030 18408 32036 18420
rect 31991 18380 32036 18408
rect 32030 18368 32036 18380
rect 32088 18368 32094 18420
rect 7392 18272 7420 18368
rect 7392 18244 7696 18272
rect 7558 18204 7564 18216
rect 7519 18176 7564 18204
rect 7558 18164 7564 18176
rect 7616 18164 7622 18216
rect 7668 18204 7696 18244
rect 14918 18232 14924 18284
rect 14976 18272 14982 18284
rect 15473 18275 15531 18281
rect 15473 18272 15485 18275
rect 14976 18244 15485 18272
rect 14976 18232 14982 18244
rect 15473 18241 15485 18244
rect 15519 18272 15531 18275
rect 15838 18272 15844 18284
rect 15519 18244 15844 18272
rect 15519 18241 15531 18244
rect 15473 18235 15531 18241
rect 15838 18232 15844 18244
rect 15896 18272 15902 18284
rect 16482 18272 16488 18284
rect 15896 18244 16488 18272
rect 15896 18232 15902 18244
rect 16482 18232 16488 18244
rect 16540 18232 16546 18284
rect 16942 18272 16948 18284
rect 16903 18244 16948 18272
rect 16942 18232 16948 18244
rect 17000 18272 17006 18284
rect 17862 18272 17868 18284
rect 17000 18244 17868 18272
rect 17000 18232 17006 18244
rect 17862 18232 17868 18244
rect 17920 18232 17926 18284
rect 18064 18281 18092 18368
rect 26697 18343 26755 18349
rect 26697 18309 26709 18343
rect 26743 18340 26755 18343
rect 27430 18340 27436 18352
rect 26743 18312 27436 18340
rect 26743 18309 26755 18312
rect 26697 18303 26755 18309
rect 27430 18300 27436 18312
rect 27488 18300 27494 18352
rect 30558 18340 30564 18352
rect 30519 18312 30564 18340
rect 30558 18300 30564 18312
rect 30616 18300 30622 18352
rect 18049 18275 18107 18281
rect 18049 18241 18061 18275
rect 18095 18241 18107 18275
rect 21818 18272 21824 18284
rect 21779 18244 21824 18272
rect 18049 18235 18107 18241
rect 21818 18232 21824 18244
rect 21876 18232 21882 18284
rect 22002 18272 22008 18284
rect 21963 18244 22008 18272
rect 22002 18232 22008 18244
rect 22060 18232 22066 18284
rect 26237 18275 26295 18281
rect 26237 18241 26249 18275
rect 26283 18272 26295 18275
rect 27249 18275 27307 18281
rect 27249 18272 27261 18275
rect 26283 18244 27261 18272
rect 26283 18241 26295 18244
rect 26237 18235 26295 18241
rect 27249 18241 27261 18244
rect 27295 18272 27307 18275
rect 27338 18272 27344 18284
rect 27295 18244 27344 18272
rect 27295 18241 27307 18244
rect 27249 18235 27307 18241
rect 27338 18232 27344 18244
rect 27396 18232 27402 18284
rect 31110 18272 31116 18284
rect 31071 18244 31116 18272
rect 31110 18232 31116 18244
rect 31168 18232 31174 18284
rect 7817 18207 7875 18213
rect 7817 18204 7829 18207
rect 7668 18176 7829 18204
rect 7817 18173 7829 18176
rect 7863 18173 7875 18207
rect 7817 18167 7875 18173
rect 14737 18207 14795 18213
rect 14737 18173 14749 18207
rect 14783 18204 14795 18207
rect 15289 18207 15347 18213
rect 15289 18204 15301 18207
rect 14783 18176 15301 18204
rect 14783 18173 14795 18176
rect 14737 18167 14795 18173
rect 15289 18173 15301 18176
rect 15335 18204 15347 18207
rect 16206 18204 16212 18216
rect 15335 18176 16212 18204
rect 15335 18173 15347 18176
rect 15289 18167 15347 18173
rect 16206 18164 16212 18176
rect 16264 18164 16270 18216
rect 16390 18164 16396 18216
rect 16448 18204 16454 18216
rect 16761 18207 16819 18213
rect 16761 18204 16773 18207
rect 16448 18176 16773 18204
rect 16448 18164 16454 18176
rect 16761 18173 16773 18176
rect 16807 18173 16819 18207
rect 16761 18167 16819 18173
rect 16850 18164 16856 18216
rect 16908 18204 16914 18216
rect 27154 18204 27160 18216
rect 16908 18176 16953 18204
rect 27115 18176 27160 18204
rect 16908 18164 16914 18176
rect 27154 18164 27160 18176
rect 27212 18164 27218 18216
rect 32048 18204 32076 18368
rect 32769 18275 32827 18281
rect 32769 18241 32781 18275
rect 32815 18272 32827 18275
rect 32950 18272 32956 18284
rect 32815 18244 32956 18272
rect 32815 18241 32827 18244
rect 32769 18235 32827 18241
rect 32493 18207 32551 18213
rect 32493 18204 32505 18207
rect 32048 18176 32505 18204
rect 32493 18173 32505 18176
rect 32539 18173 32551 18207
rect 32493 18167 32551 18173
rect 17405 18139 17463 18145
rect 17405 18136 17417 18139
rect 15212 18108 17417 18136
rect 15212 18080 15240 18108
rect 17405 18105 17417 18108
rect 17451 18136 17463 18139
rect 17494 18136 17500 18148
rect 17451 18108 17500 18136
rect 17451 18105 17463 18108
rect 17405 18099 17463 18105
rect 17494 18096 17500 18108
rect 17552 18136 17558 18148
rect 18294 18139 18352 18145
rect 18294 18136 18306 18139
rect 17552 18108 18306 18136
rect 17552 18096 17558 18108
rect 18294 18105 18306 18108
rect 18340 18105 18352 18139
rect 18294 18099 18352 18105
rect 19334 18096 19340 18148
rect 19392 18136 19398 18148
rect 19702 18136 19708 18148
rect 19392 18108 19708 18136
rect 19392 18096 19398 18108
rect 19702 18096 19708 18108
rect 19760 18136 19766 18148
rect 19981 18139 20039 18145
rect 19981 18136 19993 18139
rect 19760 18108 19993 18136
rect 19760 18096 19766 18108
rect 19981 18105 19993 18108
rect 20027 18105 20039 18139
rect 19981 18099 20039 18105
rect 26510 18096 26516 18148
rect 26568 18136 26574 18148
rect 27065 18139 27123 18145
rect 27065 18136 27077 18139
rect 26568 18108 27077 18136
rect 26568 18096 26574 18108
rect 27065 18105 27077 18108
rect 27111 18105 27123 18139
rect 27065 18099 27123 18105
rect 30469 18139 30527 18145
rect 30469 18105 30481 18139
rect 30515 18136 30527 18139
rect 30926 18136 30932 18148
rect 30515 18108 30932 18136
rect 30515 18105 30527 18108
rect 30469 18099 30527 18105
rect 30926 18096 30932 18108
rect 30984 18096 30990 18148
rect 32784 18136 32812 18235
rect 32950 18232 32956 18244
rect 33008 18232 33014 18284
rect 31588 18108 32812 18136
rect 8938 18068 8944 18080
rect 8899 18040 8944 18068
rect 8938 18028 8944 18040
rect 8996 18028 9002 18080
rect 9674 18068 9680 18080
rect 9635 18040 9680 18068
rect 9674 18028 9680 18040
rect 9732 18028 9738 18080
rect 15194 18068 15200 18080
rect 15155 18040 15200 18068
rect 15194 18028 15200 18040
rect 15252 18028 15258 18080
rect 16209 18071 16267 18077
rect 16209 18037 16221 18071
rect 16255 18068 16267 18071
rect 16298 18068 16304 18080
rect 16255 18040 16304 18068
rect 16255 18037 16267 18040
rect 16209 18031 16267 18037
rect 16298 18028 16304 18040
rect 16356 18028 16362 18080
rect 16393 18071 16451 18077
rect 16393 18037 16405 18071
rect 16439 18068 16451 18071
rect 16482 18068 16488 18080
rect 16439 18040 16488 18068
rect 16439 18037 16451 18040
rect 16393 18031 16451 18037
rect 16482 18028 16488 18040
rect 16540 18028 16546 18080
rect 21729 18071 21787 18077
rect 21729 18037 21741 18071
rect 21775 18068 21787 18071
rect 22462 18068 22468 18080
rect 21775 18040 22468 18068
rect 21775 18037 21787 18040
rect 21729 18031 21787 18037
rect 22462 18028 22468 18040
rect 22520 18028 22526 18080
rect 22830 18068 22836 18080
rect 22743 18040 22836 18068
rect 22830 18028 22836 18040
rect 22888 18068 22894 18080
rect 23382 18068 23388 18080
rect 22888 18040 23388 18068
rect 22888 18028 22894 18040
rect 23382 18028 23388 18040
rect 23440 18028 23446 18080
rect 24397 18071 24455 18077
rect 24397 18037 24409 18071
rect 24443 18068 24455 18071
rect 24670 18068 24676 18080
rect 24443 18040 24676 18068
rect 24443 18037 24455 18040
rect 24397 18031 24455 18037
rect 24670 18028 24676 18040
rect 24728 18028 24734 18080
rect 30006 18068 30012 18080
rect 29967 18040 30012 18068
rect 30006 18028 30012 18040
rect 30064 18068 30070 18080
rect 31021 18071 31079 18077
rect 31021 18068 31033 18071
rect 30064 18040 31033 18068
rect 30064 18028 30070 18040
rect 31021 18037 31033 18040
rect 31067 18037 31079 18071
rect 31021 18031 31079 18037
rect 31478 18028 31484 18080
rect 31536 18068 31542 18080
rect 31588 18077 31616 18108
rect 31573 18071 31631 18077
rect 31573 18068 31585 18071
rect 31536 18040 31585 18068
rect 31536 18028 31542 18040
rect 31573 18037 31585 18040
rect 31619 18037 31631 18071
rect 31573 18031 31631 18037
rect 32125 18071 32183 18077
rect 32125 18037 32137 18071
rect 32171 18068 32183 18071
rect 32214 18068 32220 18080
rect 32171 18040 32220 18068
rect 32171 18037 32183 18040
rect 32125 18031 32183 18037
rect 32214 18028 32220 18040
rect 32272 18028 32278 18080
rect 32585 18071 32643 18077
rect 32585 18037 32597 18071
rect 32631 18068 32643 18071
rect 32674 18068 32680 18080
rect 32631 18040 32680 18068
rect 32631 18037 32643 18040
rect 32585 18031 32643 18037
rect 32674 18028 32680 18040
rect 32732 18068 32738 18080
rect 33042 18068 33048 18080
rect 32732 18040 33048 18068
rect 32732 18028 32738 18040
rect 33042 18028 33048 18040
rect 33100 18028 33106 18080
rect 1104 17978 38824 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 38824 17978
rect 1104 17904 38824 17926
rect 14921 17867 14979 17873
rect 14921 17833 14933 17867
rect 14967 17864 14979 17867
rect 15102 17864 15108 17876
rect 14967 17836 15108 17864
rect 14967 17833 14979 17836
rect 14921 17827 14979 17833
rect 15102 17824 15108 17836
rect 15160 17824 15166 17876
rect 15565 17867 15623 17873
rect 15565 17833 15577 17867
rect 15611 17864 15623 17867
rect 15746 17864 15752 17876
rect 15611 17836 15752 17864
rect 15611 17833 15623 17836
rect 15565 17827 15623 17833
rect 15746 17824 15752 17836
rect 15804 17864 15810 17876
rect 17865 17867 17923 17873
rect 17865 17864 17877 17867
rect 15804 17836 17877 17864
rect 15804 17824 15810 17836
rect 17865 17833 17877 17836
rect 17911 17833 17923 17867
rect 17865 17827 17923 17833
rect 17954 17824 17960 17876
rect 18012 17864 18018 17876
rect 18690 17864 18696 17876
rect 18012 17836 18696 17864
rect 18012 17824 18018 17836
rect 18690 17824 18696 17836
rect 18748 17864 18754 17876
rect 18785 17867 18843 17873
rect 18785 17864 18797 17867
rect 18748 17836 18797 17864
rect 18748 17824 18754 17836
rect 18785 17833 18797 17836
rect 18831 17833 18843 17867
rect 18785 17827 18843 17833
rect 19153 17867 19211 17873
rect 19153 17833 19165 17867
rect 19199 17864 19211 17867
rect 19334 17864 19340 17876
rect 19199 17836 19340 17864
rect 19199 17833 19211 17836
rect 19153 17827 19211 17833
rect 18800 17796 18828 17827
rect 19334 17824 19340 17836
rect 19392 17824 19398 17876
rect 19426 17824 19432 17876
rect 19484 17864 19490 17876
rect 19521 17867 19579 17873
rect 19521 17864 19533 17867
rect 19484 17836 19533 17864
rect 19484 17824 19490 17836
rect 19521 17833 19533 17836
rect 19567 17833 19579 17867
rect 19521 17827 19579 17833
rect 22462 17824 22468 17876
rect 22520 17864 22526 17876
rect 23017 17867 23075 17873
rect 23017 17864 23029 17867
rect 22520 17836 23029 17864
rect 22520 17824 22526 17836
rect 23017 17833 23029 17836
rect 23063 17833 23075 17867
rect 30926 17864 30932 17876
rect 30887 17836 30932 17864
rect 23017 17827 23075 17833
rect 30926 17824 30932 17836
rect 30984 17824 30990 17876
rect 32950 17824 32956 17876
rect 33008 17864 33014 17876
rect 33505 17867 33563 17873
rect 33505 17864 33517 17867
rect 33008 17836 33517 17864
rect 33008 17824 33014 17836
rect 33505 17833 33517 17836
rect 33551 17833 33563 17867
rect 33505 17827 33563 17833
rect 20625 17799 20683 17805
rect 20625 17796 20637 17799
rect 18800 17768 20637 17796
rect 20625 17765 20637 17768
rect 20671 17796 20683 17799
rect 21542 17796 21548 17808
rect 20671 17768 21548 17796
rect 20671 17765 20683 17768
rect 20625 17759 20683 17765
rect 21542 17756 21548 17768
rect 21600 17756 21606 17808
rect 32306 17756 32312 17808
rect 32364 17805 32370 17808
rect 32364 17799 32428 17805
rect 32364 17765 32382 17799
rect 32416 17765 32428 17799
rect 32364 17759 32428 17765
rect 32364 17756 32370 17759
rect 16758 17737 16764 17740
rect 16752 17728 16764 17737
rect 16719 17700 16764 17728
rect 16752 17691 16764 17700
rect 16758 17688 16764 17691
rect 16816 17688 16822 17740
rect 18966 17728 18972 17740
rect 18927 17700 18972 17728
rect 18966 17688 18972 17700
rect 19024 17688 19030 17740
rect 20714 17688 20720 17740
rect 20772 17728 20778 17740
rect 21637 17731 21695 17737
rect 21637 17728 21649 17731
rect 20772 17700 21649 17728
rect 20772 17688 20778 17700
rect 21637 17697 21649 17700
rect 21683 17697 21695 17731
rect 22830 17728 22836 17740
rect 22791 17700 22836 17728
rect 21637 17691 21695 17697
rect 22830 17688 22836 17700
rect 22888 17688 22894 17740
rect 24118 17688 24124 17740
rect 24176 17728 24182 17740
rect 24673 17731 24731 17737
rect 24673 17728 24685 17731
rect 24176 17700 24685 17728
rect 24176 17688 24182 17700
rect 24673 17697 24685 17700
rect 24719 17697 24731 17731
rect 24673 17691 24731 17697
rect 27614 17688 27620 17740
rect 27672 17728 27678 17740
rect 28074 17728 28080 17740
rect 27672 17700 28080 17728
rect 27672 17688 27678 17700
rect 28074 17688 28080 17700
rect 28132 17728 28138 17740
rect 28308 17731 28366 17737
rect 28308 17728 28320 17731
rect 28132 17700 28320 17728
rect 28132 17688 28138 17700
rect 28308 17697 28320 17700
rect 28354 17697 28366 17731
rect 28308 17691 28366 17697
rect 28534 17688 28540 17740
rect 28592 17728 28598 17740
rect 28721 17731 28779 17737
rect 28721 17728 28733 17731
rect 28592 17700 28733 17728
rect 28592 17688 28598 17700
rect 28721 17697 28733 17700
rect 28767 17697 28779 17731
rect 35434 17728 35440 17740
rect 35395 17700 35440 17728
rect 28721 17691 28779 17697
rect 35434 17688 35440 17700
rect 35492 17688 35498 17740
rect 16298 17620 16304 17672
rect 16356 17660 16362 17672
rect 16485 17663 16543 17669
rect 16485 17660 16497 17663
rect 16356 17632 16497 17660
rect 16356 17620 16362 17632
rect 16485 17629 16497 17632
rect 16531 17629 16543 17663
rect 19978 17660 19984 17672
rect 19939 17632 19984 17660
rect 16485 17623 16543 17629
rect 19978 17620 19984 17632
rect 20036 17620 20042 17672
rect 21726 17660 21732 17672
rect 21687 17632 21732 17660
rect 21726 17620 21732 17632
rect 21784 17620 21790 17672
rect 21910 17660 21916 17672
rect 21871 17632 21916 17660
rect 21910 17620 21916 17632
rect 21968 17620 21974 17672
rect 24762 17660 24768 17672
rect 24723 17632 24768 17660
rect 24762 17620 24768 17632
rect 24820 17620 24826 17672
rect 24857 17663 24915 17669
rect 24857 17629 24869 17663
rect 24903 17629 24915 17663
rect 26602 17660 26608 17672
rect 26563 17632 26608 17660
rect 24857 17623 24915 17629
rect 7558 17552 7564 17604
rect 7616 17592 7622 17604
rect 7653 17595 7711 17601
rect 7653 17592 7665 17595
rect 7616 17564 7665 17592
rect 7616 17552 7622 17564
rect 7653 17561 7665 17564
rect 7699 17592 7711 17595
rect 8478 17592 8484 17604
rect 7699 17564 8484 17592
rect 7699 17561 7711 17564
rect 7653 17555 7711 17561
rect 8478 17552 8484 17564
rect 8536 17552 8542 17604
rect 23753 17595 23811 17601
rect 23753 17561 23765 17595
rect 23799 17592 23811 17595
rect 24026 17592 24032 17604
rect 23799 17564 24032 17592
rect 23799 17561 23811 17564
rect 23753 17555 23811 17561
rect 24026 17552 24032 17564
rect 24084 17592 24090 17604
rect 24305 17595 24363 17601
rect 24305 17592 24317 17595
rect 24084 17564 24317 17592
rect 24084 17552 24090 17564
rect 24305 17561 24317 17564
rect 24351 17561 24363 17595
rect 24305 17555 24363 17561
rect 24670 17552 24676 17604
rect 24728 17592 24734 17604
rect 24872 17592 24900 17623
rect 26602 17620 26608 17632
rect 26660 17620 26666 17672
rect 27706 17620 27712 17672
rect 27764 17660 27770 17672
rect 27985 17663 28043 17669
rect 27985 17660 27997 17663
rect 27764 17632 27997 17660
rect 27764 17620 27770 17632
rect 27985 17629 27997 17632
rect 28031 17629 28043 17663
rect 28442 17660 28448 17672
rect 28403 17632 28448 17660
rect 27985 17623 28043 17629
rect 28442 17620 28448 17632
rect 28500 17620 28506 17672
rect 32030 17620 32036 17672
rect 32088 17660 32094 17672
rect 32125 17663 32183 17669
rect 32125 17660 32137 17663
rect 32088 17632 32137 17660
rect 32088 17620 32094 17632
rect 32125 17629 32137 17632
rect 32171 17629 32183 17663
rect 32125 17623 32183 17629
rect 24728 17564 24900 17592
rect 24728 17552 24734 17564
rect 30282 17552 30288 17604
rect 30340 17592 30346 17604
rect 30745 17595 30803 17601
rect 30745 17592 30757 17595
rect 30340 17564 30757 17592
rect 30340 17552 30346 17564
rect 30745 17561 30757 17564
rect 30791 17592 30803 17595
rect 31662 17592 31668 17604
rect 30791 17564 31668 17592
rect 30791 17561 30803 17564
rect 30745 17555 30803 17561
rect 31662 17552 31668 17564
rect 31720 17552 31726 17604
rect 35618 17592 35624 17604
rect 35579 17564 35624 17592
rect 35618 17552 35624 17564
rect 35676 17552 35682 17604
rect 8294 17484 8300 17536
rect 8352 17524 8358 17536
rect 8389 17527 8447 17533
rect 8389 17524 8401 17527
rect 8352 17496 8401 17524
rect 8352 17484 8358 17496
rect 8389 17493 8401 17496
rect 8435 17493 8447 17527
rect 16206 17524 16212 17536
rect 16167 17496 16212 17524
rect 8389 17487 8447 17493
rect 16206 17484 16212 17496
rect 16264 17484 16270 17536
rect 18414 17524 18420 17536
rect 18375 17496 18420 17524
rect 18414 17484 18420 17496
rect 18472 17484 18478 17536
rect 21177 17527 21235 17533
rect 21177 17493 21189 17527
rect 21223 17524 21235 17527
rect 21269 17527 21327 17533
rect 21269 17524 21281 17527
rect 21223 17496 21281 17524
rect 21223 17493 21235 17496
rect 21177 17487 21235 17493
rect 21269 17493 21281 17496
rect 21315 17524 21327 17527
rect 21450 17524 21456 17536
rect 21315 17496 21456 17524
rect 21315 17493 21327 17496
rect 21269 17487 21327 17493
rect 21450 17484 21456 17496
rect 21508 17484 21514 17536
rect 24118 17524 24124 17536
rect 24079 17496 24124 17524
rect 24118 17484 24124 17496
rect 24176 17484 24182 17536
rect 29822 17524 29828 17536
rect 29783 17496 29828 17524
rect 29822 17484 29828 17496
rect 29880 17524 29886 17536
rect 30377 17527 30435 17533
rect 30377 17524 30389 17527
rect 29880 17496 30389 17524
rect 29880 17484 29886 17496
rect 30377 17493 30389 17496
rect 30423 17493 30435 17527
rect 30377 17487 30435 17493
rect 1104 17434 38824 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 38824 17434
rect 1104 17360 38824 17382
rect 16206 17280 16212 17332
rect 16264 17320 16270 17332
rect 16853 17323 16911 17329
rect 16853 17320 16865 17323
rect 16264 17292 16865 17320
rect 16264 17280 16270 17292
rect 16853 17289 16865 17292
rect 16899 17289 16911 17323
rect 16853 17283 16911 17289
rect 19426 17280 19432 17332
rect 19484 17320 19490 17332
rect 19797 17323 19855 17329
rect 19797 17320 19809 17323
rect 19484 17292 19809 17320
rect 19484 17280 19490 17292
rect 19797 17289 19809 17292
rect 19843 17289 19855 17323
rect 19797 17283 19855 17289
rect 21726 17280 21732 17332
rect 21784 17320 21790 17332
rect 22005 17323 22063 17329
rect 22005 17320 22017 17323
rect 21784 17292 22017 17320
rect 21784 17280 21790 17292
rect 22005 17289 22017 17292
rect 22051 17320 22063 17323
rect 22186 17320 22192 17332
rect 22051 17292 22192 17320
rect 22051 17289 22063 17292
rect 22005 17283 22063 17289
rect 22186 17280 22192 17292
rect 22244 17280 22250 17332
rect 23474 17280 23480 17332
rect 23532 17320 23538 17332
rect 23661 17323 23719 17329
rect 23661 17320 23673 17323
rect 23532 17292 23673 17320
rect 23532 17280 23538 17292
rect 23661 17289 23673 17292
rect 23707 17289 23719 17323
rect 23661 17283 23719 17289
rect 24762 17280 24768 17332
rect 24820 17320 24826 17332
rect 24949 17323 25007 17329
rect 24949 17320 24961 17323
rect 24820 17292 24961 17320
rect 24820 17280 24826 17292
rect 24949 17289 24961 17292
rect 24995 17320 25007 17323
rect 25130 17320 25136 17332
rect 24995 17292 25136 17320
rect 24995 17289 25007 17292
rect 24949 17283 25007 17289
rect 25130 17280 25136 17292
rect 25188 17320 25194 17332
rect 26973 17323 27031 17329
rect 26973 17320 26985 17323
rect 25188 17292 26985 17320
rect 25188 17280 25194 17292
rect 26973 17289 26985 17292
rect 27019 17289 27031 17323
rect 26973 17283 27031 17289
rect 28445 17323 28503 17329
rect 28445 17289 28457 17323
rect 28491 17320 28503 17323
rect 28534 17320 28540 17332
rect 28491 17292 28540 17320
rect 28491 17289 28503 17292
rect 28445 17283 28503 17289
rect 28534 17280 28540 17292
rect 28592 17280 28598 17332
rect 32122 17320 32128 17332
rect 32083 17292 32128 17320
rect 32122 17280 32128 17292
rect 32180 17320 32186 17332
rect 33045 17323 33103 17329
rect 33045 17320 33057 17323
rect 32180 17292 33057 17320
rect 32180 17280 32186 17292
rect 33045 17289 33057 17292
rect 33091 17289 33103 17323
rect 33045 17283 33103 17289
rect 18049 17255 18107 17261
rect 18049 17221 18061 17255
rect 18095 17252 18107 17255
rect 18966 17252 18972 17264
rect 18095 17224 18972 17252
rect 18095 17221 18107 17224
rect 18049 17215 18107 17221
rect 18966 17212 18972 17224
rect 19024 17252 19030 17264
rect 19061 17255 19119 17261
rect 19061 17252 19073 17255
rect 19024 17224 19073 17252
rect 19024 17212 19030 17224
rect 19061 17221 19073 17224
rect 19107 17221 19119 17255
rect 19061 17215 19119 17221
rect 23385 17255 23443 17261
rect 23385 17221 23397 17255
rect 23431 17252 23443 17255
rect 24780 17252 24808 17280
rect 25406 17252 25412 17264
rect 23431 17224 24808 17252
rect 25367 17224 25412 17252
rect 23431 17221 23443 17224
rect 23385 17215 23443 17221
rect 25406 17212 25412 17224
rect 25464 17252 25470 17264
rect 25464 17224 25636 17252
rect 25464 17212 25470 17224
rect 18690 17184 18696 17196
rect 18651 17156 18696 17184
rect 18690 17144 18696 17156
rect 18748 17144 18754 17196
rect 21450 17184 21456 17196
rect 21411 17156 21456 17184
rect 21450 17144 21456 17156
rect 21508 17144 21514 17196
rect 21542 17144 21548 17196
rect 21600 17184 21606 17196
rect 21600 17156 21645 17184
rect 21600 17144 21606 17156
rect 24026 17144 24032 17196
rect 24084 17184 24090 17196
rect 25608 17193 25636 17224
rect 27982 17212 27988 17264
rect 28040 17252 28046 17264
rect 30009 17255 30067 17261
rect 30009 17252 30021 17255
rect 28040 17224 30021 17252
rect 28040 17212 28046 17224
rect 30009 17221 30021 17224
rect 30055 17252 30067 17255
rect 30101 17255 30159 17261
rect 30101 17252 30113 17255
rect 30055 17224 30113 17252
rect 30055 17221 30067 17224
rect 30009 17215 30067 17221
rect 30101 17221 30113 17224
rect 30147 17221 30159 17255
rect 33060 17252 33088 17283
rect 33134 17280 33140 17332
rect 33192 17320 33198 17332
rect 33229 17323 33287 17329
rect 33229 17320 33241 17323
rect 33192 17292 33241 17320
rect 33192 17280 33198 17292
rect 33229 17289 33241 17292
rect 33275 17289 33287 17323
rect 35434 17320 35440 17332
rect 35395 17292 35440 17320
rect 33229 17283 33287 17289
rect 35434 17280 35440 17292
rect 35492 17280 35498 17332
rect 33060 17224 33732 17252
rect 30101 17215 30159 17221
rect 24121 17187 24179 17193
rect 24121 17184 24133 17187
rect 24084 17156 24133 17184
rect 24084 17144 24090 17156
rect 24121 17153 24133 17156
rect 24167 17153 24179 17187
rect 24121 17147 24179 17153
rect 24213 17187 24271 17193
rect 24213 17153 24225 17187
rect 24259 17153 24271 17187
rect 24213 17147 24271 17153
rect 25593 17187 25651 17193
rect 25593 17153 25605 17187
rect 25639 17153 25651 17187
rect 25593 17147 25651 17153
rect 29825 17187 29883 17193
rect 29825 17153 29837 17187
rect 29871 17184 29883 17187
rect 30745 17187 30803 17193
rect 30745 17184 30757 17187
rect 29871 17156 30757 17184
rect 29871 17153 29883 17156
rect 29825 17147 29883 17153
rect 30745 17153 30757 17156
rect 30791 17184 30803 17187
rect 33410 17184 33416 17196
rect 30791 17156 33416 17184
rect 30791 17153 30803 17156
rect 30745 17147 30803 17153
rect 8205 17119 8263 17125
rect 8205 17085 8217 17119
rect 8251 17116 8263 17119
rect 8389 17119 8447 17125
rect 8389 17116 8401 17119
rect 8251 17088 8401 17116
rect 8251 17085 8263 17088
rect 8205 17079 8263 17085
rect 8389 17085 8401 17088
rect 8435 17116 8447 17119
rect 8478 17116 8484 17128
rect 8435 17088 8484 17116
rect 8435 17085 8447 17088
rect 8389 17079 8447 17085
rect 8478 17076 8484 17088
rect 8536 17076 8542 17128
rect 15381 17119 15439 17125
rect 15381 17085 15393 17119
rect 15427 17116 15439 17119
rect 15470 17116 15476 17128
rect 15427 17088 15476 17116
rect 15427 17085 15439 17088
rect 15381 17079 15439 17085
rect 15470 17076 15476 17088
rect 15528 17076 15534 17128
rect 15746 17125 15752 17128
rect 15740 17116 15752 17125
rect 15707 17088 15752 17116
rect 15740 17079 15752 17088
rect 15746 17076 15752 17079
rect 15804 17076 15810 17128
rect 19613 17119 19671 17125
rect 19613 17085 19625 17119
rect 19659 17116 19671 17119
rect 19886 17116 19892 17128
rect 19659 17088 19892 17116
rect 19659 17085 19671 17088
rect 19613 17079 19671 17085
rect 19886 17076 19892 17088
rect 19944 17116 19950 17128
rect 20165 17119 20223 17125
rect 20165 17116 20177 17119
rect 19944 17088 20177 17116
rect 19944 17076 19950 17088
rect 20165 17085 20177 17088
rect 20211 17085 20223 17119
rect 20165 17079 20223 17085
rect 23474 17076 23480 17128
rect 23532 17116 23538 17128
rect 24228 17116 24256 17147
rect 33410 17144 33416 17156
rect 33468 17184 33474 17196
rect 33704 17193 33732 17224
rect 35250 17212 35256 17264
rect 35308 17252 35314 17264
rect 35618 17252 35624 17264
rect 35308 17224 35624 17252
rect 35308 17212 35314 17224
rect 35618 17212 35624 17224
rect 35676 17212 35682 17264
rect 33689 17187 33747 17193
rect 33468 17156 33640 17184
rect 33468 17144 33474 17156
rect 23532 17088 24256 17116
rect 23532 17076 23538 17088
rect 29730 17076 29736 17128
rect 29788 17116 29794 17128
rect 30282 17116 30288 17128
rect 29788 17088 30288 17116
rect 29788 17076 29794 17088
rect 30282 17076 30288 17088
rect 30340 17076 30346 17128
rect 31021 17119 31079 17125
rect 31021 17116 31033 17119
rect 30392 17088 31033 17116
rect 8294 17008 8300 17060
rect 8352 17048 8358 17060
rect 8634 17051 8692 17057
rect 8634 17048 8646 17051
rect 8352 17020 8646 17048
rect 8352 17008 8358 17020
rect 8634 17017 8646 17020
rect 8680 17017 8692 17051
rect 15488 17048 15516 17076
rect 16298 17048 16304 17060
rect 15488 17020 16304 17048
rect 8634 17011 8692 17017
rect 16298 17008 16304 17020
rect 16356 17008 16362 17060
rect 16574 17008 16580 17060
rect 16632 17048 16638 17060
rect 17773 17051 17831 17057
rect 17773 17048 17785 17051
rect 16632 17020 17785 17048
rect 16632 17008 16638 17020
rect 17773 17017 17785 17020
rect 17819 17048 17831 17051
rect 18509 17051 18567 17057
rect 18509 17048 18521 17051
rect 17819 17020 18521 17048
rect 17819 17017 17831 17020
rect 17773 17011 17831 17017
rect 18509 17017 18521 17020
rect 18555 17017 18567 17051
rect 18509 17011 18567 17017
rect 23109 17051 23167 17057
rect 23109 17017 23121 17051
rect 23155 17048 23167 17051
rect 23658 17048 23664 17060
rect 23155 17020 23664 17048
rect 23155 17017 23167 17020
rect 23109 17011 23167 17017
rect 23658 17008 23664 17020
rect 23716 17048 23722 17060
rect 24029 17051 24087 17057
rect 24029 17048 24041 17051
rect 23716 17020 24041 17048
rect 23716 17008 23722 17020
rect 24029 17017 24041 17020
rect 24075 17017 24087 17051
rect 24029 17011 24087 17017
rect 25682 17008 25688 17060
rect 25740 17048 25746 17060
rect 25838 17051 25896 17057
rect 25838 17048 25850 17051
rect 25740 17020 25850 17048
rect 25740 17008 25746 17020
rect 25838 17017 25850 17020
rect 25884 17017 25896 17051
rect 25838 17011 25896 17017
rect 27614 17008 27620 17060
rect 27672 17048 27678 17060
rect 28442 17048 28448 17060
rect 27672 17020 28448 17048
rect 27672 17008 27678 17020
rect 28442 17008 28448 17020
rect 28500 17048 28506 17060
rect 28721 17051 28779 17057
rect 28721 17048 28733 17051
rect 28500 17020 28733 17048
rect 28500 17008 28506 17020
rect 28721 17017 28733 17020
rect 28767 17017 28779 17051
rect 28721 17011 28779 17017
rect 29822 17008 29828 17060
rect 29880 17048 29886 17060
rect 30392 17048 30420 17088
rect 31021 17085 31033 17088
rect 31067 17085 31079 17119
rect 31662 17116 31668 17128
rect 31575 17088 31668 17116
rect 31021 17079 31079 17085
rect 31662 17076 31668 17088
rect 31720 17116 31726 17128
rect 32214 17116 32220 17128
rect 31720 17088 32220 17116
rect 31720 17076 31726 17088
rect 32214 17076 32220 17088
rect 32272 17076 32278 17128
rect 33612 17125 33640 17156
rect 33689 17153 33701 17187
rect 33735 17153 33747 17187
rect 33870 17184 33876 17196
rect 33831 17156 33876 17184
rect 33689 17147 33747 17153
rect 33870 17144 33876 17156
rect 33928 17144 33934 17196
rect 33597 17119 33655 17125
rect 33597 17085 33609 17119
rect 33643 17116 33655 17119
rect 34241 17119 34299 17125
rect 34241 17116 34253 17119
rect 33643 17088 34253 17116
rect 33643 17085 33655 17088
rect 33597 17079 33655 17085
rect 34241 17085 34253 17088
rect 34287 17085 34299 17119
rect 34241 17079 34299 17085
rect 29880 17020 30420 17048
rect 29880 17008 29886 17020
rect 8386 16940 8392 16992
rect 8444 16980 8450 16992
rect 9769 16983 9827 16989
rect 9769 16980 9781 16983
rect 8444 16952 9781 16980
rect 8444 16940 8450 16952
rect 9769 16949 9781 16952
rect 9815 16949 9827 16983
rect 9769 16943 9827 16949
rect 15378 16940 15384 16992
rect 15436 16980 15442 16992
rect 16758 16980 16764 16992
rect 15436 16952 16764 16980
rect 15436 16940 15442 16952
rect 16758 16940 16764 16952
rect 16816 16980 16822 16992
rect 17405 16983 17463 16989
rect 17405 16980 17417 16983
rect 16816 16952 17417 16980
rect 16816 16940 16822 16952
rect 17405 16949 17417 16952
rect 17451 16980 17463 16983
rect 18230 16980 18236 16992
rect 17451 16952 18236 16980
rect 17451 16949 17463 16952
rect 17405 16943 17463 16949
rect 18230 16940 18236 16952
rect 18288 16940 18294 16992
rect 18414 16980 18420 16992
rect 18375 16952 18420 16980
rect 18414 16940 18420 16952
rect 18472 16940 18478 16992
rect 20714 16940 20720 16992
rect 20772 16980 20778 16992
rect 20809 16983 20867 16989
rect 20809 16980 20821 16983
rect 20772 16952 20821 16980
rect 20772 16940 20778 16952
rect 20809 16949 20821 16952
rect 20855 16949 20867 16983
rect 20990 16980 20996 16992
rect 20951 16952 20996 16980
rect 20809 16943 20867 16949
rect 20990 16940 20996 16952
rect 21048 16940 21054 16992
rect 21266 16940 21272 16992
rect 21324 16980 21330 16992
rect 21361 16983 21419 16989
rect 21361 16980 21373 16983
rect 21324 16952 21373 16980
rect 21324 16940 21330 16952
rect 21361 16949 21373 16952
rect 21407 16980 21419 16983
rect 22373 16983 22431 16989
rect 22373 16980 22385 16983
rect 21407 16952 22385 16980
rect 21407 16949 21419 16952
rect 21361 16943 21419 16949
rect 22373 16949 22385 16952
rect 22419 16949 22431 16983
rect 27706 16980 27712 16992
rect 27667 16952 27712 16980
rect 22373 16943 22431 16949
rect 27706 16940 27712 16952
rect 27764 16940 27770 16992
rect 27982 16980 27988 16992
rect 27943 16952 27988 16980
rect 27982 16940 27988 16952
rect 28040 16940 28046 16992
rect 30009 16983 30067 16989
rect 30009 16949 30021 16983
rect 30055 16980 30067 16983
rect 30747 16983 30805 16989
rect 30747 16980 30759 16983
rect 30055 16952 30759 16980
rect 30055 16949 30067 16952
rect 30009 16943 30067 16949
rect 30747 16949 30759 16952
rect 30793 16980 30805 16983
rect 31680 16980 31708 17076
rect 30793 16952 31708 16980
rect 30793 16949 30805 16952
rect 30747 16943 30805 16949
rect 32122 16940 32128 16992
rect 32180 16980 32186 16992
rect 32769 16983 32827 16989
rect 32769 16980 32781 16983
rect 32180 16952 32781 16980
rect 32180 16940 32186 16952
rect 32769 16949 32781 16952
rect 32815 16980 32827 16983
rect 33042 16980 33048 16992
rect 32815 16952 33048 16980
rect 32815 16949 32827 16952
rect 32769 16943 32827 16949
rect 33042 16940 33048 16952
rect 33100 16940 33106 16992
rect 1104 16890 38824 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 38824 16890
rect 1104 16816 38824 16838
rect 5442 16776 5448 16788
rect 5403 16748 5448 16776
rect 5442 16736 5448 16748
rect 5500 16736 5506 16788
rect 8021 16779 8079 16785
rect 8021 16745 8033 16779
rect 8067 16776 8079 16779
rect 8110 16776 8116 16788
rect 8067 16748 8116 16776
rect 8067 16745 8079 16748
rect 8021 16739 8079 16745
rect 8110 16736 8116 16748
rect 8168 16736 8174 16788
rect 8386 16776 8392 16788
rect 8220 16748 8392 16776
rect 5905 16711 5963 16717
rect 5905 16677 5917 16711
rect 5951 16708 5963 16711
rect 5994 16708 6000 16720
rect 5951 16680 6000 16708
rect 5951 16677 5963 16680
rect 5905 16671 5963 16677
rect 5994 16668 6000 16680
rect 6052 16668 6058 16720
rect 7926 16708 7932 16720
rect 7839 16680 7932 16708
rect 7926 16668 7932 16680
rect 7984 16708 7990 16720
rect 8220 16708 8248 16748
rect 8386 16736 8392 16748
rect 8444 16736 8450 16788
rect 11054 16776 11060 16788
rect 11015 16748 11060 16776
rect 11054 16736 11060 16748
rect 11112 16736 11118 16788
rect 15286 16776 15292 16788
rect 15247 16748 15292 16776
rect 15286 16736 15292 16748
rect 15344 16736 15350 16788
rect 15657 16779 15715 16785
rect 15657 16745 15669 16779
rect 15703 16776 15715 16779
rect 15746 16776 15752 16788
rect 15703 16748 15752 16776
rect 15703 16745 15715 16748
rect 15657 16739 15715 16745
rect 15746 16736 15752 16748
rect 15804 16736 15810 16788
rect 16298 16736 16304 16788
rect 16356 16776 16362 16788
rect 16485 16779 16543 16785
rect 16485 16776 16497 16779
rect 16356 16748 16497 16776
rect 16356 16736 16362 16748
rect 16485 16745 16497 16748
rect 16531 16776 16543 16779
rect 16850 16776 16856 16788
rect 16531 16748 16856 16776
rect 16531 16745 16543 16748
rect 16485 16739 16543 16745
rect 16850 16736 16856 16748
rect 16908 16736 16914 16788
rect 18230 16776 18236 16788
rect 18191 16748 18236 16776
rect 18230 16736 18236 16748
rect 18288 16736 18294 16788
rect 20990 16736 20996 16788
rect 21048 16776 21054 16788
rect 22830 16776 22836 16788
rect 21048 16748 22836 16776
rect 21048 16736 21054 16748
rect 22830 16736 22836 16748
rect 22888 16776 22894 16788
rect 23017 16779 23075 16785
rect 23017 16776 23029 16779
rect 22888 16748 23029 16776
rect 22888 16736 22894 16748
rect 23017 16745 23029 16748
rect 23063 16745 23075 16779
rect 23474 16776 23480 16788
rect 23435 16748 23480 16776
rect 23017 16739 23075 16745
rect 23474 16736 23480 16748
rect 23532 16736 23538 16788
rect 25682 16776 25688 16788
rect 25643 16748 25688 16776
rect 25682 16736 25688 16748
rect 25740 16736 25746 16788
rect 27338 16736 27344 16788
rect 27396 16776 27402 16788
rect 27893 16779 27951 16785
rect 27893 16776 27905 16779
rect 27396 16748 27905 16776
rect 27396 16736 27402 16748
rect 27893 16745 27905 16748
rect 27939 16745 27951 16779
rect 29362 16776 29368 16788
rect 29323 16748 29368 16776
rect 27893 16739 27951 16745
rect 29362 16736 29368 16748
rect 29420 16736 29426 16788
rect 30929 16779 30987 16785
rect 30929 16745 30941 16779
rect 30975 16745 30987 16779
rect 30929 16739 30987 16745
rect 7984 16680 8248 16708
rect 7984 16668 7990 16680
rect 8294 16668 8300 16720
rect 8352 16708 8358 16720
rect 8481 16711 8539 16717
rect 8481 16708 8493 16711
rect 8352 16680 8493 16708
rect 8352 16668 8358 16680
rect 8481 16677 8493 16680
rect 8527 16708 8539 16711
rect 9582 16708 9588 16720
rect 8527 16680 9588 16708
rect 8527 16677 8539 16680
rect 8481 16671 8539 16677
rect 9582 16668 9588 16680
rect 9640 16668 9646 16720
rect 20714 16668 20720 16720
rect 20772 16708 20778 16720
rect 21330 16711 21388 16717
rect 21330 16708 21342 16711
rect 20772 16680 21342 16708
rect 20772 16668 20778 16680
rect 21330 16677 21342 16680
rect 21376 16677 21388 16711
rect 24394 16708 24400 16720
rect 21330 16671 21388 16677
rect 23584 16680 24400 16708
rect 5813 16643 5871 16649
rect 5813 16609 5825 16643
rect 5859 16640 5871 16643
rect 6270 16640 6276 16652
rect 5859 16612 6276 16640
rect 5859 16609 5871 16612
rect 5813 16603 5871 16609
rect 6270 16600 6276 16612
rect 6328 16600 6334 16652
rect 9766 16600 9772 16652
rect 9824 16640 9830 16652
rect 9944 16643 10002 16649
rect 9944 16640 9956 16643
rect 9824 16612 9956 16640
rect 9824 16600 9830 16612
rect 9944 16609 9956 16612
rect 9990 16640 10002 16643
rect 10962 16640 10968 16652
rect 9990 16612 10968 16640
rect 9990 16609 10002 16612
rect 9944 16603 10002 16609
rect 10962 16600 10968 16612
rect 11020 16600 11026 16652
rect 16758 16600 16764 16652
rect 16816 16640 16822 16652
rect 17109 16643 17167 16649
rect 17109 16640 17121 16643
rect 16816 16612 17121 16640
rect 16816 16600 16822 16612
rect 17109 16609 17121 16612
rect 17155 16609 17167 16643
rect 17109 16603 17167 16609
rect 20625 16643 20683 16649
rect 20625 16609 20637 16643
rect 20671 16640 20683 16643
rect 20806 16640 20812 16652
rect 20671 16612 20812 16640
rect 20671 16609 20683 16612
rect 20625 16603 20683 16609
rect 20806 16600 20812 16612
rect 20864 16640 20870 16652
rect 21910 16640 21916 16652
rect 20864 16612 21916 16640
rect 20864 16600 20870 16612
rect 21910 16600 21916 16612
rect 21968 16600 21974 16652
rect 23584 16649 23612 16680
rect 24394 16668 24400 16680
rect 24452 16708 24458 16720
rect 25406 16708 25412 16720
rect 24452 16680 25412 16708
rect 24452 16668 24458 16680
rect 25406 16668 25412 16680
rect 25464 16668 25470 16720
rect 29816 16711 29874 16717
rect 29816 16677 29828 16711
rect 29862 16708 29874 16711
rect 29914 16708 29920 16720
rect 29862 16680 29920 16708
rect 29862 16677 29874 16680
rect 29816 16671 29874 16677
rect 29914 16668 29920 16680
rect 29972 16668 29978 16720
rect 30282 16668 30288 16720
rect 30340 16708 30346 16720
rect 30944 16708 30972 16739
rect 31110 16736 31116 16788
rect 31168 16776 31174 16788
rect 31481 16779 31539 16785
rect 31481 16776 31493 16779
rect 31168 16748 31493 16776
rect 31168 16736 31174 16748
rect 31481 16745 31493 16748
rect 31527 16776 31539 16779
rect 31665 16779 31723 16785
rect 31665 16776 31677 16779
rect 31527 16748 31677 16776
rect 31527 16745 31539 16748
rect 31481 16739 31539 16745
rect 31665 16745 31677 16748
rect 31711 16745 31723 16779
rect 31665 16739 31723 16745
rect 31941 16779 31999 16785
rect 31941 16745 31953 16779
rect 31987 16776 31999 16779
rect 32306 16776 32312 16788
rect 31987 16748 32312 16776
rect 31987 16745 31999 16748
rect 31941 16739 31999 16745
rect 32306 16736 32312 16748
rect 32364 16776 32370 16788
rect 33870 16776 33876 16788
rect 32364 16748 33876 16776
rect 32364 16736 32370 16748
rect 33870 16736 33876 16748
rect 33928 16776 33934 16788
rect 34057 16779 34115 16785
rect 34057 16776 34069 16779
rect 33928 16748 34069 16776
rect 33928 16736 33934 16748
rect 34057 16745 34069 16748
rect 34103 16745 34115 16779
rect 34057 16739 34115 16745
rect 30340 16680 32352 16708
rect 30340 16668 30346 16680
rect 23569 16643 23627 16649
rect 23569 16609 23581 16643
rect 23615 16609 23627 16643
rect 23569 16603 23627 16609
rect 23836 16643 23894 16649
rect 23836 16609 23848 16643
rect 23882 16640 23894 16643
rect 24118 16640 24124 16652
rect 23882 16612 24124 16640
rect 23882 16609 23894 16612
rect 23836 16603 23894 16609
rect 24118 16600 24124 16612
rect 24176 16600 24182 16652
rect 4985 16575 5043 16581
rect 4985 16541 4997 16575
rect 5031 16572 5043 16575
rect 5258 16572 5264 16584
rect 5031 16544 5264 16572
rect 5031 16541 5043 16544
rect 4985 16535 5043 16541
rect 5258 16532 5264 16544
rect 5316 16532 5322 16584
rect 5997 16575 6055 16581
rect 5997 16572 6009 16575
rect 5368 16544 6009 16572
rect 5368 16448 5396 16544
rect 5997 16541 6009 16544
rect 6043 16541 6055 16575
rect 8573 16575 8631 16581
rect 8573 16572 8585 16575
rect 5997 16535 6055 16541
rect 7484 16544 8585 16572
rect 7484 16448 7512 16544
rect 8573 16541 8585 16544
rect 8619 16541 8631 16575
rect 9674 16572 9680 16584
rect 9587 16544 9680 16572
rect 8573 16535 8631 16541
rect 9674 16532 9680 16544
rect 9732 16532 9738 16584
rect 15378 16532 15384 16584
rect 15436 16572 15442 16584
rect 15749 16575 15807 16581
rect 15749 16572 15761 16575
rect 15436 16544 15761 16572
rect 15436 16532 15442 16544
rect 15749 16541 15761 16544
rect 15795 16541 15807 16575
rect 15749 16535 15807 16541
rect 15933 16575 15991 16581
rect 15933 16541 15945 16575
rect 15979 16572 15991 16575
rect 16114 16572 16120 16584
rect 15979 16544 16120 16572
rect 15979 16541 15991 16544
rect 15933 16535 15991 16541
rect 16114 16532 16120 16544
rect 16172 16572 16178 16584
rect 16666 16572 16672 16584
rect 16172 16544 16672 16572
rect 16172 16532 16178 16544
rect 16666 16532 16672 16544
rect 16724 16572 16730 16584
rect 16724 16544 16804 16572
rect 16724 16532 16730 16544
rect 8478 16464 8484 16516
rect 8536 16504 8542 16516
rect 9692 16504 9720 16532
rect 8536 16476 9720 16504
rect 8536 16464 8542 16476
rect 5350 16436 5356 16448
rect 5311 16408 5356 16436
rect 5350 16396 5356 16408
rect 5408 16396 5414 16448
rect 7190 16436 7196 16448
rect 7151 16408 7196 16436
rect 7190 16396 7196 16408
rect 7248 16396 7254 16448
rect 7466 16436 7472 16448
rect 7427 16408 7472 16436
rect 7466 16396 7472 16408
rect 7524 16396 7530 16448
rect 16776 16436 16804 16544
rect 16850 16532 16856 16584
rect 16908 16572 16914 16584
rect 21082 16572 21088 16584
rect 16908 16544 16953 16572
rect 21043 16544 21088 16572
rect 16908 16532 16914 16544
rect 21082 16532 21088 16544
rect 21140 16532 21146 16584
rect 25424 16572 25452 16668
rect 26326 16600 26332 16652
rect 26384 16640 26390 16652
rect 26769 16643 26827 16649
rect 26769 16640 26781 16643
rect 26384 16612 26781 16640
rect 26384 16600 26390 16612
rect 26769 16609 26781 16612
rect 26815 16640 26827 16643
rect 27246 16640 27252 16652
rect 26815 16612 27252 16640
rect 26815 16609 26827 16612
rect 26769 16603 26827 16609
rect 27246 16600 27252 16612
rect 27304 16600 27310 16652
rect 29546 16640 29552 16652
rect 29507 16612 29552 16640
rect 29546 16600 29552 16612
rect 29604 16640 29610 16652
rect 30374 16640 30380 16652
rect 29604 16612 30380 16640
rect 29604 16600 29610 16612
rect 30374 16600 30380 16612
rect 30432 16600 30438 16652
rect 32122 16640 32128 16652
rect 31588 16612 32128 16640
rect 26510 16572 26516 16584
rect 25424 16544 26516 16572
rect 26510 16532 26516 16544
rect 26568 16532 26574 16584
rect 30926 16532 30932 16584
rect 30984 16572 30990 16584
rect 31588 16572 31616 16612
rect 32122 16600 32128 16612
rect 32180 16600 32186 16652
rect 32324 16640 32352 16680
rect 32392 16643 32450 16649
rect 32392 16640 32404 16643
rect 32324 16612 32404 16640
rect 32392 16609 32404 16612
rect 32438 16640 32450 16643
rect 32438 16612 33180 16640
rect 32438 16609 32450 16612
rect 32392 16603 32450 16609
rect 30984 16544 31616 16572
rect 33152 16572 33180 16612
rect 33226 16572 33232 16584
rect 33152 16544 33232 16572
rect 30984 16532 30990 16544
rect 33226 16532 33232 16544
rect 33284 16532 33290 16584
rect 17034 16436 17040 16448
rect 16776 16408 17040 16436
rect 17034 16396 17040 16408
rect 17092 16396 17098 16448
rect 18782 16436 18788 16448
rect 18743 16408 18788 16436
rect 18782 16396 18788 16408
rect 18840 16396 18846 16448
rect 22094 16396 22100 16448
rect 22152 16436 22158 16448
rect 22465 16439 22523 16445
rect 22465 16436 22477 16439
rect 22152 16408 22477 16436
rect 22152 16396 22158 16408
rect 22465 16405 22477 16408
rect 22511 16405 22523 16439
rect 22465 16399 22523 16405
rect 24762 16396 24768 16448
rect 24820 16436 24826 16448
rect 24949 16439 25007 16445
rect 24949 16436 24961 16439
rect 24820 16408 24961 16436
rect 24820 16396 24826 16408
rect 24949 16405 24961 16408
rect 24995 16405 25007 16439
rect 24949 16399 25007 16405
rect 31665 16439 31723 16445
rect 31665 16405 31677 16439
rect 31711 16436 31723 16439
rect 33505 16439 33563 16445
rect 33505 16436 33517 16439
rect 31711 16408 33517 16436
rect 31711 16405 31723 16408
rect 31665 16399 31723 16405
rect 33505 16405 33517 16408
rect 33551 16405 33563 16439
rect 33505 16399 33563 16405
rect 1104 16346 38824 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 38824 16346
rect 1104 16272 38824 16294
rect 4893 16235 4951 16241
rect 4893 16201 4905 16235
rect 4939 16232 4951 16235
rect 5442 16232 5448 16244
rect 4939 16204 5448 16232
rect 4939 16201 4951 16204
rect 4893 16195 4951 16201
rect 5442 16192 5448 16204
rect 5500 16192 5506 16244
rect 8478 16232 8484 16244
rect 8439 16204 8484 16232
rect 8478 16192 8484 16204
rect 8536 16192 8542 16244
rect 9674 16192 9680 16244
rect 9732 16232 9738 16244
rect 10045 16235 10103 16241
rect 10045 16232 10057 16235
rect 9732 16204 10057 16232
rect 9732 16192 9738 16204
rect 10045 16201 10057 16204
rect 10091 16201 10103 16235
rect 10045 16195 10103 16201
rect 10689 16235 10747 16241
rect 10689 16201 10701 16235
rect 10735 16232 10747 16235
rect 10962 16232 10968 16244
rect 10735 16204 10968 16232
rect 10735 16201 10747 16204
rect 10689 16195 10747 16201
rect 10962 16192 10968 16204
rect 11020 16192 11026 16244
rect 15378 16232 15384 16244
rect 15339 16204 15384 16232
rect 15378 16192 15384 16204
rect 15436 16192 15442 16244
rect 15746 16232 15752 16244
rect 15707 16204 15752 16232
rect 15746 16192 15752 16204
rect 15804 16192 15810 16244
rect 16393 16235 16451 16241
rect 16393 16201 16405 16235
rect 16439 16232 16451 16235
rect 16482 16232 16488 16244
rect 16439 16204 16488 16232
rect 16439 16201 16451 16204
rect 16393 16195 16451 16201
rect 16482 16192 16488 16204
rect 16540 16192 16546 16244
rect 17681 16235 17739 16241
rect 17681 16201 17693 16235
rect 17727 16232 17739 16235
rect 18046 16232 18052 16244
rect 17727 16204 18052 16232
rect 17727 16201 17739 16204
rect 17681 16195 17739 16201
rect 18046 16192 18052 16204
rect 18104 16192 18110 16244
rect 20625 16235 20683 16241
rect 20625 16201 20637 16235
rect 20671 16232 20683 16235
rect 20901 16235 20959 16241
rect 20901 16232 20913 16235
rect 20671 16204 20913 16232
rect 20671 16201 20683 16204
rect 20625 16195 20683 16201
rect 20901 16201 20913 16204
rect 20947 16232 20959 16235
rect 21082 16232 21088 16244
rect 20947 16204 21088 16232
rect 20947 16201 20959 16204
rect 20901 16195 20959 16201
rect 21082 16192 21088 16204
rect 21140 16192 21146 16244
rect 22186 16192 22192 16244
rect 22244 16232 22250 16244
rect 22465 16235 22523 16241
rect 22465 16232 22477 16235
rect 22244 16204 22477 16232
rect 22244 16192 22250 16204
rect 22465 16201 22477 16204
rect 22511 16201 22523 16235
rect 22465 16195 22523 16201
rect 23474 16192 23480 16244
rect 23532 16232 23538 16244
rect 23937 16235 23995 16241
rect 23937 16232 23949 16235
rect 23532 16204 23949 16232
rect 23532 16192 23538 16204
rect 23937 16201 23949 16204
rect 23983 16201 23995 16235
rect 24394 16232 24400 16244
rect 24355 16204 24400 16232
rect 23937 16195 23995 16201
rect 24394 16192 24400 16204
rect 24452 16232 24458 16244
rect 24673 16235 24731 16241
rect 24673 16232 24685 16235
rect 24452 16204 24685 16232
rect 24452 16192 24458 16204
rect 24673 16201 24685 16204
rect 24719 16201 24731 16235
rect 26234 16232 26240 16244
rect 26195 16204 26240 16232
rect 24673 16195 24731 16201
rect 7466 16164 7472 16176
rect 6656 16136 7472 16164
rect 6656 16108 6684 16136
rect 7466 16124 7472 16136
rect 7524 16164 7530 16176
rect 15013 16167 15071 16173
rect 7524 16136 7696 16164
rect 7524 16124 7530 16136
rect 4433 16099 4491 16105
rect 4433 16065 4445 16099
rect 4479 16096 4491 16099
rect 5350 16096 5356 16108
rect 4479 16068 5356 16096
rect 4479 16065 4491 16068
rect 4433 16059 4491 16065
rect 5350 16056 5356 16068
rect 5408 16096 5414 16108
rect 5537 16099 5595 16105
rect 5537 16096 5549 16099
rect 5408 16068 5549 16096
rect 5408 16056 5414 16068
rect 5537 16065 5549 16068
rect 5583 16096 5595 16099
rect 6638 16096 6644 16108
rect 5583 16068 6644 16096
rect 5583 16065 5595 16068
rect 5537 16059 5595 16065
rect 6638 16056 6644 16068
rect 6696 16056 6702 16108
rect 7558 16096 7564 16108
rect 7519 16068 7564 16096
rect 7558 16056 7564 16068
rect 7616 16056 7622 16108
rect 7668 16105 7696 16136
rect 15013 16133 15025 16167
rect 15059 16164 15071 16167
rect 16114 16164 16120 16176
rect 15059 16136 16120 16164
rect 15059 16133 15071 16136
rect 15013 16127 15071 16133
rect 16114 16124 16120 16136
rect 16172 16124 16178 16176
rect 7653 16099 7711 16105
rect 7653 16065 7665 16099
rect 7699 16065 7711 16099
rect 7653 16059 7711 16065
rect 8205 16099 8263 16105
rect 8205 16065 8217 16099
rect 8251 16096 8263 16099
rect 17034 16096 17040 16108
rect 8251 16068 8800 16096
rect 16995 16068 17040 16096
rect 8251 16065 8263 16068
rect 8205 16059 8263 16065
rect 7190 15988 7196 16040
rect 7248 16028 7254 16040
rect 7469 16031 7527 16037
rect 7469 16028 7481 16031
rect 7248 16000 7481 16028
rect 7248 15988 7254 16000
rect 7469 15997 7481 16000
rect 7515 16028 7527 16031
rect 8220 16028 8248 16059
rect 7515 16000 8248 16028
rect 7515 15997 7527 16000
rect 7469 15991 7527 15997
rect 8478 15988 8484 16040
rect 8536 16028 8542 16040
rect 8665 16031 8723 16037
rect 8665 16028 8677 16031
rect 8536 16000 8677 16028
rect 8536 15988 8542 16000
rect 8665 15997 8677 16000
rect 8711 15997 8723 16031
rect 8772 16028 8800 16068
rect 17034 16056 17040 16068
rect 17092 16056 17098 16108
rect 18064 16105 18092 16192
rect 21100 16105 21128 16192
rect 18049 16099 18107 16105
rect 18049 16065 18061 16099
rect 18095 16065 18107 16099
rect 18049 16059 18107 16065
rect 21085 16099 21143 16105
rect 21085 16065 21097 16099
rect 21131 16065 21143 16099
rect 24688 16096 24716 16195
rect 26234 16192 26240 16204
rect 26292 16192 26298 16244
rect 26602 16192 26608 16244
rect 26660 16232 26666 16244
rect 27157 16235 27215 16241
rect 27157 16232 27169 16235
rect 26660 16204 27169 16232
rect 26660 16192 26666 16204
rect 27157 16201 27169 16204
rect 27203 16232 27215 16235
rect 29365 16235 29423 16241
rect 27203 16204 27752 16232
rect 27203 16201 27215 16204
rect 27157 16195 27215 16201
rect 26510 16124 26516 16176
rect 26568 16164 26574 16176
rect 26789 16167 26847 16173
rect 26789 16164 26801 16167
rect 26568 16136 26801 16164
rect 26568 16124 26574 16136
rect 26789 16133 26801 16136
rect 26835 16133 26847 16167
rect 26789 16127 26847 16133
rect 27341 16167 27399 16173
rect 27341 16133 27353 16167
rect 27387 16164 27399 16167
rect 27522 16164 27528 16176
rect 27387 16136 27528 16164
rect 27387 16133 27399 16136
rect 27341 16127 27399 16133
rect 27522 16124 27528 16136
rect 27580 16124 27586 16176
rect 24857 16099 24915 16105
rect 24857 16096 24869 16099
rect 24688 16068 24869 16096
rect 21085 16059 21143 16065
rect 24857 16065 24869 16068
rect 24903 16065 24915 16099
rect 24857 16059 24915 16065
rect 8932 16031 8990 16037
rect 8932 16028 8944 16031
rect 8772 16000 8944 16028
rect 8665 15991 8723 15997
rect 8932 15997 8944 16000
rect 8978 16028 8990 16031
rect 9214 16028 9220 16040
rect 8978 16000 9220 16028
rect 8978 15997 8990 16000
rect 8932 15991 8990 15997
rect 9214 15988 9220 16000
rect 9272 15988 9278 16040
rect 18316 16031 18374 16037
rect 18316 15997 18328 16031
rect 18362 16028 18374 16031
rect 18782 16028 18788 16040
rect 18362 16000 18788 16028
rect 18362 15997 18374 16000
rect 18316 15991 18374 15997
rect 18782 15988 18788 16000
rect 18840 15988 18846 16040
rect 23477 16031 23535 16037
rect 23477 15997 23489 16031
rect 23523 16028 23535 16031
rect 23750 16028 23756 16040
rect 23523 16000 23756 16028
rect 23523 15997 23535 16000
rect 23477 15991 23535 15997
rect 23750 15988 23756 16000
rect 23808 15988 23814 16040
rect 25130 16037 25136 16040
rect 25124 16028 25136 16037
rect 25091 16000 25136 16028
rect 25124 15991 25136 16000
rect 25130 15988 25136 15991
rect 25188 15988 25194 16040
rect 27724 16037 27752 16204
rect 29365 16201 29377 16235
rect 29411 16232 29423 16235
rect 30006 16232 30012 16244
rect 29411 16204 30012 16232
rect 29411 16201 29423 16204
rect 29365 16195 29423 16201
rect 30006 16192 30012 16204
rect 30064 16192 30070 16244
rect 30374 16232 30380 16244
rect 30335 16204 30380 16232
rect 30374 16192 30380 16204
rect 30432 16232 30438 16244
rect 30745 16235 30803 16241
rect 30745 16232 30757 16235
rect 30432 16204 30757 16232
rect 30432 16192 30438 16204
rect 30745 16201 30757 16204
rect 30791 16232 30803 16235
rect 32306 16232 32312 16244
rect 30791 16204 30972 16232
rect 32267 16204 32312 16232
rect 30791 16201 30803 16204
rect 30745 16195 30803 16201
rect 30944 16108 30972 16204
rect 32306 16192 32312 16204
rect 32364 16192 32370 16244
rect 33226 16232 33232 16244
rect 33187 16204 33232 16232
rect 33226 16192 33232 16204
rect 33284 16192 33290 16244
rect 27890 16096 27896 16108
rect 27851 16068 27896 16096
rect 27890 16056 27896 16068
rect 27948 16096 27954 16108
rect 28353 16099 28411 16105
rect 28353 16096 28365 16099
rect 27948 16068 28365 16096
rect 27948 16056 27954 16068
rect 28353 16065 28365 16068
rect 28399 16065 28411 16099
rect 28353 16059 28411 16065
rect 29089 16099 29147 16105
rect 29089 16065 29101 16099
rect 29135 16096 29147 16099
rect 29822 16096 29828 16108
rect 29135 16068 29828 16096
rect 29135 16065 29147 16068
rect 29089 16059 29147 16065
rect 29822 16056 29828 16068
rect 29880 16056 29886 16108
rect 30009 16099 30067 16105
rect 30009 16065 30021 16099
rect 30055 16096 30067 16099
rect 30282 16096 30288 16108
rect 30055 16068 30288 16096
rect 30055 16065 30067 16068
rect 30009 16059 30067 16065
rect 30282 16056 30288 16068
rect 30340 16056 30346 16108
rect 30926 16096 30932 16108
rect 30839 16068 30932 16096
rect 30926 16056 30932 16068
rect 30984 16056 30990 16108
rect 27709 16031 27767 16037
rect 27709 15997 27721 16031
rect 27755 15997 27767 16031
rect 27709 15991 27767 15997
rect 29362 15988 29368 16040
rect 29420 16028 29426 16040
rect 29733 16031 29791 16037
rect 29733 16028 29745 16031
rect 29420 16000 29745 16028
rect 29420 15988 29426 16000
rect 29733 15997 29745 16000
rect 29779 16028 29791 16031
rect 30190 16028 30196 16040
rect 29779 16000 30196 16028
rect 29779 15997 29791 16000
rect 29733 15991 29791 15997
rect 30190 15988 30196 16000
rect 30248 15988 30254 16040
rect 5353 15963 5411 15969
rect 5353 15960 5365 15963
rect 4816 15932 5365 15960
rect 4816 15904 4844 15932
rect 5353 15929 5365 15932
rect 5399 15929 5411 15963
rect 5353 15923 5411 15929
rect 16301 15963 16359 15969
rect 16301 15929 16313 15963
rect 16347 15960 16359 15963
rect 16853 15963 16911 15969
rect 16853 15960 16865 15963
rect 16347 15932 16865 15960
rect 16347 15929 16359 15932
rect 16301 15923 16359 15929
rect 16853 15929 16865 15932
rect 16899 15960 16911 15963
rect 17494 15960 17500 15972
rect 16899 15932 17500 15960
rect 16899 15929 16911 15932
rect 16853 15923 16911 15929
rect 17494 15920 17500 15932
rect 17552 15920 17558 15972
rect 20257 15963 20315 15969
rect 20257 15929 20269 15963
rect 20303 15960 20315 15963
rect 21330 15963 21388 15969
rect 21330 15960 21342 15963
rect 20303 15932 21342 15960
rect 20303 15929 20315 15932
rect 20257 15923 20315 15929
rect 21330 15929 21342 15932
rect 21376 15960 21388 15963
rect 22278 15960 22284 15972
rect 21376 15932 22284 15960
rect 21376 15929 21388 15932
rect 21330 15923 21388 15929
rect 22278 15920 22284 15932
rect 22336 15920 22342 15972
rect 27614 15920 27620 15972
rect 27672 15960 27678 15972
rect 27801 15963 27859 15969
rect 27801 15960 27813 15963
rect 27672 15932 27813 15960
rect 27672 15920 27678 15932
rect 27801 15929 27813 15932
rect 27847 15929 27859 15963
rect 27801 15923 27859 15929
rect 31110 15920 31116 15972
rect 31168 15969 31174 15972
rect 31168 15963 31232 15969
rect 31168 15929 31186 15963
rect 31220 15929 31232 15963
rect 31168 15923 31232 15929
rect 31168 15920 31174 15923
rect 4798 15892 4804 15904
rect 4759 15864 4804 15892
rect 4798 15852 4804 15864
rect 4856 15852 4862 15904
rect 5258 15892 5264 15904
rect 5219 15864 5264 15892
rect 5258 15852 5264 15864
rect 5316 15852 5322 15904
rect 5994 15892 6000 15904
rect 5955 15864 6000 15892
rect 5994 15852 6000 15864
rect 6052 15852 6058 15904
rect 6270 15892 6276 15904
rect 6231 15864 6276 15892
rect 6270 15852 6276 15864
rect 6328 15852 6334 15904
rect 7098 15892 7104 15904
rect 7059 15864 7104 15892
rect 7098 15852 7104 15864
rect 7156 15852 7162 15904
rect 16758 15892 16764 15904
rect 16719 15864 16764 15892
rect 16758 15852 16764 15864
rect 16816 15852 16822 15904
rect 17218 15852 17224 15904
rect 17276 15892 17282 15904
rect 17405 15895 17463 15901
rect 17405 15892 17417 15895
rect 17276 15864 17417 15892
rect 17276 15852 17282 15864
rect 17405 15861 17417 15864
rect 17451 15892 17463 15895
rect 17681 15895 17739 15901
rect 17681 15892 17693 15895
rect 17451 15864 17693 15892
rect 17451 15861 17463 15864
rect 17405 15855 17463 15861
rect 17681 15861 17693 15864
rect 17727 15892 17739 15895
rect 17773 15895 17831 15901
rect 17773 15892 17785 15895
rect 17727 15864 17785 15892
rect 17727 15861 17739 15864
rect 17681 15855 17739 15861
rect 17773 15861 17785 15864
rect 17819 15861 17831 15895
rect 19426 15892 19432 15904
rect 19387 15864 19432 15892
rect 17773 15855 17831 15861
rect 19426 15852 19432 15864
rect 19484 15852 19490 15904
rect 32953 15895 33011 15901
rect 32953 15861 32965 15895
rect 32999 15892 33011 15895
rect 33042 15892 33048 15904
rect 32999 15864 33048 15892
rect 32999 15861 33011 15864
rect 32953 15855 33011 15861
rect 33042 15852 33048 15864
rect 33100 15852 33106 15904
rect 1104 15802 38824 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 38824 15802
rect 1104 15728 38824 15750
rect 7098 15648 7104 15700
rect 7156 15688 7162 15700
rect 8018 15688 8024 15700
rect 7156 15660 8024 15688
rect 7156 15648 7162 15660
rect 8018 15648 8024 15660
rect 8076 15688 8082 15700
rect 8481 15691 8539 15697
rect 8481 15688 8493 15691
rect 8076 15660 8493 15688
rect 8076 15648 8082 15660
rect 8481 15657 8493 15660
rect 8527 15657 8539 15691
rect 8481 15651 8539 15657
rect 9766 15648 9772 15700
rect 9824 15688 9830 15700
rect 9861 15691 9919 15697
rect 9861 15688 9873 15691
rect 9824 15660 9873 15688
rect 9824 15648 9830 15660
rect 9861 15657 9873 15660
rect 9907 15657 9919 15691
rect 16114 15688 16120 15700
rect 16075 15660 16120 15688
rect 9861 15651 9919 15657
rect 16114 15648 16120 15660
rect 16172 15648 16178 15700
rect 16485 15691 16543 15697
rect 16485 15657 16497 15691
rect 16531 15688 16543 15691
rect 16758 15688 16764 15700
rect 16531 15660 16764 15688
rect 16531 15657 16543 15660
rect 16485 15651 16543 15657
rect 16758 15648 16764 15660
rect 16816 15688 16822 15700
rect 16945 15691 17003 15697
rect 16945 15688 16957 15691
rect 16816 15660 16957 15688
rect 16816 15648 16822 15660
rect 16945 15657 16957 15660
rect 16991 15688 17003 15691
rect 18601 15691 18659 15697
rect 18601 15688 18613 15691
rect 16991 15660 18613 15688
rect 16991 15657 17003 15660
rect 16945 15651 17003 15657
rect 18601 15657 18613 15660
rect 18647 15657 18659 15691
rect 20714 15688 20720 15700
rect 20675 15660 20720 15688
rect 18601 15651 18659 15657
rect 20714 15648 20720 15660
rect 20772 15688 20778 15700
rect 22465 15691 22523 15697
rect 22465 15688 22477 15691
rect 20772 15660 22477 15688
rect 20772 15648 20778 15660
rect 22465 15657 22477 15660
rect 22511 15657 22523 15691
rect 26326 15688 26332 15700
rect 26287 15660 26332 15688
rect 22465 15651 22523 15657
rect 26326 15648 26332 15660
rect 26384 15648 26390 15700
rect 27890 15688 27896 15700
rect 27851 15660 27896 15688
rect 27890 15648 27896 15660
rect 27948 15648 27954 15700
rect 30009 15691 30067 15697
rect 30009 15657 30021 15691
rect 30055 15688 30067 15691
rect 30282 15688 30288 15700
rect 30055 15660 30288 15688
rect 30055 15657 30067 15660
rect 30009 15651 30067 15657
rect 30282 15648 30288 15660
rect 30340 15648 30346 15700
rect 33410 15688 33416 15700
rect 33371 15660 33416 15688
rect 33410 15648 33416 15660
rect 33468 15648 33474 15700
rect 36538 15688 36544 15700
rect 36499 15660 36544 15688
rect 36538 15648 36544 15660
rect 36596 15648 36602 15700
rect 7193 15623 7251 15629
rect 7193 15589 7205 15623
rect 7239 15620 7251 15623
rect 7558 15620 7564 15632
rect 7239 15592 7564 15620
rect 7239 15589 7251 15592
rect 7193 15583 7251 15589
rect 7558 15580 7564 15592
rect 7616 15580 7622 15632
rect 7929 15623 7987 15629
rect 7929 15589 7941 15623
rect 7975 15620 7987 15623
rect 8202 15620 8208 15632
rect 7975 15592 8208 15620
rect 7975 15589 7987 15592
rect 7929 15583 7987 15589
rect 8202 15580 8208 15592
rect 8260 15580 8266 15632
rect 17494 15629 17500 15632
rect 17488 15620 17500 15629
rect 17455 15592 17500 15620
rect 17488 15583 17500 15592
rect 17494 15580 17500 15583
rect 17552 15580 17558 15632
rect 24394 15620 24400 15632
rect 23952 15592 24400 15620
rect 5252 15555 5310 15561
rect 5252 15521 5264 15555
rect 5298 15552 5310 15555
rect 5994 15552 6000 15564
rect 5298 15524 6000 15552
rect 5298 15521 5310 15524
rect 5252 15515 5310 15521
rect 5994 15512 6000 15524
rect 6052 15512 6058 15564
rect 8294 15512 8300 15564
rect 8352 15552 8358 15564
rect 8389 15555 8447 15561
rect 8389 15552 8401 15555
rect 8352 15524 8401 15552
rect 8352 15512 8358 15524
rect 8389 15521 8401 15524
rect 8435 15521 8447 15555
rect 8389 15515 8447 15521
rect 20714 15512 20720 15564
rect 20772 15552 20778 15564
rect 21341 15555 21399 15561
rect 21341 15552 21353 15555
rect 20772 15524 21353 15552
rect 20772 15512 20778 15524
rect 21341 15521 21353 15524
rect 21387 15552 21399 15555
rect 22186 15552 22192 15564
rect 21387 15524 22192 15552
rect 21387 15521 21399 15524
rect 21341 15515 21399 15521
rect 22186 15512 22192 15524
rect 22244 15512 22250 15564
rect 23952 15561 23980 15592
rect 24394 15580 24400 15592
rect 24452 15580 24458 15632
rect 26780 15623 26838 15629
rect 26780 15589 26792 15623
rect 26826 15620 26838 15623
rect 26970 15620 26976 15632
rect 26826 15592 26976 15620
rect 26826 15589 26838 15592
rect 26780 15583 26838 15589
rect 26970 15580 26976 15592
rect 27028 15620 27034 15632
rect 27338 15620 27344 15632
rect 27028 15592 27344 15620
rect 27028 15580 27034 15592
rect 27338 15580 27344 15592
rect 27396 15580 27402 15632
rect 23937 15555 23995 15561
rect 23937 15521 23949 15555
rect 23983 15521 23995 15555
rect 23937 15515 23995 15521
rect 24026 15512 24032 15564
rect 24084 15552 24090 15564
rect 24193 15555 24251 15561
rect 24193 15552 24205 15555
rect 24084 15524 24205 15552
rect 24084 15512 24090 15524
rect 24193 15521 24205 15524
rect 24239 15521 24251 15555
rect 26510 15552 26516 15564
rect 26471 15524 26516 15552
rect 24193 15515 24251 15521
rect 26510 15512 26516 15524
rect 26568 15512 26574 15564
rect 30558 15552 30564 15564
rect 30519 15524 30564 15552
rect 30558 15512 30564 15524
rect 30616 15512 30622 15564
rect 31297 15555 31355 15561
rect 31297 15521 31309 15555
rect 31343 15552 31355 15555
rect 31662 15552 31668 15564
rect 31343 15524 31668 15552
rect 31343 15521 31355 15524
rect 31297 15515 31355 15521
rect 31662 15512 31668 15524
rect 31720 15512 31726 15564
rect 32122 15552 32128 15564
rect 32035 15524 32128 15552
rect 32122 15512 32128 15524
rect 32180 15552 32186 15564
rect 32677 15555 32735 15561
rect 32677 15552 32689 15555
rect 32180 15524 32689 15552
rect 32180 15512 32186 15524
rect 32677 15521 32689 15524
rect 32723 15521 32735 15555
rect 33226 15552 33232 15564
rect 33187 15524 33232 15552
rect 32677 15515 32735 15521
rect 33226 15512 33232 15524
rect 33284 15512 33290 15564
rect 35069 15555 35127 15561
rect 35069 15521 35081 15555
rect 35115 15552 35127 15555
rect 35250 15552 35256 15564
rect 35115 15524 35256 15552
rect 35115 15521 35127 15524
rect 35069 15515 35127 15521
rect 35250 15512 35256 15524
rect 35308 15512 35314 15564
rect 35428 15555 35486 15561
rect 35428 15521 35440 15555
rect 35474 15552 35486 15555
rect 35894 15552 35900 15564
rect 35474 15524 35900 15552
rect 35474 15521 35486 15524
rect 35428 15515 35486 15521
rect 35894 15512 35900 15524
rect 35952 15512 35958 15564
rect 4982 15484 4988 15496
rect 4943 15456 4988 15484
rect 4982 15444 4988 15456
rect 5040 15444 5046 15496
rect 8662 15484 8668 15496
rect 8623 15456 8668 15484
rect 8662 15444 8668 15456
rect 8720 15444 8726 15496
rect 17218 15484 17224 15496
rect 17179 15456 17224 15484
rect 17218 15444 17224 15456
rect 17276 15444 17282 15496
rect 21082 15484 21088 15496
rect 21043 15456 21088 15484
rect 21082 15444 21088 15456
rect 21140 15444 21146 15496
rect 30650 15484 30656 15496
rect 30611 15456 30656 15484
rect 30650 15444 30656 15456
rect 30708 15444 30714 15496
rect 30837 15487 30895 15493
rect 30837 15453 30849 15487
rect 30883 15484 30895 15487
rect 31386 15484 31392 15496
rect 30883 15456 31392 15484
rect 30883 15453 30895 15456
rect 30837 15447 30895 15453
rect 29641 15419 29699 15425
rect 29641 15385 29653 15419
rect 29687 15416 29699 15419
rect 29914 15416 29920 15428
rect 29687 15388 29920 15416
rect 29687 15385 29699 15388
rect 29641 15379 29699 15385
rect 29914 15376 29920 15388
rect 29972 15416 29978 15428
rect 30852 15416 30880 15447
rect 31386 15444 31392 15456
rect 31444 15444 31450 15496
rect 35161 15487 35219 15493
rect 35161 15453 35173 15487
rect 35207 15453 35219 15487
rect 35161 15447 35219 15453
rect 29972 15388 30880 15416
rect 29972 15376 29978 15388
rect 4341 15351 4399 15357
rect 4341 15317 4353 15351
rect 4387 15348 4399 15351
rect 4614 15348 4620 15360
rect 4387 15320 4620 15348
rect 4387 15317 4399 15320
rect 4341 15311 4399 15317
rect 4614 15308 4620 15320
rect 4672 15348 4678 15360
rect 6270 15348 6276 15360
rect 4672 15320 6276 15348
rect 4672 15308 4678 15320
rect 6270 15308 6276 15320
rect 6328 15348 6334 15360
rect 6365 15351 6423 15357
rect 6365 15348 6377 15351
rect 6328 15320 6377 15348
rect 6328 15308 6334 15320
rect 6365 15317 6377 15320
rect 6411 15317 6423 15351
rect 6365 15311 6423 15317
rect 6638 15308 6644 15360
rect 6696 15348 6702 15360
rect 7469 15351 7527 15357
rect 7469 15348 7481 15351
rect 6696 15320 7481 15348
rect 6696 15308 6702 15320
rect 7469 15317 7481 15320
rect 7515 15317 7527 15351
rect 7469 15311 7527 15317
rect 8021 15351 8079 15357
rect 8021 15317 8033 15351
rect 8067 15348 8079 15351
rect 8294 15348 8300 15360
rect 8067 15320 8300 15348
rect 8067 15317 8079 15320
rect 8021 15311 8079 15317
rect 8294 15308 8300 15320
rect 8352 15308 8358 15360
rect 14001 15351 14059 15357
rect 14001 15317 14013 15351
rect 14047 15348 14059 15351
rect 14550 15348 14556 15360
rect 14047 15320 14556 15348
rect 14047 15317 14059 15320
rect 14001 15311 14059 15317
rect 14550 15308 14556 15320
rect 14608 15308 14614 15360
rect 23661 15351 23719 15357
rect 23661 15317 23673 15351
rect 23707 15348 23719 15351
rect 24118 15348 24124 15360
rect 23707 15320 24124 15348
rect 23707 15317 23719 15320
rect 23661 15311 23719 15317
rect 24118 15308 24124 15320
rect 24176 15348 24182 15360
rect 25317 15351 25375 15357
rect 25317 15348 25329 15351
rect 24176 15320 25329 15348
rect 24176 15308 24182 15320
rect 25317 15317 25329 15320
rect 25363 15317 25375 15351
rect 30190 15348 30196 15360
rect 30151 15320 30196 15348
rect 25317 15311 25375 15317
rect 30190 15308 30196 15320
rect 30248 15308 30254 15360
rect 31754 15308 31760 15360
rect 31812 15348 31818 15360
rect 32309 15351 32367 15357
rect 32309 15348 32321 15351
rect 31812 15320 32321 15348
rect 31812 15308 31818 15320
rect 32309 15317 32321 15320
rect 32355 15317 32367 15351
rect 32309 15311 32367 15317
rect 33686 15308 33692 15360
rect 33744 15348 33750 15360
rect 33781 15351 33839 15357
rect 33781 15348 33793 15351
rect 33744 15320 33793 15348
rect 33744 15308 33750 15320
rect 33781 15317 33793 15320
rect 33827 15317 33839 15351
rect 35176 15348 35204 15447
rect 35342 15348 35348 15360
rect 35176 15320 35348 15348
rect 33781 15311 33839 15317
rect 35342 15308 35348 15320
rect 35400 15308 35406 15360
rect 1104 15258 38824 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 38824 15258
rect 1104 15184 38824 15206
rect 7285 15147 7343 15153
rect 7285 15113 7297 15147
rect 7331 15144 7343 15147
rect 8110 15144 8116 15156
rect 7331 15116 8116 15144
rect 7331 15113 7343 15116
rect 7285 15107 7343 15113
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 17494 15104 17500 15156
rect 17552 15144 17558 15156
rect 17589 15147 17647 15153
rect 17589 15144 17601 15147
rect 17552 15116 17601 15144
rect 17552 15104 17558 15116
rect 17589 15113 17601 15116
rect 17635 15113 17647 15147
rect 20622 15144 20628 15156
rect 20583 15116 20628 15144
rect 17589 15107 17647 15113
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 20993 15147 21051 15153
rect 20993 15113 21005 15147
rect 21039 15144 21051 15147
rect 21082 15144 21088 15156
rect 21039 15116 21088 15144
rect 21039 15113 21051 15116
rect 20993 15107 21051 15113
rect 21082 15104 21088 15116
rect 21140 15104 21146 15156
rect 23658 15144 23664 15156
rect 23619 15116 23664 15144
rect 23658 15104 23664 15116
rect 23716 15104 23722 15156
rect 24394 15104 24400 15156
rect 24452 15144 24458 15156
rect 24765 15147 24823 15153
rect 24765 15144 24777 15147
rect 24452 15116 24777 15144
rect 24452 15104 24458 15116
rect 24765 15113 24777 15116
rect 24811 15113 24823 15147
rect 26050 15144 26056 15156
rect 26011 15116 26056 15144
rect 24765 15107 24823 15113
rect 26050 15104 26056 15116
rect 26108 15104 26114 15156
rect 26510 15144 26516 15156
rect 26471 15116 26516 15144
rect 26510 15104 26516 15116
rect 26568 15104 26574 15156
rect 26970 15144 26976 15156
rect 26931 15116 26976 15144
rect 26970 15104 26976 15116
rect 27028 15104 27034 15156
rect 27430 15144 27436 15156
rect 27391 15116 27436 15144
rect 27430 15104 27436 15116
rect 27488 15104 27494 15156
rect 29914 15144 29920 15156
rect 29875 15116 29920 15144
rect 29914 15104 29920 15116
rect 29972 15104 29978 15156
rect 30558 15144 30564 15156
rect 30519 15116 30564 15144
rect 30558 15104 30564 15116
rect 30616 15104 30622 15156
rect 30926 15144 30932 15156
rect 30887 15116 30932 15144
rect 30926 15104 30932 15116
rect 30984 15104 30990 15156
rect 31386 15104 31392 15156
rect 31444 15144 31450 15156
rect 32401 15147 32459 15153
rect 32401 15144 32413 15147
rect 31444 15116 32413 15144
rect 31444 15104 31450 15116
rect 32401 15113 32413 15116
rect 32447 15113 32459 15147
rect 35342 15144 35348 15156
rect 32401 15107 32459 15113
rect 35176 15116 35348 15144
rect 14550 15008 14556 15020
rect 14511 14980 14556 15008
rect 14550 14968 14556 14980
rect 14608 14968 14614 15020
rect 21100 15017 21128 15104
rect 22370 15036 22376 15088
rect 22428 15076 22434 15088
rect 24670 15076 24676 15088
rect 22428 15048 24676 15076
rect 22428 15036 22434 15048
rect 21085 15011 21143 15017
rect 21085 14977 21097 15011
rect 21131 14977 21143 15011
rect 21085 14971 21143 14977
rect 23477 15011 23535 15017
rect 23477 14977 23489 15011
rect 23523 15008 23535 15011
rect 24118 15008 24124 15020
rect 23523 14980 24124 15008
rect 23523 14977 23535 14980
rect 23477 14971 23535 14977
rect 24118 14968 24124 14980
rect 24176 14968 24182 15020
rect 24228 15017 24256 15048
rect 24670 15036 24676 15048
rect 24728 15076 24734 15088
rect 25593 15079 25651 15085
rect 25593 15076 25605 15079
rect 24728 15048 25605 15076
rect 24728 15036 24734 15048
rect 25593 15045 25605 15048
rect 25639 15045 25651 15079
rect 25593 15039 25651 15045
rect 24213 15011 24271 15017
rect 24213 14977 24225 15011
rect 24259 15008 24271 15011
rect 24302 15008 24308 15020
rect 24259 14980 24308 15008
rect 24259 14977 24271 14980
rect 24213 14971 24271 14977
rect 24302 14968 24308 14980
rect 24360 14968 24366 15020
rect 30009 15011 30067 15017
rect 30009 14977 30021 15011
rect 30055 15008 30067 15011
rect 30576 15008 30604 15104
rect 30055 14980 30604 15008
rect 30944 15008 30972 15104
rect 31021 15011 31079 15017
rect 31021 15008 31033 15011
rect 30944 14980 31033 15008
rect 30055 14977 30067 14980
rect 30009 14971 30067 14977
rect 31021 14977 31033 14980
rect 31067 14977 31079 15011
rect 31021 14971 31079 14977
rect 4157 14943 4215 14949
rect 4157 14909 4169 14943
rect 4203 14940 4215 14943
rect 4246 14940 4252 14952
rect 4203 14912 4252 14940
rect 4203 14909 4215 14912
rect 4157 14903 4215 14909
rect 4246 14900 4252 14912
rect 4304 14940 4310 14952
rect 4982 14940 4988 14952
rect 4304 14912 4988 14940
rect 4304 14900 4310 14912
rect 4982 14900 4988 14912
rect 5040 14940 5046 14952
rect 6273 14943 6331 14949
rect 6273 14940 6285 14943
rect 5040 14912 6285 14940
rect 5040 14900 5046 14912
rect 6273 14909 6285 14912
rect 6319 14940 6331 14943
rect 7653 14943 7711 14949
rect 7653 14940 7665 14943
rect 6319 14912 7665 14940
rect 6319 14909 6331 14912
rect 6273 14903 6331 14909
rect 7653 14909 7665 14912
rect 7699 14940 7711 14943
rect 7745 14943 7803 14949
rect 7745 14940 7757 14943
rect 7699 14912 7757 14940
rect 7699 14909 7711 14912
rect 7653 14903 7711 14909
rect 7745 14909 7757 14912
rect 7791 14940 7803 14943
rect 8478 14940 8484 14952
rect 7791 14912 8484 14940
rect 7791 14909 7803 14912
rect 7745 14903 7803 14909
rect 8478 14900 8484 14912
rect 8536 14900 8542 14952
rect 13449 14943 13507 14949
rect 13449 14909 13461 14943
rect 13495 14940 13507 14943
rect 13495 14912 14412 14940
rect 13495 14909 13507 14912
rect 13449 14903 13507 14909
rect 4516 14875 4574 14881
rect 4516 14841 4528 14875
rect 4562 14872 4574 14875
rect 4614 14872 4620 14884
rect 4562 14844 4620 14872
rect 4562 14841 4574 14844
rect 4516 14835 4574 14841
rect 4614 14832 4620 14844
rect 4672 14832 4678 14884
rect 5994 14832 6000 14884
rect 6052 14872 6058 14884
rect 6641 14875 6699 14881
rect 6641 14872 6653 14875
rect 6052 14844 6653 14872
rect 6052 14832 6058 14844
rect 6641 14841 6653 14844
rect 6687 14872 6699 14875
rect 6687 14844 7696 14872
rect 6687 14841 6699 14844
rect 6641 14835 6699 14841
rect 5626 14804 5632 14816
rect 5587 14776 5632 14804
rect 5626 14764 5632 14776
rect 5684 14764 5690 14816
rect 7668 14804 7696 14844
rect 7926 14832 7932 14884
rect 7984 14881 7990 14884
rect 7984 14875 8048 14881
rect 7984 14841 8002 14875
rect 8036 14841 8048 14875
rect 7984 14835 8048 14841
rect 13817 14875 13875 14881
rect 13817 14841 13829 14875
rect 13863 14872 13875 14875
rect 14090 14872 14096 14884
rect 13863 14844 14096 14872
rect 13863 14841 13875 14844
rect 13817 14835 13875 14841
rect 7984 14832 7990 14835
rect 14090 14832 14096 14844
rect 14148 14872 14154 14884
rect 14277 14875 14335 14881
rect 14277 14872 14289 14875
rect 14148 14844 14289 14872
rect 14148 14832 14154 14844
rect 14277 14841 14289 14844
rect 14323 14841 14335 14875
rect 14277 14835 14335 14841
rect 9125 14807 9183 14813
rect 9125 14804 9137 14807
rect 7668 14776 9137 14804
rect 9125 14773 9137 14776
rect 9171 14773 9183 14807
rect 13906 14804 13912 14816
rect 13867 14776 13912 14804
rect 9125 14767 9183 14773
rect 13906 14764 13912 14776
rect 13964 14764 13970 14816
rect 14384 14813 14412 14912
rect 22278 14900 22284 14952
rect 22336 14940 22342 14952
rect 23109 14943 23167 14949
rect 23109 14940 23121 14943
rect 22336 14912 23121 14940
rect 22336 14900 22342 14912
rect 23109 14909 23121 14912
rect 23155 14940 23167 14943
rect 24029 14943 24087 14949
rect 24029 14940 24041 14943
rect 23155 14912 24041 14940
rect 23155 14909 23167 14912
rect 23109 14903 23167 14909
rect 24029 14909 24041 14912
rect 24075 14940 24087 14943
rect 24762 14940 24768 14952
rect 24075 14912 24768 14940
rect 24075 14909 24087 14912
rect 24029 14903 24087 14909
rect 24762 14900 24768 14912
rect 24820 14900 24826 14952
rect 25409 14943 25467 14949
rect 25409 14909 25421 14943
rect 25455 14940 25467 14943
rect 26050 14940 26056 14952
rect 25455 14912 26056 14940
rect 25455 14909 25467 14912
rect 25409 14903 25467 14909
rect 26050 14900 26056 14912
rect 26108 14900 26114 14952
rect 31288 14943 31346 14949
rect 31288 14909 31300 14943
rect 31334 14940 31346 14943
rect 31662 14940 31668 14952
rect 31334 14912 31668 14940
rect 31334 14909 31346 14912
rect 31288 14903 31346 14909
rect 31662 14900 31668 14912
rect 31720 14900 31726 14952
rect 33686 14940 33692 14952
rect 33647 14912 33692 14940
rect 33686 14900 33692 14912
rect 33744 14900 33750 14952
rect 35176 14949 35204 15116
rect 35342 15104 35348 15116
rect 35400 15104 35406 15156
rect 35161 14943 35219 14949
rect 35161 14940 35173 14943
rect 34624 14912 35173 14940
rect 20257 14875 20315 14881
rect 20257 14841 20269 14875
rect 20303 14872 20315 14875
rect 21330 14875 21388 14881
rect 21330 14872 21342 14875
rect 20303 14844 21342 14872
rect 20303 14841 20315 14844
rect 20257 14835 20315 14841
rect 21330 14841 21342 14844
rect 21376 14872 21388 14875
rect 21726 14872 21732 14884
rect 21376 14844 21732 14872
rect 21376 14841 21388 14844
rect 21330 14835 21388 14841
rect 21726 14832 21732 14844
rect 21784 14832 21790 14884
rect 29549 14875 29607 14881
rect 29549 14841 29561 14875
rect 29595 14872 29607 14875
rect 30650 14872 30656 14884
rect 29595 14844 30656 14872
rect 29595 14841 29607 14844
rect 29549 14835 29607 14841
rect 30650 14832 30656 14844
rect 30708 14832 30714 14884
rect 33042 14832 33048 14884
rect 33100 14872 33106 14884
rect 33100 14844 34192 14872
rect 33100 14832 33106 14844
rect 34164 14816 34192 14844
rect 14369 14807 14427 14813
rect 14369 14773 14381 14807
rect 14415 14804 14427 14807
rect 15102 14804 15108 14816
rect 14415 14776 15108 14804
rect 14415 14773 14427 14776
rect 14369 14767 14427 14773
rect 15102 14764 15108 14776
rect 15160 14764 15166 14816
rect 15470 14764 15476 14816
rect 15528 14804 15534 14816
rect 17218 14804 17224 14816
rect 15528 14776 17224 14804
rect 15528 14764 15534 14776
rect 17218 14764 17224 14776
rect 17276 14764 17282 14816
rect 21634 14764 21640 14816
rect 21692 14804 21698 14816
rect 22465 14807 22523 14813
rect 22465 14804 22477 14807
rect 21692 14776 22477 14804
rect 21692 14764 21698 14776
rect 22465 14773 22477 14776
rect 22511 14773 22523 14807
rect 22465 14767 22523 14773
rect 32490 14764 32496 14816
rect 32548 14804 32554 14816
rect 33226 14804 33232 14816
rect 32548 14776 33232 14804
rect 32548 14764 32554 14776
rect 33226 14764 33232 14776
rect 33284 14764 33290 14816
rect 33870 14804 33876 14816
rect 33831 14776 33876 14804
rect 33870 14764 33876 14776
rect 33928 14764 33934 14816
rect 34146 14764 34152 14816
rect 34204 14804 34210 14816
rect 34624 14813 34652 14912
rect 35161 14909 35173 14912
rect 35207 14909 35219 14943
rect 35161 14903 35219 14909
rect 35250 14832 35256 14884
rect 35308 14872 35314 14884
rect 35406 14875 35464 14881
rect 35406 14872 35418 14875
rect 35308 14844 35418 14872
rect 35308 14832 35314 14844
rect 35406 14841 35418 14844
rect 35452 14841 35464 14875
rect 35406 14835 35464 14841
rect 34241 14807 34299 14813
rect 34241 14804 34253 14807
rect 34204 14776 34253 14804
rect 34204 14764 34210 14776
rect 34241 14773 34253 14776
rect 34287 14804 34299 14807
rect 34609 14807 34667 14813
rect 34609 14804 34621 14807
rect 34287 14776 34621 14804
rect 34287 14773 34299 14776
rect 34241 14767 34299 14773
rect 34609 14773 34621 14776
rect 34655 14773 34667 14807
rect 34609 14767 34667 14773
rect 35894 14764 35900 14816
rect 35952 14804 35958 14816
rect 36541 14807 36599 14813
rect 36541 14804 36553 14807
rect 35952 14776 36553 14804
rect 35952 14764 35958 14776
rect 36541 14773 36553 14776
rect 36587 14773 36599 14807
rect 36541 14767 36599 14773
rect 1104 14714 38824 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 38824 14714
rect 1104 14640 38824 14662
rect 7006 14560 7012 14612
rect 7064 14600 7070 14612
rect 7193 14603 7251 14609
rect 7193 14600 7205 14603
rect 7064 14572 7205 14600
rect 7064 14560 7070 14572
rect 7193 14569 7205 14572
rect 7239 14600 7251 14603
rect 7374 14600 7380 14612
rect 7239 14572 7380 14600
rect 7239 14569 7251 14572
rect 7193 14563 7251 14569
rect 7374 14560 7380 14572
rect 7432 14560 7438 14612
rect 7837 14603 7895 14609
rect 7837 14569 7849 14603
rect 7883 14600 7895 14603
rect 7926 14600 7932 14612
rect 7883 14572 7932 14600
rect 7883 14569 7895 14572
rect 7837 14563 7895 14569
rect 7926 14560 7932 14572
rect 7984 14560 7990 14612
rect 8018 14560 8024 14612
rect 8076 14600 8082 14612
rect 8113 14603 8171 14609
rect 8113 14600 8125 14603
rect 8076 14572 8125 14600
rect 8076 14560 8082 14572
rect 8113 14569 8125 14572
rect 8159 14569 8171 14603
rect 8113 14563 8171 14569
rect 8662 14560 8668 14612
rect 8720 14600 8726 14612
rect 8849 14603 8907 14609
rect 8849 14600 8861 14603
rect 8720 14572 8861 14600
rect 8720 14560 8726 14572
rect 8849 14569 8861 14572
rect 8895 14569 8907 14603
rect 8849 14563 8907 14569
rect 13906 14560 13912 14612
rect 13964 14600 13970 14612
rect 14461 14603 14519 14609
rect 14461 14600 14473 14603
rect 13964 14572 14473 14600
rect 13964 14560 13970 14572
rect 14461 14569 14473 14572
rect 14507 14600 14519 14603
rect 14918 14600 14924 14612
rect 14507 14572 14924 14600
rect 14507 14569 14519 14572
rect 14461 14563 14519 14569
rect 14918 14560 14924 14572
rect 14976 14560 14982 14612
rect 21082 14600 21088 14612
rect 21043 14572 21088 14600
rect 21082 14560 21088 14572
rect 21140 14560 21146 14612
rect 21266 14600 21272 14612
rect 21227 14572 21272 14600
rect 21266 14560 21272 14572
rect 21324 14560 21330 14612
rect 21726 14600 21732 14612
rect 21687 14572 21732 14600
rect 21726 14560 21732 14572
rect 21784 14600 21790 14612
rect 22002 14600 22008 14612
rect 21784 14572 22008 14600
rect 21784 14560 21790 14572
rect 22002 14560 22008 14572
rect 22060 14560 22066 14612
rect 24026 14600 24032 14612
rect 23987 14572 24032 14600
rect 24026 14560 24032 14572
rect 24084 14560 24090 14612
rect 24302 14600 24308 14612
rect 24263 14572 24308 14600
rect 24302 14560 24308 14572
rect 24360 14560 24366 14612
rect 30377 14603 30435 14609
rect 30377 14569 30389 14603
rect 30423 14600 30435 14603
rect 30466 14600 30472 14612
rect 30423 14572 30472 14600
rect 30423 14569 30435 14572
rect 30377 14563 30435 14569
rect 30466 14560 30472 14572
rect 30524 14560 30530 14612
rect 30558 14560 30564 14612
rect 30616 14600 30622 14612
rect 31297 14603 31355 14609
rect 31297 14600 31309 14603
rect 30616 14572 31309 14600
rect 30616 14560 30622 14572
rect 31297 14569 31309 14572
rect 31343 14600 31355 14603
rect 32122 14600 32128 14612
rect 31343 14572 31984 14600
rect 32083 14572 32128 14600
rect 31343 14569 31355 14572
rect 31297 14563 31355 14569
rect 21634 14532 21640 14544
rect 21595 14504 21640 14532
rect 21634 14492 21640 14504
rect 21692 14492 21698 14544
rect 31956 14541 31984 14572
rect 32122 14560 32128 14572
rect 32180 14560 32186 14612
rect 32490 14600 32496 14612
rect 32451 14572 32496 14600
rect 32490 14560 32496 14572
rect 32548 14560 32554 14612
rect 35894 14600 35900 14612
rect 35855 14572 35900 14600
rect 35894 14560 35900 14572
rect 35952 14560 35958 14612
rect 36814 14600 36820 14612
rect 36775 14572 36820 14600
rect 36814 14560 36820 14572
rect 36872 14560 36878 14612
rect 31941 14535 31999 14541
rect 31941 14501 31953 14535
rect 31987 14532 31999 14535
rect 33410 14532 33416 14544
rect 31987 14504 33416 14532
rect 31987 14501 31999 14504
rect 31941 14495 31999 14501
rect 33410 14492 33416 14504
rect 33468 14492 33474 14544
rect 3510 14424 3516 14476
rect 3568 14464 3574 14476
rect 4505 14467 4563 14473
rect 4505 14464 4517 14467
rect 3568 14436 4517 14464
rect 3568 14424 3574 14436
rect 4505 14433 4517 14436
rect 4551 14464 4563 14467
rect 4798 14464 4804 14476
rect 4551 14436 4804 14464
rect 4551 14433 4563 14436
rect 4505 14427 4563 14433
rect 4798 14424 4804 14436
rect 4856 14464 4862 14476
rect 5626 14464 5632 14476
rect 4856 14436 5632 14464
rect 4856 14424 4862 14436
rect 5626 14424 5632 14436
rect 5684 14424 5690 14476
rect 7098 14464 7104 14476
rect 7059 14436 7104 14464
rect 7098 14424 7104 14436
rect 7156 14424 7162 14476
rect 8294 14464 8300 14476
rect 8255 14436 8300 14464
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 9858 14464 9864 14476
rect 9819 14436 9864 14464
rect 9858 14424 9864 14436
rect 9916 14424 9922 14476
rect 11238 14424 11244 14476
rect 11296 14464 11302 14476
rect 12526 14464 12532 14476
rect 11296 14436 12532 14464
rect 11296 14424 11302 14436
rect 12526 14424 12532 14436
rect 12584 14424 12590 14476
rect 12618 14424 12624 14476
rect 12676 14464 12682 14476
rect 12785 14467 12843 14473
rect 12785 14464 12797 14467
rect 12676 14436 12797 14464
rect 12676 14424 12682 14436
rect 12785 14433 12797 14436
rect 12831 14433 12843 14467
rect 22370 14464 22376 14476
rect 12785 14427 12843 14433
rect 21928 14436 22376 14464
rect 3878 14356 3884 14408
rect 3936 14396 3942 14408
rect 4246 14396 4252 14408
rect 3936 14368 4252 14396
rect 3936 14356 3942 14368
rect 4246 14356 4252 14368
rect 4304 14356 4310 14408
rect 6270 14356 6276 14408
rect 6328 14396 6334 14408
rect 7377 14399 7435 14405
rect 7377 14396 7389 14399
rect 6328 14368 7389 14396
rect 6328 14356 6334 14368
rect 7377 14365 7389 14368
rect 7423 14396 7435 14399
rect 8662 14396 8668 14408
rect 7423 14368 8668 14396
rect 7423 14365 7435 14368
rect 7377 14359 7435 14365
rect 8662 14356 8668 14368
rect 8720 14356 8726 14408
rect 11146 14356 11152 14408
rect 11204 14396 11210 14408
rect 21928 14405 21956 14436
rect 22370 14424 22376 14436
rect 22428 14424 22434 14476
rect 29086 14424 29092 14476
rect 29144 14464 29150 14476
rect 29365 14467 29423 14473
rect 29365 14464 29377 14467
rect 29144 14436 29377 14464
rect 29144 14424 29150 14436
rect 29365 14433 29377 14436
rect 29411 14464 29423 14467
rect 30834 14464 30840 14476
rect 29411 14436 30328 14464
rect 30795 14436 30840 14464
rect 29411 14433 29423 14436
rect 29365 14427 29423 14433
rect 11517 14399 11575 14405
rect 11517 14396 11529 14399
rect 11204 14368 11529 14396
rect 11204 14356 11210 14368
rect 11517 14365 11529 14368
rect 11563 14365 11575 14399
rect 11517 14359 11575 14365
rect 21913 14399 21971 14405
rect 21913 14365 21925 14399
rect 21959 14365 21971 14399
rect 21913 14359 21971 14365
rect 5258 14220 5264 14272
rect 5316 14260 5322 14272
rect 5626 14260 5632 14272
rect 5316 14232 5632 14260
rect 5316 14220 5322 14232
rect 5626 14220 5632 14232
rect 5684 14220 5690 14272
rect 6730 14260 6736 14272
rect 6691 14232 6736 14260
rect 6730 14220 6736 14232
rect 6788 14220 6794 14272
rect 8478 14260 8484 14272
rect 8439 14232 8484 14260
rect 8478 14220 8484 14232
rect 8536 14220 8542 14272
rect 10042 14260 10048 14272
rect 10003 14232 10048 14260
rect 10042 14220 10048 14232
rect 10100 14220 10106 14272
rect 10778 14260 10784 14272
rect 10739 14232 10784 14260
rect 10778 14220 10784 14232
rect 10836 14220 10842 14272
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 13909 14263 13967 14269
rect 13909 14260 13921 14263
rect 13504 14232 13921 14260
rect 13504 14220 13510 14232
rect 13909 14229 13921 14232
rect 13955 14229 13967 14263
rect 13909 14223 13967 14229
rect 19245 14263 19303 14269
rect 19245 14229 19257 14263
rect 19291 14260 19303 14263
rect 19334 14260 19340 14272
rect 19291 14232 19340 14260
rect 19291 14229 19303 14232
rect 19245 14223 19303 14229
rect 19334 14220 19340 14232
rect 19392 14220 19398 14272
rect 26970 14260 26976 14272
rect 26931 14232 26976 14260
rect 26970 14220 26976 14232
rect 27028 14220 27034 14272
rect 29546 14260 29552 14272
rect 29507 14232 29552 14260
rect 29546 14220 29552 14232
rect 29604 14220 29610 14272
rect 30300 14260 30328 14436
rect 30834 14424 30840 14436
rect 30892 14424 30898 14476
rect 32582 14464 32588 14476
rect 32543 14436 32588 14464
rect 32582 14424 32588 14436
rect 32640 14424 32646 14476
rect 33689 14467 33747 14473
rect 33689 14433 33701 14467
rect 33735 14464 33747 14467
rect 33778 14464 33784 14476
rect 33735 14436 33784 14464
rect 33735 14433 33747 14436
rect 33689 14427 33747 14433
rect 33778 14424 33784 14436
rect 33836 14424 33842 14476
rect 34514 14424 34520 14476
rect 34572 14464 34578 14476
rect 35250 14464 35256 14476
rect 34572 14436 35256 14464
rect 34572 14424 34578 14436
rect 35250 14424 35256 14436
rect 35308 14424 35314 14476
rect 35912 14464 35940 14560
rect 36449 14535 36507 14541
rect 36449 14501 36461 14535
rect 36495 14532 36507 14535
rect 37090 14532 37096 14544
rect 36495 14504 37096 14532
rect 36495 14501 36507 14504
rect 36449 14495 36507 14501
rect 37090 14492 37096 14504
rect 37148 14492 37154 14544
rect 36538 14464 36544 14476
rect 35912 14436 36544 14464
rect 36538 14424 36544 14436
rect 36596 14464 36602 14476
rect 36633 14467 36691 14473
rect 36633 14464 36645 14467
rect 36596 14436 36645 14464
rect 36596 14424 36602 14436
rect 36633 14433 36645 14436
rect 36679 14433 36691 14467
rect 36633 14427 36691 14433
rect 30558 14356 30564 14408
rect 30616 14396 30622 14408
rect 30929 14399 30987 14405
rect 30929 14396 30941 14399
rect 30616 14368 30941 14396
rect 30616 14356 30622 14368
rect 30929 14365 30941 14368
rect 30975 14365 30987 14399
rect 30929 14359 30987 14365
rect 31113 14399 31171 14405
rect 31113 14365 31125 14399
rect 31159 14396 31171 14399
rect 31297 14399 31355 14405
rect 31297 14396 31309 14399
rect 31159 14368 31309 14396
rect 31159 14365 31171 14368
rect 31113 14359 31171 14365
rect 31297 14365 31309 14368
rect 31343 14365 31355 14399
rect 31297 14359 31355 14365
rect 31573 14399 31631 14405
rect 31573 14365 31585 14399
rect 31619 14396 31631 14399
rect 32769 14399 32827 14405
rect 32769 14396 32781 14399
rect 31619 14368 32781 14396
rect 31619 14365 31631 14368
rect 31573 14359 31631 14365
rect 32769 14365 32781 14368
rect 32815 14396 32827 14399
rect 33870 14396 33876 14408
rect 32815 14368 33876 14396
rect 32815 14365 32827 14368
rect 32769 14359 32827 14365
rect 33870 14356 33876 14368
rect 33928 14356 33934 14408
rect 34793 14399 34851 14405
rect 34793 14365 34805 14399
rect 34839 14396 34851 14399
rect 35342 14396 35348 14408
rect 34839 14368 35348 14396
rect 34839 14365 34851 14368
rect 34793 14359 34851 14365
rect 35342 14356 35348 14368
rect 35400 14356 35406 14408
rect 35437 14399 35495 14405
rect 35437 14365 35449 14399
rect 35483 14365 35495 14399
rect 35437 14359 35495 14365
rect 34514 14288 34520 14340
rect 34572 14328 34578 14340
rect 34885 14331 34943 14337
rect 34885 14328 34897 14331
rect 34572 14300 34897 14328
rect 34572 14288 34578 14300
rect 34885 14297 34897 14300
rect 34931 14297 34943 14331
rect 35452 14328 35480 14359
rect 34885 14291 34943 14297
rect 35421 14300 35480 14328
rect 35421 14272 35449 14300
rect 30469 14263 30527 14269
rect 30469 14260 30481 14263
rect 30300 14232 30481 14260
rect 30469 14229 30481 14232
rect 30515 14260 30527 14263
rect 31294 14260 31300 14272
rect 30515 14232 31300 14260
rect 30515 14229 30527 14232
rect 30469 14223 30527 14229
rect 31294 14220 31300 14232
rect 31352 14220 31358 14272
rect 33318 14260 33324 14272
rect 33279 14232 33324 14260
rect 33318 14220 33324 14232
rect 33376 14220 33382 14272
rect 33410 14220 33416 14272
rect 33468 14260 33474 14272
rect 33873 14263 33931 14269
rect 33873 14260 33885 14263
rect 33468 14232 33885 14260
rect 33468 14220 33474 14232
rect 33873 14229 33885 14232
rect 33919 14229 33931 14263
rect 33873 14223 33931 14229
rect 34054 14220 34060 14272
rect 34112 14260 34118 14272
rect 34333 14263 34391 14269
rect 34333 14260 34345 14263
rect 34112 14232 34345 14260
rect 34112 14220 34118 14232
rect 34333 14229 34345 14232
rect 34379 14260 34391 14263
rect 35421 14260 35440 14272
rect 34379 14232 35440 14260
rect 34379 14229 34391 14232
rect 34333 14223 34391 14229
rect 35434 14220 35440 14232
rect 35492 14260 35498 14272
rect 35492 14232 35554 14260
rect 35492 14220 35498 14232
rect 1104 14170 38824 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 38824 14170
rect 1104 14096 38824 14118
rect 3510 14056 3516 14068
rect 3471 14028 3516 14056
rect 3510 14016 3516 14028
rect 3568 14016 3574 14068
rect 3878 14056 3884 14068
rect 3839 14028 3884 14056
rect 3878 14016 3884 14028
rect 3936 14016 3942 14068
rect 5534 14016 5540 14068
rect 5592 14056 5598 14068
rect 6549 14059 6607 14065
rect 6549 14056 6561 14059
rect 5592 14028 6561 14056
rect 5592 14016 5598 14028
rect 6549 14025 6561 14028
rect 6595 14056 6607 14059
rect 7098 14056 7104 14068
rect 6595 14028 7104 14056
rect 6595 14025 6607 14028
rect 6549 14019 6607 14025
rect 7098 14016 7104 14028
rect 7156 14016 7162 14068
rect 7374 14056 7380 14068
rect 7335 14028 7380 14056
rect 7374 14016 7380 14028
rect 7432 14016 7438 14068
rect 8297 14059 8355 14065
rect 8297 14025 8309 14059
rect 8343 14056 8355 14059
rect 8478 14056 8484 14068
rect 8343 14028 8484 14056
rect 8343 14025 8355 14028
rect 8297 14019 8355 14025
rect 6270 13988 6276 14000
rect 6231 13960 6276 13988
rect 6270 13948 6276 13960
rect 6328 13948 6334 14000
rect 7009 13991 7067 13997
rect 7009 13957 7021 13991
rect 7055 13988 7067 13991
rect 7837 13991 7895 13997
rect 7837 13988 7849 13991
rect 7055 13960 7849 13988
rect 7055 13957 7067 13960
rect 7009 13951 7067 13957
rect 7837 13957 7849 13960
rect 7883 13957 7895 13991
rect 7837 13951 7895 13957
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13920 3203 13923
rect 3191 13892 4108 13920
rect 3191 13889 3203 13892
rect 3145 13883 3203 13889
rect 3878 13812 3884 13864
rect 3936 13852 3942 13864
rect 3973 13855 4031 13861
rect 3973 13852 3985 13855
rect 3936 13824 3985 13852
rect 3936 13812 3942 13824
rect 3973 13821 3985 13824
rect 4019 13821 4031 13855
rect 4080 13852 4108 13892
rect 4229 13855 4287 13861
rect 4229 13852 4241 13855
rect 4080 13824 4241 13852
rect 3973 13815 4031 13821
rect 4229 13821 4241 13824
rect 4275 13852 4287 13855
rect 5626 13852 5632 13864
rect 4275 13824 5632 13852
rect 4275 13821 4287 13824
rect 4229 13815 4287 13821
rect 5626 13812 5632 13824
rect 5684 13812 5690 13864
rect 6730 13812 6736 13864
rect 6788 13852 6794 13864
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6788 13824 6837 13852
rect 6788 13812 6794 13824
rect 6825 13821 6837 13824
rect 6871 13852 6883 13855
rect 6914 13852 6920 13864
rect 6871 13824 6920 13852
rect 6871 13821 6883 13824
rect 6825 13815 6883 13821
rect 6914 13812 6920 13824
rect 6972 13812 6978 13864
rect 7852 13852 7880 13951
rect 8312 13920 8340 14019
rect 8478 14016 8484 14028
rect 8536 14016 8542 14068
rect 10689 14059 10747 14065
rect 10689 14025 10701 14059
rect 10735 14056 10747 14059
rect 11146 14056 11152 14068
rect 10735 14028 11152 14056
rect 10735 14025 10747 14028
rect 10689 14019 10747 14025
rect 11146 14016 11152 14028
rect 11204 14016 11210 14068
rect 12526 14016 12532 14068
rect 12584 14056 12590 14068
rect 12621 14059 12679 14065
rect 12621 14056 12633 14059
rect 12584 14028 12633 14056
rect 12584 14016 12590 14028
rect 12621 14025 12633 14028
rect 12667 14025 12679 14059
rect 14366 14056 14372 14068
rect 12621 14019 12679 14025
rect 13280 14028 14372 14056
rect 8389 13991 8447 13997
rect 8389 13957 8401 13991
rect 8435 13988 8447 13991
rect 10781 13991 10839 13997
rect 8435 13960 9536 13988
rect 8435 13957 8447 13960
rect 8389 13951 8447 13957
rect 8849 13923 8907 13929
rect 8849 13920 8861 13923
rect 8312 13892 8861 13920
rect 8849 13889 8861 13892
rect 8895 13889 8907 13923
rect 8849 13883 8907 13889
rect 8941 13923 8999 13929
rect 8941 13889 8953 13923
rect 8987 13889 8999 13923
rect 8941 13883 8999 13889
rect 7852 13824 8248 13852
rect 8220 13784 8248 13824
rect 8662 13812 8668 13864
rect 8720 13852 8726 13864
rect 8956 13852 8984 13883
rect 9508 13864 9536 13960
rect 10781 13957 10793 13991
rect 10827 13957 10839 13991
rect 10781 13951 10839 13957
rect 9401 13855 9459 13861
rect 9401 13852 9413 13855
rect 8720 13824 9413 13852
rect 8720 13812 8726 13824
rect 9401 13821 9413 13824
rect 9447 13821 9459 13855
rect 9401 13815 9459 13821
rect 9490 13812 9496 13864
rect 9548 13852 9554 13864
rect 9858 13852 9864 13864
rect 9548 13824 9864 13852
rect 9548 13812 9554 13824
rect 9858 13812 9864 13824
rect 9916 13812 9922 13864
rect 10796 13852 10824 13951
rect 10870 13880 10876 13932
rect 10928 13920 10934 13932
rect 13280 13929 13308 14028
rect 14366 14016 14372 14028
rect 14424 14056 14430 14068
rect 16209 14059 16267 14065
rect 16209 14056 16221 14059
rect 14424 14028 16221 14056
rect 14424 14016 14430 14028
rect 16209 14025 16221 14028
rect 16255 14025 16267 14059
rect 16209 14019 16267 14025
rect 21361 14059 21419 14065
rect 21361 14025 21373 14059
rect 21407 14056 21419 14059
rect 21726 14056 21732 14068
rect 21407 14028 21732 14056
rect 21407 14025 21419 14028
rect 21361 14019 21419 14025
rect 21726 14016 21732 14028
rect 21784 14016 21790 14068
rect 22097 14059 22155 14065
rect 22097 14025 22109 14059
rect 22143 14056 22155 14059
rect 22370 14056 22376 14068
rect 22143 14028 22376 14056
rect 22143 14025 22155 14028
rect 22097 14019 22155 14025
rect 22370 14016 22376 14028
rect 22428 14016 22434 14068
rect 26694 14056 26700 14068
rect 26655 14028 26700 14056
rect 26694 14016 26700 14028
rect 26752 14016 26758 14068
rect 29086 14056 29092 14068
rect 29047 14028 29092 14056
rect 29086 14016 29092 14028
rect 29144 14016 29150 14068
rect 29457 14059 29515 14065
rect 29457 14025 29469 14059
rect 29503 14056 29515 14059
rect 30558 14056 30564 14068
rect 29503 14028 30564 14056
rect 29503 14025 29515 14028
rect 29457 14019 29515 14025
rect 30558 14016 30564 14028
rect 30616 14016 30622 14068
rect 30650 14016 30656 14068
rect 30708 14056 30714 14068
rect 31205 14059 31263 14065
rect 31205 14056 31217 14059
rect 30708 14028 31217 14056
rect 30708 14016 30714 14028
rect 31205 14025 31217 14028
rect 31251 14025 31263 14059
rect 31205 14019 31263 14025
rect 31294 14016 31300 14068
rect 31352 14056 31358 14068
rect 32309 14059 32367 14065
rect 32309 14056 32321 14059
rect 31352 14028 32321 14056
rect 31352 14016 31358 14028
rect 32309 14025 32321 14028
rect 32355 14056 32367 14059
rect 32582 14056 32588 14068
rect 32355 14028 32588 14056
rect 32355 14025 32367 14028
rect 32309 14019 32367 14025
rect 32582 14016 32588 14028
rect 32640 14016 32646 14068
rect 35250 14016 35256 14068
rect 35308 14056 35314 14068
rect 36449 14059 36507 14065
rect 36449 14056 36461 14059
rect 35308 14028 36461 14056
rect 35308 14016 35314 14028
rect 36449 14025 36461 14028
rect 36495 14025 36507 14059
rect 37090 14056 37096 14068
rect 37051 14028 37096 14056
rect 36449 14019 36507 14025
rect 37090 14016 37096 14028
rect 37148 14016 37154 14068
rect 21634 13988 21640 14000
rect 21595 13960 21640 13988
rect 21634 13948 21640 13960
rect 21692 13948 21698 14000
rect 25590 13988 25596 14000
rect 25551 13960 25596 13988
rect 25590 13948 25596 13960
rect 25648 13948 25654 14000
rect 29546 13948 29552 14000
rect 29604 13988 29610 14000
rect 31021 13991 31079 13997
rect 31021 13988 31033 13991
rect 29604 13960 31033 13988
rect 29604 13948 29610 13960
rect 31021 13957 31033 13960
rect 31067 13957 31079 13991
rect 31021 13951 31079 13957
rect 11333 13923 11391 13929
rect 11333 13920 11345 13923
rect 10928 13892 11345 13920
rect 10928 13880 10934 13892
rect 11333 13889 11345 13892
rect 11379 13920 11391 13923
rect 11793 13923 11851 13929
rect 11793 13920 11805 13923
rect 11379 13892 11805 13920
rect 11379 13889 11391 13892
rect 11333 13883 11391 13889
rect 11793 13889 11805 13892
rect 11839 13889 11851 13923
rect 11793 13883 11851 13889
rect 12253 13923 12311 13929
rect 12253 13889 12265 13923
rect 12299 13920 12311 13923
rect 13265 13923 13323 13929
rect 13265 13920 13277 13923
rect 12299 13892 13277 13920
rect 12299 13889 12311 13892
rect 12253 13883 12311 13889
rect 13265 13889 13277 13892
rect 13311 13889 13323 13923
rect 13446 13920 13452 13932
rect 13407 13892 13452 13920
rect 13265 13883 13323 13889
rect 11146 13852 11152 13864
rect 10796 13824 11008 13852
rect 11107 13824 11152 13852
rect 8757 13787 8815 13793
rect 8757 13784 8769 13787
rect 8220 13756 8769 13784
rect 8757 13753 8769 13756
rect 8803 13753 8815 13787
rect 10980 13784 11008 13824
rect 11146 13812 11152 13824
rect 11204 13812 11210 13864
rect 11808 13852 11836 13883
rect 13446 13880 13452 13892
rect 13504 13880 13510 13932
rect 14918 13929 14924 13932
rect 13909 13923 13967 13929
rect 13909 13889 13921 13923
rect 13955 13920 13967 13923
rect 14875 13923 14924 13929
rect 13955 13892 14780 13920
rect 13955 13889 13967 13892
rect 13909 13883 13967 13889
rect 12526 13852 12532 13864
rect 11808 13824 12532 13852
rect 12526 13812 12532 13824
rect 12584 13812 12590 13864
rect 14369 13855 14427 13861
rect 14369 13821 14381 13855
rect 14415 13852 14427 13855
rect 14642 13852 14648 13864
rect 14415 13824 14648 13852
rect 14415 13821 14427 13824
rect 14369 13815 14427 13821
rect 14642 13812 14648 13824
rect 14700 13812 14706 13864
rect 14752 13852 14780 13892
rect 14875 13889 14887 13923
rect 14921 13889 14924 13923
rect 14875 13883 14924 13889
rect 14918 13880 14924 13883
rect 14976 13880 14982 13932
rect 19705 13923 19763 13929
rect 19705 13920 19717 13923
rect 18616 13892 19717 13920
rect 18616 13864 18644 13892
rect 19705 13889 19717 13892
rect 19751 13889 19763 13923
rect 19705 13883 19763 13889
rect 26421 13923 26479 13929
rect 26421 13889 26433 13923
rect 26467 13920 26479 13923
rect 27430 13920 27436 13932
rect 26467 13892 27436 13920
rect 26467 13889 26479 13892
rect 26421 13883 26479 13889
rect 27430 13880 27436 13892
rect 27488 13880 27494 13932
rect 15105 13855 15163 13861
rect 15105 13852 15117 13855
rect 14752 13824 15117 13852
rect 15105 13821 15117 13824
rect 15151 13852 15163 13855
rect 18598 13852 18604 13864
rect 15151 13824 15792 13852
rect 18559 13824 18604 13852
rect 15151 13821 15163 13824
rect 15105 13815 15163 13821
rect 12434 13784 12440 13796
rect 10980 13756 12440 13784
rect 8757 13747 8815 13753
rect 12434 13744 12440 13756
rect 12492 13744 12498 13796
rect 15764 13784 15792 13824
rect 18598 13812 18604 13824
rect 18656 13812 18662 13864
rect 19061 13855 19119 13861
rect 19061 13821 19073 13855
rect 19107 13852 19119 13855
rect 19426 13852 19432 13864
rect 19107 13824 19432 13852
rect 19107 13821 19119 13824
rect 19061 13815 19119 13821
rect 19426 13812 19432 13824
rect 19484 13852 19490 13864
rect 19613 13855 19671 13861
rect 19613 13852 19625 13855
rect 19484 13824 19625 13852
rect 19484 13812 19490 13824
rect 19613 13821 19625 13824
rect 19659 13821 19671 13855
rect 19613 13815 19671 13821
rect 25777 13855 25835 13861
rect 25777 13821 25789 13855
rect 25823 13821 25835 13855
rect 25777 13815 25835 13821
rect 16114 13784 16120 13796
rect 15764 13756 16120 13784
rect 16114 13744 16120 13756
rect 16172 13744 16178 13796
rect 19334 13744 19340 13796
rect 19392 13784 19398 13796
rect 19521 13787 19579 13793
rect 19521 13784 19533 13787
rect 19392 13756 19533 13784
rect 19392 13744 19398 13756
rect 19521 13753 19533 13756
rect 19567 13753 19579 13787
rect 19521 13747 19579 13753
rect 25501 13787 25559 13793
rect 25501 13753 25513 13787
rect 25547 13784 25559 13787
rect 25682 13784 25688 13796
rect 25547 13756 25688 13784
rect 25547 13753 25559 13756
rect 25501 13747 25559 13753
rect 25682 13744 25688 13756
rect 25740 13784 25746 13796
rect 25792 13784 25820 13815
rect 26970 13812 26976 13864
rect 27028 13852 27034 13864
rect 27249 13855 27307 13861
rect 27249 13852 27261 13855
rect 27028 13824 27261 13852
rect 27028 13812 27034 13824
rect 27249 13821 27261 13824
rect 27295 13821 27307 13855
rect 27249 13815 27307 13821
rect 28721 13855 28779 13861
rect 28721 13821 28733 13855
rect 28767 13852 28779 13855
rect 28994 13852 29000 13864
rect 28767 13824 29000 13852
rect 28767 13821 28779 13824
rect 28721 13815 28779 13821
rect 28994 13812 29000 13824
rect 29052 13852 29058 13864
rect 29273 13855 29331 13861
rect 29273 13852 29285 13855
rect 29052 13824 29285 13852
rect 29052 13812 29058 13824
rect 29273 13821 29285 13824
rect 29319 13821 29331 13855
rect 29273 13815 29331 13821
rect 30193 13855 30251 13861
rect 30193 13821 30205 13855
rect 30239 13852 30251 13855
rect 30834 13852 30840 13864
rect 30239 13824 30840 13852
rect 30239 13821 30251 13824
rect 30193 13815 30251 13821
rect 30834 13812 30840 13824
rect 30892 13812 30898 13864
rect 31036 13852 31064 13951
rect 31570 13948 31576 14000
rect 31628 13988 31634 14000
rect 33870 13988 33876 14000
rect 31628 13960 31800 13988
rect 33831 13960 33876 13988
rect 31628 13948 31634 13960
rect 31662 13920 31668 13932
rect 31623 13892 31668 13920
rect 31662 13880 31668 13892
rect 31720 13880 31726 13932
rect 31772 13929 31800 13960
rect 33870 13948 33876 13960
rect 33928 13948 33934 14000
rect 31757 13923 31815 13929
rect 31757 13889 31769 13923
rect 31803 13889 31815 13923
rect 33410 13920 33416 13932
rect 33371 13892 33416 13920
rect 31757 13883 31815 13889
rect 33410 13880 33416 13892
rect 33468 13880 33474 13932
rect 34333 13923 34391 13929
rect 34333 13889 34345 13923
rect 34379 13920 34391 13923
rect 34379 13892 35204 13920
rect 34379 13889 34391 13892
rect 34333 13883 34391 13889
rect 31573 13855 31631 13861
rect 31573 13852 31585 13855
rect 31036 13824 31585 13852
rect 31573 13821 31585 13824
rect 31619 13821 31631 13855
rect 31573 13815 31631 13821
rect 34146 13812 34152 13864
rect 34204 13852 34210 13864
rect 35069 13855 35127 13861
rect 35069 13852 35081 13855
rect 34204 13824 35081 13852
rect 34204 13812 34210 13824
rect 35069 13821 35081 13824
rect 35115 13821 35127 13855
rect 35176 13852 35204 13892
rect 35342 13861 35348 13864
rect 35336 13852 35348 13861
rect 35176 13824 35348 13852
rect 35069 13815 35127 13821
rect 35336 13815 35348 13824
rect 35400 13852 35406 13864
rect 35400 13824 35848 13852
rect 25740 13756 25820 13784
rect 25740 13744 25746 13756
rect 26694 13744 26700 13796
rect 26752 13784 26758 13796
rect 27341 13787 27399 13793
rect 27341 13784 27353 13787
rect 26752 13756 27353 13784
rect 26752 13744 26758 13756
rect 27341 13753 27353 13756
rect 27387 13753 27399 13787
rect 27341 13747 27399 13753
rect 32398 13744 32404 13796
rect 32456 13784 32462 13796
rect 32677 13787 32735 13793
rect 32677 13784 32689 13787
rect 32456 13756 32689 13784
rect 32456 13744 32462 13756
rect 32677 13753 32689 13756
rect 32723 13784 32735 13787
rect 33229 13787 33287 13793
rect 33229 13784 33241 13787
rect 32723 13756 33241 13784
rect 32723 13753 32735 13756
rect 32677 13747 32735 13753
rect 33229 13753 33241 13756
rect 33275 13753 33287 13787
rect 33229 13747 33287 13753
rect 5074 13676 5080 13728
rect 5132 13716 5138 13728
rect 5353 13719 5411 13725
rect 5353 13716 5365 13719
rect 5132 13688 5365 13716
rect 5132 13676 5138 13688
rect 5353 13685 5365 13688
rect 5399 13685 5411 13719
rect 5353 13679 5411 13685
rect 9950 13676 9956 13728
rect 10008 13716 10014 13728
rect 10778 13716 10784 13728
rect 10008 13688 10784 13716
rect 10008 13676 10014 13688
rect 10778 13676 10784 13688
rect 10836 13716 10842 13728
rect 11241 13719 11299 13725
rect 11241 13716 11253 13719
rect 10836 13688 11253 13716
rect 10836 13676 10842 13688
rect 11241 13685 11253 13688
rect 11287 13685 11299 13719
rect 12802 13716 12808 13728
rect 12763 13688 12808 13716
rect 11241 13679 11299 13685
rect 12802 13676 12808 13688
rect 12860 13676 12866 13728
rect 13173 13719 13231 13725
rect 13173 13685 13185 13719
rect 13219 13716 13231 13719
rect 13262 13716 13268 13728
rect 13219 13688 13268 13716
rect 13219 13685 13231 13688
rect 13173 13679 13231 13685
rect 13262 13676 13268 13688
rect 13320 13676 13326 13728
rect 13906 13676 13912 13728
rect 13964 13716 13970 13728
rect 14185 13719 14243 13725
rect 14185 13716 14197 13719
rect 13964 13688 14197 13716
rect 13964 13676 13970 13688
rect 14185 13685 14197 13688
rect 14231 13716 14243 13719
rect 14831 13719 14889 13725
rect 14831 13716 14843 13719
rect 14231 13688 14843 13716
rect 14231 13685 14243 13688
rect 14185 13679 14243 13685
rect 14831 13685 14843 13688
rect 14877 13685 14889 13719
rect 19150 13716 19156 13728
rect 19111 13688 19156 13716
rect 14831 13679 14889 13685
rect 19150 13676 19156 13688
rect 19208 13676 19214 13728
rect 26878 13716 26884 13728
rect 26839 13688 26884 13716
rect 26878 13676 26884 13688
rect 26936 13676 26942 13728
rect 31938 13676 31944 13728
rect 31996 13716 32002 13728
rect 32490 13716 32496 13728
rect 31996 13688 32496 13716
rect 31996 13676 32002 13688
rect 32490 13676 32496 13688
rect 32548 13716 32554 13728
rect 32769 13719 32827 13725
rect 32769 13716 32781 13719
rect 32548 13688 32781 13716
rect 32548 13676 32554 13688
rect 32769 13685 32781 13688
rect 32815 13685 32827 13719
rect 33134 13716 33140 13728
rect 33095 13688 33140 13716
rect 32769 13679 32827 13685
rect 33134 13676 33140 13688
rect 33192 13676 33198 13728
rect 34701 13719 34759 13725
rect 34701 13685 34713 13719
rect 34747 13716 34759 13719
rect 35084 13716 35112 13815
rect 35342 13812 35348 13815
rect 35400 13812 35406 13824
rect 35820 13784 35848 13824
rect 35894 13784 35900 13796
rect 35820 13756 35900 13784
rect 35894 13744 35900 13756
rect 35952 13744 35958 13796
rect 35250 13716 35256 13728
rect 34747 13688 35256 13716
rect 34747 13685 34759 13688
rect 34701 13679 34759 13685
rect 35250 13676 35256 13688
rect 35308 13676 35314 13728
rect 1104 13626 38824 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 38824 13626
rect 1104 13552 38824 13574
rect 3878 13472 3884 13524
rect 3936 13512 3942 13524
rect 4249 13515 4307 13521
rect 4249 13512 4261 13515
rect 3936 13484 4261 13512
rect 3936 13472 3942 13484
rect 4249 13481 4261 13484
rect 4295 13481 4307 13515
rect 5074 13512 5080 13524
rect 5035 13484 5080 13512
rect 4249 13475 4307 13481
rect 5074 13472 5080 13484
rect 5132 13472 5138 13524
rect 6914 13512 6920 13524
rect 6875 13484 6920 13512
rect 6914 13472 6920 13484
rect 6972 13472 6978 13524
rect 8294 13512 8300 13524
rect 8255 13484 8300 13512
rect 8294 13472 8300 13484
rect 8352 13472 8358 13524
rect 9677 13515 9735 13521
rect 9677 13481 9689 13515
rect 9723 13512 9735 13515
rect 9858 13512 9864 13524
rect 9723 13484 9864 13512
rect 9723 13481 9735 13484
rect 9677 13475 9735 13481
rect 9858 13472 9864 13484
rect 9916 13472 9922 13524
rect 10042 13512 10048 13524
rect 10003 13484 10048 13512
rect 10042 13472 10048 13484
rect 10100 13472 10106 13524
rect 10870 13512 10876 13524
rect 10831 13484 10876 13512
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 12618 13512 12624 13524
rect 12579 13484 12624 13512
rect 12618 13472 12624 13484
rect 12676 13472 12682 13524
rect 13446 13472 13452 13524
rect 13504 13512 13510 13524
rect 13541 13515 13599 13521
rect 13541 13512 13553 13515
rect 13504 13484 13553 13512
rect 13504 13472 13510 13484
rect 13541 13481 13553 13484
rect 13587 13481 13599 13515
rect 14090 13512 14096 13524
rect 14051 13484 14096 13512
rect 13541 13475 13599 13481
rect 14090 13472 14096 13484
rect 14148 13472 14154 13524
rect 16666 13512 16672 13524
rect 16627 13484 16672 13512
rect 16666 13472 16672 13484
rect 16724 13472 16730 13524
rect 18509 13515 18567 13521
rect 18509 13481 18521 13515
rect 18555 13512 18567 13515
rect 18969 13515 19027 13521
rect 18969 13512 18981 13515
rect 18555 13484 18981 13512
rect 18555 13481 18567 13484
rect 18509 13475 18567 13481
rect 18969 13481 18981 13484
rect 19015 13512 19027 13515
rect 19150 13512 19156 13524
rect 19015 13484 19156 13512
rect 19015 13481 19027 13484
rect 18969 13475 19027 13481
rect 19150 13472 19156 13484
rect 19208 13472 19214 13524
rect 26970 13472 26976 13524
rect 27028 13512 27034 13524
rect 27893 13515 27951 13521
rect 27893 13512 27905 13515
rect 27028 13484 27905 13512
rect 27028 13472 27034 13484
rect 27893 13481 27905 13484
rect 27939 13481 27951 13515
rect 28994 13512 29000 13524
rect 28955 13484 29000 13512
rect 27893 13475 27951 13481
rect 28994 13472 29000 13484
rect 29052 13472 29058 13524
rect 29454 13512 29460 13524
rect 29415 13484 29460 13512
rect 29454 13472 29460 13484
rect 29512 13472 29518 13524
rect 30745 13515 30803 13521
rect 30745 13481 30757 13515
rect 30791 13512 30803 13515
rect 30834 13512 30840 13524
rect 30791 13484 30840 13512
rect 30791 13481 30803 13484
rect 30745 13475 30803 13481
rect 30834 13472 30840 13484
rect 30892 13472 30898 13524
rect 31297 13515 31355 13521
rect 31297 13481 31309 13515
rect 31343 13512 31355 13515
rect 31662 13512 31668 13524
rect 31343 13484 31668 13512
rect 31343 13481 31355 13484
rect 31297 13475 31355 13481
rect 31662 13472 31668 13484
rect 31720 13472 31726 13524
rect 31938 13512 31944 13524
rect 31899 13484 31944 13512
rect 31938 13472 31944 13484
rect 31996 13472 32002 13524
rect 32398 13512 32404 13524
rect 32359 13484 32404 13512
rect 32398 13472 32404 13484
rect 32456 13472 32462 13524
rect 32858 13512 32864 13524
rect 32771 13484 32864 13512
rect 32858 13472 32864 13484
rect 32916 13512 32922 13524
rect 33134 13512 33140 13524
rect 32916 13484 33140 13512
rect 32916 13472 32922 13484
rect 33134 13472 33140 13484
rect 33192 13472 33198 13524
rect 33410 13472 33416 13524
rect 33468 13512 33474 13524
rect 33781 13515 33839 13521
rect 33781 13512 33793 13515
rect 33468 13484 33793 13512
rect 33468 13472 33474 13484
rect 33781 13481 33793 13484
rect 33827 13512 33839 13515
rect 34885 13515 34943 13521
rect 34885 13512 34897 13515
rect 33827 13484 34897 13512
rect 33827 13481 33839 13484
rect 33781 13475 33839 13481
rect 34885 13481 34897 13484
rect 34931 13481 34943 13515
rect 36538 13512 36544 13524
rect 36499 13484 36544 13512
rect 34885 13475 34943 13481
rect 36538 13472 36544 13484
rect 36596 13472 36602 13524
rect 26694 13404 26700 13456
rect 26752 13453 26758 13456
rect 26752 13447 26816 13453
rect 26752 13413 26770 13447
rect 26804 13413 26816 13447
rect 26752 13407 26816 13413
rect 33229 13447 33287 13453
rect 33229 13413 33241 13447
rect 33275 13444 33287 13447
rect 33689 13447 33747 13453
rect 33689 13444 33701 13447
rect 33275 13416 33701 13444
rect 33275 13413 33287 13416
rect 33229 13407 33287 13413
rect 33689 13413 33701 13416
rect 33735 13444 33747 13447
rect 34422 13444 34428 13456
rect 33735 13416 34428 13444
rect 33735 13413 33747 13416
rect 33689 13407 33747 13413
rect 26752 13404 26758 13407
rect 34422 13404 34428 13416
rect 34480 13404 34486 13456
rect 4982 13376 4988 13388
rect 4943 13348 4988 13376
rect 4982 13336 4988 13348
rect 5040 13336 5046 13388
rect 8478 13376 8484 13388
rect 8439 13348 8484 13376
rect 8478 13336 8484 13348
rect 8536 13336 8542 13388
rect 9493 13379 9551 13385
rect 9493 13345 9505 13379
rect 9539 13376 9551 13379
rect 11497 13379 11555 13385
rect 11497 13376 11509 13379
rect 9539 13348 10364 13376
rect 9539 13345 9551 13348
rect 9493 13339 9551 13345
rect 5261 13311 5319 13317
rect 5261 13277 5273 13311
rect 5307 13308 5319 13311
rect 5350 13308 5356 13320
rect 5307 13280 5356 13308
rect 5307 13277 5319 13280
rect 5261 13271 5319 13277
rect 5350 13268 5356 13280
rect 5408 13268 5414 13320
rect 9398 13308 9404 13320
rect 8680 13280 9404 13308
rect 8680 13249 8708 13280
rect 9398 13268 9404 13280
rect 9456 13308 9462 13320
rect 10336 13317 10364 13348
rect 11072 13348 11509 13376
rect 11072 13320 11100 13348
rect 11497 13345 11509 13348
rect 11543 13345 11555 13379
rect 11497 13339 11555 13345
rect 15194 13336 15200 13388
rect 15252 13376 15258 13388
rect 15545 13379 15603 13385
rect 15545 13376 15557 13379
rect 15252 13348 15557 13376
rect 15252 13336 15258 13348
rect 15545 13345 15557 13348
rect 15591 13376 15603 13379
rect 16298 13376 16304 13388
rect 15591 13348 16304 13376
rect 15591 13345 15603 13348
rect 15545 13339 15603 13345
rect 16298 13336 16304 13348
rect 16356 13336 16362 13388
rect 18141 13379 18199 13385
rect 18141 13345 18153 13379
rect 18187 13376 18199 13379
rect 18187 13348 19196 13376
rect 18187 13345 18199 13348
rect 18141 13339 18199 13345
rect 19168 13320 19196 13348
rect 21082 13336 21088 13388
rect 21140 13376 21146 13388
rect 22186 13385 22192 13388
rect 21913 13379 21971 13385
rect 21913 13376 21925 13379
rect 21140 13348 21925 13376
rect 21140 13336 21146 13348
rect 21913 13345 21925 13348
rect 21959 13345 21971 13379
rect 22180 13376 22192 13385
rect 22147 13348 22192 13376
rect 21913 13339 21971 13345
rect 22180 13339 22192 13348
rect 22186 13336 22192 13339
rect 22244 13336 22250 13388
rect 26510 13376 26516 13388
rect 26471 13348 26516 13376
rect 26510 13336 26516 13348
rect 26568 13336 26574 13388
rect 29362 13376 29368 13388
rect 29323 13348 29368 13376
rect 29362 13336 29368 13348
rect 29420 13336 29426 13388
rect 30561 13379 30619 13385
rect 30561 13376 30573 13379
rect 30484 13348 30573 13376
rect 10137 13311 10195 13317
rect 10137 13308 10149 13311
rect 9456 13280 10149 13308
rect 9456 13268 9462 13280
rect 10137 13277 10149 13280
rect 10183 13277 10195 13311
rect 10137 13271 10195 13277
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13308 10379 13311
rect 11054 13308 11060 13320
rect 10367 13280 11060 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 11054 13268 11060 13280
rect 11112 13268 11118 13320
rect 11238 13268 11244 13320
rect 11296 13317 11302 13320
rect 11296 13308 11306 13317
rect 15289 13311 15347 13317
rect 11296 13280 11341 13308
rect 11296 13271 11306 13280
rect 15289 13277 15301 13311
rect 15335 13277 15347 13311
rect 15289 13271 15347 13277
rect 11296 13268 11302 13271
rect 8665 13243 8723 13249
rect 8665 13209 8677 13243
rect 8711 13209 8723 13243
rect 8665 13203 8723 13209
rect 15194 13200 15200 13252
rect 15252 13240 15258 13252
rect 15304 13240 15332 13271
rect 17954 13268 17960 13320
rect 18012 13308 18018 13320
rect 19058 13308 19064 13320
rect 18012 13280 19064 13308
rect 18012 13268 18018 13280
rect 19058 13268 19064 13280
rect 19116 13268 19122 13320
rect 19150 13268 19156 13320
rect 19208 13308 19214 13320
rect 29549 13311 29607 13317
rect 19208 13280 19301 13308
rect 19208 13268 19214 13280
rect 29549 13277 29561 13311
rect 29595 13277 29607 13311
rect 29549 13271 29607 13277
rect 15252 13212 15332 13240
rect 15252 13200 15258 13212
rect 4617 13175 4675 13181
rect 4617 13141 4629 13175
rect 4663 13172 4675 13175
rect 5442 13172 5448 13184
rect 4663 13144 5448 13172
rect 4663 13141 4675 13144
rect 4617 13135 4675 13141
rect 5442 13132 5448 13144
rect 5500 13132 5506 13184
rect 7374 13172 7380 13184
rect 7335 13144 7380 13172
rect 7374 13132 7380 13144
rect 7432 13132 7438 13184
rect 12434 13132 12440 13184
rect 12492 13172 12498 13184
rect 13262 13172 13268 13184
rect 12492 13144 13268 13172
rect 12492 13132 12498 13144
rect 13262 13132 13268 13144
rect 13320 13132 13326 13184
rect 14642 13172 14648 13184
rect 14603 13144 14648 13172
rect 14642 13132 14648 13144
rect 14700 13132 14706 13184
rect 15304 13172 15332 13212
rect 28905 13243 28963 13249
rect 28905 13209 28917 13243
rect 28951 13240 28963 13243
rect 29564 13240 29592 13271
rect 30374 13240 30380 13252
rect 28951 13212 30380 13240
rect 28951 13209 28963 13212
rect 28905 13203 28963 13209
rect 30374 13200 30380 13212
rect 30432 13200 30438 13252
rect 30484 13184 30512 13348
rect 30561 13345 30573 13348
rect 30607 13345 30619 13379
rect 32214 13376 32220 13388
rect 32175 13348 32220 13376
rect 30561 13339 30619 13345
rect 32214 13336 32220 13348
rect 32272 13336 32278 13388
rect 34330 13376 34336 13388
rect 34291 13348 34336 13376
rect 34330 13336 34336 13348
rect 34388 13336 34394 13388
rect 34793 13379 34851 13385
rect 34793 13345 34805 13379
rect 34839 13376 34851 13379
rect 35253 13379 35311 13385
rect 35253 13376 35265 13379
rect 34839 13348 35265 13376
rect 34839 13345 34851 13348
rect 34793 13339 34851 13345
rect 35253 13345 35265 13348
rect 35299 13376 35311 13379
rect 35986 13376 35992 13388
rect 35299 13348 35992 13376
rect 35299 13345 35311 13348
rect 35253 13339 35311 13345
rect 35986 13336 35992 13348
rect 36044 13336 36050 13388
rect 33965 13311 34023 13317
rect 33965 13277 33977 13311
rect 34011 13308 34023 13311
rect 34422 13308 34428 13320
rect 34011 13280 34428 13308
rect 34011 13277 34023 13280
rect 33965 13271 34023 13277
rect 34422 13268 34428 13280
rect 34480 13268 34486 13320
rect 35342 13308 35348 13320
rect 35303 13280 35348 13308
rect 35342 13268 35348 13280
rect 35400 13268 35406 13320
rect 35434 13268 35440 13320
rect 35492 13308 35498 13320
rect 35492 13280 35537 13308
rect 35492 13268 35498 13280
rect 33042 13200 33048 13252
rect 33100 13240 33106 13252
rect 33321 13243 33379 13249
rect 33321 13240 33333 13243
rect 33100 13212 33333 13240
rect 33100 13200 33106 13212
rect 33321 13209 33333 13212
rect 33367 13209 33379 13243
rect 33321 13203 33379 13209
rect 15470 13172 15476 13184
rect 15304 13144 15476 13172
rect 15470 13132 15476 13144
rect 15528 13132 15534 13184
rect 18601 13175 18659 13181
rect 18601 13141 18613 13175
rect 18647 13172 18659 13175
rect 19242 13172 19248 13184
rect 18647 13144 19248 13172
rect 18647 13141 18659 13144
rect 18601 13135 18659 13141
rect 19242 13132 19248 13144
rect 19300 13132 19306 13184
rect 21821 13175 21879 13181
rect 21821 13141 21833 13175
rect 21867 13172 21879 13175
rect 21910 13172 21916 13184
rect 21867 13144 21916 13172
rect 21867 13141 21879 13144
rect 21821 13135 21879 13141
rect 21910 13132 21916 13144
rect 21968 13132 21974 13184
rect 23290 13172 23296 13184
rect 23251 13144 23296 13172
rect 23290 13132 23296 13144
rect 23348 13132 23354 13184
rect 30466 13172 30472 13184
rect 30427 13144 30472 13172
rect 30466 13132 30472 13144
rect 30524 13132 30530 13184
rect 35986 13172 35992 13184
rect 35947 13144 35992 13172
rect 35986 13132 35992 13144
rect 36044 13132 36050 13184
rect 1104 13082 38824 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 38824 13082
rect 1104 13008 38824 13030
rect 3789 12971 3847 12977
rect 3789 12937 3801 12971
rect 3835 12968 3847 12971
rect 3878 12968 3884 12980
rect 3835 12940 3884 12968
rect 3835 12937 3847 12940
rect 3789 12931 3847 12937
rect 3878 12928 3884 12940
rect 3936 12928 3942 12980
rect 4982 12928 4988 12980
rect 5040 12968 5046 12980
rect 5261 12971 5319 12977
rect 5261 12968 5273 12971
rect 5040 12940 5273 12968
rect 5040 12928 5046 12940
rect 5261 12937 5273 12940
rect 5307 12937 5319 12971
rect 5261 12931 5319 12937
rect 6270 12928 6276 12980
rect 6328 12968 6334 12980
rect 6549 12971 6607 12977
rect 6549 12968 6561 12971
rect 6328 12940 6561 12968
rect 6328 12928 6334 12940
rect 6549 12937 6561 12940
rect 6595 12937 6607 12971
rect 6549 12931 6607 12937
rect 9033 12971 9091 12977
rect 9033 12937 9045 12971
rect 9079 12968 9091 12971
rect 10042 12968 10048 12980
rect 9079 12940 10048 12968
rect 9079 12937 9091 12940
rect 9033 12931 9091 12937
rect 3421 12835 3479 12841
rect 3421 12801 3433 12835
rect 3467 12832 3479 12835
rect 6564 12832 6592 12931
rect 10042 12928 10048 12940
rect 10100 12928 10106 12980
rect 11054 12928 11060 12980
rect 11112 12968 11118 12980
rect 11241 12971 11299 12977
rect 11241 12968 11253 12971
rect 11112 12940 11253 12968
rect 11112 12928 11118 12940
rect 11241 12937 11253 12940
rect 11287 12968 11299 12971
rect 12161 12971 12219 12977
rect 12161 12968 12173 12971
rect 11287 12940 12173 12968
rect 11287 12937 11299 12940
rect 11241 12931 11299 12937
rect 12161 12937 12173 12940
rect 12207 12937 12219 12971
rect 12161 12931 12219 12937
rect 15286 12928 15292 12980
rect 15344 12968 15350 12980
rect 15749 12971 15807 12977
rect 15749 12968 15761 12971
rect 15344 12940 15761 12968
rect 15344 12928 15350 12940
rect 15749 12937 15761 12940
rect 15795 12937 15807 12971
rect 19426 12968 19432 12980
rect 19387 12940 19432 12968
rect 15749 12931 15807 12937
rect 19426 12928 19432 12940
rect 19484 12928 19490 12980
rect 25682 12968 25688 12980
rect 25643 12940 25688 12968
rect 25682 12928 25688 12940
rect 25740 12928 25746 12980
rect 26510 12968 26516 12980
rect 26471 12940 26516 12968
rect 26510 12928 26516 12940
rect 26568 12928 26574 12980
rect 30466 12928 30472 12980
rect 30524 12968 30530 12980
rect 30837 12971 30895 12977
rect 30837 12968 30849 12971
rect 30524 12940 30849 12968
rect 30524 12928 30530 12940
rect 30837 12937 30849 12940
rect 30883 12937 30895 12971
rect 32214 12968 32220 12980
rect 32175 12940 32220 12968
rect 30837 12931 30895 12937
rect 32214 12928 32220 12940
rect 32272 12968 32278 12980
rect 32585 12971 32643 12977
rect 32585 12968 32597 12971
rect 32272 12940 32597 12968
rect 32272 12928 32278 12940
rect 32585 12937 32597 12940
rect 32631 12937 32643 12971
rect 32585 12931 32643 12937
rect 35894 12928 35900 12980
rect 35952 12968 35958 12980
rect 36541 12971 36599 12977
rect 36541 12968 36553 12971
rect 35952 12940 36553 12968
rect 35952 12928 35958 12940
rect 36541 12937 36553 12940
rect 36587 12937 36599 12971
rect 36541 12931 36599 12937
rect 9766 12900 9772 12912
rect 9727 12872 9772 12900
rect 9766 12860 9772 12872
rect 9824 12900 9830 12912
rect 9824 12872 9904 12900
rect 9824 12860 9830 12872
rect 9876 12841 9904 12872
rect 19058 12860 19064 12912
rect 19116 12900 19122 12912
rect 19981 12903 20039 12909
rect 19981 12900 19993 12903
rect 19116 12872 19993 12900
rect 19116 12860 19122 12872
rect 19981 12869 19993 12872
rect 20027 12869 20039 12903
rect 19981 12863 20039 12869
rect 7837 12835 7895 12841
rect 7837 12832 7849 12835
rect 3467 12804 4016 12832
rect 6564 12804 7849 12832
rect 3467 12801 3479 12804
rect 3421 12795 3479 12801
rect 3878 12764 3884 12776
rect 3839 12736 3884 12764
rect 3878 12724 3884 12736
rect 3936 12724 3942 12776
rect 3988 12764 4016 12804
rect 7837 12801 7849 12804
rect 7883 12801 7895 12835
rect 7837 12795 7895 12801
rect 9861 12835 9919 12841
rect 9861 12801 9873 12835
rect 9907 12801 9919 12835
rect 16298 12832 16304 12844
rect 16259 12804 16304 12832
rect 9861 12795 9919 12801
rect 4148 12767 4206 12773
rect 4148 12764 4160 12767
rect 3988 12736 4160 12764
rect 4148 12733 4160 12736
rect 4194 12764 4206 12767
rect 5074 12764 5080 12776
rect 4194 12736 5080 12764
rect 4194 12733 4206 12736
rect 4148 12727 4206 12733
rect 5074 12724 5080 12736
rect 5132 12724 5138 12776
rect 7374 12724 7380 12776
rect 7432 12764 7438 12776
rect 7653 12767 7711 12773
rect 7653 12764 7665 12767
rect 7432 12736 7665 12764
rect 7432 12724 7438 12736
rect 7653 12733 7665 12736
rect 7699 12764 7711 12767
rect 7926 12764 7932 12776
rect 7699 12736 7932 12764
rect 7699 12733 7711 12736
rect 7653 12727 7711 12733
rect 7926 12724 7932 12736
rect 7984 12724 7990 12776
rect 8478 12724 8484 12776
rect 8536 12764 8542 12776
rect 8573 12767 8631 12773
rect 8573 12764 8585 12767
rect 8536 12736 8585 12764
rect 8536 12724 8542 12736
rect 8573 12733 8585 12736
rect 8619 12764 8631 12767
rect 9582 12764 9588 12776
rect 8619 12736 9588 12764
rect 8619 12733 8631 12736
rect 8573 12727 8631 12733
rect 9582 12724 9588 12736
rect 9640 12724 9646 12776
rect 9876 12764 9904 12795
rect 16298 12792 16304 12804
rect 16356 12832 16362 12844
rect 16761 12835 16819 12841
rect 16761 12832 16773 12835
rect 16356 12804 16773 12832
rect 16356 12792 16362 12804
rect 16761 12801 16773 12804
rect 16807 12801 16819 12835
rect 16761 12795 16819 12801
rect 17770 12792 17776 12844
rect 17828 12832 17834 12844
rect 18049 12835 18107 12841
rect 18049 12832 18061 12835
rect 17828 12804 18061 12832
rect 17828 12792 17834 12804
rect 18049 12801 18061 12804
rect 18095 12801 18107 12835
rect 26528 12832 26556 12928
rect 29273 12903 29331 12909
rect 29273 12869 29285 12903
rect 29319 12900 29331 12903
rect 29362 12900 29368 12912
rect 29319 12872 29368 12900
rect 29319 12869 29331 12872
rect 29273 12863 29331 12869
rect 29362 12860 29368 12872
rect 29420 12900 29426 12912
rect 30285 12903 30343 12909
rect 30285 12900 30297 12903
rect 29420 12872 30297 12900
rect 29420 12860 29426 12872
rect 30285 12869 30297 12872
rect 30331 12869 30343 12903
rect 30285 12863 30343 12869
rect 26602 12832 26608 12844
rect 26515 12804 26608 12832
rect 18049 12795 18107 12801
rect 26602 12792 26608 12804
rect 26660 12792 26666 12844
rect 29822 12832 29828 12844
rect 29783 12804 29828 12832
rect 29822 12792 29828 12804
rect 29880 12792 29886 12844
rect 30374 12792 30380 12844
rect 30432 12832 30438 12844
rect 31389 12835 31447 12841
rect 31389 12832 31401 12835
rect 30432 12804 31401 12832
rect 30432 12792 30438 12804
rect 31389 12801 31401 12804
rect 31435 12832 31447 12835
rect 31938 12832 31944 12844
rect 31435 12804 31944 12832
rect 31435 12801 31447 12804
rect 31389 12795 31447 12801
rect 31938 12792 31944 12804
rect 31996 12832 32002 12844
rect 33229 12835 33287 12841
rect 33229 12832 33241 12835
rect 31996 12804 33241 12832
rect 31996 12792 32002 12804
rect 33229 12801 33241 12804
rect 33275 12832 33287 12835
rect 33318 12832 33324 12844
rect 33275 12804 33324 12832
rect 33275 12801 33287 12804
rect 33229 12795 33287 12801
rect 33318 12792 33324 12804
rect 33376 12832 33382 12844
rect 34422 12832 34428 12844
rect 33376 12804 34428 12832
rect 33376 12792 33382 12804
rect 34422 12792 34428 12804
rect 34480 12792 34486 12844
rect 11238 12764 11244 12776
rect 9876 12736 11244 12764
rect 11238 12724 11244 12736
rect 11296 12764 11302 12776
rect 11793 12767 11851 12773
rect 11793 12764 11805 12767
rect 11296 12736 11805 12764
rect 11296 12724 11302 12736
rect 11793 12733 11805 12736
rect 11839 12764 11851 12767
rect 13081 12767 13139 12773
rect 13081 12764 13093 12767
rect 11839 12736 13093 12764
rect 11839 12733 11851 12736
rect 11793 12727 11851 12733
rect 13081 12733 13093 12736
rect 13127 12764 13139 12767
rect 13265 12767 13323 12773
rect 13265 12764 13277 12767
rect 13127 12736 13277 12764
rect 13127 12733 13139 12736
rect 13081 12727 13139 12733
rect 13265 12733 13277 12736
rect 13311 12764 13323 12767
rect 15194 12764 15200 12776
rect 13311 12736 15200 12764
rect 13311 12733 13323 12736
rect 13265 12727 13323 12733
rect 15194 12724 15200 12736
rect 15252 12764 15258 12776
rect 15289 12767 15347 12773
rect 15289 12764 15301 12767
rect 15252 12736 15301 12764
rect 15252 12724 15258 12736
rect 15289 12733 15301 12736
rect 15335 12733 15347 12767
rect 16114 12764 16120 12776
rect 16075 12736 16120 12764
rect 15289 12727 15347 12733
rect 16114 12724 16120 12736
rect 16172 12724 16178 12776
rect 20441 12767 20499 12773
rect 20441 12733 20453 12767
rect 20487 12764 20499 12767
rect 20533 12767 20591 12773
rect 20533 12764 20545 12767
rect 20487 12736 20545 12764
rect 20487 12733 20499 12736
rect 20441 12727 20499 12733
rect 20533 12733 20545 12736
rect 20579 12764 20591 12767
rect 21082 12764 21088 12776
rect 20579 12736 21088 12764
rect 20579 12733 20591 12736
rect 20533 12727 20591 12733
rect 21082 12724 21088 12736
rect 21140 12764 21146 12776
rect 22462 12764 22468 12776
rect 21140 12736 22468 12764
rect 21140 12724 21146 12736
rect 22462 12724 22468 12736
rect 22520 12724 22526 12776
rect 35161 12767 35219 12773
rect 35161 12764 35173 12767
rect 34900 12736 35173 12764
rect 6822 12656 6828 12708
rect 6880 12696 6886 12708
rect 7193 12699 7251 12705
rect 7193 12696 7205 12699
rect 6880 12668 7205 12696
rect 6880 12656 6886 12668
rect 7193 12665 7205 12668
rect 7239 12696 7251 12699
rect 7745 12699 7803 12705
rect 7745 12696 7757 12699
rect 7239 12668 7757 12696
rect 7239 12665 7251 12668
rect 7193 12659 7251 12665
rect 7745 12665 7757 12668
rect 7791 12665 7803 12699
rect 7745 12659 7803 12665
rect 9401 12699 9459 12705
rect 9401 12665 9413 12699
rect 9447 12696 9459 12699
rect 10106 12699 10164 12705
rect 10106 12696 10118 12699
rect 9447 12668 10118 12696
rect 9447 12665 9459 12668
rect 9401 12659 9459 12665
rect 10106 12665 10118 12668
rect 10152 12696 10164 12699
rect 10410 12696 10416 12708
rect 10152 12668 10416 12696
rect 10152 12665 10164 12668
rect 10106 12659 10164 12665
rect 10410 12656 10416 12668
rect 10468 12656 10474 12708
rect 12805 12699 12863 12705
rect 12805 12665 12817 12699
rect 12851 12696 12863 12699
rect 13446 12696 13452 12708
rect 12851 12668 13452 12696
rect 12851 12665 12863 12668
rect 12805 12659 12863 12665
rect 13446 12656 13452 12668
rect 13504 12705 13510 12708
rect 13504 12699 13568 12705
rect 13504 12665 13522 12699
rect 13556 12665 13568 12699
rect 13504 12659 13568 12665
rect 13504 12656 13510 12659
rect 18230 12656 18236 12708
rect 18288 12705 18294 12708
rect 18288 12699 18352 12705
rect 18288 12665 18306 12699
rect 18340 12665 18352 12699
rect 18288 12659 18352 12665
rect 18288 12656 18294 12659
rect 19334 12656 19340 12708
rect 19392 12696 19398 12708
rect 20622 12696 20628 12708
rect 19392 12668 20628 12696
rect 19392 12656 19398 12668
rect 20622 12656 20628 12668
rect 20680 12696 20686 12708
rect 20778 12699 20836 12705
rect 20778 12696 20790 12699
rect 20680 12668 20790 12696
rect 20680 12656 20686 12668
rect 20778 12665 20790 12668
rect 20824 12665 20836 12699
rect 20778 12659 20836 12665
rect 21266 12656 21272 12708
rect 21324 12696 21330 12708
rect 22186 12696 22192 12708
rect 21324 12668 22192 12696
rect 21324 12656 21330 12668
rect 5350 12588 5356 12640
rect 5408 12628 5414 12640
rect 5813 12631 5871 12637
rect 5813 12628 5825 12631
rect 5408 12600 5825 12628
rect 5408 12588 5414 12600
rect 5813 12597 5825 12600
rect 5859 12628 5871 12631
rect 6638 12628 6644 12640
rect 5859 12600 6644 12628
rect 5859 12597 5871 12600
rect 5813 12591 5871 12597
rect 6638 12588 6644 12600
rect 6696 12628 6702 12640
rect 7098 12628 7104 12640
rect 6696 12600 7104 12628
rect 6696 12588 6702 12600
rect 7098 12588 7104 12600
rect 7156 12588 7162 12640
rect 7282 12628 7288 12640
rect 7243 12600 7288 12628
rect 7282 12588 7288 12600
rect 7340 12588 7346 12640
rect 13814 12588 13820 12640
rect 13872 12628 13878 12640
rect 14645 12631 14703 12637
rect 14645 12628 14657 12631
rect 13872 12600 14657 12628
rect 13872 12588 13878 12600
rect 14645 12597 14657 12600
rect 14691 12597 14703 12631
rect 16206 12628 16212 12640
rect 16167 12600 16212 12628
rect 14645 12591 14703 12597
rect 16206 12588 16212 12600
rect 16264 12588 16270 12640
rect 17770 12628 17776 12640
rect 17731 12600 17776 12628
rect 17770 12588 17776 12600
rect 17828 12588 17834 12640
rect 21928 12637 21956 12668
rect 22186 12656 22192 12668
rect 22244 12696 22250 12708
rect 22833 12699 22891 12705
rect 22833 12696 22845 12699
rect 22244 12668 22845 12696
rect 22244 12656 22250 12668
rect 22833 12665 22845 12668
rect 22879 12665 22891 12699
rect 22833 12659 22891 12665
rect 24305 12699 24363 12705
rect 24305 12665 24317 12699
rect 24351 12696 24363 12699
rect 24394 12696 24400 12708
rect 24351 12668 24400 12696
rect 24351 12665 24363 12668
rect 24305 12659 24363 12665
rect 24394 12656 24400 12668
rect 24452 12656 24458 12708
rect 26872 12699 26930 12705
rect 26872 12665 26884 12699
rect 26918 12696 26930 12699
rect 26970 12696 26976 12708
rect 26918 12668 26976 12696
rect 26918 12665 26930 12668
rect 26872 12659 26930 12665
rect 26970 12656 26976 12668
rect 27028 12656 27034 12708
rect 28718 12696 28724 12708
rect 28631 12668 28724 12696
rect 28718 12656 28724 12668
rect 28776 12696 28782 12708
rect 29641 12699 29699 12705
rect 29641 12696 29653 12699
rect 28776 12668 29653 12696
rect 28776 12656 28782 12668
rect 29641 12665 29653 12668
rect 29687 12665 29699 12699
rect 29641 12659 29699 12665
rect 30282 12656 30288 12708
rect 30340 12696 30346 12708
rect 30745 12699 30803 12705
rect 30745 12696 30757 12699
rect 30340 12668 30757 12696
rect 30340 12656 30346 12668
rect 30745 12665 30757 12668
rect 30791 12696 30803 12699
rect 31297 12699 31355 12705
rect 31297 12696 31309 12699
rect 30791 12668 31309 12696
rect 30791 12665 30803 12668
rect 30745 12659 30803 12665
rect 31297 12665 31309 12668
rect 31343 12665 31355 12699
rect 31297 12659 31355 12665
rect 32953 12699 33011 12705
rect 32953 12665 32965 12699
rect 32999 12696 33011 12699
rect 33594 12696 33600 12708
rect 32999 12668 33600 12696
rect 32999 12665 33011 12668
rect 32953 12659 33011 12665
rect 33594 12656 33600 12668
rect 33652 12656 33658 12708
rect 34900 12640 34928 12736
rect 35161 12733 35173 12736
rect 35207 12764 35219 12767
rect 35250 12764 35256 12776
rect 35207 12736 35256 12764
rect 35207 12733 35219 12736
rect 35161 12727 35219 12733
rect 35250 12724 35256 12736
rect 35308 12724 35314 12776
rect 35428 12767 35486 12773
rect 35428 12733 35440 12767
rect 35474 12764 35486 12767
rect 35986 12764 35992 12776
rect 35474 12736 35992 12764
rect 35474 12733 35486 12736
rect 35428 12727 35486 12733
rect 35986 12724 35992 12736
rect 36044 12724 36050 12776
rect 35710 12656 35716 12708
rect 35768 12656 35774 12708
rect 21913 12631 21971 12637
rect 21913 12597 21925 12631
rect 21959 12628 21971 12631
rect 21959 12600 21993 12628
rect 21959 12597 21971 12600
rect 21913 12591 21971 12597
rect 27614 12588 27620 12640
rect 27672 12628 27678 12640
rect 27985 12631 28043 12637
rect 27985 12628 27997 12631
rect 27672 12600 27997 12628
rect 27672 12588 27678 12600
rect 27985 12597 27997 12600
rect 28031 12628 28043 12631
rect 28997 12631 29055 12637
rect 28997 12628 29009 12631
rect 28031 12600 29009 12628
rect 28031 12597 28043 12600
rect 27985 12591 28043 12597
rect 28997 12597 29009 12600
rect 29043 12628 29055 12631
rect 29733 12631 29791 12637
rect 29733 12628 29745 12631
rect 29043 12600 29745 12628
rect 29043 12597 29055 12600
rect 28997 12591 29055 12597
rect 29733 12597 29745 12600
rect 29779 12597 29791 12631
rect 31202 12628 31208 12640
rect 31163 12600 31208 12628
rect 29733 12591 29791 12597
rect 31202 12588 31208 12600
rect 31260 12588 31266 12640
rect 31941 12631 31999 12637
rect 31941 12597 31953 12631
rect 31987 12628 31999 12631
rect 32306 12628 32312 12640
rect 31987 12600 32312 12628
rect 31987 12597 31999 12600
rect 31941 12591 31999 12597
rect 32306 12588 32312 12600
rect 32364 12628 32370 12640
rect 33045 12631 33103 12637
rect 33045 12628 33057 12631
rect 32364 12600 33057 12628
rect 32364 12588 32370 12600
rect 33045 12597 33057 12600
rect 33091 12597 33103 12631
rect 33045 12591 33103 12597
rect 34333 12631 34391 12637
rect 34333 12597 34345 12631
rect 34379 12628 34391 12631
rect 34514 12628 34520 12640
rect 34379 12600 34520 12628
rect 34379 12597 34391 12600
rect 34333 12591 34391 12597
rect 34514 12588 34520 12600
rect 34572 12588 34578 12640
rect 34701 12631 34759 12637
rect 34701 12597 34713 12631
rect 34747 12628 34759 12631
rect 34882 12628 34888 12640
rect 34747 12600 34888 12628
rect 34747 12597 34759 12600
rect 34701 12591 34759 12597
rect 34882 12588 34888 12600
rect 34940 12588 34946 12640
rect 35250 12588 35256 12640
rect 35308 12628 35314 12640
rect 35728 12628 35756 12656
rect 35308 12600 35756 12628
rect 35308 12588 35314 12600
rect 1104 12538 38824 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 38824 12538
rect 1104 12464 38824 12486
rect 4709 12427 4767 12433
rect 4709 12393 4721 12427
rect 4755 12424 4767 12427
rect 5074 12424 5080 12436
rect 4755 12396 5080 12424
rect 4755 12393 4767 12396
rect 4709 12387 4767 12393
rect 5074 12384 5080 12396
rect 5132 12384 5138 12436
rect 5442 12384 5448 12436
rect 5500 12424 5506 12436
rect 5629 12427 5687 12433
rect 5629 12424 5641 12427
rect 5500 12396 5641 12424
rect 5500 12384 5506 12396
rect 5629 12393 5641 12396
rect 5675 12393 5687 12427
rect 9398 12424 9404 12436
rect 9359 12396 9404 12424
rect 5629 12387 5687 12393
rect 9398 12384 9404 12396
rect 9456 12384 9462 12436
rect 9674 12424 9680 12436
rect 9635 12396 9680 12424
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 12713 12427 12771 12433
rect 12713 12393 12725 12427
rect 12759 12424 12771 12427
rect 12802 12424 12808 12436
rect 12759 12396 12808 12424
rect 12759 12393 12771 12396
rect 12713 12387 12771 12393
rect 12802 12384 12808 12396
rect 12860 12424 12866 12436
rect 13633 12427 13691 12433
rect 13633 12424 13645 12427
rect 12860 12396 13645 12424
rect 12860 12384 12866 12396
rect 13633 12393 13645 12396
rect 13679 12393 13691 12427
rect 16206 12424 16212 12436
rect 16167 12396 16212 12424
rect 13633 12387 13691 12393
rect 16206 12384 16212 12396
rect 16264 12384 16270 12436
rect 16669 12427 16727 12433
rect 16669 12393 16681 12427
rect 16715 12424 16727 12427
rect 17862 12424 17868 12436
rect 16715 12396 17868 12424
rect 16715 12393 16727 12396
rect 16669 12387 16727 12393
rect 17862 12384 17868 12396
rect 17920 12384 17926 12436
rect 20622 12424 20628 12436
rect 20583 12396 20628 12424
rect 20622 12384 20628 12396
rect 20680 12384 20686 12436
rect 26602 12384 26608 12436
rect 26660 12424 26666 12436
rect 26789 12427 26847 12433
rect 26789 12424 26801 12427
rect 26660 12396 26801 12424
rect 26660 12384 26666 12396
rect 26789 12393 26801 12396
rect 26835 12393 26847 12427
rect 26789 12387 26847 12393
rect 26970 12384 26976 12436
rect 27028 12424 27034 12436
rect 27433 12427 27491 12433
rect 27433 12424 27445 12427
rect 27028 12396 27445 12424
rect 27028 12384 27034 12396
rect 27433 12393 27445 12396
rect 27479 12393 27491 12427
rect 27433 12387 27491 12393
rect 29454 12384 29460 12436
rect 29512 12424 29518 12436
rect 29549 12427 29607 12433
rect 29549 12424 29561 12427
rect 29512 12396 29561 12424
rect 29512 12384 29518 12396
rect 29549 12393 29561 12396
rect 29595 12393 29607 12427
rect 29549 12387 29607 12393
rect 29822 12384 29828 12436
rect 29880 12424 29886 12436
rect 29917 12427 29975 12433
rect 29917 12424 29929 12427
rect 29880 12396 29929 12424
rect 29880 12384 29886 12396
rect 29917 12393 29929 12396
rect 29963 12393 29975 12427
rect 29917 12387 29975 12393
rect 30101 12427 30159 12433
rect 30101 12393 30113 12427
rect 30147 12424 30159 12427
rect 30282 12424 30288 12436
rect 30147 12396 30288 12424
rect 30147 12393 30159 12396
rect 30101 12387 30159 12393
rect 4982 12356 4988 12368
rect 4943 12328 4988 12356
rect 4982 12316 4988 12328
rect 5040 12316 5046 12368
rect 10410 12316 10416 12368
rect 10468 12356 10474 12368
rect 11425 12359 11483 12365
rect 11425 12356 11437 12359
rect 10468 12328 11437 12356
rect 10468 12316 10474 12328
rect 11425 12325 11437 12328
rect 11471 12325 11483 12359
rect 11425 12319 11483 12325
rect 15841 12359 15899 12365
rect 15841 12325 15853 12359
rect 15887 12356 15899 12359
rect 16114 12356 16120 12368
rect 15887 12328 16120 12356
rect 15887 12325 15899 12328
rect 15841 12319 15899 12325
rect 16114 12316 16120 12328
rect 16172 12316 16178 12368
rect 17037 12359 17095 12365
rect 17037 12325 17049 12359
rect 17083 12356 17095 12359
rect 17126 12356 17132 12368
rect 17083 12328 17132 12356
rect 17083 12325 17095 12328
rect 17037 12319 17095 12325
rect 17126 12316 17132 12328
rect 17184 12356 17190 12368
rect 18230 12356 18236 12368
rect 17184 12328 18236 12356
rect 17184 12316 17190 12328
rect 18230 12316 18236 12328
rect 18288 12316 18294 12368
rect 18500 12359 18558 12365
rect 18500 12356 18512 12359
rect 18340 12328 18512 12356
rect 4341 12291 4399 12297
rect 4341 12257 4353 12291
rect 4387 12288 4399 12291
rect 4706 12288 4712 12300
rect 4387 12260 4712 12288
rect 4387 12257 4399 12260
rect 4341 12251 4399 12257
rect 4706 12248 4712 12260
rect 4764 12288 4770 12300
rect 5537 12291 5595 12297
rect 5537 12288 5549 12291
rect 4764 12260 5549 12288
rect 4764 12248 4770 12260
rect 5537 12257 5549 12260
rect 5583 12257 5595 12291
rect 5537 12251 5595 12257
rect 6733 12291 6791 12297
rect 6733 12257 6745 12291
rect 6779 12257 6791 12291
rect 6733 12251 6791 12257
rect 5813 12223 5871 12229
rect 5813 12189 5825 12223
rect 5859 12220 5871 12223
rect 6270 12220 6276 12232
rect 5859 12192 6276 12220
rect 5859 12189 5871 12192
rect 5813 12183 5871 12189
rect 6270 12180 6276 12192
rect 6328 12180 6334 12232
rect 5169 12155 5227 12161
rect 5169 12121 5181 12155
rect 5215 12152 5227 12155
rect 6748 12152 6776 12251
rect 8294 12248 8300 12300
rect 8352 12288 8358 12300
rect 8389 12291 8447 12297
rect 8389 12288 8401 12291
rect 8352 12260 8401 12288
rect 8352 12248 8358 12260
rect 8389 12257 8401 12260
rect 8435 12257 8447 12291
rect 10045 12291 10103 12297
rect 10045 12288 10057 12291
rect 8389 12251 8447 12257
rect 9048 12260 10057 12288
rect 8478 12220 8484 12232
rect 8439 12192 8484 12220
rect 8478 12180 8484 12192
rect 8536 12180 8542 12232
rect 8662 12220 8668 12232
rect 8623 12192 8668 12220
rect 8662 12180 8668 12192
rect 8720 12180 8726 12232
rect 7285 12155 7343 12161
rect 7285 12152 7297 12155
rect 5215 12124 7297 12152
rect 5215 12121 5227 12124
rect 5169 12115 5227 12121
rect 7285 12121 7297 12124
rect 7331 12121 7343 12155
rect 7285 12115 7343 12121
rect 6914 12084 6920 12096
rect 6875 12056 6920 12084
rect 6914 12044 6920 12056
rect 6972 12044 6978 12096
rect 7098 12044 7104 12096
rect 7156 12084 7162 12096
rect 7466 12084 7472 12096
rect 7156 12056 7472 12084
rect 7156 12044 7162 12056
rect 7466 12044 7472 12056
rect 7524 12084 7530 12096
rect 9048 12093 9076 12260
rect 10045 12257 10057 12260
rect 10091 12288 10103 12291
rect 11054 12288 11060 12300
rect 10091 12260 11060 12288
rect 10091 12257 10103 12260
rect 10045 12251 10103 12257
rect 11054 12248 11060 12260
rect 11112 12248 11118 12300
rect 11238 12288 11244 12300
rect 11199 12260 11244 12288
rect 11238 12248 11244 12260
rect 11296 12248 11302 12300
rect 12710 12248 12716 12300
rect 12768 12288 12774 12300
rect 13541 12291 13599 12297
rect 13541 12288 13553 12291
rect 12768 12260 13553 12288
rect 12768 12248 12774 12260
rect 13541 12257 13553 12260
rect 13587 12288 13599 12291
rect 15289 12291 15347 12297
rect 15289 12288 15301 12291
rect 13587 12260 15301 12288
rect 13587 12257 13599 12260
rect 13541 12251 13599 12257
rect 15289 12257 15301 12260
rect 15335 12257 15347 12291
rect 18340 12288 18368 12328
rect 18500 12325 18512 12328
rect 18546 12356 18558 12359
rect 18690 12356 18696 12368
rect 18546 12328 18696 12356
rect 18546 12325 18558 12328
rect 18500 12319 18558 12325
rect 18690 12316 18696 12328
rect 18748 12316 18754 12368
rect 21453 12359 21511 12365
rect 21453 12325 21465 12359
rect 21499 12356 21511 12359
rect 22646 12356 22652 12368
rect 21499 12328 22652 12356
rect 21499 12325 21511 12328
rect 21453 12319 21511 12325
rect 22646 12316 22652 12328
rect 22704 12356 22710 12368
rect 22916 12359 22974 12365
rect 22916 12356 22928 12359
rect 22704 12328 22928 12356
rect 22704 12316 22710 12328
rect 22916 12325 22928 12328
rect 22962 12356 22974 12359
rect 23290 12356 23296 12368
rect 22962 12328 23296 12356
rect 22962 12325 22974 12328
rect 22916 12319 22974 12325
rect 23290 12316 23296 12328
rect 23348 12316 23354 12368
rect 26694 12316 26700 12368
rect 26752 12356 26758 12368
rect 27065 12359 27123 12365
rect 27065 12356 27077 12359
rect 26752 12328 27077 12356
rect 26752 12316 26758 12328
rect 27065 12325 27077 12328
rect 27111 12325 27123 12359
rect 27065 12319 27123 12325
rect 27884 12359 27942 12365
rect 27884 12325 27896 12359
rect 27930 12356 27942 12359
rect 28074 12356 28080 12368
rect 27930 12328 28080 12356
rect 27930 12325 27942 12328
rect 27884 12319 27942 12325
rect 28074 12316 28080 12328
rect 28132 12356 28138 12368
rect 28718 12356 28724 12368
rect 28132 12328 28724 12356
rect 28132 12316 28138 12328
rect 28718 12316 28724 12328
rect 28776 12316 28782 12368
rect 29932 12356 29960 12387
rect 30282 12384 30288 12396
rect 30340 12384 30346 12436
rect 31573 12427 31631 12433
rect 31573 12393 31585 12427
rect 31619 12424 31631 12427
rect 31849 12427 31907 12433
rect 31849 12424 31861 12427
rect 31619 12396 31861 12424
rect 31619 12393 31631 12396
rect 31573 12387 31631 12393
rect 31849 12393 31861 12396
rect 31895 12424 31907 12427
rect 31938 12424 31944 12436
rect 31895 12396 31944 12424
rect 31895 12393 31907 12396
rect 31849 12387 31907 12393
rect 31938 12384 31944 12396
rect 31996 12384 32002 12436
rect 32585 12427 32643 12433
rect 32585 12393 32597 12427
rect 32631 12424 32643 12427
rect 32858 12424 32864 12436
rect 32631 12396 32864 12424
rect 32631 12393 32643 12396
rect 32585 12387 32643 12393
rect 32858 12384 32864 12396
rect 32916 12384 32922 12436
rect 33042 12424 33048 12436
rect 33003 12396 33048 12424
rect 33042 12384 33048 12396
rect 33100 12384 33106 12436
rect 33410 12424 33416 12436
rect 33371 12396 33416 12424
rect 33410 12384 33416 12396
rect 33468 12384 33474 12436
rect 33505 12427 33563 12433
rect 33505 12393 33517 12427
rect 33551 12424 33563 12427
rect 33594 12424 33600 12436
rect 33551 12396 33600 12424
rect 33551 12393 33563 12396
rect 33505 12387 33563 12393
rect 33594 12384 33600 12396
rect 33652 12384 33658 12436
rect 34054 12384 34060 12436
rect 34112 12424 34118 12436
rect 34330 12424 34336 12436
rect 34112 12396 34336 12424
rect 34112 12384 34118 12396
rect 34330 12384 34336 12396
rect 34388 12424 34394 12436
rect 34609 12427 34667 12433
rect 34609 12424 34621 12427
rect 34388 12396 34621 12424
rect 34388 12384 34394 12396
rect 34609 12393 34621 12396
rect 34655 12393 34667 12427
rect 34609 12387 34667 12393
rect 35342 12384 35348 12436
rect 35400 12424 35406 12436
rect 35400 12396 35471 12424
rect 35400 12384 35406 12396
rect 29932 12328 30604 12356
rect 15289 12251 15347 12257
rect 17144 12260 18368 12288
rect 9490 12180 9496 12232
rect 9548 12220 9554 12232
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 9548 12192 10149 12220
rect 9548 12180 9554 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12220 10379 12223
rect 13081 12223 13139 12229
rect 10367 12192 10824 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 10796 12093 10824 12192
rect 13081 12189 13093 12223
rect 13127 12220 13139 12223
rect 13722 12220 13728 12232
rect 13127 12192 13728 12220
rect 13127 12189 13139 12192
rect 13081 12183 13139 12189
rect 13722 12180 13728 12192
rect 13780 12180 13786 12232
rect 16758 12180 16764 12232
rect 16816 12220 16822 12232
rect 17144 12229 17172 12260
rect 22462 12248 22468 12300
rect 22520 12288 22526 12300
rect 30466 12288 30472 12300
rect 22520 12260 22692 12288
rect 30427 12260 30472 12288
rect 22520 12248 22526 12260
rect 17129 12223 17187 12229
rect 17129 12220 17141 12223
rect 16816 12192 17141 12220
rect 16816 12180 16822 12192
rect 17129 12189 17141 12192
rect 17175 12189 17187 12223
rect 17129 12183 17187 12189
rect 17313 12223 17371 12229
rect 17313 12189 17325 12223
rect 17359 12220 17371 12223
rect 17494 12220 17500 12232
rect 17359 12192 17500 12220
rect 17359 12189 17371 12192
rect 17313 12183 17371 12189
rect 17494 12180 17500 12192
rect 17552 12180 17558 12232
rect 17770 12180 17776 12232
rect 17828 12220 17834 12232
rect 18233 12223 18291 12229
rect 18233 12220 18245 12223
rect 17828 12192 18245 12220
rect 17828 12180 17834 12192
rect 18233 12189 18245 12192
rect 18279 12189 18291 12223
rect 18233 12183 18291 12189
rect 21266 12180 21272 12232
rect 21324 12220 21330 12232
rect 22664 12229 22692 12260
rect 30466 12248 30472 12260
rect 30524 12248 30530 12300
rect 30576 12288 30604 12328
rect 32401 12291 32459 12297
rect 30576 12260 30696 12288
rect 21545 12223 21603 12229
rect 21545 12220 21557 12223
rect 21324 12192 21557 12220
rect 21324 12180 21330 12192
rect 21545 12189 21557 12192
rect 21591 12189 21603 12223
rect 21545 12183 21603 12189
rect 21729 12223 21787 12229
rect 21729 12189 21741 12223
rect 21775 12220 21787 12223
rect 22649 12223 22707 12229
rect 21775 12192 22600 12220
rect 21775 12189 21787 12192
rect 21729 12183 21787 12189
rect 22572 12096 22600 12192
rect 22649 12189 22661 12223
rect 22695 12189 22707 12223
rect 22649 12183 22707 12189
rect 26602 12180 26608 12232
rect 26660 12220 26666 12232
rect 27614 12220 27620 12232
rect 26660 12192 27620 12220
rect 26660 12180 26666 12192
rect 27614 12180 27620 12192
rect 27672 12180 27678 12232
rect 30190 12220 30196 12232
rect 29012 12192 30196 12220
rect 29012 12161 29040 12192
rect 30190 12180 30196 12192
rect 30248 12220 30254 12232
rect 30668 12229 30696 12260
rect 32401 12257 32413 12291
rect 32447 12288 32459 12291
rect 33060 12288 33088 12384
rect 34514 12316 34520 12368
rect 34572 12356 34578 12368
rect 35443 12356 35471 12396
rect 35986 12384 35992 12436
rect 36044 12424 36050 12436
rect 36541 12427 36599 12433
rect 36541 12424 36553 12427
rect 36044 12396 36553 12424
rect 36044 12384 36050 12396
rect 36541 12393 36553 12396
rect 36587 12393 36599 12427
rect 36541 12387 36599 12393
rect 34572 12328 35471 12356
rect 34572 12316 34578 12328
rect 33870 12288 33876 12300
rect 32447 12260 33088 12288
rect 33831 12260 33876 12288
rect 32447 12257 32459 12260
rect 32401 12251 32459 12257
rect 33870 12248 33876 12260
rect 33928 12248 33934 12300
rect 35443 12297 35471 12328
rect 35428 12291 35486 12297
rect 35428 12257 35440 12291
rect 35474 12288 35486 12291
rect 36262 12288 36268 12300
rect 35474 12260 36268 12288
rect 35474 12257 35486 12260
rect 35428 12251 35486 12257
rect 36262 12248 36268 12260
rect 36320 12248 36326 12300
rect 30561 12223 30619 12229
rect 30561 12220 30573 12223
rect 30248 12192 30573 12220
rect 30248 12180 30254 12192
rect 30561 12189 30573 12192
rect 30607 12189 30619 12223
rect 30561 12183 30619 12189
rect 30653 12223 30711 12229
rect 30653 12189 30665 12223
rect 30699 12220 30711 12223
rect 30834 12220 30840 12232
rect 30699 12192 30840 12220
rect 30699 12189 30711 12192
rect 30653 12183 30711 12189
rect 30834 12180 30840 12192
rect 30892 12180 30898 12232
rect 33962 12220 33968 12232
rect 33923 12192 33968 12220
rect 33962 12180 33968 12192
rect 34020 12180 34026 12232
rect 34149 12223 34207 12229
rect 34149 12189 34161 12223
rect 34195 12220 34207 12223
rect 34330 12220 34336 12232
rect 34195 12192 34336 12220
rect 34195 12189 34207 12192
rect 34149 12183 34207 12189
rect 34330 12180 34336 12192
rect 34388 12180 34394 12232
rect 34606 12220 34612 12232
rect 34440 12192 34612 12220
rect 28997 12155 29055 12161
rect 28997 12121 29009 12155
rect 29043 12121 29055 12155
rect 28997 12115 29055 12121
rect 34440 12096 34468 12192
rect 34606 12180 34612 12192
rect 34664 12180 34670 12232
rect 34882 12180 34888 12232
rect 34940 12220 34946 12232
rect 35161 12223 35219 12229
rect 35161 12220 35173 12223
rect 34940 12192 35173 12220
rect 34940 12180 34946 12192
rect 7653 12087 7711 12093
rect 7653 12084 7665 12087
rect 7524 12056 7665 12084
rect 7524 12044 7530 12056
rect 7653 12053 7665 12056
rect 7699 12053 7711 12087
rect 7653 12047 7711 12053
rect 8021 12087 8079 12093
rect 8021 12053 8033 12087
rect 8067 12084 8079 12087
rect 9033 12087 9091 12093
rect 9033 12084 9045 12087
rect 8067 12056 9045 12084
rect 8067 12053 8079 12056
rect 8021 12047 8079 12053
rect 9033 12053 9045 12056
rect 9079 12053 9091 12087
rect 9033 12047 9091 12053
rect 10781 12087 10839 12093
rect 10781 12053 10793 12087
rect 10827 12084 10839 12087
rect 10962 12084 10968 12096
rect 10827 12056 10968 12084
rect 10827 12053 10839 12056
rect 10781 12047 10839 12053
rect 10962 12044 10968 12056
rect 11020 12044 11026 12096
rect 11054 12044 11060 12096
rect 11112 12084 11118 12096
rect 11609 12087 11667 12093
rect 11609 12084 11621 12087
rect 11112 12056 11621 12084
rect 11112 12044 11118 12056
rect 11609 12053 11621 12056
rect 11655 12053 11667 12087
rect 13170 12084 13176 12096
rect 13131 12056 13176 12084
rect 11609 12047 11667 12053
rect 13170 12044 13176 12056
rect 13228 12044 13234 12096
rect 15010 12084 15016 12096
rect 14971 12056 15016 12084
rect 15010 12044 15016 12056
rect 15068 12044 15074 12096
rect 18141 12087 18199 12093
rect 18141 12053 18153 12087
rect 18187 12084 18199 12087
rect 18230 12084 18236 12096
rect 18187 12056 18236 12084
rect 18187 12053 18199 12056
rect 18141 12047 18199 12053
rect 18230 12044 18236 12056
rect 18288 12084 18294 12096
rect 19613 12087 19671 12093
rect 19613 12084 19625 12087
rect 18288 12056 19625 12084
rect 18288 12044 18294 12056
rect 19613 12053 19625 12056
rect 19659 12053 19671 12087
rect 21082 12084 21088 12096
rect 21043 12056 21088 12084
rect 19613 12047 19671 12053
rect 21082 12044 21088 12056
rect 21140 12044 21146 12096
rect 22186 12084 22192 12096
rect 22147 12056 22192 12084
rect 22186 12044 22192 12056
rect 22244 12044 22250 12096
rect 22554 12084 22560 12096
rect 22515 12056 22560 12084
rect 22554 12044 22560 12056
rect 22612 12044 22618 12096
rect 23934 12044 23940 12096
rect 23992 12084 23998 12096
rect 24029 12087 24087 12093
rect 24029 12084 24041 12087
rect 23992 12056 24041 12084
rect 23992 12044 23998 12056
rect 24029 12053 24041 12056
rect 24075 12053 24087 12087
rect 24029 12047 24087 12053
rect 30374 12044 30380 12096
rect 30432 12084 30438 12096
rect 31113 12087 31171 12093
rect 31113 12084 31125 12087
rect 30432 12056 31125 12084
rect 30432 12044 30438 12056
rect 31113 12053 31125 12056
rect 31159 12084 31171 12087
rect 31202 12084 31208 12096
rect 31159 12056 31208 12084
rect 31159 12053 31171 12056
rect 31113 12047 31171 12053
rect 31202 12044 31208 12056
rect 31260 12044 31266 12096
rect 34422 12044 34428 12096
rect 34480 12044 34486 12096
rect 34606 12044 34612 12096
rect 34664 12084 34670 12096
rect 34992 12093 35020 12192
rect 35161 12189 35173 12192
rect 35207 12189 35219 12223
rect 35161 12183 35219 12189
rect 34977 12087 35035 12093
rect 34977 12084 34989 12087
rect 34664 12056 34989 12084
rect 34664 12044 34670 12056
rect 34977 12053 34989 12056
rect 35023 12053 35035 12087
rect 34977 12047 35035 12053
rect 1104 11994 38824 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 38824 11994
rect 1104 11920 38824 11942
rect 3878 11880 3884 11892
rect 3839 11852 3884 11880
rect 3878 11840 3884 11852
rect 3936 11840 3942 11892
rect 6822 11880 6828 11892
rect 6783 11852 6828 11880
rect 6822 11840 6828 11852
rect 6880 11840 6886 11892
rect 6914 11840 6920 11892
rect 6972 11880 6978 11892
rect 8021 11883 8079 11889
rect 8021 11880 8033 11883
rect 6972 11852 8033 11880
rect 6972 11840 6978 11852
rect 8021 11849 8033 11852
rect 8067 11880 8079 11883
rect 8478 11880 8484 11892
rect 8067 11852 8484 11880
rect 8067 11849 8079 11852
rect 8021 11843 8079 11849
rect 8478 11840 8484 11852
rect 8536 11840 8542 11892
rect 8941 11883 8999 11889
rect 8941 11849 8953 11883
rect 8987 11880 8999 11883
rect 9030 11880 9036 11892
rect 8987 11852 9036 11880
rect 8987 11849 8999 11852
rect 8941 11843 8999 11849
rect 9030 11840 9036 11852
rect 9088 11880 9094 11892
rect 9766 11880 9772 11892
rect 9088 11852 9772 11880
rect 9088 11840 9094 11852
rect 9766 11840 9772 11852
rect 9824 11840 9830 11892
rect 10410 11880 10416 11892
rect 10371 11852 10416 11880
rect 10410 11840 10416 11852
rect 10468 11880 10474 11892
rect 11609 11883 11667 11889
rect 11609 11880 11621 11883
rect 10468 11852 11621 11880
rect 10468 11840 10474 11852
rect 11609 11849 11621 11852
rect 11655 11849 11667 11883
rect 12710 11880 12716 11892
rect 12671 11852 12716 11880
rect 11609 11843 11667 11849
rect 12710 11840 12716 11852
rect 12768 11840 12774 11892
rect 16758 11880 16764 11892
rect 16719 11852 16764 11880
rect 16758 11840 16764 11852
rect 16816 11840 16822 11892
rect 17126 11880 17132 11892
rect 17087 11852 17132 11880
rect 17126 11840 17132 11852
rect 17184 11840 17190 11892
rect 20622 11880 20628 11892
rect 20583 11852 20628 11880
rect 20622 11840 20628 11852
rect 20680 11840 20686 11892
rect 21266 11880 21272 11892
rect 21227 11852 21272 11880
rect 21266 11840 21272 11852
rect 21324 11840 21330 11892
rect 21726 11880 21732 11892
rect 21687 11852 21732 11880
rect 21726 11840 21732 11852
rect 21784 11840 21790 11892
rect 22462 11840 22468 11892
rect 22520 11880 22526 11892
rect 23017 11883 23075 11889
rect 23017 11880 23029 11883
rect 22520 11852 23029 11880
rect 22520 11840 22526 11852
rect 23017 11849 23029 11852
rect 23063 11880 23075 11883
rect 23385 11883 23443 11889
rect 23385 11880 23397 11883
rect 23063 11852 23397 11880
rect 23063 11849 23075 11852
rect 23017 11843 23075 11849
rect 23385 11849 23397 11852
rect 23431 11880 23443 11883
rect 26602 11880 26608 11892
rect 23431 11852 26608 11880
rect 23431 11849 23443 11852
rect 23385 11843 23443 11849
rect 3513 11747 3571 11753
rect 3513 11713 3525 11747
rect 3559 11744 3571 11747
rect 7466 11744 7472 11756
rect 3559 11716 4108 11744
rect 7427 11716 7472 11744
rect 3559 11713 3571 11716
rect 3513 11707 3571 11713
rect 3878 11636 3884 11688
rect 3936 11676 3942 11688
rect 3973 11679 4031 11685
rect 3973 11676 3985 11679
rect 3936 11648 3985 11676
rect 3936 11636 3942 11648
rect 3973 11645 3985 11648
rect 4019 11645 4031 11679
rect 4080 11676 4108 11716
rect 7466 11704 7472 11716
rect 7524 11704 7530 11756
rect 12253 11747 12311 11753
rect 12253 11713 12265 11747
rect 12299 11744 12311 11747
rect 22554 11744 22560 11756
rect 12299 11716 13308 11744
rect 22515 11716 22560 11744
rect 12299 11713 12311 11716
rect 12253 11707 12311 11713
rect 4240 11679 4298 11685
rect 4240 11676 4252 11679
rect 4080 11648 4252 11676
rect 3973 11639 4031 11645
rect 4240 11645 4252 11648
rect 4286 11676 4298 11679
rect 4982 11676 4988 11688
rect 4286 11648 4988 11676
rect 4286 11645 4298 11648
rect 4240 11639 4298 11645
rect 4982 11636 4988 11648
rect 5040 11636 5046 11688
rect 8110 11636 8116 11688
rect 8168 11676 8174 11688
rect 9030 11676 9036 11688
rect 8168 11648 9036 11676
rect 8168 11636 8174 11648
rect 9030 11636 9036 11648
rect 9088 11636 9094 11688
rect 13173 11679 13231 11685
rect 13173 11645 13185 11679
rect 13219 11645 13231 11679
rect 13280 11676 13308 11716
rect 22554 11704 22560 11716
rect 22612 11704 22618 11756
rect 23400 11744 23428 11843
rect 26602 11840 26608 11852
rect 26660 11840 26666 11892
rect 28074 11880 28080 11892
rect 28035 11852 28080 11880
rect 28074 11840 28080 11852
rect 28132 11840 28138 11892
rect 30834 11840 30840 11892
rect 30892 11880 30898 11892
rect 31389 11883 31447 11889
rect 31389 11880 31401 11883
rect 30892 11852 31401 11880
rect 30892 11840 30898 11852
rect 31389 11849 31401 11852
rect 31435 11849 31447 11883
rect 32306 11880 32312 11892
rect 32267 11852 32312 11880
rect 31389 11843 31447 11849
rect 23661 11747 23719 11753
rect 23661 11744 23673 11747
rect 23400 11716 23673 11744
rect 23661 11713 23673 11716
rect 23707 11713 23719 11747
rect 26620 11744 26648 11840
rect 26697 11747 26755 11753
rect 26697 11744 26709 11747
rect 26620 11716 26709 11744
rect 23661 11707 23719 11713
rect 26697 11713 26709 11716
rect 26743 11713 26755 11747
rect 31404 11744 31432 11843
rect 32306 11840 32312 11852
rect 32364 11840 32370 11892
rect 33597 11883 33655 11889
rect 33597 11849 33609 11883
rect 33643 11880 33655 11883
rect 33962 11880 33968 11892
rect 33643 11852 33968 11880
rect 33643 11849 33655 11852
rect 33597 11843 33655 11849
rect 33962 11840 33968 11852
rect 34020 11840 34026 11892
rect 34330 11840 34336 11892
rect 34388 11840 34394 11892
rect 36262 11880 36268 11892
rect 36175 11852 36268 11880
rect 36262 11840 36268 11852
rect 36320 11880 36326 11892
rect 36817 11883 36875 11889
rect 36817 11880 36829 11883
rect 36320 11852 36829 11880
rect 36320 11840 36326 11852
rect 36817 11849 36829 11852
rect 36863 11849 36875 11883
rect 36817 11843 36875 11849
rect 34348 11812 34376 11840
rect 32968 11784 34376 11812
rect 32968 11753 32996 11784
rect 32953 11747 33011 11753
rect 32953 11744 32965 11747
rect 31404 11716 32965 11744
rect 26697 11707 26755 11713
rect 32953 11713 32965 11716
rect 32999 11713 33011 11747
rect 32953 11707 33011 11713
rect 33870 11704 33876 11756
rect 33928 11744 33934 11756
rect 33965 11747 34023 11753
rect 33965 11744 33977 11747
rect 33928 11716 33977 11744
rect 33928 11704 33934 11716
rect 33965 11713 33977 11716
rect 34011 11744 34023 11747
rect 34333 11747 34391 11753
rect 34333 11744 34345 11747
rect 34011 11716 34345 11744
rect 34011 11713 34023 11716
rect 33965 11707 34023 11713
rect 34333 11713 34345 11716
rect 34379 11744 34391 11747
rect 34379 11716 35020 11744
rect 34379 11713 34391 11716
rect 34333 11707 34391 11713
rect 13440 11679 13498 11685
rect 13440 11676 13452 11679
rect 13280 11648 13452 11676
rect 13173 11639 13231 11645
rect 13440 11645 13452 11648
rect 13486 11676 13498 11679
rect 13722 11676 13728 11688
rect 13486 11648 13728 11676
rect 13486 11645 13498 11648
rect 13440 11639 13498 11645
rect 6638 11608 6644 11620
rect 6551 11580 6644 11608
rect 6638 11568 6644 11580
rect 6696 11608 6702 11620
rect 9306 11617 9312 11620
rect 7285 11611 7343 11617
rect 7285 11608 7297 11611
rect 6696 11580 7297 11608
rect 6696 11568 6702 11580
rect 7285 11577 7297 11580
rect 7331 11577 7343 11611
rect 9300 11608 9312 11617
rect 9267 11580 9312 11608
rect 7285 11571 7343 11577
rect 9300 11571 9312 11580
rect 9306 11568 9312 11571
rect 9364 11568 9370 11620
rect 12710 11568 12716 11620
rect 12768 11608 12774 11620
rect 12989 11611 13047 11617
rect 12989 11608 13001 11611
rect 12768 11580 13001 11608
rect 12768 11568 12774 11580
rect 12989 11577 13001 11580
rect 13035 11608 13047 11611
rect 13188 11608 13216 11639
rect 13722 11636 13728 11648
rect 13780 11636 13786 11688
rect 19245 11679 19303 11685
rect 19245 11645 19257 11679
rect 19291 11645 19303 11679
rect 21910 11676 21916 11688
rect 21871 11648 21916 11676
rect 19245 11639 19303 11645
rect 19061 11611 19119 11617
rect 19061 11608 19073 11611
rect 13035 11580 13216 11608
rect 18248 11580 19073 11608
rect 13035 11577 13047 11580
rect 12989 11571 13047 11577
rect 5166 11500 5172 11552
rect 5224 11540 5230 11552
rect 5353 11543 5411 11549
rect 5353 11540 5365 11543
rect 5224 11512 5365 11540
rect 5224 11500 5230 11512
rect 5353 11509 5365 11512
rect 5399 11509 5411 11543
rect 5353 11503 5411 11509
rect 6273 11543 6331 11549
rect 6273 11509 6285 11543
rect 6319 11540 6331 11543
rect 7193 11543 7251 11549
rect 7193 11540 7205 11543
rect 6319 11512 7205 11540
rect 6319 11509 6331 11512
rect 6273 11503 6331 11509
rect 7193 11509 7205 11512
rect 7239 11540 7251 11543
rect 7650 11540 7656 11552
rect 7239 11512 7656 11540
rect 7239 11509 7251 11512
rect 7193 11503 7251 11509
rect 7650 11500 7656 11512
rect 7708 11500 7714 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 8389 11543 8447 11549
rect 8389 11540 8401 11543
rect 8352 11512 8401 11540
rect 8352 11500 8358 11512
rect 8389 11509 8401 11512
rect 8435 11509 8447 11543
rect 8389 11503 8447 11509
rect 11238 11500 11244 11552
rect 11296 11540 11302 11552
rect 11333 11543 11391 11549
rect 11333 11540 11345 11543
rect 11296 11512 11345 11540
rect 11296 11500 11302 11512
rect 11333 11509 11345 11512
rect 11379 11540 11391 11543
rect 12894 11540 12900 11552
rect 11379 11512 12900 11540
rect 11379 11509 11391 11512
rect 11333 11503 11391 11509
rect 12894 11500 12900 11512
rect 12952 11500 12958 11552
rect 13814 11500 13820 11552
rect 13872 11540 13878 11552
rect 14553 11543 14611 11549
rect 14553 11540 14565 11543
rect 13872 11512 14565 11540
rect 13872 11500 13878 11512
rect 14553 11509 14565 11512
rect 14599 11509 14611 11543
rect 17494 11540 17500 11552
rect 17455 11512 17500 11540
rect 14553 11503 14611 11509
rect 17494 11500 17500 11512
rect 17552 11500 17558 11552
rect 17770 11500 17776 11552
rect 17828 11540 17834 11552
rect 18248 11549 18276 11580
rect 19061 11577 19073 11580
rect 19107 11608 19119 11611
rect 19260 11608 19288 11639
rect 21910 11636 21916 11648
rect 21968 11636 21974 11688
rect 23934 11685 23940 11688
rect 23928 11676 23940 11685
rect 23768 11648 23940 11676
rect 19107 11580 19288 11608
rect 19107 11577 19119 11580
rect 19061 11571 19119 11577
rect 19426 11568 19432 11620
rect 19484 11617 19490 11620
rect 19484 11611 19548 11617
rect 19484 11577 19502 11611
rect 19536 11577 19548 11611
rect 19484 11571 19548 11577
rect 21637 11611 21695 11617
rect 21637 11577 21649 11611
rect 21683 11608 21695 11611
rect 22465 11611 22523 11617
rect 22465 11608 22477 11611
rect 21683 11580 22477 11608
rect 21683 11577 21695 11580
rect 21637 11571 21695 11577
rect 22465 11577 22477 11580
rect 22511 11608 22523 11611
rect 23768 11608 23796 11648
rect 23928 11639 23940 11648
rect 23934 11636 23940 11639
rect 23992 11636 23998 11688
rect 28905 11679 28963 11685
rect 28905 11645 28917 11679
rect 28951 11676 28963 11679
rect 29273 11679 29331 11685
rect 29273 11676 29285 11679
rect 28951 11648 29285 11676
rect 28951 11645 28963 11648
rect 28905 11639 28963 11645
rect 29273 11645 29285 11648
rect 29319 11645 29331 11679
rect 34885 11679 34943 11685
rect 34885 11676 34897 11679
rect 29273 11639 29331 11645
rect 34624 11648 34897 11676
rect 22511 11580 23796 11608
rect 22511 11577 22523 11580
rect 22465 11571 22523 11577
rect 19484 11568 19490 11571
rect 26786 11568 26792 11620
rect 26844 11608 26850 11620
rect 26942 11611 27000 11617
rect 26942 11608 26954 11611
rect 26844 11580 26954 11608
rect 26844 11568 26850 11580
rect 26942 11577 26954 11580
rect 26988 11608 27000 11611
rect 27522 11608 27528 11620
rect 26988 11580 27528 11608
rect 26988 11577 27000 11580
rect 26942 11571 27000 11577
rect 27522 11568 27528 11580
rect 27580 11568 27586 11620
rect 29546 11617 29552 11620
rect 28721 11611 28779 11617
rect 28721 11577 28733 11611
rect 28767 11608 28779 11611
rect 29540 11608 29552 11617
rect 28767 11580 29552 11608
rect 28767 11577 28779 11580
rect 28721 11571 28779 11577
rect 29540 11571 29552 11580
rect 29546 11568 29552 11571
rect 29604 11568 29610 11620
rect 32217 11611 32275 11617
rect 32217 11577 32229 11611
rect 32263 11608 32275 11611
rect 32398 11608 32404 11620
rect 32263 11580 32404 11608
rect 32263 11577 32275 11580
rect 32217 11571 32275 11577
rect 32398 11568 32404 11580
rect 32456 11608 32462 11620
rect 32769 11611 32827 11617
rect 32769 11608 32781 11611
rect 32456 11580 32781 11608
rect 32456 11568 32462 11580
rect 32769 11577 32781 11580
rect 32815 11577 32827 11611
rect 32769 11571 32827 11577
rect 34624 11552 34652 11648
rect 34885 11645 34897 11648
rect 34931 11645 34943 11679
rect 34885 11639 34943 11645
rect 34992 11608 35020 11716
rect 35152 11611 35210 11617
rect 35152 11608 35164 11611
rect 34992 11580 35164 11608
rect 35152 11577 35164 11580
rect 35198 11608 35210 11611
rect 35986 11608 35992 11620
rect 35198 11580 35992 11608
rect 35198 11577 35210 11580
rect 35152 11571 35210 11577
rect 35986 11568 35992 11580
rect 36044 11568 36050 11620
rect 18233 11543 18291 11549
rect 18233 11540 18245 11543
rect 17828 11512 18245 11540
rect 17828 11500 17834 11512
rect 18233 11509 18245 11512
rect 18279 11509 18291 11543
rect 18690 11540 18696 11552
rect 18651 11512 18696 11540
rect 18233 11503 18291 11509
rect 18690 11500 18696 11512
rect 18748 11500 18754 11552
rect 22002 11540 22008 11552
rect 21963 11512 22008 11540
rect 22002 11500 22008 11512
rect 22060 11500 22066 11552
rect 22186 11500 22192 11552
rect 22244 11540 22250 11552
rect 22373 11543 22431 11549
rect 22373 11540 22385 11543
rect 22244 11512 22385 11540
rect 22244 11500 22250 11512
rect 22373 11509 22385 11512
rect 22419 11540 22431 11543
rect 22738 11540 22744 11552
rect 22419 11512 22744 11540
rect 22419 11509 22431 11512
rect 22373 11503 22431 11509
rect 22738 11500 22744 11512
rect 22796 11500 22802 11552
rect 25038 11540 25044 11552
rect 24999 11512 25044 11540
rect 25038 11500 25044 11512
rect 25096 11500 25102 11552
rect 28166 11500 28172 11552
rect 28224 11540 28230 11552
rect 28905 11543 28963 11549
rect 28905 11540 28917 11543
rect 28224 11512 28917 11540
rect 28224 11500 28230 11512
rect 28905 11509 28917 11512
rect 28951 11540 28963 11543
rect 28997 11543 29055 11549
rect 28997 11540 29009 11543
rect 28951 11512 29009 11540
rect 28951 11509 28963 11512
rect 28905 11503 28963 11509
rect 28997 11509 29009 11512
rect 29043 11509 29055 11543
rect 28997 11503 29055 11509
rect 30374 11500 30380 11552
rect 30432 11540 30438 11552
rect 30653 11543 30711 11549
rect 30653 11540 30665 11543
rect 30432 11512 30665 11540
rect 30432 11500 30438 11512
rect 30653 11509 30665 11512
rect 30699 11509 30711 11543
rect 30653 11503 30711 11509
rect 31849 11543 31907 11549
rect 31849 11509 31861 11543
rect 31895 11540 31907 11543
rect 32677 11543 32735 11549
rect 32677 11540 32689 11543
rect 31895 11512 32689 11540
rect 31895 11509 31907 11512
rect 31849 11503 31907 11509
rect 32677 11509 32689 11512
rect 32723 11540 32735 11543
rect 33502 11540 33508 11552
rect 32723 11512 33508 11540
rect 32723 11509 32735 11512
rect 32677 11503 32735 11509
rect 33502 11500 33508 11512
rect 33560 11500 33566 11552
rect 34606 11540 34612 11552
rect 34567 11512 34612 11540
rect 34606 11500 34612 11512
rect 34664 11500 34670 11552
rect 1104 11450 38824 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 38824 11450
rect 1104 11376 38824 11398
rect 4706 11336 4712 11348
rect 4667 11308 4712 11336
rect 4706 11296 4712 11308
rect 4764 11296 4770 11348
rect 5166 11336 5172 11348
rect 5127 11308 5172 11336
rect 5166 11296 5172 11308
rect 5224 11296 5230 11348
rect 5442 11296 5448 11348
rect 5500 11336 5506 11348
rect 5721 11339 5779 11345
rect 5721 11336 5733 11339
rect 5500 11308 5733 11336
rect 5500 11296 5506 11308
rect 5721 11305 5733 11308
rect 5767 11305 5779 11339
rect 5721 11299 5779 11305
rect 6181 11339 6239 11345
rect 6181 11305 6193 11339
rect 6227 11336 6239 11339
rect 6270 11336 6276 11348
rect 6227 11308 6276 11336
rect 6227 11305 6239 11308
rect 6181 11299 6239 11305
rect 6270 11296 6276 11308
rect 6328 11336 6334 11348
rect 8386 11336 8392 11348
rect 6328 11308 8392 11336
rect 6328 11296 6334 11308
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 9490 11336 9496 11348
rect 9451 11308 9496 11336
rect 9490 11296 9496 11308
rect 9548 11296 9554 11348
rect 11057 11339 11115 11345
rect 11057 11305 11069 11339
rect 11103 11305 11115 11339
rect 11057 11299 11115 11305
rect 14093 11339 14151 11345
rect 14093 11305 14105 11339
rect 14139 11336 14151 11339
rect 15010 11336 15016 11348
rect 14139 11308 15016 11336
rect 14139 11305 14151 11308
rect 14093 11299 14151 11305
rect 6540 11271 6598 11277
rect 6540 11237 6552 11271
rect 6586 11268 6598 11271
rect 6638 11268 6644 11280
rect 6586 11240 6644 11268
rect 6586 11237 6598 11240
rect 6540 11231 6598 11237
rect 6638 11228 6644 11240
rect 6696 11228 6702 11280
rect 8297 11271 8355 11277
rect 8297 11237 8309 11271
rect 8343 11268 8355 11271
rect 8478 11268 8484 11280
rect 8343 11240 8484 11268
rect 8343 11237 8355 11240
rect 8297 11231 8355 11237
rect 8478 11228 8484 11240
rect 8536 11268 8542 11280
rect 11072 11268 11100 11299
rect 15010 11296 15016 11308
rect 15068 11296 15074 11348
rect 18690 11296 18696 11348
rect 18748 11336 18754 11348
rect 19245 11339 19303 11345
rect 19245 11336 19257 11339
rect 18748 11308 19257 11336
rect 18748 11296 18754 11308
rect 19245 11305 19257 11308
rect 19291 11305 19303 11339
rect 19245 11299 19303 11305
rect 19426 11296 19432 11348
rect 19484 11336 19490 11348
rect 19797 11339 19855 11345
rect 19797 11336 19809 11339
rect 19484 11308 19809 11336
rect 19484 11296 19490 11308
rect 19797 11305 19809 11308
rect 19843 11305 19855 11339
rect 19797 11299 19855 11305
rect 21082 11296 21088 11348
rect 21140 11336 21146 11348
rect 21729 11339 21787 11345
rect 21729 11336 21741 11339
rect 21140 11308 21741 11336
rect 21140 11296 21146 11308
rect 21729 11305 21741 11308
rect 21775 11305 21787 11339
rect 22646 11336 22652 11348
rect 22607 11308 22652 11336
rect 21729 11299 21787 11305
rect 22646 11296 22652 11308
rect 22704 11296 22710 11348
rect 23385 11339 23443 11345
rect 23385 11305 23397 11339
rect 23431 11336 23443 11339
rect 23934 11336 23940 11348
rect 23431 11308 23940 11336
rect 23431 11305 23443 11308
rect 23385 11299 23443 11305
rect 23934 11296 23940 11308
rect 23992 11296 23998 11348
rect 26786 11336 26792 11348
rect 26747 11308 26792 11336
rect 26786 11296 26792 11308
rect 26844 11296 26850 11348
rect 27614 11336 27620 11348
rect 27575 11308 27620 11336
rect 27614 11296 27620 11308
rect 27672 11296 27678 11348
rect 28074 11336 28080 11348
rect 28035 11308 28080 11336
rect 28074 11296 28080 11308
rect 28132 11296 28138 11348
rect 29546 11336 29552 11348
rect 29459 11308 29552 11336
rect 29546 11296 29552 11308
rect 29604 11336 29610 11348
rect 30466 11336 30472 11348
rect 29604 11308 30472 11336
rect 29604 11296 29610 11308
rect 30466 11296 30472 11308
rect 30524 11296 30530 11348
rect 30834 11336 30840 11348
rect 30795 11308 30840 11336
rect 30834 11296 30840 11308
rect 30892 11296 30898 11348
rect 33502 11336 33508 11348
rect 33463 11308 33508 11336
rect 33502 11296 33508 11308
rect 33560 11296 33566 11348
rect 35986 11336 35992 11348
rect 35947 11308 35992 11336
rect 35986 11296 35992 11308
rect 36044 11296 36050 11348
rect 8536 11240 11100 11268
rect 8536 11228 8542 11240
rect 20990 11228 20996 11280
rect 21048 11268 21054 11280
rect 21637 11271 21695 11277
rect 21637 11268 21649 11271
rect 21048 11240 21649 11268
rect 21048 11228 21054 11240
rect 21637 11237 21649 11240
rect 21683 11268 21695 11271
rect 22002 11268 22008 11280
rect 21683 11240 22008 11268
rect 21683 11237 21695 11240
rect 21637 11231 21695 11237
rect 22002 11228 22008 11240
rect 22060 11228 22066 11280
rect 4617 11203 4675 11209
rect 4617 11169 4629 11203
rect 4663 11200 4675 11203
rect 5077 11203 5135 11209
rect 5077 11200 5089 11203
rect 4663 11172 5089 11200
rect 4663 11169 4675 11172
rect 4617 11163 4675 11169
rect 5077 11169 5089 11172
rect 5123 11200 5135 11203
rect 5442 11200 5448 11212
rect 5123 11172 5448 11200
rect 5123 11169 5135 11172
rect 5077 11163 5135 11169
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 9944 11203 10002 11209
rect 9944 11200 9956 11203
rect 8220 11172 9956 11200
rect 5261 11135 5319 11141
rect 5261 11101 5273 11135
rect 5307 11132 5319 11135
rect 5350 11132 5356 11144
rect 5307 11104 5356 11132
rect 5307 11101 5319 11104
rect 5261 11095 5319 11101
rect 5276 11064 5304 11095
rect 5350 11092 5356 11104
rect 5408 11092 5414 11144
rect 6270 11132 6276 11144
rect 6231 11104 6276 11132
rect 6270 11092 6276 11104
rect 6328 11092 6334 11144
rect 7650 11064 7656 11076
rect 4080 11036 5304 11064
rect 7563 11036 7656 11064
rect 3786 10956 3792 11008
rect 3844 10996 3850 11008
rect 4080 10996 4108 11036
rect 7650 11024 7656 11036
rect 7708 11064 7714 11076
rect 8220 11064 8248 11172
rect 9944 11169 9956 11172
rect 9990 11200 10002 11203
rect 10502 11200 10508 11212
rect 9990 11172 10508 11200
rect 9990 11169 10002 11172
rect 9944 11163 10002 11169
rect 10502 11160 10508 11172
rect 10560 11160 10566 11212
rect 12434 11160 12440 11212
rect 12492 11200 12498 11212
rect 12969 11203 13027 11209
rect 12969 11200 12981 11203
rect 12492 11172 12981 11200
rect 12492 11160 12498 11172
rect 12969 11169 12981 11172
rect 13015 11169 13027 11203
rect 12969 11163 13027 11169
rect 17770 11160 17776 11212
rect 17828 11200 17834 11212
rect 17865 11203 17923 11209
rect 17865 11200 17877 11203
rect 17828 11172 17877 11200
rect 17828 11160 17834 11172
rect 17865 11169 17877 11172
rect 17911 11169 17923 11203
rect 17865 11163 17923 11169
rect 17954 11160 17960 11212
rect 18012 11200 18018 11212
rect 18132 11203 18190 11209
rect 18132 11200 18144 11203
rect 18012 11172 18144 11200
rect 18012 11160 18018 11172
rect 18132 11169 18144 11172
rect 18178 11200 18190 11203
rect 19150 11200 19156 11212
rect 18178 11172 19156 11200
rect 18178 11169 18190 11172
rect 18132 11163 18190 11169
rect 19150 11160 19156 11172
rect 19208 11160 19214 11212
rect 21177 11203 21235 11209
rect 21177 11169 21189 11203
rect 21223 11200 21235 11203
rect 22664 11200 22692 11296
rect 22738 11228 22744 11280
rect 22796 11268 22802 11280
rect 23198 11268 23204 11280
rect 22796 11240 23204 11268
rect 22796 11228 22802 11240
rect 23198 11228 23204 11240
rect 23256 11268 23262 11280
rect 23744 11271 23802 11277
rect 23744 11268 23756 11271
rect 23256 11240 23756 11268
rect 23256 11228 23262 11240
rect 23744 11237 23756 11240
rect 23790 11268 23802 11271
rect 25038 11268 25044 11280
rect 23790 11240 25044 11268
rect 23790 11237 23802 11240
rect 23744 11231 23802 11237
rect 25038 11228 25044 11240
rect 25096 11228 25102 11280
rect 21223 11172 22692 11200
rect 27632 11200 27660 11296
rect 28436 11271 28494 11277
rect 28436 11237 28448 11271
rect 28482 11268 28494 11271
rect 28626 11268 28632 11280
rect 28482 11240 28632 11268
rect 28482 11237 28494 11240
rect 28436 11231 28494 11237
rect 28626 11228 28632 11240
rect 28684 11268 28690 11280
rect 30190 11268 30196 11280
rect 28684 11240 30196 11268
rect 28684 11228 28690 11240
rect 30190 11228 30196 11240
rect 30248 11228 30254 11280
rect 32398 11277 32404 11280
rect 32392 11268 32404 11277
rect 32359 11240 32404 11268
rect 32392 11231 32404 11240
rect 32398 11228 32404 11231
rect 32456 11228 32462 11280
rect 33962 11228 33968 11280
rect 34020 11268 34026 11280
rect 34790 11268 34796 11280
rect 34020 11240 34796 11268
rect 34020 11228 34026 11240
rect 34790 11228 34796 11240
rect 34848 11277 34854 11280
rect 34848 11271 34912 11277
rect 34848 11237 34866 11271
rect 34900 11237 34912 11271
rect 34848 11231 34912 11237
rect 34848 11228 34854 11231
rect 28166 11200 28172 11212
rect 27632 11172 28172 11200
rect 21223 11169 21235 11172
rect 21177 11163 21235 11169
rect 28166 11160 28172 11172
rect 28224 11160 28230 11212
rect 9030 11092 9036 11144
rect 9088 11132 9094 11144
rect 9677 11135 9735 11141
rect 9677 11132 9689 11135
rect 9088 11104 9689 11132
rect 9088 11092 9094 11104
rect 9677 11101 9689 11104
rect 9723 11101 9735 11135
rect 12710 11132 12716 11144
rect 12671 11104 12716 11132
rect 9677 11095 9735 11101
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 20714 11092 20720 11144
rect 20772 11132 20778 11144
rect 21821 11135 21879 11141
rect 21821 11132 21833 11135
rect 20772 11104 21833 11132
rect 20772 11092 20778 11104
rect 21821 11101 21833 11104
rect 21867 11101 21879 11135
rect 23474 11132 23480 11144
rect 23435 11104 23480 11132
rect 21821 11095 21879 11101
rect 23474 11092 23480 11104
rect 23532 11092 23538 11144
rect 32122 11132 32128 11144
rect 32083 11104 32128 11132
rect 32122 11092 32128 11104
rect 32180 11092 32186 11144
rect 34606 11132 34612 11144
rect 34567 11104 34612 11132
rect 34606 11092 34612 11104
rect 34664 11092 34670 11144
rect 8662 11064 8668 11076
rect 7708 11036 8248 11064
rect 8575 11036 8668 11064
rect 7708 11024 7714 11036
rect 8662 11024 8668 11036
rect 8720 11064 8726 11076
rect 9582 11064 9588 11076
rect 8720 11036 9588 11064
rect 8720 11024 8726 11036
rect 9582 11024 9588 11036
rect 9640 11024 9646 11076
rect 20625 11067 20683 11073
rect 20625 11033 20637 11067
rect 20671 11064 20683 11067
rect 20806 11064 20812 11076
rect 20671 11036 20812 11064
rect 20671 11033 20683 11036
rect 20625 11027 20683 11033
rect 20806 11024 20812 11036
rect 20864 11064 20870 11076
rect 22554 11064 22560 11076
rect 20864 11036 22560 11064
rect 20864 11024 20870 11036
rect 22554 11024 22560 11036
rect 22612 11024 22618 11076
rect 24854 11064 24860 11076
rect 24815 11036 24860 11064
rect 24854 11024 24860 11036
rect 24912 11024 24918 11076
rect 34149 11067 34207 11073
rect 34149 11033 34161 11067
rect 34195 11064 34207 11067
rect 34330 11064 34336 11076
rect 34195 11036 34336 11064
rect 34195 11033 34207 11036
rect 34149 11027 34207 11033
rect 34330 11024 34336 11036
rect 34388 11024 34394 11076
rect 3844 10968 4108 10996
rect 3844 10956 3850 10968
rect 8294 10956 8300 11008
rect 8352 10996 8358 11008
rect 9033 10999 9091 11005
rect 9033 10996 9045 10999
rect 8352 10968 9045 10996
rect 8352 10956 8358 10968
rect 9033 10965 9045 10968
rect 9079 10996 9091 10999
rect 9306 10996 9312 11008
rect 9079 10968 9312 10996
rect 9079 10965 9091 10968
rect 9033 10959 9091 10965
rect 9306 10956 9312 10968
rect 9364 10996 9370 11008
rect 9490 10996 9496 11008
rect 9364 10968 9496 10996
rect 9364 10956 9370 10968
rect 9490 10956 9496 10968
rect 9548 10956 9554 11008
rect 21266 10996 21272 11008
rect 21227 10968 21272 10996
rect 21266 10956 21272 10968
rect 21324 10956 21330 11008
rect 23014 10996 23020 11008
rect 22975 10968 23020 10996
rect 23014 10956 23020 10968
rect 23072 10956 23078 11008
rect 1104 10906 38824 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 38824 10906
rect 1104 10832 38824 10854
rect 3786 10792 3792 10804
rect 3747 10764 3792 10792
rect 3786 10752 3792 10764
rect 3844 10752 3850 10804
rect 3878 10752 3884 10804
rect 3936 10792 3942 10804
rect 4065 10795 4123 10801
rect 4065 10792 4077 10795
rect 3936 10764 4077 10792
rect 3936 10752 3942 10764
rect 4065 10761 4077 10764
rect 4111 10761 4123 10795
rect 4065 10755 4123 10761
rect 4080 10656 4108 10755
rect 5442 10752 5448 10804
rect 5500 10792 5506 10804
rect 5629 10795 5687 10801
rect 5629 10792 5641 10795
rect 5500 10764 5641 10792
rect 5500 10752 5506 10764
rect 5629 10761 5641 10764
rect 5675 10761 5687 10795
rect 5629 10755 5687 10761
rect 7285 10795 7343 10801
rect 7285 10761 7297 10795
rect 7331 10792 7343 10795
rect 8202 10792 8208 10804
rect 7331 10764 8208 10792
rect 7331 10761 7343 10764
rect 7285 10755 7343 10761
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 9490 10752 9496 10804
rect 9548 10792 9554 10804
rect 9585 10795 9643 10801
rect 9585 10792 9597 10795
rect 9548 10764 9597 10792
rect 9548 10752 9554 10764
rect 9585 10761 9597 10764
rect 9631 10761 9643 10795
rect 9585 10755 9643 10761
rect 9766 10752 9772 10804
rect 9824 10792 9830 10804
rect 10137 10795 10195 10801
rect 10137 10792 10149 10795
rect 9824 10764 10149 10792
rect 9824 10752 9830 10764
rect 10137 10761 10149 10764
rect 10183 10761 10195 10795
rect 10502 10792 10508 10804
rect 10463 10764 10508 10792
rect 10137 10755 10195 10761
rect 6270 10684 6276 10736
rect 6328 10724 6334 10736
rect 6365 10727 6423 10733
rect 6365 10724 6377 10727
rect 6328 10696 6377 10724
rect 6328 10684 6334 10696
rect 6365 10693 6377 10696
rect 6411 10724 6423 10727
rect 7006 10724 7012 10736
rect 6411 10696 7012 10724
rect 6411 10693 6423 10696
rect 6365 10687 6423 10693
rect 7006 10684 7012 10696
rect 7064 10724 7070 10736
rect 8110 10724 8116 10736
rect 7064 10696 8116 10724
rect 7064 10684 7070 10696
rect 8110 10684 8116 10696
rect 8168 10724 8174 10736
rect 8168 10696 8248 10724
rect 8168 10684 8174 10696
rect 4246 10656 4252 10668
rect 4080 10628 4252 10656
rect 4246 10616 4252 10628
rect 4304 10616 4310 10668
rect 8220 10665 8248 10696
rect 8205 10659 8263 10665
rect 8205 10625 8217 10659
rect 8251 10625 8263 10659
rect 10152 10656 10180 10755
rect 10502 10752 10508 10764
rect 10560 10752 10566 10804
rect 17129 10795 17187 10801
rect 17129 10761 17141 10795
rect 17175 10792 17187 10795
rect 17862 10792 17868 10804
rect 17175 10764 17868 10792
rect 17175 10761 17187 10764
rect 17129 10755 17187 10761
rect 17862 10752 17868 10764
rect 17920 10752 17926 10804
rect 19150 10752 19156 10804
rect 19208 10792 19214 10804
rect 19429 10795 19487 10801
rect 19429 10792 19441 10795
rect 19208 10764 19441 10792
rect 19208 10752 19214 10764
rect 19429 10761 19441 10764
rect 19475 10761 19487 10795
rect 20990 10792 20996 10804
rect 20951 10764 20996 10792
rect 19429 10755 19487 10761
rect 20990 10752 20996 10764
rect 21048 10752 21054 10804
rect 21082 10752 21088 10804
rect 21140 10792 21146 10804
rect 21269 10795 21327 10801
rect 21269 10792 21281 10795
rect 21140 10764 21281 10792
rect 21140 10752 21146 10764
rect 21269 10761 21281 10764
rect 21315 10761 21327 10795
rect 21269 10755 21327 10761
rect 22462 10752 22468 10804
rect 22520 10792 22526 10804
rect 23017 10795 23075 10801
rect 23017 10792 23029 10795
rect 22520 10764 23029 10792
rect 22520 10752 22526 10764
rect 23017 10761 23029 10764
rect 23063 10792 23075 10795
rect 23385 10795 23443 10801
rect 23385 10792 23397 10795
rect 23063 10764 23397 10792
rect 23063 10761 23075 10764
rect 23017 10755 23075 10761
rect 23385 10761 23397 10764
rect 23431 10792 23443 10795
rect 23474 10792 23480 10804
rect 23431 10764 23480 10792
rect 23431 10761 23443 10764
rect 23385 10755 23443 10761
rect 23474 10752 23480 10764
rect 23532 10752 23538 10804
rect 28166 10792 28172 10804
rect 28127 10764 28172 10792
rect 28166 10752 28172 10764
rect 28224 10752 28230 10804
rect 28626 10792 28632 10804
rect 28587 10764 28632 10792
rect 28626 10752 28632 10764
rect 28684 10752 28690 10804
rect 31573 10795 31631 10801
rect 31573 10792 31585 10795
rect 29656 10764 31585 10792
rect 11333 10727 11391 10733
rect 11333 10693 11345 10727
rect 11379 10724 11391 10727
rect 13173 10727 13231 10733
rect 13173 10724 13185 10727
rect 11379 10696 13185 10724
rect 11379 10693 11391 10696
rect 11333 10687 11391 10693
rect 13173 10693 13185 10696
rect 13219 10693 13231 10727
rect 28184 10724 28212 10752
rect 29457 10727 29515 10733
rect 29457 10724 29469 10727
rect 28184 10696 29469 10724
rect 13173 10687 13231 10693
rect 29457 10693 29469 10696
rect 29503 10724 29515 10727
rect 29656 10724 29684 10764
rect 31573 10761 31585 10764
rect 31619 10792 31631 10795
rect 32122 10792 32128 10804
rect 31619 10764 32128 10792
rect 31619 10761 31631 10764
rect 31573 10755 31631 10761
rect 32122 10752 32128 10764
rect 32180 10752 32186 10804
rect 32398 10752 32404 10804
rect 32456 10792 32462 10804
rect 33505 10795 33563 10801
rect 33505 10792 33517 10795
rect 32456 10764 33517 10792
rect 32456 10752 32462 10764
rect 33505 10761 33517 10764
rect 33551 10761 33563 10795
rect 34606 10792 34612 10804
rect 34567 10764 34612 10792
rect 33505 10755 33563 10761
rect 34606 10752 34612 10764
rect 34664 10752 34670 10804
rect 34790 10752 34796 10804
rect 34848 10792 34854 10804
rect 35069 10795 35127 10801
rect 35069 10792 35081 10795
rect 34848 10764 35081 10792
rect 34848 10752 34854 10764
rect 35069 10761 35081 10764
rect 35115 10761 35127 10795
rect 35069 10755 35127 10761
rect 29503 10696 29684 10724
rect 29503 10693 29515 10696
rect 29457 10687 29515 10693
rect 10594 10656 10600 10668
rect 10152 10628 10600 10656
rect 8205 10619 8263 10625
rect 10594 10616 10600 10628
rect 10652 10656 10658 10668
rect 12710 10656 12716 10668
rect 10652 10628 12716 10656
rect 10652 10616 10658 10628
rect 12710 10616 12716 10628
rect 12768 10616 12774 10668
rect 13188 10656 13216 10687
rect 13446 10656 13452 10668
rect 13188 10628 13452 10656
rect 13446 10616 13452 10628
rect 13504 10656 13510 10668
rect 14185 10659 14243 10665
rect 14185 10656 14197 10659
rect 13504 10628 14197 10656
rect 13504 10616 13510 10628
rect 14185 10625 14197 10628
rect 14231 10625 14243 10659
rect 14642 10656 14648 10668
rect 14185 10619 14243 10625
rect 14384 10628 14648 10656
rect 7101 10591 7159 10597
rect 7101 10557 7113 10591
rect 7147 10588 7159 10591
rect 7282 10588 7288 10600
rect 7147 10560 7288 10588
rect 7147 10557 7159 10560
rect 7101 10551 7159 10557
rect 7282 10548 7288 10560
rect 7340 10588 7346 10600
rect 8478 10597 8484 10600
rect 7653 10591 7711 10597
rect 7653 10588 7665 10591
rect 7340 10560 7665 10588
rect 7340 10548 7346 10560
rect 7653 10557 7665 10560
rect 7699 10557 7711 10591
rect 8472 10588 8484 10597
rect 8439 10560 8484 10588
rect 7653 10551 7711 10557
rect 8472 10551 8484 10560
rect 8478 10548 8484 10551
rect 8536 10548 8542 10600
rect 11146 10588 11152 10600
rect 11107 10560 11152 10588
rect 11146 10548 11152 10560
rect 11204 10588 11210 10600
rect 11701 10591 11759 10597
rect 11701 10588 11713 10591
rect 11204 10560 11713 10588
rect 11204 10548 11210 10560
rect 11701 10557 11713 10560
rect 11747 10557 11759 10591
rect 11701 10551 11759 10557
rect 13725 10591 13783 10597
rect 13725 10557 13737 10591
rect 13771 10588 13783 10591
rect 14384 10588 14412 10628
rect 14642 10616 14648 10628
rect 14700 10616 14706 10668
rect 22554 10656 22560 10668
rect 22515 10628 22560 10656
rect 22554 10616 22560 10628
rect 22612 10616 22618 10668
rect 23014 10616 23020 10668
rect 23072 10656 23078 10668
rect 29656 10665 29684 10696
rect 29641 10659 29699 10665
rect 23072 10628 23796 10656
rect 23072 10616 23078 10628
rect 13771 10560 14412 10588
rect 13771 10557 13783 10560
rect 13725 10551 13783 10557
rect 14458 10548 14464 10600
rect 14516 10588 14522 10600
rect 17770 10588 17776 10600
rect 14516 10560 14561 10588
rect 17420 10560 17776 10588
rect 14516 10548 14522 10560
rect 4516 10523 4574 10529
rect 4516 10489 4528 10523
rect 4562 10520 4574 10523
rect 4798 10520 4804 10532
rect 4562 10492 4804 10520
rect 4562 10489 4574 10492
rect 4516 10483 4574 10489
rect 4798 10480 4804 10492
rect 4856 10520 4862 10532
rect 5166 10520 5172 10532
rect 4856 10492 5172 10520
rect 4856 10480 4862 10492
rect 5166 10480 5172 10492
rect 5224 10480 5230 10532
rect 16850 10480 16856 10532
rect 16908 10520 16914 10532
rect 17420 10529 17448 10560
rect 17770 10548 17776 10560
rect 17828 10588 17834 10600
rect 18049 10591 18107 10597
rect 18049 10588 18061 10591
rect 17828 10560 18061 10588
rect 17828 10548 17834 10560
rect 18049 10557 18061 10560
rect 18095 10557 18107 10591
rect 18049 10551 18107 10557
rect 21913 10591 21971 10597
rect 21913 10557 21925 10591
rect 21959 10588 21971 10591
rect 22465 10591 22523 10597
rect 22465 10588 22477 10591
rect 21959 10560 22477 10588
rect 21959 10557 21971 10560
rect 21913 10551 21971 10557
rect 22465 10557 22477 10560
rect 22511 10588 22523 10591
rect 23032 10588 23060 10616
rect 22511 10560 23060 10588
rect 22511 10557 22523 10560
rect 22465 10551 22523 10557
rect 23474 10548 23480 10600
rect 23532 10588 23538 10600
rect 23661 10591 23719 10597
rect 23661 10588 23673 10591
rect 23532 10560 23673 10588
rect 23532 10548 23538 10560
rect 23661 10557 23673 10560
rect 23707 10557 23719 10591
rect 23768 10588 23796 10628
rect 29641 10625 29653 10659
rect 29687 10625 29699 10659
rect 29641 10619 29699 10625
rect 23928 10591 23986 10597
rect 23928 10588 23940 10591
rect 23768 10560 23940 10588
rect 23661 10551 23719 10557
rect 23928 10557 23940 10560
rect 23974 10588 23986 10591
rect 24762 10588 24768 10600
rect 23974 10560 24768 10588
rect 23974 10557 23986 10560
rect 23928 10551 23986 10557
rect 24762 10548 24768 10560
rect 24820 10548 24826 10600
rect 29908 10591 29966 10597
rect 29908 10588 29920 10591
rect 29840 10560 29920 10588
rect 17405 10523 17463 10529
rect 17405 10520 17417 10523
rect 16908 10492 17417 10520
rect 16908 10480 16914 10492
rect 17405 10489 17417 10492
rect 17451 10489 17463 10523
rect 17405 10483 17463 10489
rect 18230 10480 18236 10532
rect 18288 10529 18294 10532
rect 18288 10523 18352 10529
rect 18288 10489 18306 10523
rect 18340 10489 18352 10523
rect 18288 10483 18352 10489
rect 29089 10523 29147 10529
rect 29089 10489 29101 10523
rect 29135 10520 29147 10523
rect 29840 10520 29868 10560
rect 29908 10557 29920 10560
rect 29954 10588 29966 10591
rect 30282 10588 30288 10600
rect 29954 10560 30288 10588
rect 29954 10557 29966 10560
rect 29908 10551 29966 10557
rect 30282 10548 30288 10560
rect 30340 10548 30346 10600
rect 32140 10597 32168 10752
rect 34514 10684 34520 10736
rect 34572 10724 34578 10736
rect 35621 10727 35679 10733
rect 35621 10724 35633 10727
rect 34572 10696 35633 10724
rect 34572 10684 34578 10696
rect 35621 10693 35633 10696
rect 35667 10693 35679 10727
rect 35621 10687 35679 10693
rect 32125 10591 32183 10597
rect 32125 10557 32137 10591
rect 32171 10588 32183 10591
rect 35437 10591 35495 10597
rect 32171 10560 32260 10588
rect 32171 10557 32183 10560
rect 32125 10551 32183 10557
rect 29135 10492 29868 10520
rect 29135 10489 29147 10492
rect 29089 10483 29147 10489
rect 18288 10480 18294 10483
rect 12250 10452 12256 10464
rect 12211 10424 12256 10452
rect 12250 10412 12256 10424
rect 12308 10412 12314 10464
rect 13633 10455 13691 10461
rect 13633 10421 13645 10455
rect 13679 10452 13691 10455
rect 13814 10452 13820 10464
rect 13679 10424 13820 10452
rect 13679 10421 13691 10424
rect 13633 10415 13691 10421
rect 13814 10412 13820 10424
rect 13872 10452 13878 10464
rect 14187 10455 14245 10461
rect 14187 10452 14199 10455
rect 13872 10424 14199 10452
rect 13872 10412 13878 10424
rect 14187 10421 14199 10424
rect 14233 10421 14245 10455
rect 15562 10452 15568 10464
rect 15523 10424 15568 10452
rect 14187 10415 14245 10421
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 20622 10452 20628 10464
rect 20583 10424 20628 10452
rect 20622 10412 20628 10424
rect 20680 10412 20686 10464
rect 21910 10412 21916 10464
rect 21968 10452 21974 10464
rect 22005 10455 22063 10461
rect 22005 10452 22017 10455
rect 21968 10424 22017 10452
rect 21968 10412 21974 10424
rect 22005 10421 22017 10424
rect 22051 10421 22063 10455
rect 22370 10452 22376 10464
rect 22331 10424 22376 10452
rect 22005 10415 22063 10421
rect 22370 10412 22376 10424
rect 22428 10412 22434 10464
rect 25038 10452 25044 10464
rect 24999 10424 25044 10452
rect 25038 10412 25044 10424
rect 25096 10412 25102 10464
rect 30006 10412 30012 10464
rect 30064 10452 30070 10464
rect 31018 10452 31024 10464
rect 30064 10424 31024 10452
rect 30064 10412 30070 10424
rect 31018 10412 31024 10424
rect 31076 10412 31082 10464
rect 32033 10455 32091 10461
rect 32033 10421 32045 10455
rect 32079 10452 32091 10455
rect 32232 10452 32260 10560
rect 35437 10557 35449 10591
rect 35483 10588 35495 10591
rect 35618 10588 35624 10600
rect 35483 10560 35624 10588
rect 35483 10557 35495 10560
rect 35437 10551 35495 10557
rect 35618 10548 35624 10560
rect 35676 10588 35682 10600
rect 35989 10591 36047 10597
rect 35989 10588 36001 10591
rect 35676 10560 36001 10588
rect 35676 10548 35682 10560
rect 35989 10557 36001 10560
rect 36035 10557 36047 10591
rect 35989 10551 36047 10557
rect 32398 10529 32404 10532
rect 32392 10483 32404 10529
rect 32456 10520 32462 10532
rect 32456 10492 32492 10520
rect 32398 10480 32404 10483
rect 32456 10480 32462 10492
rect 32950 10452 32956 10464
rect 32079 10424 32956 10452
rect 32079 10421 32091 10424
rect 32033 10415 32091 10421
rect 32950 10412 32956 10424
rect 33008 10412 33014 10464
rect 1104 10362 38824 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 38824 10362
rect 1104 10288 38824 10310
rect 4341 10251 4399 10257
rect 4341 10217 4353 10251
rect 4387 10248 4399 10251
rect 4798 10248 4804 10260
rect 4387 10220 4804 10248
rect 4387 10217 4399 10220
rect 4341 10211 4399 10217
rect 4798 10208 4804 10220
rect 4856 10208 4862 10260
rect 6457 10251 6515 10257
rect 6457 10217 6469 10251
rect 6503 10248 6515 10251
rect 6638 10248 6644 10260
rect 6503 10220 6644 10248
rect 6503 10217 6515 10220
rect 6457 10211 6515 10217
rect 6638 10208 6644 10220
rect 6696 10248 6702 10260
rect 7009 10251 7067 10257
rect 7009 10248 7021 10251
rect 6696 10220 7021 10248
rect 6696 10208 6702 10220
rect 7009 10217 7021 10220
rect 7055 10217 7067 10251
rect 7926 10248 7932 10260
rect 7887 10220 7932 10248
rect 7009 10211 7067 10217
rect 7926 10208 7932 10220
rect 7984 10208 7990 10260
rect 8389 10251 8447 10257
rect 8389 10217 8401 10251
rect 8435 10248 8447 10251
rect 8478 10248 8484 10260
rect 8435 10220 8484 10248
rect 8435 10217 8447 10220
rect 8389 10211 8447 10217
rect 8478 10208 8484 10220
rect 8536 10208 8542 10260
rect 9582 10208 9588 10260
rect 9640 10248 9646 10260
rect 9861 10251 9919 10257
rect 9861 10248 9873 10251
rect 9640 10220 9873 10248
rect 9640 10208 9646 10220
rect 9861 10217 9873 10220
rect 9907 10217 9919 10251
rect 10962 10248 10968 10260
rect 10923 10220 10968 10248
rect 9861 10211 9919 10217
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 23198 10248 23204 10260
rect 23159 10220 23204 10248
rect 23198 10208 23204 10220
rect 23256 10208 23262 10260
rect 29641 10251 29699 10257
rect 29641 10217 29653 10251
rect 29687 10217 29699 10251
rect 29641 10211 29699 10217
rect 30101 10251 30159 10257
rect 30101 10217 30113 10251
rect 30147 10248 30159 10251
rect 30282 10248 30288 10260
rect 30147 10220 30288 10248
rect 30147 10217 30159 10220
rect 30101 10211 30159 10217
rect 5344 10183 5402 10189
rect 5344 10149 5356 10183
rect 5390 10180 5402 10183
rect 5442 10180 5448 10192
rect 5390 10152 5448 10180
rect 5390 10149 5402 10152
rect 5344 10143 5402 10149
rect 5442 10140 5448 10152
rect 5500 10140 5506 10192
rect 12980 10183 13038 10189
rect 12980 10149 12992 10183
rect 13026 10180 13038 10183
rect 13722 10180 13728 10192
rect 13026 10152 13728 10180
rect 13026 10149 13038 10152
rect 12980 10143 13038 10149
rect 13722 10140 13728 10152
rect 13780 10140 13786 10192
rect 22097 10183 22155 10189
rect 22097 10149 22109 10183
rect 22143 10180 22155 10183
rect 22370 10180 22376 10192
rect 22143 10152 22376 10180
rect 22143 10149 22155 10152
rect 22097 10143 22155 10149
rect 22370 10140 22376 10152
rect 22428 10180 22434 10192
rect 23014 10180 23020 10192
rect 22428 10152 23020 10180
rect 22428 10140 22434 10152
rect 23014 10140 23020 10152
rect 23072 10180 23078 10192
rect 23560 10183 23618 10189
rect 23560 10180 23572 10183
rect 23072 10152 23572 10180
rect 23072 10140 23078 10152
rect 23560 10149 23572 10152
rect 23606 10180 23618 10183
rect 25038 10180 25044 10192
rect 23606 10152 25044 10180
rect 23606 10149 23618 10152
rect 23560 10143 23618 10149
rect 25038 10140 25044 10152
rect 25096 10140 25102 10192
rect 29656 10180 29684 10211
rect 30282 10208 30288 10220
rect 30340 10208 30346 10260
rect 31018 10208 31024 10260
rect 31076 10248 31082 10260
rect 32398 10248 32404 10260
rect 31076 10220 32404 10248
rect 31076 10208 31082 10220
rect 32398 10208 32404 10220
rect 32456 10208 32462 10260
rect 32490 10208 32496 10260
rect 32548 10248 32554 10260
rect 32677 10251 32735 10257
rect 32677 10248 32689 10251
rect 32548 10220 32689 10248
rect 32548 10208 32554 10220
rect 32677 10217 32689 10220
rect 32723 10217 32735 10251
rect 32677 10211 32735 10217
rect 34333 10251 34391 10257
rect 34333 10217 34345 10251
rect 34379 10248 34391 10251
rect 34790 10248 34796 10260
rect 34379 10220 34796 10248
rect 34379 10217 34391 10220
rect 34333 10211 34391 10217
rect 34790 10208 34796 10220
rect 34848 10208 34854 10260
rect 30190 10180 30196 10192
rect 29656 10152 30196 10180
rect 30190 10140 30196 10152
rect 30248 10140 30254 10192
rect 33220 10183 33278 10189
rect 33220 10149 33232 10183
rect 33266 10180 33278 10183
rect 33502 10180 33508 10192
rect 33266 10152 33508 10180
rect 33266 10149 33278 10152
rect 33220 10143 33278 10149
rect 33502 10140 33508 10152
rect 33560 10140 33566 10192
rect 4246 10072 4252 10124
rect 4304 10112 4310 10124
rect 5074 10112 5080 10124
rect 4304 10084 5080 10112
rect 4304 10072 4310 10084
rect 5074 10072 5080 10084
rect 5132 10072 5138 10124
rect 8294 10112 8300 10124
rect 8255 10084 8300 10112
rect 8294 10072 8300 10084
rect 8352 10072 8358 10124
rect 9674 10112 9680 10124
rect 9635 10084 9680 10112
rect 9674 10072 9680 10084
rect 9732 10072 9738 10124
rect 10781 10115 10839 10121
rect 10781 10081 10793 10115
rect 10827 10112 10839 10115
rect 10962 10112 10968 10124
rect 10827 10084 10968 10112
rect 10827 10081 10839 10084
rect 10781 10075 10839 10081
rect 10962 10072 10968 10084
rect 11020 10072 11026 10124
rect 12710 10112 12716 10124
rect 12671 10084 12716 10112
rect 12710 10072 12716 10084
rect 12768 10072 12774 10124
rect 16666 10072 16672 10124
rect 16724 10112 16730 10124
rect 17109 10115 17167 10121
rect 17109 10112 17121 10115
rect 16724 10084 17121 10112
rect 16724 10072 16730 10084
rect 17109 10081 17121 10084
rect 17155 10081 17167 10115
rect 19334 10112 19340 10124
rect 19295 10084 19340 10112
rect 17109 10075 17167 10081
rect 19334 10072 19340 10084
rect 19392 10072 19398 10124
rect 20901 10115 20959 10121
rect 20901 10081 20913 10115
rect 20947 10112 20959 10115
rect 21266 10112 21272 10124
rect 20947 10084 21272 10112
rect 20947 10081 20959 10084
rect 20901 10075 20959 10081
rect 21266 10072 21272 10084
rect 21324 10072 21330 10124
rect 22002 10072 22008 10124
rect 22060 10112 22066 10124
rect 27982 10112 27988 10124
rect 22060 10084 27988 10112
rect 22060 10072 22066 10084
rect 27982 10072 27988 10084
rect 28040 10072 28046 10124
rect 30006 10112 30012 10124
rect 29967 10084 30012 10112
rect 30006 10072 30012 10084
rect 30064 10072 30070 10124
rect 35434 10112 35440 10124
rect 35395 10084 35440 10112
rect 35434 10072 35440 10084
rect 35492 10072 35498 10124
rect 8570 10044 8576 10056
rect 8531 10016 8576 10044
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 16298 10004 16304 10056
rect 16356 10044 16362 10056
rect 16850 10044 16856 10056
rect 16356 10016 16856 10044
rect 16356 10004 16362 10016
rect 16850 10004 16856 10016
rect 16908 10004 16914 10056
rect 23290 10044 23296 10056
rect 23251 10016 23296 10044
rect 23290 10004 23296 10016
rect 23348 10004 23354 10056
rect 30190 10044 30196 10056
rect 30151 10016 30196 10044
rect 30190 10004 30196 10016
rect 30248 10004 30254 10056
rect 32950 10044 32956 10056
rect 32911 10016 32956 10044
rect 32950 10004 32956 10016
rect 33008 10004 33014 10056
rect 34514 9936 34520 9988
rect 34572 9976 34578 9988
rect 35621 9979 35679 9985
rect 35621 9976 35633 9979
rect 34572 9948 35633 9976
rect 34572 9936 34578 9948
rect 35621 9945 35633 9948
rect 35667 9945 35679 9979
rect 35621 9939 35679 9945
rect 13814 9868 13820 9920
rect 13872 9908 13878 9920
rect 14093 9911 14151 9917
rect 14093 9908 14105 9911
rect 13872 9880 14105 9908
rect 13872 9868 13878 9880
rect 14093 9877 14105 9880
rect 14139 9877 14151 9911
rect 14642 9908 14648 9920
rect 14603 9880 14648 9908
rect 14093 9871 14151 9877
rect 14642 9868 14648 9880
rect 14700 9868 14706 9920
rect 16482 9908 16488 9920
rect 16443 9880 16488 9908
rect 16482 9868 16488 9880
rect 16540 9868 16546 9920
rect 18230 9908 18236 9920
rect 18191 9880 18236 9908
rect 18230 9868 18236 9880
rect 18288 9908 18294 9920
rect 18785 9911 18843 9917
rect 18785 9908 18797 9911
rect 18288 9880 18797 9908
rect 18288 9868 18294 9880
rect 18785 9877 18797 9880
rect 18831 9877 18843 9911
rect 18785 9871 18843 9877
rect 19334 9868 19340 9920
rect 19392 9908 19398 9920
rect 19521 9911 19579 9917
rect 19521 9908 19533 9911
rect 19392 9880 19533 9908
rect 19392 9868 19398 9880
rect 19521 9877 19533 9880
rect 19567 9877 19579 9911
rect 21082 9908 21088 9920
rect 21043 9880 21088 9908
rect 19521 9871 19579 9877
rect 21082 9868 21088 9880
rect 21140 9868 21146 9920
rect 21542 9908 21548 9920
rect 21503 9880 21548 9908
rect 21542 9868 21548 9880
rect 21600 9868 21606 9920
rect 22465 9911 22523 9917
rect 22465 9877 22477 9911
rect 22511 9908 22523 9911
rect 22554 9908 22560 9920
rect 22511 9880 22560 9908
rect 22511 9877 22523 9880
rect 22465 9871 22523 9877
rect 22554 9868 22560 9880
rect 22612 9908 22618 9920
rect 23198 9908 23204 9920
rect 22612 9880 23204 9908
rect 22612 9868 22618 9880
rect 23198 9868 23204 9880
rect 23256 9868 23262 9920
rect 24670 9908 24676 9920
rect 24631 9880 24676 9908
rect 24670 9868 24676 9880
rect 24728 9868 24734 9920
rect 1104 9818 38824 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 38824 9818
rect 1104 9744 38824 9766
rect 5074 9704 5080 9716
rect 5035 9676 5080 9704
rect 5074 9664 5080 9676
rect 5132 9664 5138 9716
rect 5442 9704 5448 9716
rect 5403 9676 5448 9704
rect 5442 9664 5448 9676
rect 5500 9664 5506 9716
rect 8478 9704 8484 9716
rect 8220 9676 8484 9704
rect 7101 9639 7159 9645
rect 7101 9605 7113 9639
rect 7147 9636 7159 9639
rect 8110 9636 8116 9648
rect 7147 9608 8116 9636
rect 7147 9605 7159 9608
rect 7101 9599 7159 9605
rect 8110 9596 8116 9608
rect 8168 9596 8174 9648
rect 8220 9645 8248 9676
rect 8478 9664 8484 9676
rect 8536 9664 8542 9716
rect 8570 9664 8576 9716
rect 8628 9704 8634 9716
rect 9217 9707 9275 9713
rect 9217 9704 9229 9707
rect 8628 9676 9229 9704
rect 8628 9664 8634 9676
rect 9217 9673 9229 9676
rect 9263 9673 9275 9707
rect 9217 9667 9275 9673
rect 10873 9707 10931 9713
rect 10873 9673 10885 9707
rect 10919 9704 10931 9707
rect 10962 9704 10968 9716
rect 10919 9676 10968 9704
rect 10919 9673 10931 9676
rect 10873 9667 10931 9673
rect 10962 9664 10968 9676
rect 11020 9664 11026 9716
rect 12710 9704 12716 9716
rect 12671 9676 12716 9704
rect 12710 9664 12716 9676
rect 12768 9664 12774 9716
rect 14001 9707 14059 9713
rect 14001 9673 14013 9707
rect 14047 9704 14059 9707
rect 14458 9704 14464 9716
rect 14047 9676 14464 9704
rect 14047 9673 14059 9676
rect 14001 9667 14059 9673
rect 14458 9664 14464 9676
rect 14516 9664 14522 9716
rect 16850 9664 16856 9716
rect 16908 9704 16914 9716
rect 17405 9707 17463 9713
rect 17405 9704 17417 9707
rect 16908 9676 17417 9704
rect 16908 9664 16914 9676
rect 17405 9673 17417 9676
rect 17451 9673 17463 9707
rect 19426 9704 19432 9716
rect 19387 9676 19432 9704
rect 17405 9667 17463 9673
rect 19426 9664 19432 9676
rect 19484 9664 19490 9716
rect 20993 9707 21051 9713
rect 20993 9673 21005 9707
rect 21039 9704 21051 9707
rect 21266 9704 21272 9716
rect 21039 9676 21272 9704
rect 21039 9673 21051 9676
rect 20993 9667 21051 9673
rect 21266 9664 21272 9676
rect 21324 9664 21330 9716
rect 23014 9704 23020 9716
rect 22975 9676 23020 9704
rect 23014 9664 23020 9676
rect 23072 9664 23078 9716
rect 24670 9704 24676 9716
rect 24136 9676 24676 9704
rect 8205 9639 8263 9645
rect 8205 9605 8217 9639
rect 8251 9605 8263 9639
rect 8205 9599 8263 9605
rect 12161 9639 12219 9645
rect 12161 9605 12173 9639
rect 12207 9636 12219 9639
rect 12250 9636 12256 9648
rect 12207 9608 12256 9636
rect 12207 9605 12219 9608
rect 12161 9599 12219 9605
rect 12250 9596 12256 9608
rect 12308 9596 12314 9648
rect 16301 9639 16359 9645
rect 16301 9605 16313 9639
rect 16347 9636 16359 9639
rect 16666 9636 16672 9648
rect 16347 9608 16672 9636
rect 16347 9605 16359 9608
rect 16301 9599 16359 9605
rect 16666 9596 16672 9608
rect 16724 9596 16730 9648
rect 23658 9636 23664 9648
rect 20824 9608 22048 9636
rect 23619 9608 23664 9636
rect 7193 9503 7251 9509
rect 7193 9469 7205 9503
rect 7239 9500 7251 9503
rect 7834 9500 7840 9512
rect 7239 9472 7840 9500
rect 7239 9469 7251 9472
rect 7193 9463 7251 9469
rect 7834 9460 7840 9472
rect 7892 9460 7898 9512
rect 8297 9503 8355 9509
rect 8297 9469 8309 9503
rect 8343 9500 8355 9503
rect 12268 9500 12296 9596
rect 13449 9571 13507 9577
rect 13449 9568 13461 9571
rect 12912 9540 13461 9568
rect 12912 9500 12940 9540
rect 13449 9537 13461 9540
rect 13495 9568 13507 9571
rect 13722 9568 13728 9580
rect 13495 9540 13728 9568
rect 13495 9537 13507 9540
rect 13449 9531 13507 9537
rect 13722 9528 13728 9540
rect 13780 9528 13786 9580
rect 15565 9571 15623 9577
rect 15565 9537 15577 9571
rect 15611 9568 15623 9571
rect 17034 9568 17040 9580
rect 15611 9540 17040 9568
rect 15611 9537 15623 9540
rect 15565 9531 15623 9537
rect 17034 9528 17040 9540
rect 17092 9528 17098 9580
rect 17865 9571 17923 9577
rect 17865 9537 17877 9571
rect 17911 9568 17923 9571
rect 18230 9568 18236 9580
rect 17911 9540 18236 9568
rect 17911 9537 17923 9540
rect 17865 9531 17923 9537
rect 18230 9528 18236 9540
rect 18288 9568 18294 9580
rect 18509 9571 18567 9577
rect 18509 9568 18521 9571
rect 18288 9540 18521 9568
rect 18288 9528 18294 9540
rect 18509 9537 18521 9540
rect 18555 9537 18567 9571
rect 18690 9568 18696 9580
rect 18651 9540 18696 9568
rect 18509 9531 18567 9537
rect 18690 9528 18696 9540
rect 18748 9528 18754 9580
rect 20824 9512 20852 9608
rect 21361 9571 21419 9577
rect 21361 9537 21373 9571
rect 21407 9568 21419 9571
rect 21910 9568 21916 9580
rect 21407 9540 21916 9568
rect 21407 9537 21419 9540
rect 21361 9531 21419 9537
rect 21910 9528 21916 9540
rect 21968 9528 21974 9580
rect 22020 9577 22048 9608
rect 23658 9596 23664 9608
rect 23716 9596 23722 9648
rect 24136 9580 24164 9676
rect 24670 9664 24676 9676
rect 24728 9664 24734 9716
rect 30006 9704 30012 9716
rect 29967 9676 30012 9704
rect 30006 9664 30012 9676
rect 30064 9664 30070 9716
rect 30190 9664 30196 9716
rect 30248 9704 30254 9716
rect 32950 9704 32956 9716
rect 30248 9676 30420 9704
rect 32911 9676 32956 9704
rect 30248 9664 30254 9676
rect 29733 9639 29791 9645
rect 29733 9605 29745 9639
rect 29779 9636 29791 9639
rect 30282 9636 30288 9648
rect 29779 9608 30288 9636
rect 29779 9605 29791 9608
rect 29733 9599 29791 9605
rect 30282 9596 30288 9608
rect 30340 9596 30346 9648
rect 30392 9636 30420 9676
rect 32950 9664 32956 9676
rect 33008 9664 33014 9716
rect 33413 9707 33471 9713
rect 33413 9673 33425 9707
rect 33459 9704 33471 9707
rect 33502 9704 33508 9716
rect 33459 9676 33508 9704
rect 33459 9673 33471 9676
rect 33413 9667 33471 9673
rect 33502 9664 33508 9676
rect 33560 9664 33566 9716
rect 35434 9704 35440 9716
rect 35395 9676 35440 9704
rect 35434 9664 35440 9676
rect 35492 9664 35498 9716
rect 30469 9639 30527 9645
rect 30469 9636 30481 9639
rect 30392 9608 30481 9636
rect 30469 9605 30481 9608
rect 30515 9636 30527 9639
rect 30834 9636 30840 9648
rect 30515 9608 30840 9636
rect 30515 9605 30527 9608
rect 30469 9599 30527 9605
rect 30834 9596 30840 9608
rect 30892 9596 30898 9648
rect 22005 9571 22063 9577
rect 22005 9537 22017 9571
rect 22051 9537 22063 9571
rect 24118 9568 24124 9580
rect 24031 9540 24124 9568
rect 22005 9531 22063 9537
rect 24118 9528 24124 9540
rect 24176 9528 24182 9580
rect 24305 9571 24363 9577
rect 24305 9537 24317 9571
rect 24351 9568 24363 9571
rect 25409 9571 25467 9577
rect 25409 9568 25421 9571
rect 24351 9540 25421 9568
rect 24351 9537 24363 9540
rect 24305 9531 24363 9537
rect 25409 9537 25421 9540
rect 25455 9537 25467 9571
rect 25409 9531 25467 9537
rect 8343 9472 8984 9500
rect 12268 9472 12940 9500
rect 8343 9469 8355 9472
rect 8297 9463 8355 9469
rect 7466 9432 7472 9444
rect 7379 9404 7472 9432
rect 7392 9373 7420 9404
rect 7466 9392 7472 9404
rect 7524 9432 7530 9444
rect 8570 9432 8576 9444
rect 7524 9404 8576 9432
rect 7524 9392 7530 9404
rect 8570 9392 8576 9404
rect 8628 9392 8634 9444
rect 8956 9376 8984 9472
rect 12986 9460 12992 9512
rect 13044 9500 13050 9512
rect 13265 9503 13323 9509
rect 13265 9500 13277 9503
rect 13044 9472 13277 9500
rect 13044 9460 13050 9472
rect 13265 9469 13277 9472
rect 13311 9500 13323 9503
rect 14461 9503 14519 9509
rect 14461 9500 14473 9503
rect 13311 9472 14473 9500
rect 13311 9469 13323 9472
rect 13265 9463 13323 9469
rect 14461 9469 14473 9472
rect 14507 9469 14519 9503
rect 16758 9500 16764 9512
rect 14461 9463 14519 9469
rect 16592 9472 16764 9500
rect 11885 9435 11943 9441
rect 11885 9401 11897 9435
rect 11931 9432 11943 9435
rect 11931 9404 13032 9432
rect 11931 9401 11943 9404
rect 11885 9395 11943 9401
rect 7377 9367 7435 9373
rect 7377 9333 7389 9367
rect 7423 9333 7435 9367
rect 7834 9364 7840 9376
rect 7795 9336 7840 9364
rect 7377 9327 7435 9333
rect 7834 9324 7840 9336
rect 7892 9324 7898 9376
rect 8386 9324 8392 9376
rect 8444 9364 8450 9376
rect 8481 9367 8539 9373
rect 8481 9364 8493 9367
rect 8444 9336 8493 9364
rect 8444 9324 8450 9336
rect 8481 9333 8493 9336
rect 8527 9333 8539 9367
rect 8938 9364 8944 9376
rect 8899 9336 8944 9364
rect 8481 9327 8539 9333
rect 8938 9324 8944 9336
rect 8996 9324 9002 9376
rect 9674 9324 9680 9376
rect 9732 9364 9738 9376
rect 9769 9367 9827 9373
rect 9769 9364 9781 9367
rect 9732 9336 9781 9364
rect 9732 9324 9738 9336
rect 9769 9333 9781 9336
rect 9815 9364 9827 9367
rect 11606 9364 11612 9376
rect 9815 9336 11612 9364
rect 9815 9333 9827 9336
rect 9769 9327 9827 9333
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 12802 9324 12808 9376
rect 12860 9364 12866 9376
rect 12897 9367 12955 9373
rect 12897 9364 12909 9367
rect 12860 9336 12909 9364
rect 12860 9324 12866 9336
rect 12897 9333 12909 9336
rect 12943 9333 12955 9367
rect 13004 9364 13032 9404
rect 13078 9392 13084 9444
rect 13136 9432 13142 9444
rect 13357 9435 13415 9441
rect 13357 9432 13369 9435
rect 13136 9404 13369 9432
rect 13136 9392 13142 9404
rect 13357 9401 13369 9404
rect 13403 9432 13415 9435
rect 14277 9435 14335 9441
rect 14277 9432 14289 9435
rect 13403 9404 14289 9432
rect 13403 9401 13415 9404
rect 13357 9395 13415 9401
rect 14277 9401 14289 9404
rect 14323 9401 14335 9435
rect 14277 9395 14335 9401
rect 15933 9435 15991 9441
rect 15933 9401 15945 9435
rect 15979 9432 15991 9435
rect 16592 9432 16620 9472
rect 16758 9460 16764 9472
rect 16816 9460 16822 9512
rect 18414 9500 18420 9512
rect 18327 9472 18420 9500
rect 18414 9460 18420 9472
rect 18472 9500 18478 9512
rect 19150 9500 19156 9512
rect 18472 9472 19156 9500
rect 18472 9460 18478 9472
rect 19150 9460 19156 9472
rect 19208 9460 19214 9512
rect 20622 9500 20628 9512
rect 20535 9472 20628 9500
rect 20622 9460 20628 9472
rect 20680 9500 20686 9512
rect 20806 9500 20812 9512
rect 20680 9472 20812 9500
rect 20680 9460 20686 9472
rect 20806 9460 20812 9472
rect 20864 9460 20870 9512
rect 21542 9460 21548 9512
rect 21600 9500 21606 9512
rect 21821 9503 21879 9509
rect 21821 9500 21833 9503
rect 21600 9472 21833 9500
rect 21600 9460 21606 9472
rect 21821 9469 21833 9472
rect 21867 9469 21879 9503
rect 21821 9463 21879 9469
rect 23198 9460 23204 9512
rect 23256 9500 23262 9512
rect 24320 9500 24348 9531
rect 23256 9472 24348 9500
rect 23256 9460 23262 9472
rect 16853 9435 16911 9441
rect 16853 9432 16865 9435
rect 15979 9404 16620 9432
rect 16684 9404 16865 9432
rect 15979 9401 15991 9404
rect 15933 9395 15991 9401
rect 13630 9364 13636 9376
rect 13004 9336 13636 9364
rect 12897 9327 12955 9333
rect 13630 9324 13636 9336
rect 13688 9324 13694 9376
rect 16390 9364 16396 9376
rect 16351 9336 16396 9364
rect 16390 9324 16396 9336
rect 16448 9324 16454 9376
rect 16482 9324 16488 9376
rect 16540 9364 16546 9376
rect 16574 9364 16580 9376
rect 16540 9336 16580 9364
rect 16540 9324 16546 9336
rect 16574 9324 16580 9336
rect 16632 9364 16638 9376
rect 16684 9364 16712 9404
rect 16853 9401 16865 9404
rect 16899 9401 16911 9435
rect 16853 9395 16911 9401
rect 17124 9404 18092 9432
rect 16632 9336 16725 9364
rect 16632 9324 16638 9336
rect 16758 9324 16764 9376
rect 16816 9364 16822 9376
rect 17124 9364 17152 9404
rect 18064 9373 18092 9404
rect 16816 9336 17152 9364
rect 18049 9367 18107 9373
rect 16816 9324 16822 9336
rect 18049 9333 18061 9367
rect 18095 9333 18107 9367
rect 18049 9327 18107 9333
rect 20622 9324 20628 9376
rect 20680 9364 20686 9376
rect 21453 9367 21511 9373
rect 21453 9364 21465 9367
rect 20680 9336 21465 9364
rect 20680 9324 20686 9336
rect 21453 9333 21465 9336
rect 21499 9333 21511 9367
rect 21453 9327 21511 9333
rect 22646 9324 22652 9376
rect 22704 9364 22710 9376
rect 23290 9364 23296 9376
rect 22704 9336 23296 9364
rect 22704 9324 22710 9336
rect 23290 9324 23296 9336
rect 23348 9324 23354 9376
rect 24026 9364 24032 9376
rect 23939 9336 24032 9364
rect 24026 9324 24032 9336
rect 24084 9364 24090 9376
rect 25041 9367 25099 9373
rect 25041 9364 25053 9367
rect 24084 9336 25053 9364
rect 24084 9324 24090 9336
rect 25041 9333 25053 9336
rect 25087 9333 25099 9367
rect 25041 9327 25099 9333
rect 1104 9274 38824 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 38824 9274
rect 1104 9200 38824 9222
rect 13078 9160 13084 9172
rect 13039 9132 13084 9160
rect 13078 9120 13084 9132
rect 13136 9120 13142 9172
rect 13446 9160 13452 9172
rect 13407 9132 13452 9160
rect 13446 9120 13452 9132
rect 13504 9120 13510 9172
rect 13538 9120 13544 9172
rect 13596 9160 13602 9172
rect 13596 9132 13641 9160
rect 13596 9120 13602 9132
rect 16758 9120 16764 9172
rect 16816 9160 16822 9172
rect 17402 9160 17408 9172
rect 16816 9132 17408 9160
rect 16816 9120 16822 9132
rect 17402 9120 17408 9132
rect 17460 9160 17466 9172
rect 17589 9163 17647 9169
rect 17589 9160 17601 9163
rect 17460 9132 17601 9160
rect 17460 9120 17466 9132
rect 17589 9129 17601 9132
rect 17635 9129 17647 9163
rect 17589 9123 17647 9129
rect 18233 9163 18291 9169
rect 18233 9129 18245 9163
rect 18279 9160 18291 9163
rect 18414 9160 18420 9172
rect 18279 9132 18420 9160
rect 18279 9129 18291 9132
rect 18233 9123 18291 9129
rect 18414 9120 18420 9132
rect 18472 9120 18478 9172
rect 18601 9163 18659 9169
rect 18601 9129 18613 9163
rect 18647 9160 18659 9163
rect 18690 9160 18696 9172
rect 18647 9132 18696 9160
rect 18647 9129 18659 9132
rect 18601 9123 18659 9129
rect 18690 9120 18696 9132
rect 18748 9120 18754 9172
rect 19245 9163 19303 9169
rect 19245 9129 19257 9163
rect 19291 9160 19303 9163
rect 19334 9160 19340 9172
rect 19291 9132 19340 9160
rect 19291 9129 19303 9132
rect 19245 9123 19303 9129
rect 19334 9120 19340 9132
rect 19392 9120 19398 9172
rect 21082 9120 21088 9172
rect 21140 9160 21146 9172
rect 21361 9163 21419 9169
rect 21361 9160 21373 9163
rect 21140 9132 21373 9160
rect 21140 9120 21146 9132
rect 21361 9129 21373 9132
rect 21407 9129 21419 9163
rect 24026 9160 24032 9172
rect 23987 9132 24032 9160
rect 21361 9123 21419 9129
rect 24026 9120 24032 9132
rect 24084 9120 24090 9172
rect 28166 9160 28172 9172
rect 28000 9132 28172 9160
rect 12986 9092 12992 9104
rect 12947 9064 12992 9092
rect 12986 9052 12992 9064
rect 13044 9052 13050 9104
rect 16476 9095 16534 9101
rect 16476 9061 16488 9095
rect 16522 9092 16534 9095
rect 16666 9092 16672 9104
rect 16522 9064 16672 9092
rect 16522 9061 16534 9064
rect 16476 9055 16534 9061
rect 16666 9052 16672 9064
rect 16724 9052 16730 9104
rect 22916 9095 22974 9101
rect 22916 9061 22928 9095
rect 22962 9092 22974 9095
rect 23106 9092 23112 9104
rect 22962 9064 23112 9092
rect 22962 9061 22974 9064
rect 22916 9055 22974 9061
rect 23106 9052 23112 9064
rect 23164 9092 23170 9104
rect 24118 9092 24124 9104
rect 23164 9064 24124 9092
rect 23164 9052 23170 9064
rect 24118 9052 24124 9064
rect 24176 9052 24182 9104
rect 7282 9033 7288 9036
rect 7276 9024 7288 9033
rect 7243 8996 7288 9024
rect 7276 8987 7288 8996
rect 7282 8984 7288 8987
rect 7340 8984 7346 9036
rect 10870 9033 10876 9036
rect 10505 9027 10563 9033
rect 10505 8993 10517 9027
rect 10551 9024 10563 9027
rect 10864 9024 10876 9033
rect 10551 8996 10876 9024
rect 10551 8993 10563 8996
rect 10505 8987 10563 8993
rect 10864 8987 10876 8996
rect 10870 8984 10876 8987
rect 10928 8984 10934 9036
rect 12710 8984 12716 9036
rect 12768 9024 12774 9036
rect 16209 9027 16267 9033
rect 16209 9024 16221 9027
rect 12768 8996 16221 9024
rect 12768 8984 12774 8996
rect 16209 8993 16221 8996
rect 16255 9024 16267 9027
rect 16298 9024 16304 9036
rect 16255 8996 16304 9024
rect 16255 8993 16267 8996
rect 16209 8987 16267 8993
rect 16298 8984 16304 8996
rect 16356 8984 16362 9036
rect 21269 9027 21327 9033
rect 21269 8993 21281 9027
rect 21315 9024 21327 9027
rect 21358 9024 21364 9036
rect 21315 8996 21364 9024
rect 21315 8993 21327 8996
rect 21269 8987 21327 8993
rect 21358 8984 21364 8996
rect 21416 8984 21422 9036
rect 26602 8984 26608 9036
rect 26660 9024 26666 9036
rect 28000 9033 28028 9132
rect 28166 9120 28172 9132
rect 28224 9120 28230 9172
rect 27985 9027 28043 9033
rect 27985 9024 27997 9027
rect 26660 8996 27997 9024
rect 26660 8984 26666 8996
rect 27985 8993 27997 8996
rect 28031 8993 28043 9027
rect 27985 8987 28043 8993
rect 28074 8984 28080 9036
rect 28132 9024 28138 9036
rect 28241 9027 28299 9033
rect 28241 9024 28253 9027
rect 28132 8996 28253 9024
rect 28132 8984 28138 8996
rect 28241 8993 28253 8996
rect 28287 8993 28299 9027
rect 28241 8987 28299 8993
rect 6822 8916 6828 8968
rect 6880 8956 6886 8968
rect 7006 8956 7012 8968
rect 6880 8928 7012 8956
rect 6880 8916 6886 8928
rect 7006 8916 7012 8928
rect 7064 8916 7070 8968
rect 10594 8956 10600 8968
rect 10555 8928 10600 8956
rect 10594 8916 10600 8928
rect 10652 8916 10658 8968
rect 13630 8956 13636 8968
rect 13591 8928 13636 8956
rect 13630 8916 13636 8928
rect 13688 8916 13694 8968
rect 18966 8916 18972 8968
rect 19024 8956 19030 8968
rect 19337 8959 19395 8965
rect 19337 8956 19349 8959
rect 19024 8928 19349 8956
rect 19024 8916 19030 8928
rect 19337 8925 19349 8928
rect 19383 8925 19395 8959
rect 19518 8956 19524 8968
rect 19479 8928 19524 8956
rect 19337 8919 19395 8925
rect 19518 8916 19524 8928
rect 19576 8916 19582 8968
rect 21450 8956 21456 8968
rect 21411 8928 21456 8956
rect 21450 8916 21456 8928
rect 21508 8916 21514 8968
rect 22646 8956 22652 8968
rect 22607 8928 22652 8956
rect 22646 8916 22652 8928
rect 22704 8916 22710 8968
rect 6914 8820 6920 8832
rect 6875 8792 6920 8820
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 8386 8820 8392 8832
rect 8347 8792 8392 8820
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 10778 8780 10784 8832
rect 10836 8820 10842 8832
rect 11977 8823 12035 8829
rect 11977 8820 11989 8823
rect 10836 8792 11989 8820
rect 10836 8780 10842 8792
rect 11977 8789 11989 8792
rect 12023 8789 12035 8823
rect 18874 8820 18880 8832
rect 18835 8792 18880 8820
rect 11977 8783 12035 8789
rect 18874 8780 18880 8792
rect 18932 8780 18938 8832
rect 19981 8823 20039 8829
rect 19981 8789 19993 8823
rect 20027 8820 20039 8823
rect 20530 8820 20536 8832
rect 20027 8792 20536 8820
rect 20027 8789 20039 8792
rect 19981 8783 20039 8789
rect 20530 8780 20536 8792
rect 20588 8780 20594 8832
rect 20714 8780 20720 8832
rect 20772 8820 20778 8832
rect 20901 8823 20959 8829
rect 20901 8820 20913 8823
rect 20772 8792 20913 8820
rect 20772 8780 20778 8792
rect 20901 8789 20913 8792
rect 20947 8789 20959 8823
rect 20901 8783 20959 8789
rect 25225 8823 25283 8829
rect 25225 8789 25237 8823
rect 25271 8820 25283 8823
rect 25498 8820 25504 8832
rect 25271 8792 25504 8820
rect 25271 8789 25283 8792
rect 25225 8783 25283 8789
rect 25498 8780 25504 8792
rect 25556 8780 25562 8832
rect 29362 8820 29368 8832
rect 29323 8792 29368 8820
rect 29362 8780 29368 8792
rect 29420 8780 29426 8832
rect 1104 8730 38824 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 38824 8730
rect 1104 8656 38824 8678
rect 10594 8576 10600 8628
rect 10652 8616 10658 8628
rect 11425 8619 11483 8625
rect 11425 8616 11437 8619
rect 10652 8588 11437 8616
rect 10652 8576 10658 8588
rect 11425 8585 11437 8588
rect 11471 8616 11483 8619
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 11471 8588 12173 8616
rect 11471 8585 11483 8588
rect 11425 8579 11483 8585
rect 12161 8585 12173 8588
rect 12207 8585 12219 8619
rect 12161 8579 12219 8585
rect 7834 8508 7840 8560
rect 7892 8548 7898 8560
rect 8205 8551 8263 8557
rect 8205 8548 8217 8551
rect 7892 8520 8217 8548
rect 7892 8508 7898 8520
rect 8205 8517 8217 8520
rect 8251 8517 8263 8551
rect 8205 8511 8263 8517
rect 10318 8508 10324 8560
rect 10376 8548 10382 8560
rect 10413 8551 10471 8557
rect 10413 8548 10425 8551
rect 10376 8520 10425 8548
rect 10376 8508 10382 8520
rect 10413 8517 10425 8520
rect 10459 8517 10471 8551
rect 10413 8511 10471 8517
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8480 10287 8483
rect 10870 8480 10876 8492
rect 10275 8452 10876 8480
rect 10275 8449 10287 8452
rect 10229 8443 10287 8449
rect 10870 8440 10876 8452
rect 10928 8440 10934 8492
rect 10965 8483 11023 8489
rect 10965 8449 10977 8483
rect 11011 8449 11023 8483
rect 12176 8480 12204 8579
rect 13630 8576 13636 8628
rect 13688 8616 13694 8628
rect 14369 8619 14427 8625
rect 14369 8616 14381 8619
rect 13688 8588 14381 8616
rect 13688 8576 13694 8588
rect 14369 8585 14381 8588
rect 14415 8585 14427 8619
rect 14369 8579 14427 8585
rect 16393 8619 16451 8625
rect 16393 8585 16405 8619
rect 16439 8616 16451 8619
rect 16574 8616 16580 8628
rect 16439 8588 16580 8616
rect 16439 8585 16451 8588
rect 16393 8579 16451 8585
rect 16574 8576 16580 8588
rect 16632 8576 16638 8628
rect 17402 8616 17408 8628
rect 17363 8588 17408 8616
rect 17402 8576 17408 8588
rect 17460 8576 17466 8628
rect 18233 8619 18291 8625
rect 18233 8585 18245 8619
rect 18279 8616 18291 8619
rect 18966 8616 18972 8628
rect 18279 8588 18972 8616
rect 18279 8585 18291 8588
rect 18233 8579 18291 8585
rect 18966 8576 18972 8588
rect 19024 8576 19030 8628
rect 19334 8616 19340 8628
rect 19295 8588 19340 8616
rect 19334 8576 19340 8588
rect 19392 8576 19398 8628
rect 20622 8616 20628 8628
rect 20583 8588 20628 8616
rect 20622 8576 20628 8588
rect 20680 8576 20686 8628
rect 21082 8576 21088 8628
rect 21140 8616 21146 8628
rect 21269 8619 21327 8625
rect 21269 8616 21281 8619
rect 21140 8588 21281 8616
rect 21140 8576 21146 8588
rect 21269 8585 21281 8588
rect 21315 8585 21327 8619
rect 23106 8616 23112 8628
rect 23067 8588 23112 8616
rect 21269 8579 21327 8585
rect 23106 8576 23112 8588
rect 23164 8576 23170 8628
rect 26602 8616 26608 8628
rect 26563 8588 26608 8616
rect 26602 8576 26608 8588
rect 26660 8576 26666 8628
rect 28074 8616 28080 8628
rect 28035 8588 28080 8616
rect 28074 8576 28080 8588
rect 28132 8576 28138 8628
rect 28166 8576 28172 8628
rect 28224 8616 28230 8628
rect 28629 8619 28687 8625
rect 28629 8616 28641 8619
rect 28224 8588 28641 8616
rect 28224 8576 28230 8588
rect 28629 8585 28641 8588
rect 28675 8616 28687 8619
rect 28718 8616 28724 8628
rect 28675 8588 28724 8616
rect 28675 8585 28687 8588
rect 28629 8579 28687 8585
rect 28718 8576 28724 8588
rect 28776 8576 28782 8628
rect 13814 8548 13820 8560
rect 13775 8520 13820 8548
rect 13814 8508 13820 8520
rect 13872 8508 13878 8560
rect 19613 8551 19671 8557
rect 19613 8517 19625 8551
rect 19659 8548 19671 8551
rect 19886 8548 19892 8560
rect 19659 8520 19892 8548
rect 19659 8517 19671 8520
rect 19613 8511 19671 8517
rect 19886 8508 19892 8520
rect 19944 8508 19950 8560
rect 20901 8551 20959 8557
rect 20901 8517 20913 8551
rect 20947 8548 20959 8551
rect 21358 8548 21364 8560
rect 20947 8520 21364 8548
rect 20947 8517 20959 8520
rect 20901 8511 20959 8517
rect 21358 8508 21364 8520
rect 21416 8548 21422 8560
rect 21637 8551 21695 8557
rect 21637 8548 21649 8551
rect 21416 8520 21649 8548
rect 21416 8508 21422 8520
rect 21637 8517 21649 8520
rect 21683 8517 21695 8551
rect 21637 8511 21695 8517
rect 12437 8483 12495 8489
rect 12437 8480 12449 8483
rect 12176 8452 12449 8480
rect 10965 8443 11023 8449
rect 12437 8449 12449 8452
rect 12483 8449 12495 8483
rect 12437 8443 12495 8449
rect 17037 8483 17095 8489
rect 17037 8449 17049 8483
rect 17083 8480 17095 8483
rect 17310 8480 17316 8492
rect 17083 8452 17316 8480
rect 17083 8449 17095 8452
rect 17037 8443 17095 8449
rect 6822 8412 6828 8424
rect 6564 8384 6828 8412
rect 6178 8276 6184 8288
rect 6139 8248 6184 8276
rect 6178 8236 6184 8248
rect 6236 8276 6242 8288
rect 6564 8285 6592 8384
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 9953 8415 10011 8421
rect 9953 8381 9965 8415
rect 9999 8412 10011 8415
rect 10594 8412 10600 8424
rect 9999 8384 10600 8412
rect 9999 8381 10011 8384
rect 9953 8375 10011 8381
rect 10594 8372 10600 8384
rect 10652 8412 10658 8424
rect 10778 8412 10784 8424
rect 10652 8384 10784 8412
rect 10652 8372 10658 8384
rect 10778 8372 10784 8384
rect 10836 8372 10842 8424
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 7092 8347 7150 8353
rect 7092 8344 7104 8347
rect 6972 8316 7104 8344
rect 6972 8304 6978 8316
rect 7092 8313 7104 8316
rect 7138 8344 7150 8347
rect 8202 8344 8208 8356
rect 7138 8316 8208 8344
rect 7138 8313 7150 8316
rect 7092 8307 7150 8313
rect 8202 8304 8208 8316
rect 8260 8304 8266 8356
rect 10980 8344 11008 8443
rect 17310 8440 17316 8452
rect 17368 8480 17374 8492
rect 18690 8480 18696 8492
rect 17368 8452 18696 8480
rect 17368 8440 17374 8452
rect 18690 8440 18696 8452
rect 18748 8440 18754 8492
rect 24673 8483 24731 8489
rect 24673 8449 24685 8483
rect 24719 8480 24731 8483
rect 25590 8480 25596 8492
rect 24719 8452 25596 8480
rect 24719 8449 24731 8452
rect 24673 8443 24731 8449
rect 25590 8440 25596 8452
rect 25648 8480 25654 8492
rect 25685 8483 25743 8489
rect 25685 8480 25697 8483
rect 25648 8452 25697 8480
rect 25648 8440 25654 8452
rect 25685 8449 25697 8452
rect 25731 8449 25743 8483
rect 26620 8480 26648 8576
rect 26697 8483 26755 8489
rect 26697 8480 26709 8483
rect 26620 8452 26709 8480
rect 25685 8443 25743 8449
rect 26697 8449 26709 8452
rect 26743 8449 26755 8483
rect 26697 8443 26755 8449
rect 13998 8412 14004 8424
rect 13188 8384 14004 8412
rect 9508 8316 11100 8344
rect 6549 8279 6607 8285
rect 6549 8276 6561 8279
rect 6236 8248 6561 8276
rect 6236 8236 6242 8248
rect 6549 8245 6561 8248
rect 6595 8245 6607 8279
rect 6549 8239 6607 8245
rect 8754 8236 8760 8288
rect 8812 8276 8818 8288
rect 9508 8285 9536 8316
rect 9493 8279 9551 8285
rect 9493 8276 9505 8279
rect 8812 8248 9505 8276
rect 8812 8236 8818 8248
rect 9493 8245 9505 8248
rect 9539 8245 9551 8279
rect 11072 8276 11100 8316
rect 12526 8304 12532 8356
rect 12584 8344 12590 8356
rect 12682 8347 12740 8353
rect 12682 8344 12694 8347
rect 12584 8316 12694 8344
rect 12584 8304 12590 8316
rect 12682 8313 12694 8316
rect 12728 8344 12740 8347
rect 13188 8344 13216 8384
rect 13998 8372 14004 8384
rect 14056 8372 14062 8424
rect 16390 8372 16396 8424
rect 16448 8412 16454 8424
rect 17773 8415 17831 8421
rect 17773 8412 17785 8415
rect 16448 8384 17785 8412
rect 16448 8372 16454 8384
rect 17773 8381 17785 8384
rect 17819 8412 17831 8415
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 17819 8384 18061 8412
rect 17819 8381 17831 8384
rect 17773 8375 17831 8381
rect 18049 8381 18061 8384
rect 18095 8381 18107 8415
rect 18049 8375 18107 8381
rect 19429 8415 19487 8421
rect 19429 8381 19441 8415
rect 19475 8412 19487 8415
rect 20530 8412 20536 8424
rect 19475 8384 20536 8412
rect 19475 8381 19487 8384
rect 19429 8375 19487 8381
rect 20530 8372 20536 8384
rect 20588 8372 20594 8424
rect 20622 8372 20628 8424
rect 20680 8412 20686 8424
rect 20717 8415 20775 8421
rect 20717 8412 20729 8415
rect 20680 8384 20729 8412
rect 20680 8372 20686 8384
rect 20717 8381 20729 8384
rect 20763 8381 20775 8415
rect 25498 8412 25504 8424
rect 25459 8384 25504 8412
rect 20717 8375 20775 8381
rect 25498 8372 25504 8384
rect 25556 8412 25562 8424
rect 26234 8412 26240 8424
rect 25556 8384 26240 8412
rect 25556 8372 25562 8384
rect 26234 8372 26240 8384
rect 26292 8372 26298 8424
rect 12728 8316 13216 8344
rect 12728 8313 12740 8316
rect 12682 8307 12740 8313
rect 13262 8304 13268 8356
rect 13320 8344 13326 8356
rect 14921 8347 14979 8353
rect 14921 8344 14933 8347
rect 13320 8316 14933 8344
rect 13320 8304 13326 8316
rect 14921 8313 14933 8316
rect 14967 8313 14979 8347
rect 14921 8307 14979 8313
rect 15565 8347 15623 8353
rect 15565 8313 15577 8347
rect 15611 8344 15623 8347
rect 15841 8347 15899 8353
rect 15841 8344 15853 8347
rect 15611 8316 15853 8344
rect 15611 8313 15623 8316
rect 15565 8307 15623 8313
rect 15841 8313 15853 8316
rect 15887 8344 15899 8347
rect 16666 8344 16672 8356
rect 15887 8316 16672 8344
rect 15887 8313 15899 8316
rect 15841 8307 15899 8313
rect 16666 8304 16672 8316
rect 16724 8344 16730 8356
rect 16853 8347 16911 8353
rect 16853 8344 16865 8347
rect 16724 8316 16865 8344
rect 16724 8304 16730 8316
rect 16853 8313 16865 8316
rect 16899 8313 16911 8347
rect 16853 8307 16911 8313
rect 19518 8304 19524 8356
rect 19576 8344 19582 8356
rect 20073 8347 20131 8353
rect 20073 8344 20085 8347
rect 19576 8316 20085 8344
rect 19576 8304 19582 8316
rect 20073 8313 20085 8316
rect 20119 8344 20131 8347
rect 20162 8344 20168 8356
rect 20119 8316 20168 8344
rect 20119 8313 20131 8316
rect 20073 8307 20131 8313
rect 20162 8304 20168 8316
rect 20220 8344 20226 8356
rect 21450 8344 21456 8356
rect 20220 8316 21456 8344
rect 20220 8304 20226 8316
rect 21450 8304 21456 8316
rect 21508 8304 21514 8356
rect 25041 8347 25099 8353
rect 25041 8313 25053 8347
rect 25087 8344 25099 8347
rect 25593 8347 25651 8353
rect 25593 8344 25605 8347
rect 25087 8316 25605 8344
rect 25087 8313 25099 8316
rect 25041 8307 25099 8313
rect 25593 8313 25605 8316
rect 25639 8344 25651 8347
rect 26142 8344 26148 8356
rect 25639 8316 26148 8344
rect 25639 8313 25651 8316
rect 25593 8307 25651 8313
rect 26142 8304 26148 8316
rect 26200 8304 26206 8356
rect 26786 8304 26792 8356
rect 26844 8344 26850 8356
rect 26942 8347 27000 8353
rect 26942 8344 26954 8347
rect 26844 8316 26954 8344
rect 26844 8304 26850 8316
rect 26942 8313 26954 8316
rect 26988 8313 27000 8347
rect 26942 8307 27000 8313
rect 11238 8276 11244 8288
rect 11072 8248 11244 8276
rect 9493 8239 9551 8245
rect 11238 8236 11244 8248
rect 11296 8236 11302 8288
rect 16298 8276 16304 8288
rect 16259 8248 16304 8276
rect 16298 8236 16304 8248
rect 16356 8236 16362 8288
rect 16758 8276 16764 8288
rect 16719 8248 16764 8276
rect 16758 8236 16764 8248
rect 16816 8236 16822 8288
rect 22646 8236 22652 8288
rect 22704 8276 22710 8288
rect 22741 8279 22799 8285
rect 22741 8276 22753 8279
rect 22704 8248 22753 8276
rect 22704 8236 22710 8248
rect 22741 8245 22753 8248
rect 22787 8276 22799 8279
rect 22922 8276 22928 8288
rect 22787 8248 22928 8276
rect 22787 8245 22799 8248
rect 22741 8239 22799 8245
rect 22922 8236 22928 8248
rect 22980 8236 22986 8288
rect 25130 8276 25136 8288
rect 25091 8248 25136 8276
rect 25130 8236 25136 8248
rect 25188 8236 25194 8288
rect 1104 8186 38824 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 38824 8186
rect 1104 8112 38824 8134
rect 8297 8075 8355 8081
rect 8297 8041 8309 8075
rect 8343 8072 8355 8075
rect 8386 8072 8392 8084
rect 8343 8044 8392 8072
rect 8343 8041 8355 8044
rect 8297 8035 8355 8041
rect 8386 8032 8392 8044
rect 8444 8032 8450 8084
rect 12526 8072 12532 8084
rect 12487 8044 12532 8072
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 13446 8032 13452 8084
rect 13504 8072 13510 8084
rect 13541 8075 13599 8081
rect 13541 8072 13553 8075
rect 13504 8044 13553 8072
rect 13504 8032 13510 8044
rect 13541 8041 13553 8044
rect 13587 8041 13599 8075
rect 16666 8072 16672 8084
rect 16627 8044 16672 8072
rect 13541 8035 13599 8041
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 17310 8072 17316 8084
rect 17271 8044 17316 8072
rect 17310 8032 17316 8044
rect 17368 8072 17374 8084
rect 17957 8075 18015 8081
rect 17957 8072 17969 8075
rect 17368 8044 17969 8072
rect 17368 8032 17374 8044
rect 17957 8041 17969 8044
rect 18003 8041 18015 8075
rect 17957 8035 18015 8041
rect 19613 8075 19671 8081
rect 19613 8041 19625 8075
rect 19659 8072 19671 8075
rect 19978 8072 19984 8084
rect 19659 8044 19984 8072
rect 19659 8041 19671 8044
rect 19613 8035 19671 8041
rect 19978 8032 19984 8044
rect 20036 8072 20042 8084
rect 20622 8072 20628 8084
rect 20036 8044 20628 8072
rect 20036 8032 20042 8044
rect 20622 8032 20628 8044
rect 20680 8032 20686 8084
rect 21177 8075 21235 8081
rect 21177 8041 21189 8075
rect 21223 8072 21235 8075
rect 21450 8072 21456 8084
rect 21223 8044 21456 8072
rect 21223 8041 21235 8044
rect 21177 8035 21235 8041
rect 21450 8032 21456 8044
rect 21508 8032 21514 8084
rect 26234 8032 26240 8084
rect 26292 8072 26298 8084
rect 26881 8075 26939 8081
rect 26881 8072 26893 8075
rect 26292 8044 26893 8072
rect 26292 8032 26298 8044
rect 26881 8041 26893 8044
rect 26927 8041 26939 8075
rect 26881 8035 26939 8041
rect 27249 8075 27307 8081
rect 27249 8041 27261 8075
rect 27295 8072 27307 8075
rect 27614 8072 27620 8084
rect 27295 8044 27620 8072
rect 27295 8041 27307 8044
rect 27249 8035 27307 8041
rect 27614 8032 27620 8044
rect 27672 8072 27678 8084
rect 28074 8072 28080 8084
rect 27672 8044 28080 8072
rect 27672 8032 27678 8044
rect 28074 8032 28080 8044
rect 28132 8032 28138 8084
rect 5261 8007 5319 8013
rect 5261 7973 5273 8007
rect 5307 8004 5319 8007
rect 5534 8004 5540 8016
rect 5307 7976 5540 8004
rect 5307 7973 5319 7976
rect 5261 7967 5319 7973
rect 5534 7964 5540 7976
rect 5592 8004 5598 8016
rect 5712 8007 5770 8013
rect 5712 8004 5724 8007
rect 5592 7976 5724 8004
rect 5592 7964 5598 7976
rect 5712 7973 5724 7976
rect 5758 8004 5770 8007
rect 7834 8004 7840 8016
rect 5758 7976 7840 8004
rect 5758 7973 5770 7976
rect 5712 7967 5770 7973
rect 7834 7964 7840 7976
rect 7892 7964 7898 8016
rect 12713 8007 12771 8013
rect 12713 7973 12725 8007
rect 12759 8004 12771 8007
rect 13722 8004 13728 8016
rect 12759 7976 13728 8004
rect 12759 7973 12771 7976
rect 12713 7967 12771 7973
rect 13722 7964 13728 7976
rect 13780 7964 13786 8016
rect 16298 8004 16304 8016
rect 15304 7976 16304 8004
rect 5445 7939 5503 7945
rect 5445 7905 5457 7939
rect 5491 7936 5503 7939
rect 6178 7936 6184 7948
rect 5491 7908 6184 7936
rect 5491 7905 5503 7908
rect 5445 7899 5503 7905
rect 6178 7896 6184 7908
rect 6236 7896 6242 7948
rect 10220 7939 10278 7945
rect 10220 7905 10232 7939
rect 10266 7936 10278 7939
rect 10502 7936 10508 7948
rect 10266 7908 10508 7936
rect 10266 7905 10278 7908
rect 10220 7899 10278 7905
rect 10502 7896 10508 7908
rect 10560 7896 10566 7948
rect 13265 7939 13323 7945
rect 13265 7905 13277 7939
rect 13311 7936 13323 7939
rect 13538 7936 13544 7948
rect 13311 7908 13544 7936
rect 13311 7905 13323 7908
rect 13265 7899 13323 7905
rect 13538 7896 13544 7908
rect 13596 7896 13602 7948
rect 15304 7945 15332 7976
rect 16298 7964 16304 7976
rect 16356 7964 16362 8016
rect 21726 8013 21732 8016
rect 21720 8004 21732 8013
rect 21687 7976 21732 8004
rect 21720 7967 21732 7976
rect 21726 7964 21732 7967
rect 21784 7964 21790 8016
rect 23845 8007 23903 8013
rect 23845 7973 23857 8007
rect 23891 8004 23903 8007
rect 24182 8007 24240 8013
rect 24182 8004 24194 8007
rect 23891 7976 24194 8004
rect 23891 7973 23903 7976
rect 23845 7967 23903 7973
rect 24182 7973 24194 7976
rect 24228 8004 24240 8007
rect 25314 8004 25320 8016
rect 24228 7976 25320 8004
rect 24228 7973 24240 7976
rect 24182 7967 24240 7973
rect 25314 7964 25320 7976
rect 25372 7964 25378 8016
rect 26786 8004 26792 8016
rect 26747 7976 26792 8004
rect 26786 7964 26792 7976
rect 26844 8004 26850 8016
rect 27341 8007 27399 8013
rect 27341 8004 27353 8007
rect 26844 7976 27353 8004
rect 26844 7964 26850 7976
rect 27341 7973 27353 7976
rect 27387 8004 27399 8007
rect 27798 8004 27804 8016
rect 27387 7976 27804 8004
rect 27387 7973 27399 7976
rect 27341 7967 27399 7973
rect 27798 7964 27804 7976
rect 27856 7964 27862 8016
rect 28810 7964 28816 8016
rect 28868 8004 28874 8016
rect 28988 8007 29046 8013
rect 28988 8004 29000 8007
rect 28868 7976 29000 8004
rect 28868 7964 28874 7976
rect 28988 7973 29000 7976
rect 29034 8004 29046 8007
rect 29362 8004 29368 8016
rect 29034 7976 29368 8004
rect 29034 7973 29046 7976
rect 28988 7967 29046 7973
rect 29362 7964 29368 7976
rect 29420 7964 29426 8016
rect 15289 7939 15347 7945
rect 15289 7905 15301 7939
rect 15335 7905 15347 7939
rect 15545 7939 15603 7945
rect 15545 7936 15557 7939
rect 15289 7899 15347 7905
rect 15396 7908 15557 7936
rect 7282 7828 7288 7880
rect 7340 7868 7346 7880
rect 7469 7871 7527 7877
rect 7469 7868 7481 7871
rect 7340 7840 7481 7868
rect 7340 7828 7346 7840
rect 7469 7837 7481 7840
rect 7515 7868 7527 7871
rect 8386 7868 8392 7880
rect 7515 7840 8392 7868
rect 7515 7837 7527 7840
rect 7469 7831 7527 7837
rect 8386 7828 8392 7840
rect 8444 7828 8450 7880
rect 8573 7871 8631 7877
rect 8573 7837 8585 7871
rect 8619 7868 8631 7871
rect 8754 7868 8760 7880
rect 8619 7840 8760 7868
rect 8619 7837 8631 7840
rect 8573 7831 8631 7837
rect 8754 7828 8760 7840
rect 8812 7828 8818 7880
rect 9950 7868 9956 7880
rect 9911 7840 9956 7868
rect 9950 7828 9956 7840
rect 10008 7828 10014 7880
rect 13725 7871 13783 7877
rect 13725 7837 13737 7871
rect 13771 7868 13783 7871
rect 13998 7868 14004 7880
rect 13771 7840 14004 7868
rect 13771 7837 13783 7840
rect 13725 7831 13783 7837
rect 13998 7828 14004 7840
rect 14056 7828 14062 7880
rect 15194 7828 15200 7880
rect 15252 7868 15258 7880
rect 15396 7868 15424 7908
rect 15545 7905 15557 7908
rect 15591 7905 15603 7939
rect 17770 7936 17776 7948
rect 17731 7908 17776 7936
rect 15545 7899 15603 7905
rect 17770 7896 17776 7908
rect 17828 7896 17834 7948
rect 28718 7936 28724 7948
rect 28679 7908 28724 7936
rect 28718 7896 28724 7908
rect 28776 7896 28782 7948
rect 15252 7840 15424 7868
rect 15252 7828 15258 7840
rect 18138 7828 18144 7880
rect 18196 7868 18202 7880
rect 18874 7868 18880 7880
rect 18196 7840 18880 7868
rect 18196 7828 18202 7840
rect 18874 7828 18880 7840
rect 18932 7868 18938 7880
rect 19705 7871 19763 7877
rect 19705 7868 19717 7871
rect 18932 7840 19717 7868
rect 18932 7828 18938 7840
rect 19705 7837 19717 7840
rect 19751 7837 19763 7871
rect 19886 7868 19892 7880
rect 19847 7840 19892 7868
rect 19705 7831 19763 7837
rect 19886 7828 19892 7840
rect 19944 7828 19950 7880
rect 21450 7868 21456 7880
rect 21411 7840 21456 7868
rect 21450 7828 21456 7840
rect 21508 7828 21514 7880
rect 23934 7868 23940 7880
rect 23895 7840 23940 7868
rect 23934 7828 23940 7840
rect 23992 7828 23998 7880
rect 26694 7828 26700 7880
rect 26752 7868 26758 7880
rect 27433 7871 27491 7877
rect 27433 7868 27445 7871
rect 26752 7840 27445 7868
rect 26752 7828 26758 7840
rect 27433 7837 27445 7840
rect 27479 7837 27491 7871
rect 27433 7831 27491 7837
rect 18969 7803 19027 7809
rect 18969 7769 18981 7803
rect 19015 7800 19027 7803
rect 19150 7800 19156 7812
rect 19015 7772 19156 7800
rect 19015 7769 19027 7772
rect 18969 7763 19027 7769
rect 19150 7760 19156 7772
rect 19208 7760 19214 7812
rect 6822 7732 6828 7744
rect 6783 7704 6828 7732
rect 6822 7692 6828 7704
rect 6880 7692 6886 7744
rect 7926 7732 7932 7744
rect 7887 7704 7932 7732
rect 7926 7692 7932 7704
rect 7984 7692 7990 7744
rect 11330 7732 11336 7744
rect 11291 7704 11336 7732
rect 11330 7692 11336 7704
rect 11388 7692 11394 7744
rect 19242 7732 19248 7744
rect 19203 7704 19248 7732
rect 19242 7692 19248 7704
rect 19300 7692 19306 7744
rect 21082 7692 21088 7744
rect 21140 7732 21146 7744
rect 22833 7735 22891 7741
rect 22833 7732 22845 7735
rect 21140 7704 22845 7732
rect 21140 7692 21146 7704
rect 22833 7701 22845 7704
rect 22879 7701 22891 7735
rect 22833 7695 22891 7701
rect 25317 7735 25375 7741
rect 25317 7701 25329 7735
rect 25363 7732 25375 7735
rect 25958 7732 25964 7744
rect 25363 7704 25964 7732
rect 25363 7701 25375 7704
rect 25317 7695 25375 7701
rect 25958 7692 25964 7704
rect 26016 7692 26022 7744
rect 30098 7732 30104 7744
rect 30059 7704 30104 7732
rect 30098 7692 30104 7704
rect 30156 7692 30162 7744
rect 1104 7642 38824 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 38824 7642
rect 1104 7568 38824 7590
rect 7377 7531 7435 7537
rect 7377 7497 7389 7531
rect 7423 7528 7435 7531
rect 8386 7528 8392 7540
rect 7423 7500 8392 7528
rect 7423 7497 7435 7500
rect 7377 7491 7435 7497
rect 8386 7488 8392 7500
rect 8444 7528 8450 7540
rect 9585 7531 9643 7537
rect 9585 7528 9597 7531
rect 8444 7500 9597 7528
rect 8444 7488 8450 7500
rect 9585 7497 9597 7500
rect 9631 7497 9643 7531
rect 9585 7491 9643 7497
rect 9950 7488 9956 7540
rect 10008 7528 10014 7540
rect 10137 7531 10195 7537
rect 10137 7528 10149 7531
rect 10008 7500 10149 7528
rect 10008 7488 10014 7500
rect 10137 7497 10149 7500
rect 10183 7497 10195 7531
rect 10502 7528 10508 7540
rect 10463 7500 10508 7528
rect 10137 7491 10195 7497
rect 10502 7488 10508 7500
rect 10560 7488 10566 7540
rect 17497 7531 17555 7537
rect 17497 7497 17509 7531
rect 17543 7528 17555 7531
rect 19242 7528 19248 7540
rect 17543 7500 19248 7528
rect 17543 7497 17555 7500
rect 17497 7491 17555 7497
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7392 5135 7395
rect 5810 7392 5816 7404
rect 5123 7364 5672 7392
rect 5771 7364 5816 7392
rect 5123 7361 5135 7364
rect 5077 7355 5135 7361
rect 4709 7327 4767 7333
rect 4709 7293 4721 7327
rect 4755 7324 4767 7327
rect 5534 7324 5540 7336
rect 4755 7296 5540 7324
rect 4755 7293 4767 7296
rect 4709 7287 4767 7293
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 5644 7333 5672 7364
rect 5810 7352 5816 7364
rect 5868 7352 5874 7404
rect 10520 7392 10548 7488
rect 11149 7395 11207 7401
rect 11149 7392 11161 7395
rect 10520 7364 11161 7392
rect 11149 7361 11161 7364
rect 11195 7361 11207 7395
rect 11149 7355 11207 7361
rect 5629 7327 5687 7333
rect 5629 7293 5641 7327
rect 5675 7324 5687 7327
rect 6730 7324 6736 7336
rect 5675 7296 6736 7324
rect 5675 7293 5687 7296
rect 5629 7287 5687 7293
rect 6730 7284 6736 7296
rect 6788 7284 6794 7336
rect 7929 7327 7987 7333
rect 7929 7293 7941 7327
rect 7975 7324 7987 7327
rect 8205 7327 8263 7333
rect 8205 7324 8217 7327
rect 7975 7296 8217 7324
rect 7975 7293 7987 7296
rect 7929 7287 7987 7293
rect 8205 7293 8217 7296
rect 8251 7293 8263 7327
rect 11164 7324 11192 7355
rect 11238 7352 11244 7404
rect 11296 7392 11302 7404
rect 11296 7364 11341 7392
rect 11296 7352 11302 7364
rect 11698 7324 11704 7336
rect 11164 7296 11704 7324
rect 8205 7287 8263 7293
rect 11698 7284 11704 7296
rect 11756 7284 11762 7336
rect 12437 7327 12495 7333
rect 12437 7293 12449 7327
rect 12483 7324 12495 7327
rect 12526 7324 12532 7336
rect 12483 7296 12532 7324
rect 12483 7293 12495 7296
rect 12437 7287 12495 7293
rect 12526 7284 12532 7296
rect 12584 7324 12590 7336
rect 12989 7327 13047 7333
rect 12989 7324 13001 7327
rect 12584 7296 13001 7324
rect 12584 7284 12590 7296
rect 12989 7293 13001 7296
rect 13035 7293 13047 7327
rect 12989 7287 13047 7293
rect 13817 7327 13875 7333
rect 13817 7293 13829 7327
rect 13863 7324 13875 7327
rect 13909 7327 13967 7333
rect 13909 7324 13921 7327
rect 13863 7296 13921 7324
rect 13863 7293 13875 7296
rect 13817 7287 13875 7293
rect 13909 7293 13921 7296
rect 13955 7324 13967 7327
rect 16853 7327 16911 7333
rect 13955 7296 15976 7324
rect 13955 7293 13967 7296
rect 13909 7287 13967 7293
rect 4341 7259 4399 7265
rect 4341 7225 4353 7259
rect 4387 7256 4399 7259
rect 5810 7256 5816 7268
rect 4387 7228 5816 7256
rect 4387 7225 4399 7228
rect 4341 7219 4399 7225
rect 5810 7216 5816 7228
rect 5868 7216 5874 7268
rect 7745 7259 7803 7265
rect 7745 7225 7757 7259
rect 7791 7256 7803 7259
rect 8450 7259 8508 7265
rect 8450 7256 8462 7259
rect 7791 7228 8462 7256
rect 7791 7225 7803 7228
rect 7745 7219 7803 7225
rect 8450 7225 8462 7228
rect 8496 7256 8508 7259
rect 11057 7259 11115 7265
rect 11057 7256 11069 7259
rect 8496 7228 11069 7256
rect 8496 7225 8508 7228
rect 8450 7219 8508 7225
rect 11057 7225 11069 7228
rect 11103 7256 11115 7259
rect 11330 7256 11336 7268
rect 11103 7228 11336 7256
rect 11103 7225 11115 7228
rect 11057 7219 11115 7225
rect 11330 7216 11336 7228
rect 11388 7256 11394 7268
rect 12069 7259 12127 7265
rect 12069 7256 12081 7259
rect 11388 7228 12081 7256
rect 11388 7216 11394 7228
rect 12069 7225 12081 7228
rect 12115 7225 12127 7259
rect 12069 7219 12127 7225
rect 13354 7216 13360 7268
rect 13412 7256 13418 7268
rect 15948 7265 15976 7296
rect 16853 7293 16865 7327
rect 16899 7324 16911 7327
rect 17512 7324 17540 7491
rect 19242 7488 19248 7500
rect 19300 7488 19306 7540
rect 19886 7488 19892 7540
rect 19944 7528 19950 7540
rect 20809 7531 20867 7537
rect 20809 7528 20821 7531
rect 19944 7500 20821 7528
rect 19944 7488 19950 7500
rect 20809 7497 20821 7500
rect 20855 7497 20867 7531
rect 20809 7491 20867 7497
rect 21726 7488 21732 7540
rect 21784 7528 21790 7540
rect 21821 7531 21879 7537
rect 21821 7528 21833 7531
rect 21784 7500 21833 7528
rect 21784 7488 21790 7500
rect 21821 7497 21833 7500
rect 21867 7497 21879 7531
rect 25314 7528 25320 7540
rect 25275 7500 25320 7528
rect 21821 7491 21879 7497
rect 25314 7488 25320 7500
rect 25372 7488 25378 7540
rect 25958 7528 25964 7540
rect 25919 7500 25964 7528
rect 25958 7488 25964 7500
rect 26016 7488 26022 7540
rect 26329 7531 26387 7537
rect 26329 7497 26341 7531
rect 26375 7528 26387 7531
rect 26418 7528 26424 7540
rect 26375 7500 26424 7528
rect 26375 7497 26387 7500
rect 26329 7491 26387 7497
rect 26418 7488 26424 7500
rect 26476 7528 26482 7540
rect 26602 7528 26608 7540
rect 26476 7500 26608 7528
rect 26476 7488 26482 7500
rect 26602 7488 26608 7500
rect 26660 7488 26666 7540
rect 27798 7528 27804 7540
rect 27759 7500 27804 7528
rect 27798 7488 27804 7500
rect 27856 7488 27862 7540
rect 28445 7531 28503 7537
rect 28445 7497 28457 7531
rect 28491 7528 28503 7531
rect 28718 7528 28724 7540
rect 28491 7500 28724 7528
rect 28491 7497 28503 7500
rect 28445 7491 28503 7497
rect 28718 7488 28724 7500
rect 28776 7488 28782 7540
rect 35250 7488 35256 7540
rect 35308 7528 35314 7540
rect 35526 7528 35532 7540
rect 35308 7500 35532 7528
rect 35308 7488 35314 7500
rect 35526 7488 35532 7500
rect 35584 7488 35590 7540
rect 25976 7392 26004 7488
rect 28736 7392 28764 7488
rect 29270 7392 29276 7404
rect 25976 7364 26556 7392
rect 28736 7364 29276 7392
rect 26528 7336 26556 7364
rect 29270 7352 29276 7364
rect 29328 7352 29334 7404
rect 16899 7296 17540 7324
rect 16899 7293 16911 7296
rect 16853 7287 16911 7293
rect 18046 7284 18052 7336
rect 18104 7324 18110 7336
rect 19150 7333 19156 7336
rect 18693 7327 18751 7333
rect 18693 7324 18705 7327
rect 18104 7296 18705 7324
rect 18104 7284 18110 7296
rect 18693 7293 18705 7296
rect 18739 7324 18751 7327
rect 18877 7327 18935 7333
rect 18877 7324 18889 7327
rect 18739 7296 18889 7324
rect 18739 7293 18751 7296
rect 18693 7287 18751 7293
rect 18877 7293 18889 7296
rect 18923 7293 18935 7327
rect 19144 7324 19156 7333
rect 19111 7296 19156 7324
rect 18877 7287 18935 7293
rect 19144 7287 19156 7296
rect 19150 7284 19156 7287
rect 19208 7284 19214 7336
rect 21450 7284 21456 7336
rect 21508 7324 21514 7336
rect 21545 7327 21603 7333
rect 21545 7324 21557 7327
rect 21508 7296 21557 7324
rect 21508 7284 21514 7296
rect 21545 7293 21557 7296
rect 21591 7324 21603 7327
rect 22922 7324 22928 7336
rect 21591 7296 22928 7324
rect 21591 7293 21603 7296
rect 21545 7287 21603 7293
rect 22922 7284 22928 7296
rect 22980 7324 22986 7336
rect 23109 7327 23167 7333
rect 23109 7324 23121 7327
rect 22980 7296 23121 7324
rect 22980 7284 22986 7296
rect 23109 7293 23121 7296
rect 23155 7324 23167 7327
rect 23477 7327 23535 7333
rect 23477 7324 23489 7327
rect 23155 7296 23489 7324
rect 23155 7293 23167 7296
rect 23109 7287 23167 7293
rect 23477 7293 23489 7296
rect 23523 7324 23535 7327
rect 23934 7324 23940 7336
rect 23523 7296 23940 7324
rect 23523 7293 23535 7296
rect 23477 7287 23535 7293
rect 23934 7284 23940 7296
rect 23992 7324 23998 7336
rect 26418 7324 26424 7336
rect 23992 7296 26424 7324
rect 23992 7284 23998 7296
rect 26418 7284 26424 7296
rect 26476 7284 26482 7336
rect 26510 7284 26516 7336
rect 26568 7324 26574 7336
rect 26677 7327 26735 7333
rect 26677 7324 26689 7327
rect 26568 7296 26689 7324
rect 26568 7284 26574 7296
rect 26677 7293 26689 7296
rect 26723 7293 26735 7327
rect 26677 7287 26735 7293
rect 29362 7284 29368 7336
rect 29420 7324 29426 7336
rect 29540 7327 29598 7333
rect 29540 7324 29552 7327
rect 29420 7296 29552 7324
rect 29420 7284 29426 7296
rect 29540 7293 29552 7296
rect 29586 7324 29598 7327
rect 30098 7324 30104 7336
rect 29586 7296 30104 7324
rect 29586 7293 29598 7296
rect 29540 7287 29598 7293
rect 30098 7284 30104 7296
rect 30156 7284 30162 7336
rect 13449 7259 13507 7265
rect 13449 7256 13461 7259
rect 13412 7228 13461 7256
rect 13412 7216 13418 7228
rect 13449 7225 13461 7228
rect 13495 7256 13507 7259
rect 14154 7259 14212 7265
rect 14154 7256 14166 7259
rect 13495 7228 14166 7256
rect 13495 7225 13507 7228
rect 13449 7219 13507 7225
rect 14154 7225 14166 7228
rect 14200 7225 14212 7259
rect 14154 7219 14212 7225
rect 15933 7259 15991 7265
rect 15933 7225 15945 7259
rect 15979 7256 15991 7259
rect 16298 7256 16304 7268
rect 15979 7228 16304 7256
rect 15979 7225 15991 7228
rect 15933 7219 15991 7225
rect 16298 7216 16304 7228
rect 16356 7256 16362 7268
rect 18064 7256 18092 7284
rect 16356 7228 18092 7256
rect 16356 7216 16362 7228
rect 18138 7216 18144 7268
rect 18196 7256 18202 7268
rect 24210 7265 24216 7268
rect 18325 7259 18383 7265
rect 18325 7256 18337 7259
rect 18196 7228 18337 7256
rect 18196 7216 18202 7228
rect 18325 7225 18337 7228
rect 18371 7225 18383 7259
rect 24204 7256 24216 7265
rect 24171 7228 24216 7256
rect 18325 7219 18383 7225
rect 24204 7219 24216 7228
rect 24210 7216 24216 7219
rect 24268 7216 24274 7268
rect 5166 7188 5172 7200
rect 5127 7160 5172 7188
rect 5166 7148 5172 7160
rect 5224 7148 5230 7200
rect 6178 7188 6184 7200
rect 6139 7160 6184 7188
rect 6178 7148 6184 7160
rect 6236 7188 6242 7200
rect 7929 7191 7987 7197
rect 7929 7188 7941 7191
rect 6236 7160 7941 7188
rect 6236 7148 6242 7160
rect 7929 7157 7941 7160
rect 7975 7188 7987 7191
rect 8021 7191 8079 7197
rect 8021 7188 8033 7191
rect 7975 7160 8033 7188
rect 7975 7157 7987 7160
rect 7929 7151 7987 7157
rect 8021 7157 8033 7160
rect 8067 7157 8079 7191
rect 10686 7188 10692 7200
rect 10647 7160 10692 7188
rect 8021 7151 8079 7157
rect 10686 7148 10692 7160
rect 10744 7148 10750 7200
rect 12621 7191 12679 7197
rect 12621 7157 12633 7191
rect 12667 7188 12679 7191
rect 12894 7188 12900 7200
rect 12667 7160 12900 7188
rect 12667 7157 12679 7160
rect 12621 7151 12679 7157
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 15194 7148 15200 7200
rect 15252 7188 15258 7200
rect 15289 7191 15347 7197
rect 15289 7188 15301 7191
rect 15252 7160 15301 7188
rect 15252 7148 15258 7160
rect 15289 7157 15301 7160
rect 15335 7157 15347 7191
rect 17034 7188 17040 7200
rect 16995 7160 17040 7188
rect 15289 7151 15347 7157
rect 17034 7148 17040 7160
rect 17092 7148 17098 7200
rect 17770 7148 17776 7200
rect 17828 7188 17834 7200
rect 17865 7191 17923 7197
rect 17865 7188 17877 7191
rect 17828 7160 17877 7188
rect 17828 7148 17834 7160
rect 17865 7157 17877 7160
rect 17911 7188 17923 7191
rect 18230 7188 18236 7200
rect 17911 7160 18236 7188
rect 17911 7157 17923 7160
rect 17865 7151 17923 7157
rect 18230 7148 18236 7160
rect 18288 7148 18294 7200
rect 20254 7188 20260 7200
rect 20215 7160 20260 7188
rect 20254 7148 20260 7160
rect 20312 7148 20318 7200
rect 30374 7148 30380 7200
rect 30432 7188 30438 7200
rect 30653 7191 30711 7197
rect 30653 7188 30665 7191
rect 30432 7160 30665 7188
rect 30432 7148 30438 7160
rect 30653 7157 30665 7160
rect 30699 7157 30711 7191
rect 30653 7151 30711 7157
rect 1104 7098 38824 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 38824 7098
rect 1104 7024 38824 7046
rect 7742 6984 7748 6996
rect 7703 6956 7748 6984
rect 7742 6944 7748 6956
rect 7800 6944 7806 6996
rect 7837 6987 7895 6993
rect 7837 6953 7849 6987
rect 7883 6984 7895 6987
rect 7926 6984 7932 6996
rect 7883 6956 7932 6984
rect 7883 6953 7895 6956
rect 7837 6947 7895 6953
rect 7926 6944 7932 6956
rect 7984 6944 7990 6996
rect 8478 6984 8484 6996
rect 8439 6956 8484 6984
rect 8478 6944 8484 6956
rect 8536 6944 8542 6996
rect 11698 6984 11704 6996
rect 11659 6956 11704 6984
rect 11698 6944 11704 6956
rect 11756 6944 11762 6996
rect 13446 6944 13452 6996
rect 13504 6984 13510 6996
rect 13998 6984 14004 6996
rect 13504 6956 14004 6984
rect 13504 6944 13510 6956
rect 13998 6944 14004 6956
rect 14056 6944 14062 6996
rect 19978 6984 19984 6996
rect 19939 6956 19984 6984
rect 19978 6944 19984 6956
rect 20036 6944 20042 6996
rect 27249 6987 27307 6993
rect 27249 6953 27261 6987
rect 27295 6984 27307 6987
rect 27798 6984 27804 6996
rect 27295 6956 27804 6984
rect 27295 6953 27307 6956
rect 27249 6947 27307 6953
rect 27798 6944 27804 6956
rect 27856 6944 27862 6996
rect 29181 6987 29239 6993
rect 29181 6984 29193 6987
rect 28092 6956 29193 6984
rect 18138 6916 18144 6928
rect 17880 6888 18144 6916
rect 5160 6851 5218 6857
rect 5160 6817 5172 6851
rect 5206 6848 5218 6851
rect 5442 6848 5448 6860
rect 5206 6820 5448 6848
rect 5206 6817 5218 6820
rect 5160 6811 5218 6817
rect 5442 6808 5448 6820
rect 5500 6848 5506 6860
rect 6822 6848 6828 6860
rect 5500 6820 6828 6848
rect 5500 6808 5506 6820
rect 6822 6808 6828 6820
rect 6880 6808 6886 6860
rect 9950 6808 9956 6860
rect 10008 6848 10014 6860
rect 10594 6857 10600 6860
rect 10321 6851 10379 6857
rect 10321 6848 10333 6851
rect 10008 6820 10333 6848
rect 10008 6808 10014 6820
rect 10321 6817 10333 6820
rect 10367 6817 10379 6851
rect 10588 6848 10600 6857
rect 10555 6820 10600 6848
rect 10321 6811 10379 6817
rect 10588 6811 10600 6820
rect 10594 6808 10600 6811
rect 10652 6808 10658 6860
rect 16850 6808 16856 6860
rect 16908 6848 16914 6860
rect 16945 6851 17003 6857
rect 16945 6848 16957 6851
rect 16908 6820 16957 6848
rect 16908 6808 16914 6820
rect 16945 6817 16957 6820
rect 16991 6848 17003 6851
rect 17880 6848 17908 6888
rect 18138 6876 18144 6888
rect 18196 6876 18202 6928
rect 24029 6919 24087 6925
rect 24029 6916 24041 6919
rect 23939 6888 24041 6916
rect 24029 6885 24041 6888
rect 24075 6916 24087 6919
rect 24210 6916 24216 6928
rect 24075 6888 24216 6916
rect 24075 6885 24087 6888
rect 24029 6879 24087 6885
rect 16991 6820 17908 6848
rect 17957 6851 18015 6857
rect 16991 6817 17003 6820
rect 16945 6811 17003 6817
rect 17957 6817 17969 6851
rect 18003 6848 18015 6851
rect 18305 6851 18363 6857
rect 18305 6848 18317 6851
rect 18003 6820 18317 6848
rect 18003 6817 18015 6820
rect 17957 6811 18015 6817
rect 18305 6817 18317 6820
rect 18351 6848 18363 6851
rect 20254 6848 20260 6860
rect 18351 6820 20260 6848
rect 18351 6817 18363 6820
rect 18305 6811 18363 6817
rect 20254 6808 20260 6820
rect 20312 6808 20318 6860
rect 20898 6848 20904 6860
rect 20859 6820 20904 6848
rect 20898 6808 20904 6820
rect 20956 6808 20962 6860
rect 21082 6848 21088 6860
rect 21043 6820 21088 6848
rect 21082 6808 21088 6820
rect 21140 6808 21146 6860
rect 23201 6851 23259 6857
rect 23201 6817 23213 6851
rect 23247 6848 23259 6851
rect 24044 6848 24072 6879
rect 24210 6876 24216 6888
rect 24268 6916 24274 6928
rect 24762 6916 24768 6928
rect 24268 6888 24768 6916
rect 24268 6876 24274 6888
rect 24762 6876 24768 6888
rect 24820 6876 24826 6928
rect 27614 6916 27620 6928
rect 27575 6888 27620 6916
rect 27614 6876 27620 6888
rect 27672 6876 27678 6928
rect 28092 6860 28120 6956
rect 29181 6953 29193 6956
rect 29227 6984 29239 6987
rect 29362 6984 29368 6996
rect 29227 6956 29368 6984
rect 29227 6953 29239 6956
rect 29181 6947 29239 6953
rect 29362 6944 29368 6956
rect 29420 6944 29426 6996
rect 23247 6820 24072 6848
rect 24121 6851 24179 6857
rect 23247 6817 23259 6820
rect 23201 6811 23259 6817
rect 24121 6817 24133 6851
rect 24167 6848 24179 6851
rect 24394 6848 24400 6860
rect 24167 6820 24400 6848
rect 24167 6817 24179 6820
rect 24121 6811 24179 6817
rect 4890 6780 4896 6792
rect 4851 6752 4896 6780
rect 4890 6740 4896 6752
rect 4948 6740 4954 6792
rect 8018 6780 8024 6792
rect 7979 6752 8024 6780
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 13541 6783 13599 6789
rect 13541 6749 13553 6783
rect 13587 6780 13599 6783
rect 13630 6780 13636 6792
rect 13587 6752 13636 6780
rect 13587 6749 13599 6752
rect 13541 6743 13599 6749
rect 13630 6740 13636 6752
rect 13688 6780 13694 6792
rect 14093 6783 14151 6789
rect 14093 6780 14105 6783
rect 13688 6752 14105 6780
rect 13688 6740 13694 6752
rect 14093 6749 14105 6752
rect 14139 6749 14151 6783
rect 14093 6743 14151 6749
rect 14182 6740 14188 6792
rect 14240 6780 14246 6792
rect 15194 6780 15200 6792
rect 14240 6752 15200 6780
rect 14240 6740 14246 6752
rect 15194 6740 15200 6752
rect 15252 6780 15258 6792
rect 15473 6783 15531 6789
rect 15473 6780 15485 6783
rect 15252 6752 15485 6780
rect 15252 6740 15258 6752
rect 15473 6749 15485 6752
rect 15519 6749 15531 6783
rect 15473 6743 15531 6749
rect 15933 6783 15991 6789
rect 15933 6749 15945 6783
rect 15979 6780 15991 6783
rect 17402 6780 17408 6792
rect 15979 6752 17408 6780
rect 15979 6749 15991 6752
rect 15933 6743 15991 6749
rect 17402 6740 17408 6752
rect 17460 6740 17466 6792
rect 18046 6780 18052 6792
rect 18007 6752 18052 6780
rect 18046 6740 18052 6752
rect 18104 6740 18110 6792
rect 20714 6740 20720 6792
rect 20772 6780 20778 6792
rect 21269 6783 21327 6789
rect 21269 6780 21281 6783
rect 20772 6752 21281 6780
rect 20772 6740 20778 6752
rect 21269 6749 21281 6752
rect 21315 6749 21327 6783
rect 21269 6743 21327 6749
rect 23569 6783 23627 6789
rect 23569 6749 23581 6783
rect 23615 6780 23627 6783
rect 24136 6780 24164 6811
rect 24394 6808 24400 6820
rect 24452 6808 24458 6860
rect 25130 6808 25136 6860
rect 25188 6848 25194 6860
rect 25317 6851 25375 6857
rect 25317 6848 25329 6851
rect 25188 6820 25329 6848
rect 25188 6808 25194 6820
rect 25317 6817 25329 6820
rect 25363 6848 25375 6851
rect 25406 6848 25412 6860
rect 25363 6820 25412 6848
rect 25363 6817 25375 6820
rect 25317 6811 25375 6817
rect 25406 6808 25412 6820
rect 25464 6808 25470 6860
rect 26605 6851 26663 6857
rect 26605 6817 26617 6851
rect 26651 6848 26663 6851
rect 27246 6848 27252 6860
rect 26651 6820 27252 6848
rect 26651 6817 26663 6820
rect 26605 6811 26663 6817
rect 27246 6808 27252 6820
rect 27304 6808 27310 6860
rect 28074 6808 28080 6860
rect 28132 6848 28138 6860
rect 28810 6848 28816 6860
rect 28132 6820 28177 6848
rect 28771 6820 28816 6848
rect 28132 6808 28138 6820
rect 28810 6808 28816 6820
rect 28868 6808 28874 6860
rect 29270 6848 29276 6860
rect 29231 6820 29276 6848
rect 29270 6808 29276 6820
rect 29328 6808 29334 6860
rect 29540 6851 29598 6857
rect 29540 6817 29552 6851
rect 29586 6848 29598 6851
rect 30374 6848 30380 6860
rect 29586 6820 30380 6848
rect 29586 6817 29598 6820
rect 29540 6811 29598 6817
rect 30374 6808 30380 6820
rect 30432 6808 30438 6860
rect 23615 6752 24164 6780
rect 24305 6783 24363 6789
rect 23615 6749 23627 6752
rect 23569 6743 23627 6749
rect 24305 6749 24317 6783
rect 24351 6749 24363 6783
rect 24305 6743 24363 6749
rect 28169 6783 28227 6789
rect 28169 6749 28181 6783
rect 28215 6749 28227 6783
rect 28169 6743 28227 6749
rect 28261 6783 28319 6789
rect 28261 6749 28273 6783
rect 28307 6780 28319 6783
rect 28442 6780 28448 6792
rect 28307 6752 28448 6780
rect 28307 6749 28319 6752
rect 28261 6743 28319 6749
rect 13906 6672 13912 6724
rect 13964 6712 13970 6724
rect 13964 6684 14688 6712
rect 13964 6672 13970 6684
rect 14660 6656 14688 6684
rect 22094 6672 22100 6724
rect 22152 6712 22158 6724
rect 22833 6715 22891 6721
rect 22833 6712 22845 6715
rect 22152 6684 22845 6712
rect 22152 6672 22158 6684
rect 22833 6681 22845 6684
rect 22879 6712 22891 6715
rect 24320 6712 24348 6743
rect 25866 6712 25872 6724
rect 22879 6684 25872 6712
rect 22879 6681 22891 6684
rect 22833 6675 22891 6681
rect 25866 6672 25872 6684
rect 25924 6712 25930 6724
rect 25961 6715 26019 6721
rect 25961 6712 25973 6715
rect 25924 6684 25973 6712
rect 25924 6672 25930 6684
rect 25961 6681 25973 6684
rect 26007 6712 26019 6715
rect 26329 6715 26387 6721
rect 26329 6712 26341 6715
rect 26007 6684 26341 6712
rect 26007 6681 26019 6684
rect 25961 6675 26019 6681
rect 26329 6681 26341 6684
rect 26375 6712 26387 6715
rect 26694 6712 26700 6724
rect 26375 6684 26700 6712
rect 26375 6681 26387 6684
rect 26329 6675 26387 6681
rect 26694 6672 26700 6684
rect 26752 6672 26758 6724
rect 28184 6712 28212 6743
rect 28442 6740 28448 6752
rect 28500 6740 28506 6792
rect 28350 6712 28356 6724
rect 28184 6684 28356 6712
rect 28350 6672 28356 6684
rect 28408 6712 28414 6724
rect 28828 6712 28856 6808
rect 28408 6684 28856 6712
rect 28408 6672 28414 6684
rect 6270 6644 6276 6656
rect 6231 6616 6276 6644
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 7374 6644 7380 6656
rect 7335 6616 7380 6644
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 8754 6644 8760 6656
rect 8715 6616 8760 6644
rect 8754 6604 8760 6616
rect 8812 6644 8818 6656
rect 10137 6647 10195 6653
rect 10137 6644 10149 6647
rect 8812 6616 10149 6644
rect 8812 6604 8818 6616
rect 10137 6613 10149 6616
rect 10183 6613 10195 6647
rect 10137 6607 10195 6613
rect 13633 6647 13691 6653
rect 13633 6613 13645 6647
rect 13679 6644 13691 6647
rect 14366 6644 14372 6656
rect 13679 6616 14372 6644
rect 13679 6613 13691 6616
rect 13633 6607 13691 6613
rect 14366 6604 14372 6616
rect 14424 6604 14430 6656
rect 14642 6604 14648 6656
rect 14700 6644 14706 6656
rect 14737 6647 14795 6653
rect 14737 6644 14749 6647
rect 14700 6616 14749 6644
rect 14700 6604 14706 6616
rect 14737 6613 14749 6616
rect 14783 6644 14795 6647
rect 14826 6644 14832 6656
rect 14783 6616 14832 6644
rect 14783 6613 14795 6616
rect 14737 6607 14795 6613
rect 14826 6604 14832 6616
rect 14884 6604 14890 6656
rect 17126 6644 17132 6656
rect 17087 6616 17132 6644
rect 17126 6604 17132 6616
rect 17184 6604 17190 6656
rect 17586 6644 17592 6656
rect 17547 6616 17592 6644
rect 17586 6604 17592 6616
rect 17644 6604 17650 6656
rect 19150 6604 19156 6656
rect 19208 6644 19214 6656
rect 19429 6647 19487 6653
rect 19429 6644 19441 6647
rect 19208 6616 19441 6644
rect 19208 6604 19214 6616
rect 19429 6613 19441 6616
rect 19475 6613 19487 6647
rect 23658 6644 23664 6656
rect 23619 6616 23664 6644
rect 19429 6607 19487 6613
rect 23658 6604 23664 6616
rect 23716 6604 23722 6656
rect 24762 6644 24768 6656
rect 24723 6616 24768 6644
rect 24762 6604 24768 6616
rect 24820 6604 24826 6656
rect 25498 6644 25504 6656
rect 25459 6616 25504 6644
rect 25498 6604 25504 6616
rect 25556 6604 25562 6656
rect 26789 6647 26847 6653
rect 26789 6613 26801 6647
rect 26835 6644 26847 6647
rect 27338 6644 27344 6656
rect 26835 6616 27344 6644
rect 26835 6613 26847 6616
rect 26789 6607 26847 6613
rect 27338 6604 27344 6616
rect 27396 6604 27402 6656
rect 27706 6644 27712 6656
rect 27667 6616 27712 6644
rect 27706 6604 27712 6616
rect 27764 6604 27770 6656
rect 30650 6644 30656 6656
rect 30611 6616 30656 6644
rect 30650 6604 30656 6616
rect 30708 6604 30714 6656
rect 1104 6554 38824 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 38824 6554
rect 1104 6480 38824 6502
rect 4890 6440 4896 6452
rect 4851 6412 4896 6440
rect 4890 6400 4896 6412
rect 4948 6400 4954 6452
rect 5353 6443 5411 6449
rect 5353 6409 5365 6443
rect 5399 6440 5411 6443
rect 5442 6440 5448 6452
rect 5399 6412 5448 6440
rect 5399 6409 5411 6412
rect 5353 6403 5411 6409
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 8202 6440 8208 6452
rect 8163 6412 8208 6440
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 9950 6400 9956 6452
rect 10008 6440 10014 6452
rect 10873 6443 10931 6449
rect 10873 6440 10885 6443
rect 10008 6412 10885 6440
rect 10008 6400 10014 6412
rect 10873 6409 10885 6412
rect 10919 6440 10931 6443
rect 11054 6440 11060 6452
rect 10919 6412 11060 6440
rect 10919 6409 10931 6412
rect 10873 6403 10931 6409
rect 11054 6400 11060 6412
rect 11112 6400 11118 6452
rect 13446 6440 13452 6452
rect 13407 6412 13452 6440
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 16850 6440 16856 6452
rect 16811 6412 16856 6440
rect 16850 6400 16856 6412
rect 16908 6400 16914 6452
rect 17402 6440 17408 6452
rect 17363 6412 17408 6440
rect 17402 6400 17408 6412
rect 17460 6400 17466 6452
rect 19150 6440 19156 6452
rect 19111 6412 19156 6440
rect 19150 6400 19156 6412
rect 19208 6400 19214 6452
rect 19426 6440 19432 6452
rect 19387 6412 19432 6440
rect 19426 6400 19432 6412
rect 19484 6400 19490 6452
rect 21082 6400 21088 6452
rect 21140 6440 21146 6452
rect 21729 6443 21787 6449
rect 21729 6440 21741 6443
rect 21140 6412 21741 6440
rect 21140 6400 21146 6412
rect 21729 6409 21741 6412
rect 21775 6409 21787 6443
rect 21729 6403 21787 6409
rect 24762 6400 24768 6452
rect 24820 6440 24826 6452
rect 25041 6443 25099 6449
rect 25041 6440 25053 6443
rect 24820 6412 25053 6440
rect 24820 6400 24826 6412
rect 25041 6409 25053 6412
rect 25087 6409 25099 6443
rect 25041 6403 25099 6409
rect 25406 6400 25412 6452
rect 25464 6440 25470 6452
rect 25593 6443 25651 6449
rect 25593 6440 25605 6443
rect 25464 6412 25605 6440
rect 25464 6400 25470 6412
rect 25593 6409 25605 6412
rect 25639 6409 25651 6443
rect 26142 6440 26148 6452
rect 26103 6412 26148 6440
rect 25593 6403 25651 6409
rect 26142 6400 26148 6412
rect 26200 6400 26206 6452
rect 27617 6443 27675 6449
rect 27617 6409 27629 6443
rect 27663 6440 27675 6443
rect 28074 6440 28080 6452
rect 27663 6412 28080 6440
rect 27663 6409 27675 6412
rect 27617 6403 27675 6409
rect 28074 6400 28080 6412
rect 28132 6400 28138 6452
rect 28350 6440 28356 6452
rect 28311 6412 28356 6440
rect 28350 6400 28356 6412
rect 28408 6400 28414 6452
rect 28721 6443 28779 6449
rect 28721 6409 28733 6443
rect 28767 6440 28779 6443
rect 30374 6440 30380 6452
rect 28767 6412 30380 6440
rect 28767 6409 28779 6412
rect 28721 6403 28779 6409
rect 4908 6372 4936 6400
rect 6178 6372 6184 6384
rect 4908 6344 6184 6372
rect 6178 6332 6184 6344
rect 6236 6372 6242 6384
rect 6549 6375 6607 6381
rect 6549 6372 6561 6375
rect 6236 6344 6561 6372
rect 6236 6332 6242 6344
rect 6549 6341 6561 6344
rect 6595 6372 6607 6375
rect 13081 6375 13139 6381
rect 6595 6344 6868 6372
rect 6595 6341 6607 6344
rect 6549 6335 6607 6341
rect 6840 6313 6868 6344
rect 13081 6341 13093 6375
rect 13127 6372 13139 6375
rect 13538 6372 13544 6384
rect 13127 6344 13544 6372
rect 13127 6341 13139 6344
rect 13081 6335 13139 6341
rect 13538 6332 13544 6344
rect 13596 6332 13602 6384
rect 19613 6375 19671 6381
rect 19613 6372 19625 6375
rect 18524 6344 19625 6372
rect 6825 6307 6883 6313
rect 6825 6273 6837 6307
rect 6871 6273 6883 6307
rect 6825 6267 6883 6273
rect 9769 6307 9827 6313
rect 9769 6273 9781 6307
rect 9815 6304 9827 6307
rect 10318 6304 10324 6316
rect 9815 6276 10324 6304
rect 9815 6273 9827 6276
rect 9769 6267 9827 6273
rect 10318 6264 10324 6276
rect 10376 6264 10382 6316
rect 10502 6304 10508 6316
rect 10463 6276 10508 6304
rect 10502 6264 10508 6276
rect 10560 6264 10566 6316
rect 13556 6304 13584 6332
rect 14366 6304 14372 6316
rect 13556 6276 14044 6304
rect 14327 6276 14372 6304
rect 6914 6196 6920 6248
rect 6972 6236 6978 6248
rect 7092 6239 7150 6245
rect 7092 6236 7104 6239
rect 6972 6208 7104 6236
rect 6972 6196 6978 6208
rect 7092 6205 7104 6208
rect 7138 6236 7150 6239
rect 8478 6236 8484 6248
rect 7138 6208 8484 6236
rect 7138 6205 7150 6208
rect 7092 6199 7150 6205
rect 8478 6196 8484 6208
rect 8536 6196 8542 6248
rect 9950 6196 9956 6248
rect 10008 6236 10014 6248
rect 10229 6239 10287 6245
rect 10229 6236 10241 6239
rect 10008 6208 10241 6236
rect 10008 6196 10014 6208
rect 10229 6205 10241 6208
rect 10275 6236 10287 6239
rect 10686 6236 10692 6248
rect 10275 6208 10692 6236
rect 10275 6205 10287 6208
rect 10229 6199 10287 6205
rect 10686 6196 10692 6208
rect 10744 6196 10750 6248
rect 12437 6239 12495 6245
rect 12437 6205 12449 6239
rect 12483 6205 12495 6239
rect 13906 6236 13912 6248
rect 13867 6208 13912 6236
rect 12437 6199 12495 6205
rect 8018 6128 8024 6180
rect 8076 6168 8082 6180
rect 8849 6171 8907 6177
rect 8849 6168 8861 6171
rect 8076 6140 8861 6168
rect 8076 6128 8082 6140
rect 8849 6137 8861 6140
rect 8895 6168 8907 6171
rect 9401 6171 9459 6177
rect 9401 6168 9413 6171
rect 8895 6140 9413 6168
rect 8895 6137 8907 6140
rect 8849 6131 8907 6137
rect 9401 6137 9413 6140
rect 9447 6168 9459 6171
rect 10502 6168 10508 6180
rect 9447 6140 10508 6168
rect 9447 6137 9459 6140
rect 9401 6131 9459 6137
rect 10502 6128 10508 6140
rect 10560 6128 10566 6180
rect 12452 6168 12480 6199
rect 13906 6196 13912 6208
rect 13964 6196 13970 6248
rect 14016 6236 14044 6276
rect 14366 6264 14372 6276
rect 14424 6264 14430 6316
rect 17862 6264 17868 6316
rect 17920 6304 17926 6316
rect 18524 6313 18552 6344
rect 19613 6341 19625 6344
rect 19659 6341 19671 6375
rect 19613 6335 19671 6341
rect 19978 6332 19984 6384
rect 20036 6372 20042 6384
rect 20036 6344 21220 6372
rect 20036 6332 20042 6344
rect 18509 6307 18567 6313
rect 18509 6304 18521 6307
rect 17920 6276 18521 6304
rect 17920 6264 17926 6276
rect 18509 6273 18521 6276
rect 18555 6273 18567 6307
rect 18690 6304 18696 6316
rect 18603 6276 18696 6304
rect 18509 6267 18567 6273
rect 18690 6264 18696 6276
rect 18748 6304 18754 6316
rect 19150 6304 19156 6316
rect 18748 6276 19156 6304
rect 18748 6264 18754 6276
rect 19150 6264 19156 6276
rect 19208 6264 19214 6316
rect 20070 6304 20076 6316
rect 20031 6276 20076 6304
rect 20070 6264 20076 6276
rect 20128 6264 20134 6316
rect 20254 6304 20260 6316
rect 20215 6276 20260 6304
rect 20254 6264 20260 6276
rect 20312 6264 20318 6316
rect 14645 6239 14703 6245
rect 14645 6236 14657 6239
rect 14016 6208 14657 6236
rect 14645 6205 14657 6208
rect 14691 6205 14703 6239
rect 14645 6199 14703 6205
rect 17402 6196 17408 6248
rect 17460 6236 17466 6248
rect 18417 6239 18475 6245
rect 18417 6236 18429 6239
rect 17460 6208 18429 6236
rect 17460 6196 17466 6208
rect 18417 6205 18429 6208
rect 18463 6205 18475 6239
rect 18417 6199 18475 6205
rect 19426 6196 19432 6248
rect 19484 6236 19490 6248
rect 21192 6245 21220 6344
rect 25314 6332 25320 6384
rect 25372 6372 25378 6384
rect 25961 6375 26019 6381
rect 25961 6372 25973 6375
rect 25372 6344 25973 6372
rect 25372 6332 25378 6344
rect 25961 6341 25973 6344
rect 26007 6372 26019 6375
rect 29089 6375 29147 6381
rect 26007 6344 26648 6372
rect 26007 6341 26019 6344
rect 25961 6335 26019 6341
rect 26620 6313 26648 6344
rect 29089 6341 29101 6375
rect 29135 6372 29147 6375
rect 29270 6372 29276 6384
rect 29135 6344 29276 6372
rect 29135 6341 29147 6344
rect 29089 6335 29147 6341
rect 29270 6332 29276 6344
rect 29328 6332 29334 6384
rect 26605 6307 26663 6313
rect 26605 6273 26617 6307
rect 26651 6273 26663 6307
rect 26605 6267 26663 6273
rect 26694 6264 26700 6316
rect 26752 6304 26758 6316
rect 26789 6307 26847 6313
rect 26789 6304 26801 6307
rect 26752 6276 26801 6304
rect 26752 6264 26758 6276
rect 26789 6273 26801 6276
rect 26835 6304 26847 6307
rect 28442 6304 28448 6316
rect 26835 6276 28448 6304
rect 26835 6273 26847 6276
rect 26789 6267 26847 6273
rect 28442 6264 28448 6276
rect 28500 6264 28506 6316
rect 29748 6313 29776 6412
rect 30374 6400 30380 6412
rect 30432 6400 30438 6452
rect 30650 6440 30656 6452
rect 30611 6412 30656 6440
rect 30650 6400 30656 6412
rect 30708 6400 30714 6452
rect 29733 6307 29791 6313
rect 29733 6273 29745 6307
rect 29779 6273 29791 6307
rect 29914 6304 29920 6316
rect 29827 6276 29920 6304
rect 29733 6267 29791 6273
rect 29914 6264 29920 6276
rect 29972 6304 29978 6316
rect 29972 6276 31156 6304
rect 29972 6264 29978 6276
rect 19981 6239 20039 6245
rect 19981 6236 19993 6239
rect 19484 6208 19993 6236
rect 19484 6196 19490 6208
rect 19981 6205 19993 6208
rect 20027 6205 20039 6239
rect 19981 6199 20039 6205
rect 21177 6239 21235 6245
rect 21177 6205 21189 6239
rect 21223 6236 21235 6239
rect 21358 6236 21364 6248
rect 21223 6208 21364 6236
rect 21223 6205 21235 6208
rect 21177 6199 21235 6205
rect 21358 6196 21364 6208
rect 21416 6196 21422 6248
rect 22373 6239 22431 6245
rect 22373 6205 22385 6239
rect 22419 6236 22431 6239
rect 22465 6239 22523 6245
rect 22465 6236 22477 6239
rect 22419 6208 22477 6236
rect 22419 6205 22431 6208
rect 22373 6199 22431 6205
rect 22465 6205 22477 6208
rect 22511 6236 22523 6239
rect 23290 6236 23296 6248
rect 22511 6208 23296 6236
rect 22511 6205 22523 6208
rect 22465 6199 22523 6205
rect 23290 6196 23296 6208
rect 23348 6196 23354 6248
rect 23566 6196 23572 6248
rect 23624 6236 23630 6248
rect 23661 6239 23719 6245
rect 23661 6236 23673 6239
rect 23624 6208 23673 6236
rect 23624 6196 23630 6208
rect 23661 6205 23673 6208
rect 23707 6205 23719 6239
rect 26510 6236 26516 6248
rect 26471 6208 26516 6236
rect 23661 6199 23719 6205
rect 26510 6196 26516 6208
rect 26568 6196 26574 6248
rect 27709 6239 27767 6245
rect 27709 6205 27721 6239
rect 27755 6236 27767 6239
rect 28350 6236 28356 6248
rect 27755 6208 28356 6236
rect 27755 6205 27767 6208
rect 27709 6199 27767 6205
rect 28350 6196 28356 6208
rect 28408 6196 28414 6248
rect 29638 6236 29644 6248
rect 29551 6208 29644 6236
rect 29638 6196 29644 6208
rect 29696 6236 29702 6248
rect 30650 6236 30656 6248
rect 29696 6208 30656 6236
rect 29696 6196 29702 6208
rect 30650 6196 30656 6208
rect 30708 6196 30714 6248
rect 12176 6140 12480 6168
rect 12176 6109 12204 6140
rect 20898 6128 20904 6180
rect 20956 6168 20962 6180
rect 20993 6171 21051 6177
rect 20993 6168 21005 6171
rect 20956 6140 21005 6168
rect 20956 6128 20962 6140
rect 20993 6137 21005 6140
rect 21039 6168 21051 6171
rect 21634 6168 21640 6180
rect 21039 6140 21640 6168
rect 21039 6137 21051 6140
rect 20993 6131 21051 6137
rect 21634 6128 21640 6140
rect 21692 6128 21698 6180
rect 23109 6171 23167 6177
rect 23109 6137 23121 6171
rect 23155 6168 23167 6171
rect 23928 6171 23986 6177
rect 23928 6168 23940 6171
rect 23155 6140 23940 6168
rect 23155 6137 23167 6140
rect 23109 6131 23167 6137
rect 23928 6137 23940 6140
rect 23974 6168 23986 6171
rect 24394 6168 24400 6180
rect 23974 6140 24400 6168
rect 23974 6137 23986 6140
rect 23928 6131 23986 6137
rect 24394 6128 24400 6140
rect 24452 6128 24458 6180
rect 9861 6103 9919 6109
rect 9861 6069 9873 6103
rect 9907 6100 9919 6103
rect 12161 6103 12219 6109
rect 12161 6100 12173 6103
rect 9907 6072 12173 6100
rect 9907 6069 9919 6072
rect 9861 6063 9919 6069
rect 12161 6069 12173 6072
rect 12207 6069 12219 6103
rect 12618 6100 12624 6112
rect 12579 6072 12624 6100
rect 12161 6063 12219 6069
rect 12618 6060 12624 6072
rect 12676 6060 12682 6112
rect 13814 6100 13820 6112
rect 13727 6072 13820 6100
rect 13814 6060 13820 6072
rect 13872 6100 13878 6112
rect 14371 6103 14429 6109
rect 14371 6100 14383 6103
rect 13872 6072 14383 6100
rect 13872 6060 13878 6072
rect 14371 6069 14383 6072
rect 14417 6100 14429 6103
rect 14642 6100 14648 6112
rect 14417 6072 14648 6100
rect 14417 6069 14429 6072
rect 14371 6063 14429 6069
rect 14642 6060 14648 6072
rect 14700 6060 14706 6112
rect 15562 6060 15568 6112
rect 15620 6100 15626 6112
rect 15749 6103 15807 6109
rect 15749 6100 15761 6103
rect 15620 6072 15761 6100
rect 15620 6060 15626 6072
rect 15749 6069 15761 6072
rect 15795 6069 15807 6103
rect 16942 6100 16948 6112
rect 16903 6072 16948 6100
rect 15749 6063 15807 6069
rect 16942 6060 16948 6072
rect 17000 6060 17006 6112
rect 17865 6103 17923 6109
rect 17865 6069 17877 6103
rect 17911 6100 17923 6103
rect 17954 6100 17960 6112
rect 17911 6072 17960 6100
rect 17911 6069 17923 6072
rect 17865 6063 17923 6069
rect 17954 6060 17960 6072
rect 18012 6060 18018 6112
rect 18049 6103 18107 6109
rect 18049 6069 18061 6103
rect 18095 6100 18107 6103
rect 18506 6100 18512 6112
rect 18095 6072 18512 6100
rect 18095 6069 18107 6072
rect 18049 6063 18107 6069
rect 18506 6060 18512 6072
rect 18564 6060 18570 6112
rect 21361 6103 21419 6109
rect 21361 6069 21373 6103
rect 21407 6100 21419 6103
rect 21450 6100 21456 6112
rect 21407 6072 21456 6100
rect 21407 6069 21419 6072
rect 21361 6063 21419 6069
rect 21450 6060 21456 6072
rect 21508 6060 21514 6112
rect 22646 6100 22652 6112
rect 22607 6072 22652 6100
rect 22646 6060 22652 6072
rect 22704 6060 22710 6112
rect 22922 6060 22928 6112
rect 22980 6100 22986 6112
rect 23385 6103 23443 6109
rect 23385 6100 23397 6103
rect 22980 6072 23397 6100
rect 22980 6060 22986 6072
rect 23385 6069 23397 6072
rect 23431 6100 23443 6103
rect 23566 6100 23572 6112
rect 23431 6072 23572 6100
rect 23431 6069 23443 6072
rect 23385 6063 23443 6069
rect 23566 6060 23572 6072
rect 23624 6060 23630 6112
rect 27246 6100 27252 6112
rect 27207 6072 27252 6100
rect 27246 6060 27252 6072
rect 27304 6060 27310 6112
rect 27522 6060 27528 6112
rect 27580 6100 27586 6112
rect 27893 6103 27951 6109
rect 27893 6100 27905 6103
rect 27580 6072 27905 6100
rect 27580 6060 27586 6072
rect 27893 6069 27905 6072
rect 27939 6069 27951 6103
rect 29270 6100 29276 6112
rect 29231 6072 29276 6100
rect 27893 6063 27951 6069
rect 29270 6060 29276 6072
rect 29328 6060 29334 6112
rect 31128 6109 31156 6276
rect 31113 6103 31171 6109
rect 31113 6069 31125 6103
rect 31159 6100 31171 6103
rect 31386 6100 31392 6112
rect 31159 6072 31392 6100
rect 31159 6069 31171 6072
rect 31113 6063 31171 6069
rect 31386 6060 31392 6072
rect 31444 6060 31450 6112
rect 33318 6100 33324 6112
rect 33279 6072 33324 6100
rect 33318 6060 33324 6072
rect 33376 6060 33382 6112
rect 1104 6010 38824 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 38824 6010
rect 1104 5936 38824 5958
rect 4341 5899 4399 5905
rect 4341 5865 4353 5899
rect 4387 5896 4399 5899
rect 4614 5896 4620 5908
rect 4387 5868 4620 5896
rect 4387 5865 4399 5868
rect 4341 5859 4399 5865
rect 4614 5856 4620 5868
rect 4672 5896 4678 5908
rect 5997 5899 6055 5905
rect 5997 5896 6009 5899
rect 4672 5868 6009 5896
rect 4672 5856 4678 5868
rect 5997 5865 6009 5868
rect 6043 5896 6055 5899
rect 6270 5896 6276 5908
rect 6043 5868 6276 5896
rect 6043 5865 6055 5868
rect 5997 5859 6055 5865
rect 6270 5856 6276 5868
rect 6328 5856 6334 5908
rect 6914 5896 6920 5908
rect 6875 5868 6920 5896
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 7745 5899 7803 5905
rect 7745 5865 7757 5899
rect 7791 5896 7803 5899
rect 7926 5896 7932 5908
rect 7791 5868 7932 5896
rect 7791 5865 7803 5868
rect 7745 5859 7803 5865
rect 7926 5856 7932 5868
rect 7984 5856 7990 5908
rect 9950 5896 9956 5908
rect 9911 5868 9956 5896
rect 9950 5856 9956 5868
rect 10008 5856 10014 5908
rect 10413 5899 10471 5905
rect 10413 5865 10425 5899
rect 10459 5896 10471 5899
rect 10594 5896 10600 5908
rect 10459 5868 10600 5896
rect 10459 5865 10471 5868
rect 10413 5859 10471 5865
rect 10594 5856 10600 5868
rect 10652 5856 10658 5908
rect 11238 5856 11244 5908
rect 11296 5896 11302 5908
rect 11793 5899 11851 5905
rect 11793 5896 11805 5899
rect 11296 5868 11805 5896
rect 11296 5856 11302 5868
rect 11793 5865 11805 5868
rect 11839 5865 11851 5899
rect 13630 5896 13636 5908
rect 13591 5868 13636 5896
rect 11793 5859 11851 5865
rect 13630 5856 13636 5868
rect 13688 5856 13694 5908
rect 14366 5856 14372 5908
rect 14424 5896 14430 5908
rect 14645 5899 14703 5905
rect 14645 5896 14657 5899
rect 14424 5868 14657 5896
rect 14424 5856 14430 5868
rect 14645 5865 14657 5868
rect 14691 5865 14703 5899
rect 14645 5859 14703 5865
rect 15562 5856 15568 5908
rect 15620 5896 15626 5908
rect 15749 5899 15807 5905
rect 15749 5896 15761 5899
rect 15620 5868 15761 5896
rect 15620 5856 15626 5868
rect 15749 5865 15761 5868
rect 15795 5865 15807 5899
rect 17586 5896 17592 5908
rect 15749 5859 15807 5865
rect 16408 5868 17592 5896
rect 5442 5788 5448 5840
rect 5500 5828 5506 5840
rect 6089 5831 6147 5837
rect 6089 5828 6101 5831
rect 5500 5800 6101 5828
rect 5500 5788 5506 5800
rect 6089 5797 6101 5800
rect 6135 5828 6147 5831
rect 6178 5828 6184 5840
rect 6135 5800 6184 5828
rect 6135 5797 6147 5800
rect 6089 5791 6147 5797
rect 6178 5788 6184 5800
rect 6236 5788 6242 5840
rect 13541 5831 13599 5837
rect 13541 5797 13553 5831
rect 13587 5828 13599 5831
rect 14182 5828 14188 5840
rect 13587 5800 14188 5828
rect 13587 5797 13599 5800
rect 13541 5791 13599 5797
rect 14182 5788 14188 5800
rect 14240 5788 14246 5840
rect 7374 5720 7380 5772
rect 7432 5760 7438 5772
rect 8205 5763 8263 5769
rect 8205 5760 8217 5763
rect 7432 5732 8217 5760
rect 7432 5720 7438 5732
rect 8205 5729 8217 5732
rect 8251 5760 8263 5763
rect 8294 5760 8300 5772
rect 8251 5732 8300 5760
rect 8251 5729 8263 5732
rect 8205 5723 8263 5729
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 10505 5763 10563 5769
rect 10505 5729 10517 5763
rect 10551 5760 10563 5763
rect 10594 5760 10600 5772
rect 10551 5732 10600 5760
rect 10551 5729 10563 5732
rect 10505 5723 10563 5729
rect 10594 5720 10600 5732
rect 10652 5720 10658 5772
rect 11609 5763 11667 5769
rect 11609 5729 11621 5763
rect 11655 5760 11667 5763
rect 11698 5760 11704 5772
rect 11655 5732 11704 5760
rect 11655 5729 11667 5732
rect 11609 5723 11667 5729
rect 11698 5720 11704 5732
rect 11756 5720 11762 5772
rect 13630 5720 13636 5772
rect 13688 5760 13694 5772
rect 14001 5763 14059 5769
rect 14001 5760 14013 5763
rect 13688 5732 14013 5760
rect 13688 5720 13694 5732
rect 14001 5729 14013 5732
rect 14047 5729 14059 5763
rect 15657 5763 15715 5769
rect 15657 5760 15669 5763
rect 14001 5723 14059 5729
rect 14108 5732 15669 5760
rect 14108 5704 14136 5732
rect 15657 5729 15669 5732
rect 15703 5760 15715 5763
rect 16206 5760 16212 5772
rect 15703 5732 16212 5760
rect 15703 5729 15715 5732
rect 15657 5723 15715 5729
rect 16206 5720 16212 5732
rect 16264 5720 16270 5772
rect 16408 5760 16436 5868
rect 17586 5856 17592 5868
rect 17644 5856 17650 5908
rect 17862 5896 17868 5908
rect 17823 5868 17868 5896
rect 17862 5856 17868 5868
rect 17920 5856 17926 5908
rect 19981 5899 20039 5905
rect 19981 5865 19993 5899
rect 20027 5896 20039 5899
rect 20070 5896 20076 5908
rect 20027 5868 20076 5896
rect 20027 5865 20039 5868
rect 19981 5859 20039 5865
rect 20070 5856 20076 5868
rect 20128 5856 20134 5908
rect 20254 5896 20260 5908
rect 20215 5868 20260 5896
rect 20254 5856 20260 5868
rect 20312 5856 20318 5908
rect 21358 5896 21364 5908
rect 21319 5868 21364 5896
rect 21358 5856 21364 5868
rect 21416 5856 21422 5908
rect 21821 5899 21879 5905
rect 21821 5865 21833 5899
rect 21867 5896 21879 5899
rect 22094 5896 22100 5908
rect 21867 5868 22100 5896
rect 21867 5865 21879 5868
rect 21821 5859 21879 5865
rect 22094 5856 22100 5868
rect 22152 5856 22158 5908
rect 24394 5896 24400 5908
rect 24355 5868 24400 5896
rect 24394 5856 24400 5868
rect 24452 5856 24458 5908
rect 26237 5899 26295 5905
rect 26237 5865 26249 5899
rect 26283 5896 26295 5899
rect 26510 5896 26516 5908
rect 26283 5868 26516 5896
rect 26283 5865 26295 5868
rect 26237 5859 26295 5865
rect 26510 5856 26516 5868
rect 26568 5856 26574 5908
rect 27249 5899 27307 5905
rect 27249 5865 27261 5899
rect 27295 5896 27307 5899
rect 27706 5896 27712 5908
rect 27295 5868 27712 5896
rect 27295 5865 27307 5868
rect 27249 5859 27307 5865
rect 27706 5856 27712 5868
rect 27764 5896 27770 5908
rect 27801 5899 27859 5905
rect 27801 5896 27813 5899
rect 27764 5868 27813 5896
rect 27764 5856 27770 5868
rect 27801 5865 27813 5868
rect 27847 5865 27859 5899
rect 28350 5896 28356 5908
rect 28311 5868 28356 5896
rect 27801 5859 27859 5865
rect 28350 5856 28356 5868
rect 28408 5856 28414 5908
rect 28442 5856 28448 5908
rect 28500 5896 28506 5908
rect 28813 5899 28871 5905
rect 28813 5896 28825 5899
rect 28500 5868 28825 5896
rect 28500 5856 28506 5868
rect 28813 5865 28825 5868
rect 28859 5896 28871 5899
rect 29914 5896 29920 5908
rect 28859 5868 29920 5896
rect 28859 5865 28871 5868
rect 28813 5859 28871 5865
rect 29914 5856 29920 5868
rect 29972 5856 29978 5908
rect 18224 5831 18282 5837
rect 18224 5797 18236 5831
rect 18270 5828 18282 5831
rect 18690 5828 18696 5840
rect 18270 5800 18696 5828
rect 18270 5797 18282 5800
rect 18224 5791 18282 5797
rect 18690 5788 18696 5800
rect 18748 5788 18754 5840
rect 23014 5788 23020 5840
rect 23072 5828 23078 5840
rect 23262 5831 23320 5837
rect 23262 5828 23274 5831
rect 23072 5800 23274 5828
rect 23072 5788 23078 5800
rect 23262 5797 23274 5800
rect 23308 5797 23320 5831
rect 23262 5791 23320 5797
rect 29448 5831 29506 5837
rect 29448 5797 29460 5831
rect 29494 5828 29506 5831
rect 29638 5828 29644 5840
rect 29494 5800 29644 5828
rect 29494 5797 29506 5800
rect 29448 5791 29506 5797
rect 29638 5788 29644 5800
rect 29696 5788 29702 5840
rect 16316 5732 16436 5760
rect 17957 5763 18015 5769
rect 5810 5652 5816 5704
rect 5868 5692 5874 5704
rect 6181 5695 6239 5701
rect 6181 5692 6193 5695
rect 5868 5664 6193 5692
rect 5868 5652 5874 5664
rect 6181 5661 6193 5664
rect 6227 5661 6239 5695
rect 7190 5692 7196 5704
rect 7151 5664 7196 5692
rect 6181 5655 6239 5661
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 7742 5652 7748 5704
rect 7800 5692 7806 5704
rect 8021 5695 8079 5701
rect 8021 5692 8033 5695
rect 7800 5664 8033 5692
rect 7800 5652 7806 5664
rect 8021 5661 8033 5664
rect 8067 5661 8079 5695
rect 14090 5692 14096 5704
rect 14051 5664 14096 5692
rect 8021 5655 8079 5661
rect 14090 5652 14096 5664
rect 14148 5652 14154 5704
rect 14277 5695 14335 5701
rect 14277 5661 14289 5695
rect 14323 5692 14335 5695
rect 15102 5692 15108 5704
rect 14323 5664 15108 5692
rect 14323 5661 14335 5664
rect 14277 5655 14335 5661
rect 9030 5584 9036 5636
rect 9088 5624 9094 5636
rect 9493 5627 9551 5633
rect 9493 5624 9505 5627
rect 9088 5596 9505 5624
rect 9088 5584 9094 5596
rect 9493 5593 9505 5596
rect 9539 5624 9551 5627
rect 12805 5627 12863 5633
rect 9539 5596 10732 5624
rect 9539 5593 9551 5596
rect 9493 5587 9551 5593
rect 10704 5568 10732 5596
rect 12805 5593 12817 5627
rect 12851 5624 12863 5627
rect 13354 5624 13360 5636
rect 12851 5596 13360 5624
rect 12851 5593 12863 5596
rect 12805 5587 12863 5593
rect 13354 5584 13360 5596
rect 13412 5624 13418 5636
rect 14292 5624 14320 5655
rect 15102 5652 15108 5664
rect 15160 5652 15166 5704
rect 15838 5692 15844 5704
rect 15799 5664 15844 5692
rect 15838 5652 15844 5664
rect 15896 5652 15902 5704
rect 13412 5596 14320 5624
rect 13412 5584 13418 5596
rect 14826 5584 14832 5636
rect 14884 5624 14890 5636
rect 16316 5633 16344 5732
rect 17957 5729 17969 5763
rect 18003 5760 18015 5763
rect 18046 5760 18052 5772
rect 18003 5732 18052 5760
rect 18003 5729 18015 5732
rect 17957 5723 18015 5729
rect 18046 5720 18052 5732
rect 18104 5720 18110 5772
rect 21910 5760 21916 5772
rect 21871 5732 21916 5760
rect 21910 5720 21916 5732
rect 21968 5720 21974 5772
rect 26881 5763 26939 5769
rect 26881 5729 26893 5763
rect 26927 5760 26939 5763
rect 27709 5763 27767 5769
rect 27709 5760 27721 5763
rect 26927 5732 27721 5760
rect 26927 5729 26939 5732
rect 26881 5723 26939 5729
rect 27709 5729 27721 5732
rect 27755 5760 27767 5763
rect 29270 5760 29276 5772
rect 27755 5732 29276 5760
rect 27755 5729 27767 5732
rect 27709 5723 27767 5729
rect 29270 5720 29276 5732
rect 29328 5720 29334 5772
rect 34330 5760 34336 5772
rect 34291 5732 34336 5760
rect 34330 5720 34336 5732
rect 34388 5720 34394 5772
rect 16945 5695 17003 5701
rect 16945 5661 16957 5695
rect 16991 5692 17003 5695
rect 17862 5692 17868 5704
rect 16991 5664 17868 5692
rect 16991 5661 17003 5664
rect 16945 5655 17003 5661
rect 17862 5652 17868 5664
rect 17920 5652 17926 5704
rect 20898 5692 20904 5704
rect 20859 5664 20904 5692
rect 20898 5652 20904 5664
rect 20956 5652 20962 5704
rect 22922 5652 22928 5704
rect 22980 5692 22986 5704
rect 23017 5695 23075 5701
rect 23017 5692 23029 5695
rect 22980 5664 23029 5692
rect 22980 5652 22986 5664
rect 23017 5661 23029 5664
rect 23063 5661 23075 5695
rect 23017 5655 23075 5661
rect 26786 5652 26792 5704
rect 26844 5692 26850 5704
rect 27893 5695 27951 5701
rect 27893 5692 27905 5695
rect 26844 5664 27905 5692
rect 26844 5652 26850 5664
rect 27893 5661 27905 5664
rect 27939 5661 27951 5695
rect 29178 5692 29184 5704
rect 29139 5664 29184 5692
rect 27893 5655 27951 5661
rect 29178 5652 29184 5664
rect 29236 5652 29242 5704
rect 32674 5692 32680 5704
rect 32635 5664 32680 5692
rect 32674 5652 32680 5664
rect 32732 5652 32738 5704
rect 33962 5652 33968 5704
rect 34020 5692 34026 5704
rect 34425 5695 34483 5701
rect 34425 5692 34437 5695
rect 34020 5664 34437 5692
rect 34020 5652 34026 5664
rect 34425 5661 34437 5664
rect 34471 5661 34483 5695
rect 34425 5655 34483 5661
rect 34517 5695 34575 5701
rect 34517 5661 34529 5695
rect 34563 5661 34575 5695
rect 34517 5655 34575 5661
rect 16301 5627 16359 5633
rect 16301 5624 16313 5627
rect 14884 5596 16313 5624
rect 14884 5584 14890 5596
rect 16301 5593 16313 5596
rect 16347 5593 16359 5627
rect 16301 5587 16359 5593
rect 16853 5627 16911 5633
rect 16853 5593 16865 5627
rect 16899 5624 16911 5627
rect 27341 5627 27399 5633
rect 16899 5596 17908 5624
rect 16899 5593 16911 5596
rect 16853 5587 16911 5593
rect 5626 5556 5632 5568
rect 5587 5528 5632 5556
rect 5626 5516 5632 5528
rect 5684 5516 5690 5568
rect 8389 5559 8447 5565
rect 8389 5525 8401 5559
rect 8435 5556 8447 5559
rect 9306 5556 9312 5568
rect 8435 5528 9312 5556
rect 8435 5525 8447 5528
rect 8389 5519 8447 5525
rect 9306 5516 9312 5528
rect 9364 5516 9370 5568
rect 10686 5556 10692 5568
rect 10647 5528 10692 5556
rect 10686 5516 10692 5528
rect 10744 5516 10750 5568
rect 10962 5516 10968 5568
rect 11020 5556 11026 5568
rect 11057 5559 11115 5565
rect 11057 5556 11069 5559
rect 11020 5528 11069 5556
rect 11020 5516 11026 5528
rect 11057 5525 11069 5528
rect 11103 5525 11115 5559
rect 11057 5519 11115 5525
rect 13173 5559 13231 5565
rect 13173 5525 13185 5559
rect 13219 5556 13231 5559
rect 13814 5556 13820 5568
rect 13219 5528 13820 5556
rect 13219 5525 13231 5528
rect 13173 5519 13231 5525
rect 13814 5516 13820 5528
rect 13872 5516 13878 5568
rect 15010 5556 15016 5568
rect 14971 5528 15016 5556
rect 15010 5516 15016 5528
rect 15068 5516 15074 5568
rect 15102 5516 15108 5568
rect 15160 5556 15166 5568
rect 15289 5559 15347 5565
rect 15289 5556 15301 5559
rect 15160 5528 15301 5556
rect 15160 5516 15166 5528
rect 15289 5525 15301 5528
rect 15335 5525 15347 5559
rect 15289 5519 15347 5525
rect 17497 5559 17555 5565
rect 17497 5525 17509 5559
rect 17543 5556 17555 5559
rect 17678 5556 17684 5568
rect 17543 5528 17684 5556
rect 17543 5525 17555 5528
rect 17497 5519 17555 5525
rect 17678 5516 17684 5528
rect 17736 5516 17742 5568
rect 17880 5556 17908 5596
rect 27341 5593 27353 5627
rect 27387 5624 27399 5627
rect 28350 5624 28356 5636
rect 27387 5596 28356 5624
rect 27387 5593 27399 5596
rect 27341 5587 27399 5593
rect 28350 5584 28356 5596
rect 28408 5584 28414 5636
rect 31938 5624 31944 5636
rect 31851 5596 31944 5624
rect 31938 5584 31944 5596
rect 31996 5624 32002 5636
rect 32490 5624 32496 5636
rect 31996 5596 32496 5624
rect 31996 5584 32002 5596
rect 32490 5584 32496 5596
rect 32548 5584 32554 5636
rect 34238 5584 34244 5636
rect 34296 5624 34302 5636
rect 34532 5624 34560 5655
rect 34296 5596 34560 5624
rect 34296 5584 34302 5596
rect 17954 5556 17960 5568
rect 17880 5528 17960 5556
rect 17954 5516 17960 5528
rect 18012 5516 18018 5568
rect 19334 5556 19340 5568
rect 19295 5528 19340 5556
rect 19334 5516 19340 5528
rect 19392 5516 19398 5568
rect 22462 5556 22468 5568
rect 22423 5528 22468 5556
rect 22462 5516 22468 5528
rect 22520 5516 22526 5568
rect 22925 5559 22983 5565
rect 22925 5525 22937 5559
rect 22971 5556 22983 5559
rect 23014 5556 23020 5568
rect 22971 5528 23020 5556
rect 22971 5525 22983 5528
rect 22925 5519 22983 5525
rect 23014 5516 23020 5528
rect 23072 5516 23078 5568
rect 24946 5556 24952 5568
rect 24907 5528 24952 5556
rect 24946 5516 24952 5528
rect 25004 5516 25010 5568
rect 30558 5556 30564 5568
rect 30519 5528 30564 5556
rect 30558 5516 30564 5528
rect 30616 5516 30622 5568
rect 31202 5556 31208 5568
rect 31163 5528 31208 5556
rect 31202 5516 31208 5528
rect 31260 5516 31266 5568
rect 32306 5556 32312 5568
rect 32267 5528 32312 5556
rect 32306 5516 32312 5528
rect 32364 5516 32370 5568
rect 33134 5556 33140 5568
rect 33095 5528 33140 5556
rect 33134 5516 33140 5528
rect 33192 5516 33198 5568
rect 33965 5559 34023 5565
rect 33965 5525 33977 5559
rect 34011 5556 34023 5559
rect 34514 5556 34520 5568
rect 34011 5528 34520 5556
rect 34011 5525 34023 5528
rect 33965 5519 34023 5525
rect 34514 5516 34520 5528
rect 34572 5516 34578 5568
rect 1104 5466 38824 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 38824 5466
rect 1104 5392 38824 5414
rect 4157 5355 4215 5361
rect 4157 5321 4169 5355
rect 4203 5352 4215 5355
rect 4890 5352 4896 5364
rect 4203 5324 4896 5352
rect 4203 5321 4215 5324
rect 4157 5315 4215 5321
rect 4062 5176 4068 5228
rect 4120 5216 4126 5228
rect 4264 5225 4292 5324
rect 4890 5312 4896 5324
rect 4948 5312 4954 5364
rect 6178 5352 6184 5364
rect 6139 5324 6184 5352
rect 6178 5312 6184 5324
rect 6236 5312 6242 5364
rect 7837 5355 7895 5361
rect 7837 5321 7849 5355
rect 7883 5352 7895 5355
rect 8018 5352 8024 5364
rect 7883 5324 8024 5352
rect 7883 5321 7895 5324
rect 7837 5315 7895 5321
rect 8018 5312 8024 5324
rect 8076 5312 8082 5364
rect 8294 5312 8300 5364
rect 8352 5352 8358 5364
rect 8849 5355 8907 5361
rect 8849 5352 8861 5355
rect 8352 5324 8861 5352
rect 8352 5312 8358 5324
rect 8849 5321 8861 5324
rect 8895 5321 8907 5355
rect 10594 5352 10600 5364
rect 10555 5324 10600 5352
rect 8849 5315 8907 5321
rect 10594 5312 10600 5324
rect 10652 5312 10658 5364
rect 12434 5312 12440 5364
rect 12492 5352 12498 5364
rect 12621 5355 12679 5361
rect 12621 5352 12633 5355
rect 12492 5324 12633 5352
rect 12492 5312 12498 5324
rect 12621 5321 12633 5324
rect 12667 5321 12679 5355
rect 12621 5315 12679 5321
rect 13449 5355 13507 5361
rect 13449 5321 13461 5355
rect 13495 5352 13507 5355
rect 13538 5352 13544 5364
rect 13495 5324 13544 5352
rect 13495 5321 13507 5324
rect 13449 5315 13507 5321
rect 13538 5312 13544 5324
rect 13596 5312 13602 5364
rect 15194 5312 15200 5364
rect 15252 5352 15258 5364
rect 15289 5355 15347 5361
rect 15289 5352 15301 5355
rect 15252 5324 15301 5352
rect 15252 5312 15258 5324
rect 15289 5321 15301 5324
rect 15335 5321 15347 5355
rect 16206 5352 16212 5364
rect 16167 5324 16212 5352
rect 15289 5315 15347 5321
rect 16206 5312 16212 5324
rect 16264 5312 16270 5364
rect 17954 5312 17960 5364
rect 18012 5352 18018 5364
rect 18049 5355 18107 5361
rect 18049 5352 18061 5355
rect 18012 5324 18061 5352
rect 18012 5312 18018 5324
rect 18049 5321 18061 5324
rect 18095 5321 18107 5355
rect 18049 5315 18107 5321
rect 18690 5312 18696 5364
rect 18748 5352 18754 5364
rect 19061 5355 19119 5361
rect 19061 5352 19073 5355
rect 18748 5324 19073 5352
rect 18748 5312 18754 5324
rect 19061 5321 19073 5324
rect 19107 5321 19119 5355
rect 19061 5315 19119 5321
rect 19334 5312 19340 5364
rect 19392 5352 19398 5364
rect 19429 5355 19487 5361
rect 19429 5352 19441 5355
rect 19392 5324 19441 5352
rect 19392 5312 19398 5324
rect 19429 5321 19441 5324
rect 19475 5321 19487 5355
rect 19429 5315 19487 5321
rect 19797 5355 19855 5361
rect 19797 5321 19809 5355
rect 19843 5352 19855 5355
rect 20162 5352 20168 5364
rect 19843 5324 20168 5352
rect 19843 5321 19855 5324
rect 19797 5315 19855 5321
rect 20162 5312 20168 5324
rect 20220 5312 20226 5364
rect 20622 5352 20628 5364
rect 20583 5324 20628 5352
rect 20622 5312 20628 5324
rect 20680 5312 20686 5364
rect 20806 5312 20812 5364
rect 20864 5352 20870 5364
rect 20901 5355 20959 5361
rect 20901 5352 20913 5355
rect 20864 5324 20913 5352
rect 20864 5312 20870 5324
rect 20901 5321 20913 5324
rect 20947 5321 20959 5355
rect 20901 5315 20959 5321
rect 20990 5312 20996 5364
rect 21048 5352 21054 5364
rect 22922 5352 22928 5364
rect 21048 5324 22928 5352
rect 21048 5312 21054 5324
rect 22922 5312 22928 5324
rect 22980 5352 22986 5364
rect 23017 5355 23075 5361
rect 23017 5352 23029 5355
rect 22980 5324 23029 5352
rect 22980 5312 22986 5324
rect 23017 5321 23029 5324
rect 23063 5352 23075 5355
rect 23385 5355 23443 5361
rect 23385 5352 23397 5355
rect 23063 5324 23397 5352
rect 23063 5321 23075 5324
rect 23017 5315 23075 5321
rect 23385 5321 23397 5324
rect 23431 5321 23443 5355
rect 25590 5352 25596 5364
rect 25551 5324 25596 5352
rect 23385 5315 23443 5321
rect 22094 5244 22100 5296
rect 22152 5284 22158 5296
rect 22152 5256 22600 5284
rect 22152 5244 22158 5256
rect 4249 5219 4307 5225
rect 4249 5216 4261 5219
rect 4120 5188 4261 5216
rect 4120 5176 4126 5188
rect 4249 5185 4261 5188
rect 4295 5185 4307 5219
rect 4249 5179 4307 5185
rect 9309 5219 9367 5225
rect 9309 5185 9321 5219
rect 9355 5216 9367 5219
rect 9858 5216 9864 5228
rect 9355 5188 9864 5216
rect 9355 5185 9367 5188
rect 9309 5179 9367 5185
rect 9858 5176 9864 5188
rect 9916 5176 9922 5228
rect 10045 5219 10103 5225
rect 10045 5185 10057 5219
rect 10091 5216 10103 5219
rect 10686 5216 10692 5228
rect 10091 5188 10692 5216
rect 10091 5185 10103 5188
rect 10045 5179 10103 5185
rect 10686 5176 10692 5188
rect 10744 5176 10750 5228
rect 13814 5176 13820 5228
rect 13872 5216 13878 5228
rect 13872 5188 14044 5216
rect 13872 5176 13878 5188
rect 6825 5151 6883 5157
rect 6825 5117 6837 5151
rect 6871 5117 6883 5151
rect 7926 5148 7932 5160
rect 7887 5120 7932 5148
rect 6825 5111 6883 5117
rect 4516 5083 4574 5089
rect 4516 5049 4528 5083
rect 4562 5080 4574 5083
rect 4614 5080 4620 5092
rect 4562 5052 4620 5080
rect 4562 5049 4574 5052
rect 4516 5043 4574 5049
rect 4614 5040 4620 5052
rect 4672 5040 4678 5092
rect 6840 5080 6868 5111
rect 7926 5108 7932 5120
rect 7984 5148 7990 5160
rect 8481 5151 8539 5157
rect 8481 5148 8493 5151
rect 7984 5120 8493 5148
rect 7984 5108 7990 5120
rect 8481 5117 8493 5120
rect 8527 5117 8539 5151
rect 10962 5148 10968 5160
rect 10923 5120 10968 5148
rect 8481 5111 8539 5117
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5148 12495 5151
rect 13078 5148 13084 5160
rect 12483 5120 13084 5148
rect 12483 5117 12495 5120
rect 12437 5111 12495 5117
rect 13078 5108 13084 5120
rect 13136 5108 13142 5160
rect 13909 5151 13967 5157
rect 13909 5117 13921 5151
rect 13955 5117 13967 5151
rect 14016 5148 14044 5188
rect 17678 5176 17684 5228
rect 17736 5216 17742 5228
rect 18693 5219 18751 5225
rect 18693 5216 18705 5219
rect 17736 5188 18705 5216
rect 17736 5176 17742 5188
rect 18693 5185 18705 5188
rect 18739 5216 18751 5219
rect 18874 5216 18880 5228
rect 18739 5188 18880 5216
rect 18739 5185 18751 5188
rect 18693 5179 18751 5185
rect 18874 5176 18880 5188
rect 18932 5176 18938 5228
rect 22462 5216 22468 5228
rect 22423 5188 22468 5216
rect 22462 5176 22468 5188
rect 22520 5176 22526 5228
rect 22572 5225 22600 5256
rect 22557 5219 22615 5225
rect 22557 5185 22569 5219
rect 22603 5185 22615 5219
rect 23400 5216 23428 5315
rect 25590 5312 25596 5324
rect 25648 5352 25654 5364
rect 25961 5355 26019 5361
rect 25961 5352 25973 5355
rect 25648 5324 25973 5352
rect 25648 5312 25654 5324
rect 25961 5321 25973 5324
rect 26007 5352 26019 5355
rect 26234 5352 26240 5364
rect 26007 5324 26240 5352
rect 26007 5321 26019 5324
rect 25961 5315 26019 5321
rect 26234 5312 26240 5324
rect 26292 5352 26298 5364
rect 26786 5352 26792 5364
rect 26292 5324 26792 5352
rect 26292 5312 26298 5324
rect 26786 5312 26792 5324
rect 26844 5312 26850 5364
rect 29089 5355 29147 5361
rect 29089 5321 29101 5355
rect 29135 5352 29147 5355
rect 29178 5352 29184 5364
rect 29135 5324 29184 5352
rect 29135 5321 29147 5324
rect 29089 5315 29147 5321
rect 29178 5312 29184 5324
rect 29236 5312 29242 5364
rect 30377 5355 30435 5361
rect 30377 5321 30389 5355
rect 30423 5352 30435 5355
rect 30650 5352 30656 5364
rect 30423 5324 30656 5352
rect 30423 5321 30435 5324
rect 30377 5315 30435 5321
rect 30650 5312 30656 5324
rect 30708 5312 30714 5364
rect 32493 5355 32551 5361
rect 32493 5321 32505 5355
rect 32539 5352 32551 5355
rect 32674 5352 32680 5364
rect 32539 5324 32680 5352
rect 32539 5321 32551 5324
rect 32493 5315 32551 5321
rect 32674 5312 32680 5324
rect 32732 5312 32738 5364
rect 33962 5352 33968 5364
rect 33923 5324 33968 5352
rect 33962 5312 33968 5324
rect 34020 5312 34026 5364
rect 34330 5352 34336 5364
rect 34291 5324 34336 5352
rect 34330 5312 34336 5324
rect 34388 5312 34394 5364
rect 33226 5244 33232 5296
rect 33284 5284 33290 5296
rect 34348 5284 34376 5312
rect 33284 5256 34376 5284
rect 33284 5244 33290 5256
rect 23661 5219 23719 5225
rect 23661 5216 23673 5219
rect 23400 5188 23673 5216
rect 22557 5179 22615 5185
rect 23661 5185 23673 5188
rect 23707 5185 23719 5219
rect 28258 5216 28264 5228
rect 28219 5188 28264 5216
rect 23661 5179 23719 5185
rect 14165 5151 14223 5157
rect 14165 5148 14177 5151
rect 14016 5120 14177 5148
rect 13909 5111 13967 5117
rect 14165 5117 14177 5120
rect 14211 5117 14223 5151
rect 16390 5148 16396 5160
rect 16303 5120 16396 5148
rect 14165 5111 14223 5117
rect 7466 5080 7472 5092
rect 6840 5052 7472 5080
rect 7466 5040 7472 5052
rect 7524 5040 7530 5092
rect 9306 5040 9312 5092
rect 9364 5080 9370 5092
rect 9769 5083 9827 5089
rect 9769 5080 9781 5083
rect 9364 5052 9781 5080
rect 9364 5040 9370 5052
rect 9769 5049 9781 5052
rect 9815 5049 9827 5083
rect 9769 5043 9827 5049
rect 11054 5040 11060 5092
rect 11112 5080 11118 5092
rect 13725 5083 13783 5089
rect 13725 5080 13737 5083
rect 11112 5052 13737 5080
rect 11112 5040 11118 5052
rect 13725 5049 13737 5052
rect 13771 5080 13783 5083
rect 13924 5080 13952 5111
rect 16390 5108 16396 5120
rect 16448 5148 16454 5160
rect 16945 5151 17003 5157
rect 16945 5148 16957 5151
rect 16448 5120 16957 5148
rect 16448 5108 16454 5120
rect 16945 5117 16957 5120
rect 16991 5117 17003 5151
rect 16945 5111 17003 5117
rect 19613 5151 19671 5157
rect 19613 5117 19625 5151
rect 19659 5148 19671 5151
rect 20257 5151 20315 5157
rect 20257 5148 20269 5151
rect 19659 5120 20269 5148
rect 19659 5117 19671 5120
rect 19613 5111 19671 5117
rect 20257 5117 20269 5120
rect 20303 5148 20315 5151
rect 20530 5148 20536 5160
rect 20303 5120 20536 5148
rect 20303 5117 20315 5120
rect 20257 5111 20315 5117
rect 20530 5108 20536 5120
rect 20588 5108 20594 5160
rect 20714 5148 20720 5160
rect 20675 5120 20720 5148
rect 20714 5108 20720 5120
rect 20772 5148 20778 5160
rect 21269 5151 21327 5157
rect 21269 5148 21281 5151
rect 20772 5120 21281 5148
rect 20772 5108 20778 5120
rect 21269 5117 21281 5120
rect 21315 5117 21327 5151
rect 21269 5111 21327 5117
rect 22373 5151 22431 5157
rect 22373 5117 22385 5151
rect 22419 5148 22431 5151
rect 23014 5148 23020 5160
rect 22419 5120 23020 5148
rect 22419 5117 22431 5120
rect 22373 5111 22431 5117
rect 23014 5108 23020 5120
rect 23072 5108 23078 5160
rect 23676 5148 23704 5179
rect 28258 5176 28264 5188
rect 28316 5176 28322 5228
rect 29914 5216 29920 5228
rect 29875 5188 29920 5216
rect 29914 5176 29920 5188
rect 29972 5176 29978 5228
rect 31386 5216 31392 5228
rect 31347 5188 31392 5216
rect 31386 5176 31392 5188
rect 31444 5176 31450 5228
rect 32125 5219 32183 5225
rect 32125 5185 32137 5219
rect 32171 5216 32183 5219
rect 33042 5216 33048 5228
rect 32171 5188 33048 5216
rect 32171 5185 32183 5188
rect 32125 5179 32183 5185
rect 33042 5176 33048 5188
rect 33100 5216 33106 5228
rect 33137 5219 33195 5225
rect 33137 5216 33149 5219
rect 33100 5188 33149 5216
rect 33100 5176 33106 5188
rect 33137 5185 33149 5188
rect 33183 5185 33195 5219
rect 33137 5179 33195 5185
rect 24762 5148 24768 5160
rect 23676 5120 24768 5148
rect 24762 5108 24768 5120
rect 24820 5108 24826 5160
rect 24854 5108 24860 5160
rect 24912 5148 24918 5160
rect 26145 5151 26203 5157
rect 26145 5148 26157 5151
rect 24912 5120 26157 5148
rect 24912 5108 24918 5120
rect 26145 5117 26157 5120
rect 26191 5148 26203 5151
rect 26697 5151 26755 5157
rect 26697 5148 26709 5151
rect 26191 5120 26709 5148
rect 26191 5117 26203 5120
rect 26145 5111 26203 5117
rect 26697 5117 26709 5120
rect 26743 5117 26755 5151
rect 27154 5148 27160 5160
rect 27067 5120 27160 5148
rect 26697 5111 26755 5117
rect 27154 5108 27160 5120
rect 27212 5148 27218 5160
rect 27982 5148 27988 5160
rect 27212 5120 27988 5148
rect 27212 5108 27218 5120
rect 27982 5108 27988 5120
rect 28040 5108 28046 5160
rect 32674 5108 32680 5160
rect 32732 5148 32738 5160
rect 32953 5151 33011 5157
rect 32953 5148 32965 5151
rect 32732 5120 32965 5148
rect 32732 5108 32738 5120
rect 32953 5117 32965 5120
rect 32999 5117 33011 5151
rect 32953 5111 33011 5117
rect 13998 5080 14004 5092
rect 13771 5052 14004 5080
rect 13771 5049 13783 5052
rect 13725 5043 13783 5049
rect 13998 5040 14004 5052
rect 14056 5040 14062 5092
rect 17865 5083 17923 5089
rect 17865 5049 17877 5083
rect 17911 5080 17923 5083
rect 18046 5080 18052 5092
rect 17911 5052 18052 5080
rect 17911 5049 17923 5052
rect 17865 5043 17923 5049
rect 18046 5040 18052 5052
rect 18104 5040 18110 5092
rect 21910 5080 21916 5092
rect 21823 5052 21916 5080
rect 21910 5040 21916 5052
rect 21968 5080 21974 5092
rect 22738 5080 22744 5092
rect 21968 5052 22744 5080
rect 21968 5040 21974 5052
rect 22738 5040 22744 5052
rect 22796 5040 22802 5092
rect 23934 5089 23940 5092
rect 23928 5080 23940 5089
rect 23895 5052 23940 5080
rect 23928 5043 23940 5052
rect 23934 5040 23940 5043
rect 23992 5040 23998 5092
rect 28077 5083 28135 5089
rect 28077 5080 28089 5083
rect 27448 5052 28089 5080
rect 27448 5024 27476 5052
rect 28077 5049 28089 5052
rect 28123 5049 28135 5083
rect 28077 5043 28135 5049
rect 28721 5083 28779 5089
rect 28721 5049 28733 5083
rect 28767 5080 28779 5083
rect 29454 5080 29460 5092
rect 28767 5052 29460 5080
rect 28767 5049 28779 5052
rect 28721 5043 28779 5049
rect 29454 5040 29460 5052
rect 29512 5080 29518 5092
rect 29641 5083 29699 5089
rect 29641 5080 29653 5083
rect 29512 5052 29653 5080
rect 29512 5040 29518 5052
rect 29641 5049 29653 5052
rect 29687 5049 29699 5083
rect 31297 5083 31355 5089
rect 31297 5080 31309 5083
rect 29641 5043 29699 5049
rect 30668 5052 31309 5080
rect 30668 5024 30696 5052
rect 31297 5049 31309 5052
rect 31343 5049 31355 5083
rect 31297 5043 31355 5049
rect 31754 5040 31760 5092
rect 31812 5080 31818 5092
rect 33045 5083 33103 5089
rect 33045 5080 33057 5083
rect 31812 5052 33057 5080
rect 31812 5040 31818 5052
rect 33045 5049 33057 5052
rect 33091 5080 33103 5083
rect 33134 5080 33140 5092
rect 33091 5052 33140 5080
rect 33091 5049 33103 5052
rect 33045 5043 33103 5049
rect 33134 5040 33140 5052
rect 33192 5040 33198 5092
rect 33689 5083 33747 5089
rect 33689 5049 33701 5083
rect 33735 5080 33747 5083
rect 34238 5080 34244 5092
rect 33735 5052 34244 5080
rect 33735 5049 33747 5052
rect 33689 5043 33747 5049
rect 34238 5040 34244 5052
rect 34296 5040 34302 5092
rect 4982 4972 4988 5024
rect 5040 5012 5046 5024
rect 5629 5015 5687 5021
rect 5629 5012 5641 5015
rect 5040 4984 5641 5012
rect 5040 4972 5046 4984
rect 5629 4981 5641 4984
rect 5675 4981 5687 5015
rect 5629 4975 5687 4981
rect 5810 4972 5816 5024
rect 5868 5012 5874 5024
rect 6549 5015 6607 5021
rect 6549 5012 6561 5015
rect 5868 4984 6561 5012
rect 5868 4972 5874 4984
rect 6549 4981 6561 4984
rect 6595 4981 6607 5015
rect 6549 4975 6607 4981
rect 7009 5015 7067 5021
rect 7009 4981 7021 5015
rect 7055 5012 7067 5015
rect 7190 5012 7196 5024
rect 7055 4984 7196 5012
rect 7055 4981 7067 4984
rect 7009 4975 7067 4981
rect 7190 4972 7196 4984
rect 7248 4972 7254 5024
rect 8113 5015 8171 5021
rect 8113 4981 8125 5015
rect 8159 5012 8171 5015
rect 8386 5012 8392 5024
rect 8159 4984 8392 5012
rect 8159 4981 8171 4984
rect 8113 4975 8171 4981
rect 8386 4972 8392 4984
rect 8444 4972 8450 5024
rect 9401 5015 9459 5021
rect 9401 4981 9413 5015
rect 9447 5012 9459 5015
rect 10502 5012 10508 5024
rect 9447 4984 10508 5012
rect 9447 4981 9459 4984
rect 9401 4975 9459 4981
rect 10502 4972 10508 4984
rect 10560 4972 10566 5024
rect 11146 5012 11152 5024
rect 11107 4984 11152 5012
rect 11146 4972 11152 4984
rect 11204 4972 11210 5024
rect 11698 5012 11704 5024
rect 11659 4984 11704 5012
rect 11698 4972 11704 4984
rect 11756 4972 11762 5024
rect 12250 5012 12256 5024
rect 12211 4984 12256 5012
rect 12250 4972 12256 4984
rect 12308 4972 12314 5024
rect 13078 5012 13084 5024
rect 13039 4984 13084 5012
rect 13078 4972 13084 4984
rect 13136 4972 13142 5024
rect 15562 4972 15568 5024
rect 15620 5012 15626 5024
rect 15841 5015 15899 5021
rect 15841 5012 15853 5015
rect 15620 4984 15853 5012
rect 15620 4972 15626 4984
rect 15841 4981 15853 4984
rect 15887 4981 15899 5015
rect 15841 4975 15899 4981
rect 16574 4972 16580 5024
rect 16632 5012 16638 5024
rect 17494 5012 17500 5024
rect 16632 4984 16677 5012
rect 17407 4984 17500 5012
rect 16632 4972 16638 4984
rect 17494 4972 17500 4984
rect 17552 5012 17558 5024
rect 18138 5012 18144 5024
rect 17552 4984 18144 5012
rect 17552 4972 17558 4984
rect 18138 4972 18144 4984
rect 18196 5012 18202 5024
rect 18417 5015 18475 5021
rect 18417 5012 18429 5015
rect 18196 4984 18429 5012
rect 18196 4972 18202 4984
rect 18417 4981 18429 4984
rect 18463 4981 18475 5015
rect 18417 4975 18475 4981
rect 18506 4972 18512 5024
rect 18564 5012 18570 5024
rect 18690 5012 18696 5024
rect 18564 4984 18696 5012
rect 18564 4972 18570 4984
rect 18690 4972 18696 4984
rect 18748 4972 18754 5024
rect 22002 5012 22008 5024
rect 21963 4984 22008 5012
rect 22002 4972 22008 4984
rect 22060 4972 22066 5024
rect 25038 5012 25044 5024
rect 24999 4984 25044 5012
rect 25038 4972 25044 4984
rect 25096 4972 25102 5024
rect 26326 5012 26332 5024
rect 26287 4984 26332 5012
rect 26326 4972 26332 4984
rect 26384 4972 26390 5024
rect 27430 5012 27436 5024
rect 27391 4984 27436 5012
rect 27430 4972 27436 4984
rect 27488 4972 27494 5024
rect 27614 5012 27620 5024
rect 27575 4984 27620 5012
rect 27614 4972 27620 4984
rect 27672 4972 27678 5024
rect 27982 5012 27988 5024
rect 27943 4984 27988 5012
rect 27982 4972 27988 4984
rect 28040 4972 28046 5024
rect 29270 5012 29276 5024
rect 29231 4984 29276 5012
rect 29270 4972 29276 4984
rect 29328 4972 29334 5024
rect 29730 4972 29736 5024
rect 29788 5012 29794 5024
rect 30650 5012 30656 5024
rect 29788 4984 29833 5012
rect 30611 4984 30656 5012
rect 29788 4972 29794 4984
rect 30650 4972 30656 4984
rect 30708 4972 30714 5024
rect 30834 5012 30840 5024
rect 30795 4984 30840 5012
rect 30834 4972 30840 4984
rect 30892 4972 30898 5024
rect 31202 5012 31208 5024
rect 31163 4984 31208 5012
rect 31202 4972 31208 4984
rect 31260 4972 31266 5024
rect 32585 5015 32643 5021
rect 32585 4981 32597 5015
rect 32631 5012 32643 5015
rect 32674 5012 32680 5024
rect 32631 4984 32680 5012
rect 32631 4981 32643 4984
rect 32585 4975 32643 4981
rect 32674 4972 32680 4984
rect 32732 4972 32738 5024
rect 34698 4972 34704 5024
rect 34756 5012 34762 5024
rect 34885 5015 34943 5021
rect 34885 5012 34897 5015
rect 34756 4984 34897 5012
rect 34756 4972 34762 4984
rect 34885 4981 34897 4984
rect 34931 4981 34943 5015
rect 34885 4975 34943 4981
rect 1104 4922 38824 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 38824 4922
rect 1104 4848 38824 4870
rect 4525 4811 4583 4817
rect 4525 4777 4537 4811
rect 4571 4777 4583 4811
rect 4982 4808 4988 4820
rect 4943 4780 4988 4808
rect 4525 4771 4583 4777
rect 4540 4740 4568 4771
rect 4982 4768 4988 4780
rect 5040 4768 5046 4820
rect 5626 4768 5632 4820
rect 5684 4808 5690 4820
rect 6178 4808 6184 4820
rect 5684 4780 6184 4808
rect 5684 4768 5690 4780
rect 6178 4768 6184 4780
rect 6236 4808 6242 4820
rect 6549 4811 6607 4817
rect 6549 4808 6561 4811
rect 6236 4780 6561 4808
rect 6236 4768 6242 4780
rect 6549 4777 6561 4780
rect 6595 4777 6607 4811
rect 8386 4808 8392 4820
rect 8347 4780 8392 4808
rect 6549 4771 6607 4777
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 9306 4768 9312 4820
rect 9364 4808 9370 4820
rect 9401 4811 9459 4817
rect 9401 4808 9413 4811
rect 9364 4780 9413 4808
rect 9364 4768 9370 4780
rect 9401 4777 9413 4780
rect 9447 4777 9459 4811
rect 9401 4771 9459 4777
rect 10137 4811 10195 4817
rect 10137 4777 10149 4811
rect 10183 4808 10195 4811
rect 10962 4808 10968 4820
rect 10183 4780 10968 4808
rect 10183 4777 10195 4780
rect 10137 4771 10195 4777
rect 10962 4768 10968 4780
rect 11020 4768 11026 4820
rect 13814 4808 13820 4820
rect 13775 4780 13820 4808
rect 13814 4768 13820 4780
rect 13872 4768 13878 4820
rect 13909 4811 13967 4817
rect 13909 4777 13921 4811
rect 13955 4808 13967 4811
rect 15102 4808 15108 4820
rect 13955 4780 15108 4808
rect 13955 4777 13967 4780
rect 13909 4771 13967 4777
rect 6454 4740 6460 4752
rect 4540 4712 6460 4740
rect 6454 4700 6460 4712
rect 6512 4700 6518 4752
rect 8018 4700 8024 4752
rect 8076 4740 8082 4752
rect 8757 4743 8815 4749
rect 8757 4740 8769 4743
rect 8076 4712 8769 4740
rect 8076 4700 8082 4712
rect 8757 4709 8769 4712
rect 8803 4709 8815 4743
rect 10502 4740 10508 4752
rect 10463 4712 10508 4740
rect 8757 4703 8815 4709
rect 10502 4700 10508 4712
rect 10560 4700 10566 4752
rect 10778 4740 10784 4752
rect 10739 4712 10784 4740
rect 10778 4700 10784 4712
rect 10836 4700 10842 4752
rect 12250 4700 12256 4752
rect 12308 4740 12314 4752
rect 13924 4740 13952 4771
rect 15102 4768 15108 4780
rect 15160 4768 15166 4820
rect 15749 4811 15807 4817
rect 15749 4777 15761 4811
rect 15795 4808 15807 4811
rect 17034 4808 17040 4820
rect 15795 4780 17040 4808
rect 15795 4777 15807 4780
rect 15749 4771 15807 4777
rect 17034 4768 17040 4780
rect 17092 4808 17098 4820
rect 17494 4808 17500 4820
rect 17092 4780 17500 4808
rect 17092 4768 17098 4780
rect 17494 4768 17500 4780
rect 17552 4768 17558 4820
rect 17954 4768 17960 4820
rect 18012 4808 18018 4820
rect 18141 4811 18199 4817
rect 18141 4808 18153 4811
rect 18012 4780 18153 4808
rect 18012 4768 18018 4780
rect 18141 4777 18153 4780
rect 18187 4777 18199 4811
rect 18141 4771 18199 4777
rect 19426 4768 19432 4820
rect 19484 4808 19490 4820
rect 19613 4811 19671 4817
rect 19613 4808 19625 4811
rect 19484 4780 19625 4808
rect 19484 4768 19490 4780
rect 19613 4777 19625 4780
rect 19659 4808 19671 4811
rect 19978 4808 19984 4820
rect 19659 4780 19984 4808
rect 19659 4777 19671 4780
rect 19613 4771 19671 4777
rect 19978 4768 19984 4780
rect 20036 4768 20042 4820
rect 22281 4811 22339 4817
rect 22281 4777 22293 4811
rect 22327 4808 22339 4811
rect 22462 4808 22468 4820
rect 22327 4780 22468 4808
rect 22327 4777 22339 4780
rect 22281 4771 22339 4777
rect 22462 4768 22468 4780
rect 22520 4808 22526 4820
rect 23934 4808 23940 4820
rect 22520 4780 23940 4808
rect 22520 4768 22526 4780
rect 23934 4768 23940 4780
rect 23992 4768 23998 4820
rect 24302 4808 24308 4820
rect 24263 4780 24308 4808
rect 24302 4768 24308 4780
rect 24360 4768 24366 4820
rect 24765 4811 24823 4817
rect 24765 4777 24777 4811
rect 24811 4808 24823 4811
rect 25225 4811 25283 4817
rect 25225 4808 25237 4811
rect 24811 4780 25237 4808
rect 24811 4777 24823 4780
rect 24765 4771 24823 4777
rect 25225 4777 25237 4780
rect 25271 4808 25283 4811
rect 25498 4808 25504 4820
rect 25271 4780 25504 4808
rect 25271 4777 25283 4780
rect 25225 4771 25283 4777
rect 25498 4768 25504 4780
rect 25556 4768 25562 4820
rect 25866 4808 25872 4820
rect 25827 4780 25872 4808
rect 25866 4768 25872 4780
rect 25924 4768 25930 4820
rect 26234 4768 26240 4820
rect 26292 4808 26298 4820
rect 26292 4780 26337 4808
rect 26292 4768 26298 4780
rect 28258 4768 28264 4820
rect 28316 4808 28322 4820
rect 28445 4811 28503 4817
rect 28445 4808 28457 4811
rect 28316 4780 28457 4808
rect 28316 4768 28322 4780
rect 28445 4777 28457 4780
rect 28491 4777 28503 4811
rect 28445 4771 28503 4777
rect 29181 4811 29239 4817
rect 29181 4777 29193 4811
rect 29227 4808 29239 4811
rect 29641 4811 29699 4817
rect 29641 4808 29653 4811
rect 29227 4780 29653 4808
rect 29227 4777 29239 4780
rect 29181 4771 29239 4777
rect 29641 4777 29653 4780
rect 29687 4808 29699 4811
rect 29730 4808 29736 4820
rect 29687 4780 29736 4808
rect 29687 4777 29699 4780
rect 29641 4771 29699 4777
rect 29730 4768 29736 4780
rect 29788 4768 29794 4820
rect 29914 4808 29920 4820
rect 29875 4780 29920 4808
rect 29914 4768 29920 4780
rect 29972 4768 29978 4820
rect 31386 4808 31392 4820
rect 31347 4780 31392 4808
rect 31386 4768 31392 4780
rect 31444 4768 31450 4820
rect 31754 4768 31760 4820
rect 31812 4808 31818 4820
rect 32306 4808 32312 4820
rect 31812 4780 32312 4808
rect 31812 4768 31818 4780
rect 32306 4768 32312 4780
rect 32364 4768 32370 4820
rect 33045 4811 33103 4817
rect 33045 4777 33057 4811
rect 33091 4808 33103 4811
rect 33318 4808 33324 4820
rect 33091 4780 33324 4808
rect 33091 4777 33103 4780
rect 33045 4771 33103 4777
rect 33318 4768 33324 4780
rect 33376 4808 33382 4820
rect 33505 4811 33563 4817
rect 33505 4808 33517 4811
rect 33376 4780 33517 4808
rect 33376 4768 33382 4780
rect 33505 4777 33517 4780
rect 33551 4777 33563 4811
rect 34514 4808 34520 4820
rect 34475 4780 34520 4808
rect 33505 4771 33563 4777
rect 34514 4768 34520 4780
rect 34572 4808 34578 4820
rect 35161 4811 35219 4817
rect 35161 4808 35173 4811
rect 34572 4780 35173 4808
rect 34572 4768 34578 4780
rect 35161 4777 35173 4780
rect 35207 4777 35219 4811
rect 35161 4771 35219 4777
rect 12308 4712 13952 4740
rect 12308 4700 12314 4712
rect 16390 4700 16396 4752
rect 16448 4740 16454 4752
rect 16758 4740 16764 4752
rect 16448 4712 16764 4740
rect 16448 4700 16454 4712
rect 16758 4700 16764 4712
rect 16816 4700 16822 4752
rect 23106 4740 23112 4752
rect 23067 4712 23112 4740
rect 23106 4700 23112 4712
rect 23164 4700 23170 4752
rect 24578 4700 24584 4752
rect 24636 4740 24642 4752
rect 25884 4740 25912 4768
rect 24636 4712 25912 4740
rect 26780 4743 26838 4749
rect 24636 4700 24642 4712
rect 26780 4709 26792 4743
rect 26826 4740 26838 4743
rect 27706 4740 27712 4752
rect 26826 4712 27712 4740
rect 26826 4709 26838 4712
rect 26780 4703 26838 4709
rect 27706 4700 27712 4712
rect 27764 4700 27770 4752
rect 29270 4700 29276 4752
rect 29328 4740 29334 4752
rect 30745 4743 30803 4749
rect 30745 4740 30757 4743
rect 29328 4712 30757 4740
rect 29328 4700 29334 4712
rect 30745 4709 30757 4712
rect 30791 4740 30803 4743
rect 31478 4740 31484 4752
rect 30791 4712 31484 4740
rect 30791 4709 30803 4712
rect 30745 4703 30803 4709
rect 31478 4700 31484 4712
rect 31536 4700 31542 4752
rect 4890 4672 4896 4684
rect 4851 4644 4896 4672
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 5721 4675 5779 4681
rect 5721 4641 5733 4675
rect 5767 4672 5779 4675
rect 6270 4672 6276 4684
rect 5767 4644 6276 4672
rect 5767 4641 5779 4644
rect 5721 4635 5779 4641
rect 6270 4632 6276 4644
rect 6328 4632 6334 4684
rect 7745 4675 7803 4681
rect 7745 4641 7757 4675
rect 7791 4672 7803 4675
rect 7834 4672 7840 4684
rect 7791 4644 7840 4672
rect 7791 4641 7803 4644
rect 7745 4635 7803 4641
rect 7834 4632 7840 4644
rect 7892 4632 7898 4684
rect 9766 4672 9772 4684
rect 9727 4644 9772 4672
rect 9766 4632 9772 4644
rect 9824 4632 9830 4684
rect 9858 4632 9864 4684
rect 9916 4672 9922 4684
rect 9953 4675 10011 4681
rect 9953 4672 9965 4675
rect 9916 4644 9965 4672
rect 9916 4632 9922 4644
rect 9953 4641 9965 4644
rect 9999 4641 10011 4675
rect 9953 4635 10011 4641
rect 10965 4675 11023 4681
rect 10965 4641 10977 4675
rect 11011 4672 11023 4675
rect 11054 4672 11060 4684
rect 11011 4644 11060 4672
rect 11011 4641 11023 4644
rect 10965 4635 11023 4641
rect 11054 4632 11060 4644
rect 11112 4632 11118 4684
rect 11238 4681 11244 4684
rect 11232 4635 11244 4681
rect 11296 4672 11302 4684
rect 15654 4672 15660 4684
rect 11296 4644 11332 4672
rect 15615 4644 15660 4672
rect 11238 4632 11244 4635
rect 11296 4632 11302 4644
rect 15654 4632 15660 4644
rect 15712 4632 15718 4684
rect 17954 4632 17960 4684
rect 18012 4672 18018 4684
rect 18049 4675 18107 4681
rect 18049 4672 18061 4675
rect 18012 4644 18061 4672
rect 18012 4632 18018 4644
rect 18049 4641 18061 4644
rect 18095 4641 18107 4675
rect 20625 4675 20683 4681
rect 20625 4672 20637 4675
rect 18049 4635 18107 4641
rect 19720 4644 20637 4672
rect 19720 4616 19748 4644
rect 20625 4641 20637 4644
rect 20671 4641 20683 4675
rect 20625 4635 20683 4641
rect 20901 4675 20959 4681
rect 20901 4641 20913 4675
rect 20947 4672 20959 4675
rect 20990 4672 20996 4684
rect 20947 4644 20996 4672
rect 20947 4641 20959 4644
rect 20901 4635 20959 4641
rect 20990 4632 20996 4644
rect 21048 4632 21054 4684
rect 21174 4681 21180 4684
rect 21168 4672 21180 4681
rect 21135 4644 21180 4672
rect 21168 4635 21180 4644
rect 21174 4632 21180 4635
rect 21232 4632 21238 4684
rect 23385 4675 23443 4681
rect 23385 4641 23397 4675
rect 23431 4672 23443 4675
rect 23842 4672 23848 4684
rect 23431 4644 23848 4672
rect 23431 4641 23443 4644
rect 23385 4635 23443 4641
rect 23842 4632 23848 4644
rect 23900 4632 23906 4684
rect 27614 4632 27620 4684
rect 27672 4672 27678 4684
rect 28626 4672 28632 4684
rect 27672 4644 28632 4672
rect 27672 4632 27678 4644
rect 28626 4632 28632 4644
rect 28684 4672 28690 4684
rect 28997 4675 29055 4681
rect 28997 4672 29009 4675
rect 28684 4644 29009 4672
rect 28684 4632 28690 4644
rect 28997 4641 29009 4644
rect 29043 4641 29055 4675
rect 28997 4635 29055 4641
rect 30374 4632 30380 4684
rect 30432 4672 30438 4684
rect 30653 4675 30711 4681
rect 30653 4672 30665 4675
rect 30432 4644 30665 4672
rect 30432 4632 30438 4644
rect 30653 4641 30665 4644
rect 30699 4672 30711 4675
rect 32125 4675 32183 4681
rect 32125 4672 32137 4675
rect 30699 4644 32137 4672
rect 30699 4641 30711 4644
rect 30653 4635 30711 4641
rect 32125 4641 32137 4644
rect 32171 4641 32183 4675
rect 32125 4635 32183 4641
rect 34698 4632 34704 4684
rect 34756 4672 34762 4684
rect 35069 4675 35127 4681
rect 35069 4672 35081 4675
rect 34756 4644 35081 4672
rect 34756 4632 34762 4644
rect 35069 4641 35081 4644
rect 35115 4641 35127 4675
rect 35069 4635 35127 4641
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4604 4399 4607
rect 4982 4604 4988 4616
rect 4387 4576 4988 4604
rect 4387 4573 4399 4576
rect 4341 4567 4399 4573
rect 4982 4564 4988 4576
rect 5040 4564 5046 4616
rect 5077 4607 5135 4613
rect 5077 4573 5089 4607
rect 5123 4573 5135 4607
rect 5077 4567 5135 4573
rect 6733 4607 6791 4613
rect 6733 4573 6745 4607
rect 6779 4604 6791 4607
rect 8018 4604 8024 4616
rect 6779 4576 8024 4604
rect 6779 4573 6791 4576
rect 6733 4567 6791 4573
rect 4614 4496 4620 4548
rect 4672 4536 4678 4548
rect 5092 4536 5120 4567
rect 8018 4564 8024 4576
rect 8076 4564 8082 4616
rect 13357 4607 13415 4613
rect 13357 4573 13369 4607
rect 13403 4604 13415 4607
rect 14001 4607 14059 4613
rect 14001 4604 14013 4607
rect 13403 4576 14013 4604
rect 13403 4573 13415 4576
rect 13357 4567 13415 4573
rect 14001 4573 14013 4576
rect 14047 4604 14059 4607
rect 14274 4604 14280 4616
rect 14047 4576 14280 4604
rect 14047 4573 14059 4576
rect 14001 4567 14059 4573
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 15194 4564 15200 4616
rect 15252 4604 15258 4616
rect 15841 4607 15899 4613
rect 15841 4604 15853 4607
rect 15252 4576 15853 4604
rect 15252 4564 15258 4576
rect 15841 4573 15853 4576
rect 15887 4604 15899 4607
rect 16482 4604 16488 4616
rect 15887 4576 16488 4604
rect 15887 4573 15899 4576
rect 15841 4567 15899 4573
rect 16482 4564 16488 4576
rect 16540 4564 16546 4616
rect 17589 4607 17647 4613
rect 17589 4573 17601 4607
rect 17635 4604 17647 4607
rect 18325 4607 18383 4613
rect 18325 4604 18337 4607
rect 17635 4576 18337 4604
rect 17635 4573 17647 4576
rect 17589 4567 17647 4573
rect 18325 4573 18337 4576
rect 18371 4604 18383 4607
rect 18414 4604 18420 4616
rect 18371 4576 18420 4604
rect 18371 4573 18383 4576
rect 18325 4567 18383 4573
rect 18414 4564 18420 4576
rect 18472 4564 18478 4616
rect 18690 4604 18696 4616
rect 18651 4576 18696 4604
rect 18690 4564 18696 4576
rect 18748 4564 18754 4616
rect 19702 4604 19708 4616
rect 19663 4576 19708 4604
rect 19702 4564 19708 4576
rect 19760 4564 19766 4616
rect 19797 4607 19855 4613
rect 19797 4573 19809 4607
rect 19843 4573 19855 4607
rect 19797 4567 19855 4573
rect 5810 4536 5816 4548
rect 4672 4508 5816 4536
rect 4672 4496 4678 4508
rect 5810 4496 5816 4508
rect 5868 4496 5874 4548
rect 14182 4496 14188 4548
rect 14240 4536 14246 4548
rect 15013 4539 15071 4545
rect 15013 4536 15025 4539
rect 14240 4508 15025 4536
rect 14240 4496 14246 4508
rect 15013 4505 15025 4508
rect 15059 4536 15071 4539
rect 15746 4536 15752 4548
rect 15059 4508 15752 4536
rect 15059 4505 15071 4508
rect 15013 4499 15071 4505
rect 15746 4496 15752 4508
rect 15804 4496 15810 4548
rect 16298 4536 16304 4548
rect 16259 4508 16304 4536
rect 16298 4496 16304 4508
rect 16356 4496 16362 4548
rect 17221 4539 17279 4545
rect 17221 4505 17233 4539
rect 17267 4536 17279 4539
rect 17681 4539 17739 4545
rect 17681 4536 17693 4539
rect 17267 4508 17693 4536
rect 17267 4505 17279 4508
rect 17221 4499 17279 4505
rect 17681 4505 17693 4508
rect 17727 4536 17739 4539
rect 17862 4536 17868 4548
rect 17727 4508 17868 4536
rect 17727 4505 17739 4508
rect 17681 4499 17739 4505
rect 17862 4496 17868 4508
rect 17920 4496 17926 4548
rect 19153 4539 19211 4545
rect 19153 4505 19165 4539
rect 19199 4536 19211 4539
rect 19334 4536 19340 4548
rect 19199 4508 19340 4536
rect 19199 4505 19211 4508
rect 19153 4499 19211 4505
rect 19334 4496 19340 4508
rect 19392 4536 19398 4548
rect 19812 4536 19840 4567
rect 24670 4564 24676 4616
rect 24728 4604 24734 4616
rect 25317 4607 25375 4613
rect 25317 4604 25329 4607
rect 24728 4576 25329 4604
rect 24728 4564 24734 4576
rect 25317 4573 25329 4576
rect 25363 4573 25375 4607
rect 25317 4567 25375 4573
rect 25409 4607 25467 4613
rect 25409 4573 25421 4607
rect 25455 4573 25467 4607
rect 26510 4604 26516 4616
rect 26471 4576 26516 4604
rect 25409 4567 25467 4573
rect 19392 4508 19840 4536
rect 19392 4496 19398 4508
rect 24946 4496 24952 4548
rect 25004 4536 25010 4548
rect 25424 4536 25452 4567
rect 26510 4564 26516 4576
rect 26568 4564 26574 4616
rect 30834 4564 30840 4616
rect 30892 4604 30898 4616
rect 33597 4607 33655 4613
rect 30892 4576 30937 4604
rect 30892 4564 30898 4576
rect 33597 4573 33609 4607
rect 33643 4573 33655 4607
rect 33778 4604 33784 4616
rect 33739 4576 33784 4604
rect 33597 4567 33655 4573
rect 26142 4536 26148 4548
rect 25004 4508 26148 4536
rect 25004 4496 25010 4508
rect 26142 4496 26148 4508
rect 26200 4496 26206 4548
rect 27890 4536 27896 4548
rect 27851 4508 27896 4536
rect 27890 4496 27896 4508
rect 27948 4496 27954 4548
rect 32677 4539 32735 4545
rect 32677 4505 32689 4539
rect 32723 4536 32735 4539
rect 33042 4536 33048 4548
rect 32723 4508 33048 4536
rect 32723 4505 32735 4508
rect 32677 4499 32735 4505
rect 33042 4496 33048 4508
rect 33100 4536 33106 4548
rect 33137 4539 33195 4545
rect 33137 4536 33149 4539
rect 33100 4508 33149 4536
rect 33100 4496 33106 4508
rect 33137 4505 33149 4508
rect 33183 4505 33195 4539
rect 33137 4499 33195 4505
rect 6086 4468 6092 4480
rect 6047 4440 6092 4468
rect 6086 4428 6092 4440
rect 6144 4428 6150 4480
rect 7193 4471 7251 4477
rect 7193 4437 7205 4471
rect 7239 4468 7251 4471
rect 7282 4468 7288 4480
rect 7239 4440 7288 4468
rect 7239 4437 7251 4440
rect 7193 4431 7251 4437
rect 7282 4428 7288 4440
rect 7340 4428 7346 4480
rect 7466 4468 7472 4480
rect 7427 4440 7472 4468
rect 7466 4428 7472 4440
rect 7524 4428 7530 4480
rect 7929 4471 7987 4477
rect 7929 4437 7941 4471
rect 7975 4468 7987 4471
rect 8294 4468 8300 4480
rect 7975 4440 8300 4468
rect 7975 4437 7987 4440
rect 7929 4431 7987 4437
rect 8294 4428 8300 4440
rect 8352 4428 8358 4480
rect 12342 4468 12348 4480
rect 12303 4440 12348 4468
rect 12342 4428 12348 4440
rect 12400 4428 12406 4480
rect 12894 4468 12900 4480
rect 12855 4440 12900 4468
rect 12894 4428 12900 4440
rect 12952 4428 12958 4480
rect 13354 4428 13360 4480
rect 13412 4468 13418 4480
rect 13449 4471 13507 4477
rect 13449 4468 13461 4471
rect 13412 4440 13461 4468
rect 13412 4428 13418 4440
rect 13449 4437 13461 4440
rect 13495 4437 13507 4471
rect 13449 4431 13507 4437
rect 13814 4428 13820 4480
rect 13872 4468 13878 4480
rect 14090 4468 14096 4480
rect 13872 4440 14096 4468
rect 13872 4428 13878 4440
rect 14090 4428 14096 4440
rect 14148 4468 14154 4480
rect 14461 4471 14519 4477
rect 14461 4468 14473 4471
rect 14148 4440 14473 4468
rect 14148 4428 14154 4440
rect 14461 4437 14473 4440
rect 14507 4437 14519 4471
rect 15286 4468 15292 4480
rect 15247 4440 15292 4468
rect 14461 4431 14519 4437
rect 15286 4428 15292 4440
rect 15344 4428 15350 4480
rect 19242 4468 19248 4480
rect 19203 4440 19248 4468
rect 19242 4428 19248 4440
rect 19300 4428 19306 4480
rect 20346 4468 20352 4480
rect 20307 4440 20352 4468
rect 20346 4428 20352 4440
rect 20404 4428 20410 4480
rect 23566 4468 23572 4480
rect 23527 4440 23572 4468
rect 23566 4428 23572 4440
rect 23624 4428 23630 4480
rect 24857 4471 24915 4477
rect 24857 4437 24869 4471
rect 24903 4468 24915 4471
rect 27430 4468 27436 4480
rect 24903 4440 27436 4468
rect 24903 4437 24915 4440
rect 24857 4431 24915 4437
rect 27430 4428 27436 4440
rect 27488 4468 27494 4480
rect 28994 4468 29000 4480
rect 27488 4440 29000 4468
rect 27488 4428 27494 4440
rect 28994 4428 29000 4440
rect 29052 4428 29058 4480
rect 30282 4468 30288 4480
rect 30243 4440 30288 4468
rect 30282 4428 30288 4440
rect 30340 4428 30346 4480
rect 33612 4468 33640 4567
rect 33778 4564 33784 4576
rect 33836 4564 33842 4616
rect 35345 4607 35403 4613
rect 35345 4573 35357 4607
rect 35391 4604 35403 4607
rect 35434 4604 35440 4616
rect 35391 4576 35440 4604
rect 35391 4573 35403 4576
rect 35345 4567 35403 4573
rect 35434 4564 35440 4576
rect 35492 4564 35498 4616
rect 34701 4539 34759 4545
rect 34701 4505 34713 4539
rect 34747 4536 34759 4539
rect 34790 4536 34796 4548
rect 34747 4508 34796 4536
rect 34747 4505 34759 4508
rect 34701 4499 34759 4505
rect 34790 4496 34796 4508
rect 34848 4536 34854 4548
rect 36078 4536 36084 4548
rect 34848 4508 36084 4536
rect 34848 4496 34854 4508
rect 36078 4496 36084 4508
rect 36136 4496 36142 4548
rect 34241 4471 34299 4477
rect 34241 4468 34253 4471
rect 33612 4440 34253 4468
rect 34241 4437 34253 4440
rect 34287 4468 34299 4471
rect 34422 4468 34428 4480
rect 34287 4440 34428 4468
rect 34287 4437 34299 4440
rect 34241 4431 34299 4437
rect 34422 4428 34428 4440
rect 34480 4428 34486 4480
rect 35710 4468 35716 4480
rect 35671 4440 35716 4468
rect 35710 4428 35716 4440
rect 35768 4428 35774 4480
rect 1104 4378 38824 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 38824 4378
rect 1104 4304 38824 4326
rect 4062 4264 4068 4276
rect 4023 4236 4068 4264
rect 4062 4224 4068 4236
rect 4120 4224 4126 4276
rect 6178 4264 6184 4276
rect 6139 4236 6184 4264
rect 6178 4224 6184 4236
rect 6236 4224 6242 4276
rect 6454 4224 6460 4276
rect 6512 4264 6518 4276
rect 6549 4267 6607 4273
rect 6549 4264 6561 4267
rect 6512 4236 6561 4264
rect 6512 4224 6518 4236
rect 6549 4233 6561 4236
rect 6595 4233 6607 4267
rect 6549 4227 6607 4233
rect 6825 4267 6883 4273
rect 6825 4233 6837 4267
rect 6871 4264 6883 4267
rect 7926 4264 7932 4276
rect 6871 4236 7932 4264
rect 6871 4233 6883 4236
rect 6825 4227 6883 4233
rect 7926 4224 7932 4236
rect 7984 4224 7990 4276
rect 11054 4264 11060 4276
rect 11015 4236 11060 4264
rect 11054 4224 11060 4236
rect 11112 4224 11118 4276
rect 11146 4224 11152 4276
rect 11204 4264 11210 4276
rect 11333 4267 11391 4273
rect 11333 4264 11345 4267
rect 11204 4236 11345 4264
rect 11204 4224 11210 4236
rect 11333 4233 11345 4236
rect 11379 4233 11391 4267
rect 11333 4227 11391 4233
rect 13998 4224 14004 4276
rect 14056 4264 14062 4276
rect 14093 4267 14151 4273
rect 14093 4264 14105 4267
rect 14056 4236 14105 4264
rect 14056 4224 14062 4236
rect 14093 4233 14105 4236
rect 14139 4233 14151 4267
rect 14093 4227 14151 4233
rect 8018 4196 8024 4208
rect 7392 4168 8024 4196
rect 3050 4128 3056 4140
rect 3011 4100 3056 4128
rect 3050 4088 3056 4100
rect 3108 4128 3114 4140
rect 7392 4137 7420 4168
rect 8018 4156 8024 4168
rect 8076 4156 8082 4208
rect 11164 4196 11192 4224
rect 10612 4168 11192 4196
rect 3789 4131 3847 4137
rect 3108 4100 3188 4128
rect 3108 4088 3114 4100
rect 3160 4069 3188 4100
rect 3789 4097 3801 4131
rect 3835 4128 3847 4131
rect 7377 4131 7435 4137
rect 3835 4100 4384 4128
rect 3835 4097 3847 4100
rect 3789 4091 3847 4097
rect 3145 4063 3203 4069
rect 3145 4029 3157 4063
rect 3191 4029 3203 4063
rect 3145 4023 3203 4029
rect 4062 4020 4068 4072
rect 4120 4060 4126 4072
rect 4249 4063 4307 4069
rect 4249 4060 4261 4063
rect 4120 4032 4261 4060
rect 4120 4020 4126 4032
rect 4249 4029 4261 4032
rect 4295 4029 4307 4063
rect 4356 4060 4384 4100
rect 7377 4097 7389 4131
rect 7423 4097 7435 4131
rect 7926 4128 7932 4140
rect 7887 4100 7932 4128
rect 7377 4091 7435 4097
rect 7926 4088 7932 4100
rect 7984 4088 7990 4140
rect 9030 4128 9036 4140
rect 8991 4100 9036 4128
rect 9030 4088 9036 4100
rect 9088 4088 9094 4140
rect 10413 4131 10471 4137
rect 10413 4097 10425 4131
rect 10459 4128 10471 4131
rect 10502 4128 10508 4140
rect 10459 4100 10508 4128
rect 10459 4097 10471 4100
rect 10413 4091 10471 4097
rect 10502 4088 10508 4100
rect 10560 4088 10566 4140
rect 10612 4137 10640 4168
rect 10597 4131 10655 4137
rect 10597 4097 10609 4131
rect 10643 4097 10655 4131
rect 10597 4091 10655 4097
rect 11882 4088 11888 4140
rect 11940 4128 11946 4140
rect 12342 4128 12348 4140
rect 11940 4100 12348 4128
rect 11940 4088 11946 4100
rect 12342 4088 12348 4100
rect 12400 4128 12406 4140
rect 12989 4131 13047 4137
rect 12989 4128 13001 4131
rect 12400 4100 13001 4128
rect 12400 4088 12406 4100
rect 12989 4097 13001 4100
rect 13035 4097 13047 4131
rect 12989 4091 13047 4097
rect 13541 4131 13599 4137
rect 13541 4097 13553 4131
rect 13587 4128 13599 4131
rect 13722 4128 13728 4140
rect 13587 4100 13728 4128
rect 13587 4097 13599 4100
rect 13541 4091 13599 4097
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 14108 4128 14136 4227
rect 15654 4224 15660 4276
rect 15712 4264 15718 4276
rect 16209 4267 16267 4273
rect 16209 4264 16221 4267
rect 15712 4236 16221 4264
rect 15712 4224 15718 4236
rect 16209 4233 16221 4236
rect 16255 4233 16267 4267
rect 16209 4227 16267 4233
rect 18414 4224 18420 4276
rect 18472 4264 18478 4276
rect 19981 4267 20039 4273
rect 19981 4264 19993 4267
rect 18472 4236 19993 4264
rect 18472 4224 18478 4236
rect 19981 4233 19993 4236
rect 20027 4264 20039 4267
rect 21174 4264 21180 4276
rect 20027 4236 21180 4264
rect 20027 4233 20039 4236
rect 19981 4227 20039 4233
rect 21174 4224 21180 4236
rect 21232 4264 21238 4276
rect 22097 4267 22155 4273
rect 22097 4264 22109 4267
rect 21232 4236 22109 4264
rect 21232 4224 21238 4236
rect 22097 4233 22109 4236
rect 22143 4233 22155 4267
rect 22097 4227 22155 4233
rect 26510 4224 26516 4276
rect 26568 4264 26574 4276
rect 27525 4267 27583 4273
rect 27525 4264 27537 4267
rect 26568 4236 27537 4264
rect 26568 4224 26574 4236
rect 27525 4233 27537 4236
rect 27571 4233 27583 4267
rect 28258 4264 28264 4276
rect 28219 4236 28264 4264
rect 27525 4227 27583 4233
rect 28258 4224 28264 4236
rect 28316 4224 28322 4276
rect 28626 4264 28632 4276
rect 28587 4236 28632 4264
rect 28626 4224 28632 4236
rect 28684 4224 28690 4276
rect 29454 4264 29460 4276
rect 29415 4236 29460 4264
rect 29454 4224 29460 4236
rect 29512 4224 29518 4276
rect 30374 4264 30380 4276
rect 30335 4236 30380 4264
rect 30374 4224 30380 4236
rect 30432 4224 30438 4276
rect 34698 4264 34704 4276
rect 34659 4236 34704 4264
rect 34698 4224 34704 4236
rect 34756 4224 34762 4276
rect 20346 4196 20352 4208
rect 19628 4168 20352 4196
rect 14277 4131 14335 4137
rect 14277 4128 14289 4131
rect 14108 4100 14289 4128
rect 14277 4097 14289 4100
rect 14323 4097 14335 4131
rect 17770 4128 17776 4140
rect 17731 4100 17776 4128
rect 14277 4091 14335 4097
rect 17770 4088 17776 4100
rect 17828 4088 17834 4140
rect 4516 4063 4574 4069
rect 4516 4060 4528 4063
rect 4356 4032 4528 4060
rect 4249 4023 4307 4029
rect 4516 4029 4528 4032
rect 4562 4060 4574 4063
rect 4982 4060 4988 4072
rect 4562 4032 4988 4060
rect 4562 4029 4574 4032
rect 4516 4023 4574 4029
rect 4982 4020 4988 4032
rect 5040 4020 5046 4072
rect 7193 4063 7251 4069
rect 7193 4029 7205 4063
rect 7239 4060 7251 4063
rect 7466 4060 7472 4072
rect 7239 4032 7472 4060
rect 7239 4029 7251 4032
rect 7193 4023 7251 4029
rect 7466 4020 7472 4032
rect 7524 4020 7530 4072
rect 8386 4020 8392 4072
rect 8444 4060 8450 4072
rect 8757 4063 8815 4069
rect 8757 4060 8769 4063
rect 8444 4032 8769 4060
rect 8444 4020 8450 4032
rect 8757 4029 8769 4032
rect 8803 4029 8815 4063
rect 10321 4063 10379 4069
rect 10321 4060 10333 4063
rect 8757 4023 8815 4029
rect 9416 4032 10333 4060
rect 8297 3995 8355 4001
rect 8297 3961 8309 3995
rect 8343 3992 8355 3995
rect 8478 3992 8484 4004
rect 8343 3964 8484 3992
rect 8343 3961 8355 3964
rect 8297 3955 8355 3961
rect 8478 3952 8484 3964
rect 8536 3992 8542 4004
rect 8849 3995 8907 4001
rect 8849 3992 8861 3995
rect 8536 3964 8861 3992
rect 8536 3952 8542 3964
rect 8849 3961 8861 3964
rect 8895 3961 8907 3995
rect 8849 3955 8907 3961
rect 3326 3924 3332 3936
rect 3287 3896 3332 3924
rect 3326 3884 3332 3896
rect 3384 3884 3390 3936
rect 4890 3884 4896 3936
rect 4948 3924 4954 3936
rect 5629 3927 5687 3933
rect 5629 3924 5641 3927
rect 4948 3896 5641 3924
rect 4948 3884 4954 3896
rect 5629 3893 5641 3896
rect 5675 3893 5687 3927
rect 7282 3924 7288 3936
rect 7243 3896 7288 3924
rect 5629 3887 5687 3893
rect 7282 3884 7288 3896
rect 7340 3884 7346 3936
rect 8389 3927 8447 3933
rect 8389 3893 8401 3927
rect 8435 3924 8447 3927
rect 9416 3924 9444 4032
rect 10321 4029 10333 4032
rect 10367 4060 10379 4063
rect 10778 4060 10784 4072
rect 10367 4032 10784 4060
rect 10367 4029 10379 4032
rect 10321 4023 10379 4029
rect 10778 4020 10784 4032
rect 10836 4020 10842 4072
rect 12158 4060 12164 4072
rect 12119 4032 12164 4060
rect 12158 4020 12164 4032
rect 12216 4060 12222 4072
rect 12805 4063 12863 4069
rect 12805 4060 12817 4063
rect 12216 4032 12817 4060
rect 12216 4020 12222 4032
rect 12805 4029 12817 4032
rect 12851 4029 12863 4063
rect 12805 4023 12863 4029
rect 14544 4063 14602 4069
rect 14544 4029 14556 4063
rect 14590 4060 14602 4063
rect 15010 4060 15016 4072
rect 14590 4032 15016 4060
rect 14590 4029 14602 4032
rect 14544 4023 14602 4029
rect 15010 4020 15016 4032
rect 15068 4020 15074 4072
rect 16758 4060 16764 4072
rect 16671 4032 16764 4060
rect 16758 4020 16764 4032
rect 16816 4060 16822 4072
rect 18874 4069 18880 4072
rect 17313 4063 17371 4069
rect 17313 4060 17325 4063
rect 16816 4032 17325 4060
rect 16816 4020 16822 4032
rect 17313 4029 17325 4032
rect 17359 4029 17371 4063
rect 18601 4063 18659 4069
rect 18601 4060 18613 4063
rect 17313 4023 17371 4029
rect 18432 4032 18613 4060
rect 9493 3995 9551 4001
rect 9493 3961 9505 3995
rect 9539 3992 9551 3995
rect 9858 3992 9864 4004
rect 9539 3964 9864 3992
rect 9539 3961 9551 3964
rect 9493 3955 9551 3961
rect 9858 3952 9864 3964
rect 9916 3952 9922 4004
rect 13722 3992 13728 4004
rect 12452 3964 13728 3992
rect 9766 3924 9772 3936
rect 8435 3896 9444 3924
rect 9727 3896 9772 3924
rect 8435 3893 8447 3896
rect 8389 3887 8447 3893
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 9950 3924 9956 3936
rect 9911 3896 9956 3924
rect 9950 3884 9956 3896
rect 10008 3884 10014 3936
rect 11882 3924 11888 3936
rect 11843 3896 11888 3924
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 12452 3933 12480 3964
rect 13722 3952 13728 3964
rect 13780 3952 13786 4004
rect 12437 3927 12495 3933
rect 12437 3893 12449 3927
rect 12483 3893 12495 3927
rect 12894 3924 12900 3936
rect 12855 3896 12900 3924
rect 12437 3887 12495 3893
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 15654 3924 15660 3936
rect 15615 3896 15660 3924
rect 15654 3884 15660 3896
rect 15712 3884 15718 3936
rect 16666 3924 16672 3936
rect 16627 3896 16672 3924
rect 16666 3884 16672 3896
rect 16724 3884 16730 3936
rect 16942 3924 16948 3936
rect 16903 3896 16948 3924
rect 16942 3884 16948 3896
rect 17000 3884 17006 3936
rect 18046 3884 18052 3936
rect 18104 3924 18110 3936
rect 18432 3933 18460 4032
rect 18601 4029 18613 4032
rect 18647 4029 18659 4063
rect 18868 4060 18880 4069
rect 18787 4032 18880 4060
rect 18601 4023 18659 4029
rect 18868 4023 18880 4032
rect 18932 4060 18938 4072
rect 19628 4060 19656 4168
rect 20346 4156 20352 4168
rect 20404 4156 20410 4208
rect 23566 4156 23572 4208
rect 23624 4196 23630 4208
rect 25590 4196 25596 4208
rect 23624 4168 25596 4196
rect 23624 4156 23630 4168
rect 21542 4088 21548 4140
rect 21600 4128 21606 4140
rect 21637 4131 21695 4137
rect 21637 4128 21649 4131
rect 21600 4100 21649 4128
rect 21600 4088 21606 4100
rect 21637 4097 21649 4100
rect 21683 4128 21695 4131
rect 22830 4128 22836 4140
rect 21683 4100 22836 4128
rect 21683 4097 21695 4100
rect 21637 4091 21695 4097
rect 22830 4088 22836 4100
rect 22888 4088 22894 4140
rect 24228 4137 24256 4168
rect 25590 4156 25596 4168
rect 25648 4156 25654 4208
rect 30834 4196 30840 4208
rect 30392 4168 30840 4196
rect 24213 4131 24271 4137
rect 24213 4097 24225 4131
rect 24259 4097 24271 4131
rect 24670 4128 24676 4140
rect 24631 4100 24676 4128
rect 24213 4091 24271 4097
rect 24670 4088 24676 4100
rect 24728 4088 24734 4140
rect 25133 4131 25191 4137
rect 25133 4097 25145 4131
rect 25179 4128 25191 4131
rect 25179 4100 25728 4128
rect 25179 4097 25191 4100
rect 25133 4091 25191 4097
rect 20990 4060 20996 4072
rect 18932 4032 19656 4060
rect 20951 4032 20996 4060
rect 18874 4020 18880 4023
rect 18932 4020 18938 4032
rect 20990 4020 20996 4032
rect 21048 4020 21054 4072
rect 21450 4060 21456 4072
rect 21411 4032 21456 4060
rect 21450 4020 21456 4032
rect 21508 4060 21514 4072
rect 22465 4063 22523 4069
rect 22465 4060 22477 4063
rect 21508 4032 22477 4060
rect 21508 4020 21514 4032
rect 22465 4029 22477 4032
rect 22511 4029 22523 4063
rect 22465 4023 22523 4029
rect 23658 4020 23664 4072
rect 23716 4060 23722 4072
rect 24029 4063 24087 4069
rect 24029 4060 24041 4063
rect 23716 4032 24041 4060
rect 23716 4020 23722 4032
rect 24029 4029 24041 4032
rect 24075 4029 24087 4063
rect 24029 4023 24087 4029
rect 24121 4063 24179 4069
rect 24121 4029 24133 4063
rect 24167 4060 24179 4063
rect 24302 4060 24308 4072
rect 24167 4032 24308 4060
rect 24167 4029 24179 4032
rect 24121 4023 24179 4029
rect 24302 4020 24308 4032
rect 24360 4020 24366 4072
rect 24762 4020 24768 4072
rect 24820 4060 24826 4072
rect 25409 4063 25467 4069
rect 25409 4060 25421 4063
rect 24820 4032 25421 4060
rect 24820 4020 24826 4032
rect 25409 4029 25421 4032
rect 25455 4060 25467 4063
rect 25498 4060 25504 4072
rect 25455 4032 25504 4060
rect 25455 4029 25467 4032
rect 25409 4023 25467 4029
rect 25498 4020 25504 4032
rect 25556 4060 25562 4072
rect 25593 4063 25651 4069
rect 25593 4060 25605 4063
rect 25556 4032 25605 4060
rect 25556 4020 25562 4032
rect 25593 4029 25605 4032
rect 25639 4029 25651 4063
rect 25700 4060 25728 4100
rect 27706 4088 27712 4140
rect 27764 4128 27770 4140
rect 27893 4131 27951 4137
rect 27893 4128 27905 4131
rect 27764 4100 27905 4128
rect 27764 4088 27770 4100
rect 27893 4097 27905 4100
rect 27939 4097 27951 4131
rect 27893 4091 27951 4097
rect 28994 4088 29000 4140
rect 29052 4128 29058 4140
rect 30006 4128 30012 4140
rect 29052 4100 29097 4128
rect 29919 4100 30012 4128
rect 29052 4088 29058 4100
rect 30006 4088 30012 4100
rect 30064 4128 30070 4140
rect 30392 4128 30420 4168
rect 30834 4156 30840 4168
rect 30892 4156 30898 4208
rect 30064 4100 30420 4128
rect 30064 4088 30070 4100
rect 30742 4088 30748 4140
rect 30800 4128 30806 4140
rect 31389 4131 31447 4137
rect 31389 4128 31401 4131
rect 30800 4100 31401 4128
rect 30800 4088 30806 4100
rect 31389 4097 31401 4100
rect 31435 4128 31447 4131
rect 31754 4128 31760 4140
rect 31435 4100 31760 4128
rect 31435 4097 31447 4100
rect 31389 4091 31447 4097
rect 31754 4088 31760 4100
rect 31812 4128 31818 4140
rect 31812 4100 32444 4128
rect 31812 4088 31818 4100
rect 25866 4069 25872 4072
rect 25860 4060 25872 4069
rect 25700 4032 25872 4060
rect 25593 4023 25651 4029
rect 25860 4023 25872 4032
rect 20625 3995 20683 4001
rect 20625 3961 20637 3995
rect 20671 3992 20683 3995
rect 23477 3995 23535 4001
rect 20671 3964 21588 3992
rect 20671 3961 20683 3964
rect 20625 3955 20683 3961
rect 18417 3927 18475 3933
rect 18417 3924 18429 3927
rect 18104 3896 18429 3924
rect 18104 3884 18110 3896
rect 18417 3893 18429 3896
rect 18463 3893 18475 3927
rect 21082 3924 21088 3936
rect 21043 3896 21088 3924
rect 18417 3887 18475 3893
rect 21082 3884 21088 3896
rect 21140 3884 21146 3936
rect 21560 3933 21588 3964
rect 23477 3961 23489 3995
rect 23523 3992 23535 3995
rect 23842 3992 23848 4004
rect 23523 3964 23848 3992
rect 23523 3961 23535 3964
rect 23477 3955 23535 3961
rect 23842 3952 23848 3964
rect 23900 3952 23906 4004
rect 25608 3992 25636 4023
rect 25866 4020 25872 4023
rect 25924 4020 25930 4072
rect 28077 4063 28135 4069
rect 28077 4029 28089 4063
rect 28123 4060 28135 4063
rect 28258 4060 28264 4072
rect 28123 4032 28264 4060
rect 28123 4029 28135 4032
rect 28077 4023 28135 4029
rect 28258 4020 28264 4032
rect 28316 4020 28322 4072
rect 29012 4060 29040 4088
rect 29273 4063 29331 4069
rect 29273 4060 29285 4063
rect 29012 4032 29285 4060
rect 29273 4029 29285 4032
rect 29319 4029 29331 4063
rect 29273 4023 29331 4029
rect 30374 4020 30380 4072
rect 30432 4060 30438 4072
rect 31113 4063 31171 4069
rect 31113 4060 31125 4063
rect 30432 4032 31125 4060
rect 30432 4020 30438 4032
rect 31113 4029 31125 4032
rect 31159 4060 31171 4063
rect 32309 4063 32367 4069
rect 32309 4060 32321 4063
rect 31159 4032 31892 4060
rect 31159 4029 31171 4032
rect 31113 4023 31171 4029
rect 26510 3992 26516 4004
rect 25608 3964 26516 3992
rect 26510 3952 26516 3964
rect 26568 3952 26574 4004
rect 31662 3992 31668 4004
rect 30760 3964 31668 3992
rect 21545 3927 21603 3933
rect 21545 3893 21557 3927
rect 21591 3924 21603 3927
rect 22370 3924 22376 3936
rect 21591 3896 22376 3924
rect 21591 3893 21603 3896
rect 21545 3887 21603 3893
rect 22370 3884 22376 3896
rect 22428 3884 22434 3936
rect 23290 3884 23296 3936
rect 23348 3924 23354 3936
rect 23661 3927 23719 3933
rect 23661 3924 23673 3927
rect 23348 3896 23673 3924
rect 23348 3884 23354 3896
rect 23661 3893 23673 3896
rect 23707 3893 23719 3927
rect 26970 3924 26976 3936
rect 26931 3896 26976 3924
rect 23661 3887 23719 3893
rect 26970 3884 26976 3896
rect 27028 3884 27034 3936
rect 30760 3933 30788 3964
rect 31662 3952 31668 3964
rect 31720 3952 31726 4004
rect 31864 3936 31892 4032
rect 32140 4032 32321 4060
rect 32140 3936 32168 4032
rect 32309 4029 32321 4032
rect 32355 4029 32367 4063
rect 32416 4060 32444 4100
rect 32565 4063 32623 4069
rect 32565 4060 32577 4063
rect 32416 4032 32577 4060
rect 32309 4023 32367 4029
rect 32565 4029 32577 4032
rect 32611 4029 32623 4063
rect 32565 4023 32623 4029
rect 35158 4020 35164 4072
rect 35216 4060 35222 4072
rect 35710 4069 35716 4072
rect 35345 4063 35403 4069
rect 35345 4060 35357 4063
rect 35216 4032 35357 4060
rect 35216 4020 35222 4032
rect 35345 4029 35357 4032
rect 35391 4060 35403 4063
rect 35437 4063 35495 4069
rect 35437 4060 35449 4063
rect 35391 4032 35449 4060
rect 35391 4029 35403 4032
rect 35345 4023 35403 4029
rect 35437 4029 35449 4032
rect 35483 4029 35495 4063
rect 35704 4060 35716 4069
rect 35671 4032 35716 4060
rect 35437 4023 35495 4029
rect 35704 4023 35716 4032
rect 35710 4020 35716 4023
rect 35768 4020 35774 4072
rect 35250 3952 35256 4004
rect 35308 3992 35314 4004
rect 35526 3992 35532 4004
rect 35308 3964 35532 3992
rect 35308 3952 35314 3964
rect 35526 3952 35532 3964
rect 35584 3952 35590 4004
rect 30745 3927 30803 3933
rect 30745 3893 30757 3927
rect 30791 3893 30803 3927
rect 30745 3887 30803 3893
rect 31202 3884 31208 3936
rect 31260 3924 31266 3936
rect 31846 3924 31852 3936
rect 31260 3896 31305 3924
rect 31807 3896 31852 3924
rect 31260 3884 31266 3896
rect 31846 3884 31852 3896
rect 31904 3884 31910 3936
rect 32122 3924 32128 3936
rect 32083 3896 32128 3924
rect 32122 3884 32128 3896
rect 32180 3884 32186 3936
rect 32950 3884 32956 3936
rect 33008 3924 33014 3936
rect 33686 3924 33692 3936
rect 33008 3896 33692 3924
rect 33008 3884 33014 3896
rect 33686 3884 33692 3896
rect 33744 3884 33750 3936
rect 33778 3884 33784 3936
rect 33836 3924 33842 3936
rect 34333 3927 34391 3933
rect 34333 3924 34345 3927
rect 33836 3896 34345 3924
rect 33836 3884 33842 3896
rect 34333 3893 34345 3896
rect 34379 3924 34391 3927
rect 35894 3924 35900 3936
rect 34379 3896 35900 3924
rect 34379 3893 34391 3896
rect 34333 3887 34391 3893
rect 35894 3884 35900 3896
rect 35952 3924 35958 3936
rect 36817 3927 36875 3933
rect 36817 3924 36829 3927
rect 35952 3896 36829 3924
rect 35952 3884 35958 3896
rect 36817 3893 36829 3896
rect 36863 3893 36875 3927
rect 36817 3887 36875 3893
rect 1104 3834 38824 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 38824 3834
rect 1104 3760 38824 3782
rect 4062 3680 4068 3732
rect 4120 3720 4126 3732
rect 4801 3723 4859 3729
rect 4801 3720 4813 3723
rect 4120 3692 4813 3720
rect 4120 3680 4126 3692
rect 4801 3689 4813 3692
rect 4847 3689 4859 3723
rect 4801 3683 4859 3689
rect 4249 3587 4307 3593
rect 4249 3553 4261 3587
rect 4295 3584 4307 3587
rect 4706 3584 4712 3596
rect 4295 3556 4712 3584
rect 4295 3553 4307 3556
rect 4249 3547 4307 3553
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 4816 3584 4844 3683
rect 4890 3680 4896 3732
rect 4948 3720 4954 3732
rect 5169 3723 5227 3729
rect 5169 3720 5181 3723
rect 4948 3692 5181 3720
rect 4948 3680 4954 3692
rect 5169 3689 5181 3692
rect 5215 3689 5227 3723
rect 5169 3683 5227 3689
rect 7466 3680 7472 3732
rect 7524 3720 7530 3732
rect 7837 3723 7895 3729
rect 7837 3720 7849 3723
rect 7524 3692 7849 3720
rect 7524 3680 7530 3692
rect 7837 3689 7849 3692
rect 7883 3689 7895 3723
rect 7837 3683 7895 3689
rect 9030 3680 9036 3732
rect 9088 3720 9094 3732
rect 9217 3723 9275 3729
rect 9217 3720 9229 3723
rect 9088 3692 9229 3720
rect 9088 3680 9094 3692
rect 9217 3689 9229 3692
rect 9263 3689 9275 3723
rect 10502 3720 10508 3732
rect 10463 3692 10508 3720
rect 9217 3683 9275 3689
rect 10502 3680 10508 3692
rect 10560 3680 10566 3732
rect 10870 3720 10876 3732
rect 10831 3692 10876 3720
rect 10870 3680 10876 3692
rect 10928 3680 10934 3732
rect 13906 3680 13912 3732
rect 13964 3720 13970 3732
rect 14921 3723 14979 3729
rect 14921 3720 14933 3723
rect 13964 3692 14933 3720
rect 13964 3680 13970 3692
rect 14921 3689 14933 3692
rect 14967 3720 14979 3723
rect 15654 3720 15660 3732
rect 14967 3692 15660 3720
rect 14967 3689 14979 3692
rect 14921 3683 14979 3689
rect 15654 3680 15660 3692
rect 15712 3680 15718 3732
rect 15838 3720 15844 3732
rect 15799 3692 15844 3720
rect 15838 3680 15844 3692
rect 15896 3680 15902 3732
rect 16209 3723 16267 3729
rect 16209 3689 16221 3723
rect 16255 3720 16267 3723
rect 16298 3720 16304 3732
rect 16255 3692 16304 3720
rect 16255 3689 16267 3692
rect 16209 3683 16267 3689
rect 16298 3680 16304 3692
rect 16356 3680 16362 3732
rect 16850 3720 16856 3732
rect 16811 3692 16856 3720
rect 16850 3680 16856 3692
rect 16908 3680 16914 3732
rect 17494 3680 17500 3732
rect 17552 3720 17558 3732
rect 17867 3723 17925 3729
rect 17867 3720 17879 3723
rect 17552 3692 17879 3720
rect 17552 3680 17558 3692
rect 17867 3689 17879 3692
rect 17913 3689 17925 3723
rect 17867 3683 17925 3689
rect 19889 3723 19947 3729
rect 19889 3689 19901 3723
rect 19935 3720 19947 3723
rect 19978 3720 19984 3732
rect 19935 3692 19984 3720
rect 19935 3689 19947 3692
rect 19889 3683 19947 3689
rect 19978 3680 19984 3692
rect 20036 3680 20042 3732
rect 23290 3720 23296 3732
rect 23251 3692 23296 3720
rect 23290 3680 23296 3692
rect 23348 3680 23354 3732
rect 23658 3720 23664 3732
rect 23619 3692 23664 3720
rect 23658 3680 23664 3692
rect 23716 3680 23722 3732
rect 23937 3723 23995 3729
rect 23937 3689 23949 3723
rect 23983 3689 23995 3723
rect 24854 3720 24860 3732
rect 24815 3692 24860 3720
rect 23937 3683 23995 3689
rect 5534 3612 5540 3664
rect 5592 3661 5598 3664
rect 5592 3655 5656 3661
rect 5592 3621 5610 3655
rect 5644 3621 5656 3655
rect 5592 3615 5656 3621
rect 10413 3655 10471 3661
rect 10413 3621 10425 3655
rect 10459 3652 10471 3655
rect 10888 3652 10916 3680
rect 10459 3624 10916 3652
rect 10459 3621 10471 3624
rect 10413 3615 10471 3621
rect 5592 3612 5598 3615
rect 11882 3612 11888 3664
rect 11940 3652 11946 3664
rect 12590 3655 12648 3661
rect 12590 3652 12602 3655
rect 11940 3624 12602 3652
rect 11940 3612 11946 3624
rect 12590 3621 12602 3624
rect 12636 3621 12648 3655
rect 12590 3615 12648 3621
rect 14458 3612 14464 3664
rect 14516 3652 14522 3664
rect 14553 3655 14611 3661
rect 14553 3652 14565 3655
rect 14516 3624 14565 3652
rect 14516 3612 14522 3624
rect 14553 3621 14565 3624
rect 14599 3652 14611 3655
rect 15102 3652 15108 3664
rect 14599 3624 15108 3652
rect 14599 3621 14611 3624
rect 14553 3615 14611 3621
rect 15102 3612 15108 3624
rect 15160 3612 15166 3664
rect 19426 3612 19432 3664
rect 19484 3652 19490 3664
rect 20622 3652 20628 3664
rect 19484 3624 20628 3652
rect 19484 3612 19490 3624
rect 20622 3612 20628 3624
rect 20680 3612 20686 3664
rect 23952 3652 23980 3683
rect 24854 3680 24860 3692
rect 24912 3680 24918 3732
rect 25314 3720 25320 3732
rect 25275 3692 25320 3720
rect 25314 3680 25320 3692
rect 25372 3680 25378 3732
rect 25961 3723 26019 3729
rect 25961 3689 25973 3723
rect 26007 3720 26019 3723
rect 26326 3720 26332 3732
rect 26007 3692 26332 3720
rect 26007 3689 26019 3692
rect 25961 3683 26019 3689
rect 26326 3680 26332 3692
rect 26384 3720 26390 3732
rect 26881 3723 26939 3729
rect 26881 3720 26893 3723
rect 26384 3692 26893 3720
rect 26384 3680 26390 3692
rect 26881 3689 26893 3692
rect 26927 3689 26939 3723
rect 26881 3683 26939 3689
rect 26973 3723 27031 3729
rect 26973 3689 26985 3723
rect 27019 3720 27031 3723
rect 27062 3720 27068 3732
rect 27019 3692 27068 3720
rect 27019 3689 27031 3692
rect 26973 3683 27031 3689
rect 27062 3680 27068 3692
rect 27120 3720 27126 3732
rect 27522 3720 27528 3732
rect 27120 3692 27528 3720
rect 27120 3680 27126 3692
rect 27522 3680 27528 3692
rect 27580 3680 27586 3732
rect 29825 3723 29883 3729
rect 29825 3689 29837 3723
rect 29871 3720 29883 3723
rect 29914 3720 29920 3732
rect 29871 3692 29920 3720
rect 29871 3689 29883 3692
rect 29825 3683 29883 3689
rect 29914 3680 29920 3692
rect 29972 3720 29978 3732
rect 30377 3723 30435 3729
rect 30377 3720 30389 3723
rect 29972 3692 30389 3720
rect 29972 3680 29978 3692
rect 30377 3689 30389 3692
rect 30423 3689 30435 3723
rect 31478 3720 31484 3732
rect 31439 3692 31484 3720
rect 30377 3683 30435 3689
rect 31478 3680 31484 3692
rect 31536 3680 31542 3732
rect 34514 3680 34520 3732
rect 34572 3720 34578 3732
rect 35437 3723 35495 3729
rect 35437 3720 35449 3723
rect 34572 3692 35449 3720
rect 34572 3680 34578 3692
rect 35437 3689 35449 3692
rect 35483 3689 35495 3723
rect 35437 3683 35495 3689
rect 24946 3652 24952 3664
rect 23952 3624 24952 3652
rect 24946 3612 24952 3624
rect 25004 3612 25010 3664
rect 27617 3655 27675 3661
rect 27617 3652 27629 3655
rect 26252 3624 27629 3652
rect 5353 3587 5411 3593
rect 5353 3584 5365 3587
rect 4816 3556 5365 3584
rect 5353 3553 5365 3556
rect 5399 3584 5411 3587
rect 6178 3584 6184 3596
rect 5399 3556 6184 3584
rect 5399 3553 5411 3556
rect 5353 3547 5411 3553
rect 6178 3544 6184 3556
rect 6236 3544 6242 3596
rect 7745 3587 7803 3593
rect 7745 3553 7757 3587
rect 7791 3584 7803 3587
rect 8202 3584 8208 3596
rect 7791 3556 8208 3584
rect 7791 3553 7803 3556
rect 7745 3547 7803 3553
rect 8202 3544 8208 3556
rect 8260 3544 8266 3596
rect 10962 3544 10968 3596
rect 11020 3584 11026 3596
rect 16301 3587 16359 3593
rect 11020 3556 11065 3584
rect 11020 3544 11026 3556
rect 16301 3553 16313 3587
rect 16347 3584 16359 3587
rect 17221 3587 17279 3593
rect 17221 3584 17233 3587
rect 16347 3556 17233 3584
rect 16347 3553 16359 3556
rect 16301 3547 16359 3553
rect 17221 3553 17233 3556
rect 17267 3584 17279 3587
rect 17267 3556 19288 3584
rect 17267 3553 17279 3556
rect 17221 3547 17279 3553
rect 8110 3476 8116 3528
rect 8168 3516 8174 3528
rect 8297 3519 8355 3525
rect 8297 3516 8309 3519
rect 8168 3488 8309 3516
rect 8168 3476 8174 3488
rect 8297 3485 8309 3488
rect 8343 3485 8355 3519
rect 8297 3479 8355 3485
rect 8386 3476 8392 3528
rect 8444 3516 8450 3528
rect 8754 3516 8760 3528
rect 8444 3488 8760 3516
rect 8444 3476 8450 3488
rect 8754 3476 8760 3488
rect 8812 3516 8818 3528
rect 8849 3519 8907 3525
rect 8849 3516 8861 3519
rect 8812 3488 8861 3516
rect 8812 3476 8818 3488
rect 8849 3485 8861 3488
rect 8895 3485 8907 3519
rect 8849 3479 8907 3485
rect 11149 3519 11207 3525
rect 11149 3485 11161 3519
rect 11195 3516 11207 3519
rect 11238 3516 11244 3528
rect 11195 3488 11244 3516
rect 11195 3485 11207 3488
rect 11149 3479 11207 3485
rect 11238 3476 11244 3488
rect 11296 3516 11302 3528
rect 11517 3519 11575 3525
rect 11517 3516 11529 3519
rect 11296 3488 11529 3516
rect 11296 3476 11302 3488
rect 11517 3485 11529 3488
rect 11563 3516 11575 3519
rect 11885 3519 11943 3525
rect 11885 3516 11897 3519
rect 11563 3488 11897 3516
rect 11563 3485 11575 3488
rect 11517 3479 11575 3485
rect 11885 3485 11897 3488
rect 11931 3485 11943 3519
rect 12342 3516 12348 3528
rect 12303 3488 12348 3516
rect 11885 3479 11943 3485
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 16390 3516 16396 3528
rect 16351 3488 16396 3516
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 17405 3519 17463 3525
rect 17405 3485 17417 3519
rect 17451 3516 17463 3519
rect 17586 3516 17592 3528
rect 17451 3488 17592 3516
rect 17451 3485 17463 3488
rect 17405 3479 17463 3485
rect 17586 3476 17592 3488
rect 17644 3476 17650 3528
rect 17862 3516 17868 3528
rect 17823 3488 17868 3516
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 18138 3516 18144 3528
rect 18099 3488 18144 3516
rect 18138 3476 18144 3488
rect 18196 3476 18202 3528
rect 19260 3525 19288 3556
rect 20806 3544 20812 3596
rect 20864 3584 20870 3596
rect 21249 3587 21307 3593
rect 21249 3584 21261 3587
rect 20864 3556 21261 3584
rect 20864 3544 20870 3556
rect 21249 3553 21261 3556
rect 21295 3584 21307 3587
rect 21542 3584 21548 3596
rect 21295 3556 21548 3584
rect 21295 3553 21307 3556
rect 21249 3547 21307 3553
rect 21542 3544 21548 3556
rect 21600 3544 21606 3596
rect 23750 3584 23756 3596
rect 23711 3556 23756 3584
rect 23750 3544 23756 3556
rect 23808 3544 23814 3596
rect 25222 3584 25228 3596
rect 25183 3556 25228 3584
rect 25222 3544 25228 3556
rect 25280 3584 25286 3596
rect 26252 3584 26280 3624
rect 27617 3621 27629 3624
rect 27663 3621 27675 3655
rect 27617 3615 27675 3621
rect 34606 3612 34612 3664
rect 34664 3652 34670 3664
rect 35345 3655 35403 3661
rect 35345 3652 35357 3655
rect 34664 3624 35357 3652
rect 34664 3612 34670 3624
rect 35345 3621 35357 3624
rect 35391 3652 35403 3655
rect 35897 3655 35955 3661
rect 35897 3652 35909 3655
rect 35391 3624 35909 3652
rect 35391 3621 35403 3624
rect 35345 3615 35403 3621
rect 35897 3621 35909 3624
rect 35943 3621 35955 3655
rect 35897 3615 35955 3621
rect 25280 3556 26280 3584
rect 26329 3587 26387 3593
rect 25280 3544 25286 3556
rect 26329 3553 26341 3587
rect 26375 3584 26387 3587
rect 27062 3584 27068 3596
rect 26375 3556 27068 3584
rect 26375 3553 26387 3556
rect 26329 3547 26387 3553
rect 27062 3544 27068 3556
rect 27120 3544 27126 3596
rect 28166 3544 28172 3596
rect 28224 3584 28230 3596
rect 28701 3587 28759 3593
rect 28701 3584 28713 3587
rect 28224 3556 28713 3584
rect 28224 3544 28230 3556
rect 28701 3553 28713 3556
rect 28747 3553 28759 3587
rect 28701 3547 28759 3553
rect 30929 3587 30987 3593
rect 30929 3553 30941 3587
rect 30975 3584 30987 3587
rect 31294 3584 31300 3596
rect 30975 3556 31300 3584
rect 30975 3553 30987 3556
rect 30929 3547 30987 3553
rect 31294 3544 31300 3556
rect 31352 3544 31358 3596
rect 32306 3544 32312 3596
rect 32364 3584 32370 3596
rect 33226 3584 33232 3596
rect 32364 3556 33232 3584
rect 32364 3544 32370 3556
rect 33226 3544 33232 3556
rect 33284 3544 33290 3596
rect 34790 3544 34796 3596
rect 34848 3584 34854 3596
rect 35805 3587 35863 3593
rect 35805 3584 35817 3587
rect 34848 3556 35817 3584
rect 34848 3544 34854 3556
rect 35805 3553 35817 3556
rect 35851 3553 35863 3587
rect 35805 3547 35863 3553
rect 19245 3519 19303 3525
rect 19245 3485 19257 3519
rect 19291 3516 19303 3519
rect 19978 3516 19984 3528
rect 19291 3488 19984 3516
rect 19291 3485 19303 3488
rect 19245 3479 19303 3485
rect 19978 3476 19984 3488
rect 20036 3476 20042 3528
rect 20990 3516 20996 3528
rect 20951 3488 20996 3516
rect 20990 3476 20996 3488
rect 21048 3476 21054 3528
rect 25501 3519 25559 3525
rect 25501 3485 25513 3519
rect 25547 3516 25559 3519
rect 25590 3516 25596 3528
rect 25547 3488 25596 3516
rect 25547 3485 25559 3488
rect 25501 3479 25559 3485
rect 25590 3476 25596 3488
rect 25648 3476 25654 3528
rect 26142 3476 26148 3528
rect 26200 3516 26206 3528
rect 27157 3519 27215 3525
rect 27157 3516 27169 3519
rect 26200 3488 27169 3516
rect 26200 3476 26206 3488
rect 27157 3485 27169 3488
rect 27203 3516 27215 3519
rect 27893 3519 27951 3525
rect 27893 3516 27905 3519
rect 27203 3488 27905 3516
rect 27203 3485 27215 3488
rect 27157 3479 27215 3485
rect 27893 3485 27905 3488
rect 27939 3485 27951 3519
rect 28442 3516 28448 3528
rect 28403 3488 28448 3516
rect 27893 3479 27951 3485
rect 28442 3476 28448 3488
rect 28500 3476 28506 3528
rect 32490 3516 32496 3528
rect 32451 3488 32496 3516
rect 32490 3476 32496 3488
rect 32548 3476 32554 3528
rect 32674 3476 32680 3528
rect 32732 3516 32738 3528
rect 32816 3519 32874 3525
rect 32816 3516 32828 3519
rect 32732 3488 32828 3516
rect 32732 3476 32738 3488
rect 32816 3485 32828 3488
rect 32862 3485 32874 3519
rect 32816 3479 32874 3485
rect 32953 3519 33011 3525
rect 32953 3485 32965 3519
rect 32999 3516 33011 3519
rect 33042 3516 33048 3528
rect 32999 3488 33048 3516
rect 32999 3485 33011 3488
rect 32953 3479 33011 3485
rect 33042 3476 33048 3488
rect 33100 3476 33106 3528
rect 35989 3519 36047 3525
rect 35989 3485 36001 3519
rect 36035 3516 36047 3519
rect 36814 3516 36820 3528
rect 36035 3488 36820 3516
rect 36035 3485 36047 3488
rect 35989 3479 36047 3485
rect 4433 3451 4491 3457
rect 4433 3417 4445 3451
rect 4479 3448 4491 3451
rect 4479 3420 5396 3448
rect 4479 3417 4491 3420
rect 4433 3411 4491 3417
rect 2774 3340 2780 3392
rect 2832 3380 2838 3392
rect 3789 3383 3847 3389
rect 3789 3380 3801 3383
rect 2832 3352 3801 3380
rect 2832 3340 2838 3352
rect 3789 3349 3801 3352
rect 3835 3380 3847 3383
rect 4614 3380 4620 3392
rect 3835 3352 4620 3380
rect 3835 3349 3847 3352
rect 3789 3343 3847 3349
rect 4614 3340 4620 3352
rect 4672 3340 4678 3392
rect 5368 3380 5396 3420
rect 19334 3408 19340 3460
rect 19392 3448 19398 3460
rect 20165 3451 20223 3457
rect 20165 3448 20177 3451
rect 19392 3420 20177 3448
rect 19392 3408 19398 3420
rect 20165 3417 20177 3420
rect 20211 3417 20223 3451
rect 20165 3411 20223 3417
rect 20717 3451 20775 3457
rect 20717 3417 20729 3451
rect 20763 3448 20775 3451
rect 21008 3448 21036 3476
rect 20763 3420 21036 3448
rect 30837 3451 30895 3457
rect 20763 3417 20775 3420
rect 20717 3411 20775 3417
rect 30837 3417 30849 3451
rect 30883 3448 30895 3451
rect 31202 3448 31208 3460
rect 30883 3420 31208 3448
rect 30883 3417 30895 3420
rect 30837 3411 30895 3417
rect 31202 3408 31208 3420
rect 31260 3448 31266 3460
rect 31941 3451 31999 3457
rect 31941 3448 31953 3451
rect 31260 3420 31953 3448
rect 31260 3408 31266 3420
rect 31941 3417 31953 3420
rect 31987 3448 31999 3451
rect 32398 3448 32404 3460
rect 31987 3420 32404 3448
rect 31987 3417 31999 3420
rect 31941 3411 31999 3417
rect 32398 3408 32404 3420
rect 32456 3408 32462 3460
rect 34977 3451 35035 3457
rect 34977 3417 34989 3451
rect 35023 3448 35035 3451
rect 35434 3448 35440 3460
rect 35023 3420 35440 3448
rect 35023 3417 35035 3420
rect 34977 3411 35035 3417
rect 35434 3408 35440 3420
rect 35492 3448 35498 3460
rect 35492 3420 35664 3448
rect 35492 3408 35498 3420
rect 6086 3380 6092 3392
rect 5368 3352 6092 3380
rect 6086 3340 6092 3352
rect 6144 3340 6150 3392
rect 6730 3380 6736 3392
rect 6691 3352 6736 3380
rect 6730 3340 6736 3352
rect 6788 3380 6794 3392
rect 7285 3383 7343 3389
rect 7285 3380 7297 3383
rect 6788 3352 7297 3380
rect 6788 3340 6794 3352
rect 7285 3349 7297 3352
rect 7331 3349 7343 3383
rect 9950 3380 9956 3392
rect 9911 3352 9956 3380
rect 7285 3343 7343 3349
rect 9950 3340 9956 3352
rect 10008 3340 10014 3392
rect 13722 3380 13728 3392
rect 13683 3352 13728 3380
rect 13722 3340 13728 3352
rect 13780 3380 13786 3392
rect 14182 3380 14188 3392
rect 13780 3352 14188 3380
rect 13780 3340 13786 3352
rect 14182 3340 14188 3352
rect 14240 3340 14246 3392
rect 15565 3383 15623 3389
rect 15565 3349 15577 3383
rect 15611 3380 15623 3383
rect 15746 3380 15752 3392
rect 15611 3352 15752 3380
rect 15611 3349 15623 3352
rect 15565 3343 15623 3349
rect 15746 3340 15752 3352
rect 15804 3340 15810 3392
rect 22094 3340 22100 3392
rect 22152 3380 22158 3392
rect 22373 3383 22431 3389
rect 22373 3380 22385 3383
rect 22152 3352 22385 3380
rect 22152 3340 22158 3352
rect 22373 3349 22385 3352
rect 22419 3380 22431 3383
rect 23382 3380 23388 3392
rect 22419 3352 23388 3380
rect 22419 3349 22431 3352
rect 22373 3343 22431 3349
rect 23382 3340 23388 3352
rect 23440 3340 23446 3392
rect 24394 3380 24400 3392
rect 24355 3352 24400 3380
rect 24394 3340 24400 3352
rect 24452 3340 24458 3392
rect 24762 3380 24768 3392
rect 24723 3352 24768 3380
rect 24762 3340 24768 3352
rect 24820 3340 24826 3392
rect 26513 3383 26571 3389
rect 26513 3349 26525 3383
rect 26559 3380 26571 3383
rect 27154 3380 27160 3392
rect 26559 3352 27160 3380
rect 26559 3349 26571 3352
rect 26513 3343 26571 3349
rect 27154 3340 27160 3352
rect 27212 3340 27218 3392
rect 28258 3380 28264 3392
rect 28219 3352 28264 3380
rect 28258 3340 28264 3352
rect 28316 3340 28322 3392
rect 31113 3383 31171 3389
rect 31113 3349 31125 3383
rect 31159 3380 31171 3383
rect 31846 3380 31852 3392
rect 31159 3352 31852 3380
rect 31159 3349 31171 3352
rect 31113 3343 31171 3349
rect 31846 3340 31852 3352
rect 31904 3340 31910 3392
rect 32306 3380 32312 3392
rect 32267 3352 32312 3380
rect 32306 3340 32312 3352
rect 32364 3340 32370 3392
rect 34330 3380 34336 3392
rect 34291 3352 34336 3380
rect 34330 3340 34336 3352
rect 34388 3340 34394 3392
rect 35636 3380 35664 3420
rect 35710 3408 35716 3460
rect 35768 3448 35774 3460
rect 36004 3448 36032 3479
rect 36814 3476 36820 3488
rect 36872 3476 36878 3528
rect 35768 3420 36032 3448
rect 35768 3408 35774 3420
rect 36538 3380 36544 3392
rect 35636 3352 36544 3380
rect 36538 3340 36544 3352
rect 36596 3340 36602 3392
rect 1104 3290 38824 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 38824 3290
rect 1104 3216 38824 3238
rect 2038 3176 2044 3188
rect 1999 3148 2044 3176
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 3786 3176 3792 3188
rect 3747 3148 3792 3176
rect 3786 3136 3792 3148
rect 3844 3136 3850 3188
rect 6178 3176 6184 3188
rect 6139 3148 6184 3176
rect 6178 3136 6184 3148
rect 6236 3176 6242 3188
rect 6549 3179 6607 3185
rect 6549 3176 6561 3179
rect 6236 3148 6561 3176
rect 6236 3136 6242 3148
rect 6549 3145 6561 3148
rect 6595 3145 6607 3179
rect 6549 3139 6607 3145
rect 3329 3111 3387 3117
rect 3329 3077 3341 3111
rect 3375 3108 3387 3111
rect 3878 3108 3884 3120
rect 3375 3080 3884 3108
rect 3375 3077 3387 3080
rect 3329 3071 3387 3077
rect 3878 3068 3884 3080
rect 3936 3068 3942 3120
rect 4154 3108 4160 3120
rect 4115 3080 4160 3108
rect 4154 3068 4160 3080
rect 4212 3068 4218 3120
rect 4062 3000 4068 3052
rect 4120 3040 4126 3052
rect 4249 3043 4307 3049
rect 4249 3040 4261 3043
rect 4120 3012 4261 3040
rect 4120 3000 4126 3012
rect 4249 3009 4261 3012
rect 4295 3009 4307 3043
rect 6564 3040 6592 3139
rect 8110 3136 8116 3188
rect 8168 3176 8174 3188
rect 8205 3179 8263 3185
rect 8205 3176 8217 3179
rect 8168 3148 8217 3176
rect 8168 3136 8174 3148
rect 8205 3145 8217 3148
rect 8251 3176 8263 3179
rect 8386 3176 8392 3188
rect 8251 3148 8392 3176
rect 8251 3145 8263 3148
rect 8205 3139 8263 3145
rect 8386 3136 8392 3148
rect 8444 3176 8450 3188
rect 8757 3179 8815 3185
rect 8757 3176 8769 3179
rect 8444 3148 8769 3176
rect 8444 3136 8450 3148
rect 8757 3145 8769 3148
rect 8803 3176 8815 3179
rect 8846 3176 8852 3188
rect 8803 3148 8852 3176
rect 8803 3145 8815 3148
rect 8757 3139 8815 3145
rect 8846 3136 8852 3148
rect 8904 3136 8910 3188
rect 9401 3179 9459 3185
rect 9401 3145 9413 3179
rect 9447 3176 9459 3179
rect 10962 3176 10968 3188
rect 9447 3148 10968 3176
rect 9447 3145 9459 3148
rect 9401 3139 9459 3145
rect 10962 3136 10968 3148
rect 11020 3136 11026 3188
rect 11238 3176 11244 3188
rect 11199 3148 11244 3176
rect 11238 3136 11244 3148
rect 11296 3136 11302 3188
rect 11882 3176 11888 3188
rect 11843 3148 11888 3176
rect 11882 3136 11888 3148
rect 11940 3136 11946 3188
rect 15746 3136 15752 3188
rect 15804 3176 15810 3188
rect 16393 3179 16451 3185
rect 16393 3176 16405 3179
rect 15804 3148 16405 3176
rect 15804 3136 15810 3148
rect 16393 3145 16405 3148
rect 16439 3176 16451 3179
rect 17034 3176 17040 3188
rect 16439 3148 17040 3176
rect 16439 3145 16451 3148
rect 16393 3139 16451 3145
rect 17034 3136 17040 3148
rect 17092 3136 17098 3188
rect 17494 3176 17500 3188
rect 17455 3148 17500 3176
rect 17494 3136 17500 3148
rect 17552 3136 17558 3188
rect 19978 3176 19984 3188
rect 19939 3148 19984 3176
rect 19978 3136 19984 3148
rect 20036 3136 20042 3188
rect 22830 3136 22836 3188
rect 22888 3176 22894 3188
rect 23293 3179 23351 3185
rect 23293 3176 23305 3179
rect 22888 3148 23305 3176
rect 22888 3136 22894 3148
rect 23293 3145 23305 3148
rect 23339 3145 23351 3179
rect 23293 3139 23351 3145
rect 24213 3179 24271 3185
rect 24213 3145 24225 3179
rect 24259 3176 24271 3179
rect 25222 3176 25228 3188
rect 24259 3148 25228 3176
rect 24259 3145 24271 3148
rect 24213 3139 24271 3145
rect 25222 3136 25228 3148
rect 25280 3136 25286 3188
rect 25498 3136 25504 3188
rect 25556 3176 25562 3188
rect 25593 3179 25651 3185
rect 25593 3176 25605 3179
rect 25556 3148 25605 3176
rect 25556 3136 25562 3148
rect 25593 3145 25605 3148
rect 25639 3145 25651 3179
rect 27154 3176 27160 3188
rect 27115 3148 27160 3176
rect 25593 3139 25651 3145
rect 6638 3040 6644 3052
rect 6551 3012 6644 3040
rect 4249 3003 4307 3009
rect 6638 3000 6644 3012
rect 6696 3040 6702 3052
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 6696 3012 6837 3040
rect 6696 3000 6702 3012
rect 6825 3009 6837 3012
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 12342 3040 12348 3052
rect 11112 3012 12348 3040
rect 11112 3000 11118 3012
rect 12342 3000 12348 3012
rect 12400 3040 12406 3052
rect 12621 3043 12679 3049
rect 12621 3040 12633 3043
rect 12400 3012 12633 3040
rect 12400 3000 12406 3012
rect 12621 3009 12633 3012
rect 12667 3009 12679 3043
rect 13446 3040 13452 3052
rect 13407 3012 13452 3040
rect 12621 3003 12679 3009
rect 13446 3000 13452 3012
rect 13504 3000 13510 3052
rect 13633 3043 13691 3049
rect 13633 3009 13645 3043
rect 13679 3040 13691 3043
rect 13906 3040 13912 3052
rect 13679 3012 13912 3040
rect 13679 3009 13691 3012
rect 13633 3003 13691 3009
rect 13906 3000 13912 3012
rect 13964 3000 13970 3052
rect 14093 3043 14151 3049
rect 14093 3009 14105 3043
rect 14139 3040 14151 3043
rect 15013 3043 15071 3049
rect 14139 3012 14964 3040
rect 14139 3009 14151 3012
rect 14093 3003 14151 3009
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2972 1455 2975
rect 2038 2972 2044 2984
rect 1443 2944 2044 2972
rect 1443 2941 1455 2944
rect 1397 2935 1455 2941
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 3145 2975 3203 2981
rect 3145 2941 3157 2975
rect 3191 2972 3203 2975
rect 3786 2972 3792 2984
rect 3191 2944 3792 2972
rect 3191 2941 3203 2944
rect 3145 2935 3203 2941
rect 3786 2932 3792 2944
rect 3844 2932 3850 2984
rect 4516 2975 4574 2981
rect 4516 2941 4528 2975
rect 4562 2972 4574 2975
rect 4890 2972 4896 2984
rect 4562 2944 4896 2972
rect 4562 2941 4574 2944
rect 4516 2935 4574 2941
rect 4890 2932 4896 2944
rect 4948 2932 4954 2984
rect 9766 2972 9772 2984
rect 9679 2944 9772 2972
rect 9766 2932 9772 2944
rect 9824 2972 9830 2984
rect 9861 2975 9919 2981
rect 9861 2972 9873 2975
rect 9824 2944 9873 2972
rect 9824 2932 9830 2944
rect 9861 2941 9873 2944
rect 9907 2972 9919 2975
rect 11072 2972 11100 3000
rect 9907 2944 11100 2972
rect 12253 2975 12311 2981
rect 9907 2941 9919 2944
rect 9861 2935 9919 2941
rect 12253 2941 12265 2975
rect 12299 2972 12311 2975
rect 13262 2972 13268 2984
rect 12299 2944 13268 2972
rect 12299 2941 12311 2944
rect 12253 2935 12311 2941
rect 13262 2932 13268 2944
rect 13320 2972 13326 2984
rect 13357 2975 13415 2981
rect 13357 2972 13369 2975
rect 13320 2944 13369 2972
rect 13320 2932 13326 2944
rect 13357 2941 13369 2944
rect 13403 2941 13415 2975
rect 13357 2935 13415 2941
rect 14553 2975 14611 2981
rect 14553 2941 14565 2975
rect 14599 2972 14611 2975
rect 14826 2972 14832 2984
rect 14599 2944 14832 2972
rect 14599 2941 14611 2944
rect 14553 2935 14611 2941
rect 14826 2932 14832 2944
rect 14884 2932 14890 2984
rect 14936 2972 14964 3012
rect 15013 3009 15025 3043
rect 15059 3040 15071 3043
rect 15102 3040 15108 3052
rect 15059 3012 15108 3040
rect 15059 3009 15071 3012
rect 15013 3003 15071 3009
rect 15102 3000 15108 3012
rect 15160 3000 15166 3052
rect 19996 3040 20024 3136
rect 24578 3068 24584 3120
rect 24636 3108 24642 3120
rect 24636 3080 24808 3108
rect 24636 3068 24642 3080
rect 19996 3012 20668 3040
rect 15289 2975 15347 2981
rect 15289 2972 15301 2975
rect 14936 2944 15301 2972
rect 15289 2941 15301 2944
rect 15335 2972 15347 2975
rect 15562 2972 15568 2984
rect 15335 2944 15568 2972
rect 15335 2941 15347 2944
rect 15289 2935 15347 2941
rect 15562 2932 15568 2944
rect 15620 2932 15626 2984
rect 17865 2975 17923 2981
rect 17865 2941 17877 2975
rect 17911 2972 17923 2975
rect 18046 2972 18052 2984
rect 17911 2944 18052 2972
rect 17911 2941 17923 2944
rect 17865 2935 17923 2941
rect 18046 2932 18052 2944
rect 18104 2932 18110 2984
rect 20438 2932 20444 2984
rect 20496 2972 20502 2984
rect 20533 2975 20591 2981
rect 20533 2972 20545 2975
rect 20496 2944 20545 2972
rect 20496 2932 20502 2944
rect 20533 2941 20545 2944
rect 20579 2941 20591 2975
rect 20640 2972 20668 3012
rect 20714 3000 20720 3052
rect 20772 3040 20778 3052
rect 20993 3043 21051 3049
rect 20993 3040 21005 3043
rect 20772 3012 21005 3040
rect 20772 3000 20778 3012
rect 20993 3009 21005 3012
rect 21039 3040 21051 3043
rect 21450 3040 21456 3052
rect 21039 3012 21456 3040
rect 21039 3009 21051 3012
rect 20993 3003 21051 3009
rect 21450 3000 21456 3012
rect 21508 3000 21514 3052
rect 24394 3000 24400 3052
rect 24452 3040 24458 3052
rect 24780 3049 24808 3080
rect 24673 3043 24731 3049
rect 24673 3040 24685 3043
rect 24452 3012 24685 3040
rect 24452 3000 24458 3012
rect 24673 3009 24685 3012
rect 24719 3009 24731 3043
rect 24673 3003 24731 3009
rect 24765 3043 24823 3049
rect 24765 3009 24777 3043
rect 24811 3009 24823 3043
rect 25608 3040 25636 3139
rect 27154 3136 27160 3148
rect 27212 3176 27218 3188
rect 27709 3179 27767 3185
rect 27709 3176 27721 3179
rect 27212 3148 27721 3176
rect 27212 3136 27218 3148
rect 27709 3145 27721 3148
rect 27755 3145 27767 3179
rect 27709 3139 27767 3145
rect 28442 3136 28448 3188
rect 28500 3176 28506 3188
rect 28537 3179 28595 3185
rect 28537 3176 28549 3179
rect 28500 3148 28549 3176
rect 28500 3136 28506 3148
rect 28537 3145 28549 3148
rect 28583 3176 28595 3179
rect 29089 3179 29147 3185
rect 29089 3176 29101 3179
rect 28583 3148 29101 3176
rect 28583 3145 28595 3148
rect 28537 3139 28595 3145
rect 29089 3145 29101 3148
rect 29135 3176 29147 3179
rect 29178 3176 29184 3188
rect 29135 3148 29184 3176
rect 29135 3145 29147 3148
rect 29089 3139 29147 3145
rect 29178 3136 29184 3148
rect 29236 3136 29242 3188
rect 30742 3176 30748 3188
rect 30703 3148 30748 3176
rect 30742 3136 30748 3148
rect 30800 3136 30806 3188
rect 31294 3176 31300 3188
rect 31255 3148 31300 3176
rect 31294 3136 31300 3148
rect 31352 3136 31358 3188
rect 32490 3176 32496 3188
rect 31864 3148 32496 3176
rect 25777 3043 25835 3049
rect 25777 3040 25789 3043
rect 25608 3012 25789 3040
rect 24765 3003 24823 3009
rect 25777 3009 25789 3012
rect 25823 3009 25835 3043
rect 29196 3040 29224 3136
rect 31864 3049 31892 3148
rect 32490 3136 32496 3148
rect 32548 3136 32554 3188
rect 33226 3136 33232 3188
rect 33284 3176 33290 3188
rect 34609 3179 34667 3185
rect 34609 3176 34621 3179
rect 33284 3148 34621 3176
rect 33284 3136 33290 3148
rect 34609 3145 34621 3148
rect 34655 3176 34667 3179
rect 34790 3176 34796 3188
rect 34655 3148 34796 3176
rect 34655 3145 34667 3148
rect 34609 3139 34667 3145
rect 34790 3136 34796 3148
rect 34848 3136 34854 3188
rect 35250 3176 35256 3188
rect 35211 3148 35256 3176
rect 35250 3136 35256 3148
rect 35308 3136 35314 3188
rect 36814 3176 36820 3188
rect 36775 3148 36820 3176
rect 36814 3136 36820 3148
rect 36872 3136 36878 3188
rect 37366 3176 37372 3188
rect 37327 3148 37372 3176
rect 37366 3136 37372 3148
rect 37424 3136 37430 3188
rect 33689 3111 33747 3117
rect 33689 3077 33701 3111
rect 33735 3108 33747 3111
rect 33962 3108 33968 3120
rect 33735 3080 33968 3108
rect 33735 3077 33747 3080
rect 33689 3071 33747 3077
rect 33962 3068 33968 3080
rect 34020 3068 34026 3120
rect 29365 3043 29423 3049
rect 29365 3040 29377 3043
rect 29196 3012 29377 3040
rect 25777 3003 25835 3009
rect 29365 3009 29377 3012
rect 29411 3009 29423 3043
rect 29365 3003 29423 3009
rect 31849 3043 31907 3049
rect 31849 3009 31861 3043
rect 31895 3009 31907 3043
rect 31849 3003 31907 3009
rect 32309 3043 32367 3049
rect 32309 3009 32321 3043
rect 32355 3009 32367 3043
rect 32309 3003 32367 3009
rect 21269 2975 21327 2981
rect 21269 2972 21281 2975
rect 20640 2944 21281 2972
rect 20533 2935 20591 2941
rect 21269 2941 21281 2944
rect 21315 2941 21327 2975
rect 24688 2972 24716 3003
rect 25225 2975 25283 2981
rect 25225 2972 25237 2975
rect 24688 2944 25237 2972
rect 21269 2935 21327 2941
rect 25225 2941 25237 2944
rect 25271 2941 25283 2975
rect 26970 2972 26976 2984
rect 25225 2935 25283 2941
rect 26068 2944 26976 2972
rect 5902 2864 5908 2916
rect 5960 2904 5966 2916
rect 6730 2904 6736 2916
rect 5960 2876 6736 2904
rect 5960 2864 5966 2876
rect 6730 2864 6736 2876
rect 6788 2904 6794 2916
rect 7070 2907 7128 2913
rect 7070 2904 7082 2907
rect 6788 2876 7082 2904
rect 6788 2864 6794 2876
rect 7070 2873 7082 2876
rect 7116 2873 7128 2907
rect 7070 2867 7128 2873
rect 9950 2864 9956 2916
rect 10008 2904 10014 2916
rect 10128 2907 10186 2913
rect 10128 2904 10140 2907
rect 10008 2876 10140 2904
rect 10008 2864 10014 2876
rect 10128 2873 10140 2876
rect 10174 2904 10186 2907
rect 10962 2904 10968 2916
rect 10174 2876 10968 2904
rect 10174 2873 10186 2876
rect 10128 2867 10186 2873
rect 10962 2864 10968 2876
rect 11020 2864 11026 2916
rect 18230 2864 18236 2916
rect 18288 2913 18294 2916
rect 18288 2907 18352 2913
rect 18288 2873 18306 2907
rect 18340 2873 18352 2907
rect 18288 2867 18352 2873
rect 18288 2864 18294 2867
rect 23750 2864 23756 2916
rect 23808 2904 23814 2916
rect 23937 2907 23995 2913
rect 23937 2904 23949 2907
rect 23808 2876 23949 2904
rect 23808 2864 23814 2876
rect 23937 2873 23949 2876
rect 23983 2904 23995 2907
rect 24581 2907 24639 2913
rect 23983 2876 24348 2904
rect 23983 2873 23995 2876
rect 23937 2867 23995 2873
rect 1581 2839 1639 2845
rect 1581 2805 1593 2839
rect 1627 2836 1639 2839
rect 1670 2836 1676 2848
rect 1627 2808 1676 2836
rect 1627 2805 1639 2808
rect 1581 2799 1639 2805
rect 1670 2796 1676 2808
rect 1728 2796 1734 2848
rect 5534 2796 5540 2848
rect 5592 2836 5598 2848
rect 5629 2839 5687 2845
rect 5629 2836 5641 2839
rect 5592 2808 5641 2836
rect 5592 2796 5598 2808
rect 5629 2805 5641 2808
rect 5675 2805 5687 2839
rect 12986 2836 12992 2848
rect 12947 2808 12992 2836
rect 5629 2799 5687 2805
rect 12986 2796 12992 2808
rect 13044 2796 13050 2848
rect 14461 2839 14519 2845
rect 14461 2805 14473 2839
rect 14507 2836 14519 2839
rect 14642 2836 14648 2848
rect 14507 2808 14648 2836
rect 14507 2805 14519 2808
rect 14461 2799 14519 2805
rect 14642 2796 14648 2808
rect 14700 2836 14706 2848
rect 15015 2839 15073 2845
rect 15015 2836 15027 2839
rect 14700 2808 15027 2836
rect 14700 2796 14706 2808
rect 15015 2805 15027 2808
rect 15061 2836 15073 2839
rect 17494 2836 17500 2848
rect 15061 2808 17500 2836
rect 15061 2805 15073 2808
rect 15015 2799 15073 2805
rect 17494 2796 17500 2808
rect 17552 2796 17558 2848
rect 19334 2796 19340 2848
rect 19392 2836 19398 2848
rect 19429 2839 19487 2845
rect 19429 2836 19441 2839
rect 19392 2808 19441 2836
rect 19392 2796 19398 2808
rect 19429 2805 19441 2808
rect 19475 2805 19487 2839
rect 19429 2799 19487 2805
rect 20070 2796 20076 2848
rect 20128 2836 20134 2848
rect 20441 2839 20499 2845
rect 20441 2836 20453 2839
rect 20128 2808 20453 2836
rect 20128 2796 20134 2808
rect 20441 2805 20453 2808
rect 20487 2836 20499 2839
rect 20995 2839 21053 2845
rect 20995 2836 21007 2839
rect 20487 2808 21007 2836
rect 20487 2805 20499 2808
rect 20441 2799 20499 2805
rect 20995 2805 21007 2808
rect 21041 2836 21053 2839
rect 21910 2836 21916 2848
rect 21041 2808 21916 2836
rect 21041 2805 21053 2808
rect 20995 2799 21053 2805
rect 21910 2796 21916 2808
rect 21968 2796 21974 2848
rect 22370 2836 22376 2848
rect 22331 2808 22376 2836
rect 22370 2796 22376 2808
rect 22428 2796 22434 2848
rect 23017 2839 23075 2845
rect 23017 2805 23029 2839
rect 23063 2836 23075 2839
rect 23382 2836 23388 2848
rect 23063 2808 23388 2836
rect 23063 2805 23075 2808
rect 23017 2799 23075 2805
rect 23382 2796 23388 2808
rect 23440 2796 23446 2848
rect 24320 2836 24348 2876
rect 24581 2873 24593 2907
rect 24627 2904 24639 2907
rect 24762 2904 24768 2916
rect 24627 2876 24768 2904
rect 24627 2873 24639 2876
rect 24581 2867 24639 2873
rect 24762 2864 24768 2876
rect 24820 2864 24826 2916
rect 25240 2904 25268 2935
rect 26068 2913 26096 2944
rect 26970 2932 26976 2944
rect 27028 2932 27034 2984
rect 29632 2975 29690 2981
rect 29632 2941 29644 2975
rect 29678 2972 29690 2975
rect 30006 2972 30012 2984
rect 29678 2944 30012 2972
rect 29678 2941 29690 2944
rect 29632 2935 29690 2941
rect 30006 2932 30012 2944
rect 30064 2932 30070 2984
rect 31938 2932 31944 2984
rect 31996 2972 32002 2984
rect 32324 2972 32352 3003
rect 32398 3000 32404 3052
rect 32456 3040 32462 3052
rect 32585 3043 32643 3049
rect 32585 3040 32597 3043
rect 32456 3012 32597 3040
rect 32456 3000 32462 3012
rect 32585 3009 32597 3012
rect 32631 3040 32643 3043
rect 34330 3040 34336 3052
rect 32631 3012 34336 3040
rect 32631 3009 32643 3012
rect 32585 3003 32643 3009
rect 34330 3000 34336 3012
rect 34388 3000 34394 3052
rect 35268 3040 35296 3136
rect 35437 3043 35495 3049
rect 35437 3040 35449 3043
rect 35268 3012 35449 3040
rect 35437 3009 35449 3012
rect 35483 3009 35495 3043
rect 35437 3003 35495 3009
rect 33042 2972 33048 2984
rect 31996 2944 33048 2972
rect 31996 2932 32002 2944
rect 33042 2932 33048 2944
rect 33100 2932 33106 2984
rect 35704 2975 35762 2981
rect 35704 2941 35716 2975
rect 35750 2972 35762 2975
rect 36538 2972 36544 2984
rect 35750 2944 36544 2972
rect 35750 2941 35762 2944
rect 35704 2935 35762 2941
rect 36538 2932 36544 2944
rect 36596 2932 36602 2984
rect 26022 2907 26096 2913
rect 26022 2904 26034 2907
rect 25240 2876 26034 2904
rect 26022 2873 26034 2876
rect 26068 2876 26096 2907
rect 26068 2873 26080 2876
rect 26022 2867 26080 2873
rect 24946 2836 24952 2848
rect 24320 2808 24952 2836
rect 24946 2796 24952 2808
rect 25004 2796 25010 2848
rect 28166 2836 28172 2848
rect 28127 2808 28172 2836
rect 28166 2796 28172 2808
rect 28224 2796 28230 2848
rect 31757 2839 31815 2845
rect 31757 2805 31769 2839
rect 31803 2836 31815 2839
rect 32311 2839 32369 2845
rect 32311 2836 32323 2839
rect 31803 2808 32323 2836
rect 31803 2805 31815 2808
rect 31757 2799 31815 2805
rect 32311 2805 32323 2808
rect 32357 2836 32369 2839
rect 32674 2836 32680 2848
rect 32357 2808 32680 2836
rect 32357 2805 32369 2808
rect 32311 2799 32369 2805
rect 32674 2796 32680 2808
rect 32732 2836 32738 2848
rect 34241 2839 34299 2845
rect 34241 2836 34253 2839
rect 32732 2808 34253 2836
rect 32732 2796 32738 2808
rect 34241 2805 34253 2808
rect 34287 2836 34299 2839
rect 34422 2836 34428 2848
rect 34287 2808 34428 2836
rect 34287 2805 34299 2808
rect 34241 2799 34299 2805
rect 34422 2796 34428 2808
rect 34480 2796 34486 2848
rect 1104 2746 38824 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 38824 2746
rect 1104 2672 38824 2694
rect 2409 2635 2467 2641
rect 2409 2601 2421 2635
rect 2455 2632 2467 2635
rect 2682 2632 2688 2644
rect 2455 2604 2688 2632
rect 2455 2601 2467 2604
rect 2409 2595 2467 2601
rect 2682 2592 2688 2604
rect 2740 2592 2746 2644
rect 3142 2632 3148 2644
rect 3103 2604 3148 2632
rect 3142 2592 3148 2604
rect 3200 2592 3206 2644
rect 4890 2592 4896 2644
rect 4948 2632 4954 2644
rect 5077 2635 5135 2641
rect 5077 2632 5089 2635
rect 4948 2604 5089 2632
rect 4948 2592 4954 2604
rect 5077 2601 5089 2604
rect 5123 2601 5135 2635
rect 5258 2632 5264 2644
rect 5219 2604 5264 2632
rect 5077 2595 5135 2601
rect 5258 2592 5264 2604
rect 5316 2592 5322 2644
rect 6638 2632 6644 2644
rect 6599 2604 6644 2632
rect 6638 2592 6644 2604
rect 6696 2592 6702 2644
rect 8202 2592 8208 2644
rect 8260 2632 8266 2644
rect 8573 2635 8631 2641
rect 8573 2632 8585 2635
rect 8260 2604 8585 2632
rect 8260 2592 8266 2604
rect 8573 2601 8585 2604
rect 8619 2601 8631 2635
rect 8573 2595 8631 2601
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2496 1455 2499
rect 2038 2496 2044 2508
rect 1443 2468 2044 2496
rect 1443 2465 1455 2468
rect 1397 2459 1455 2465
rect 2038 2456 2044 2468
rect 2096 2456 2102 2508
rect 2501 2499 2559 2505
rect 2501 2465 2513 2499
rect 2547 2496 2559 2499
rect 3160 2496 3188 2592
rect 3881 2567 3939 2573
rect 3881 2533 3893 2567
rect 3927 2564 3939 2567
rect 5534 2564 5540 2576
rect 3927 2536 5540 2564
rect 3927 2533 3939 2536
rect 3881 2527 3939 2533
rect 5534 2524 5540 2536
rect 5592 2564 5598 2576
rect 5721 2567 5779 2573
rect 5721 2564 5733 2567
rect 5592 2536 5733 2564
rect 5592 2524 5598 2536
rect 5721 2533 5733 2536
rect 5767 2564 5779 2567
rect 6273 2567 6331 2573
rect 6273 2564 6285 2567
rect 5767 2536 6285 2564
rect 5767 2533 5779 2536
rect 5721 2527 5779 2533
rect 6273 2533 6285 2536
rect 6319 2533 6331 2567
rect 6273 2527 6331 2533
rect 2547 2468 3188 2496
rect 4157 2499 4215 2505
rect 2547 2465 2559 2468
rect 2501 2459 2559 2465
rect 4157 2465 4169 2499
rect 4203 2496 4215 2499
rect 4798 2496 4804 2508
rect 4203 2468 4804 2496
rect 4203 2465 4215 2468
rect 4157 2459 4215 2465
rect 4798 2456 4804 2468
rect 4856 2456 4862 2508
rect 5629 2499 5687 2505
rect 5629 2465 5641 2499
rect 5675 2496 5687 2499
rect 5902 2496 5908 2508
rect 5675 2468 5908 2496
rect 5675 2465 5687 2468
rect 5629 2459 5687 2465
rect 3513 2431 3571 2437
rect 3513 2397 3525 2431
rect 3559 2428 3571 2431
rect 5644 2428 5672 2459
rect 5902 2456 5908 2468
rect 5960 2456 5966 2508
rect 6656 2496 6684 2592
rect 7460 2567 7518 2573
rect 7460 2533 7472 2567
rect 7506 2564 7518 2567
rect 8386 2564 8392 2576
rect 7506 2536 8392 2564
rect 7506 2533 7518 2536
rect 7460 2527 7518 2533
rect 8386 2524 8392 2536
rect 8444 2524 8450 2576
rect 8588 2564 8616 2595
rect 8846 2592 8852 2644
rect 8904 2632 8910 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 8904 2604 9137 2632
rect 8904 2592 8910 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 9125 2595 9183 2601
rect 11054 2592 11060 2644
rect 11112 2632 11118 2644
rect 11149 2635 11207 2641
rect 11149 2632 11161 2635
rect 11112 2604 11161 2632
rect 11112 2592 11118 2604
rect 11149 2601 11161 2604
rect 11195 2601 11207 2635
rect 12342 2632 12348 2644
rect 12303 2604 12348 2632
rect 11149 2595 11207 2601
rect 12342 2592 12348 2604
rect 12400 2592 12406 2644
rect 14274 2632 14280 2644
rect 14235 2604 14280 2632
rect 14274 2592 14280 2604
rect 14332 2632 14338 2644
rect 14829 2635 14887 2641
rect 14829 2632 14841 2635
rect 14332 2604 14841 2632
rect 14332 2592 14338 2604
rect 14829 2601 14841 2604
rect 14875 2601 14887 2635
rect 14829 2595 14887 2601
rect 10036 2567 10094 2573
rect 10036 2564 10048 2567
rect 8588 2536 10048 2564
rect 10036 2533 10048 2536
rect 10082 2564 10094 2567
rect 11701 2567 11759 2573
rect 11701 2564 11713 2567
rect 10082 2536 11713 2564
rect 10082 2533 10094 2536
rect 10036 2527 10094 2533
rect 11701 2533 11713 2536
rect 11747 2533 11759 2567
rect 11701 2527 11759 2533
rect 7193 2499 7251 2505
rect 7193 2496 7205 2499
rect 6656 2468 7205 2496
rect 7193 2465 7205 2468
rect 7239 2496 7251 2499
rect 9493 2499 9551 2505
rect 9493 2496 9505 2499
rect 7239 2468 9505 2496
rect 7239 2465 7251 2468
rect 7193 2459 7251 2465
rect 9493 2465 9505 2468
rect 9539 2496 9551 2499
rect 9766 2496 9772 2508
rect 9539 2468 9772 2496
rect 9539 2465 9551 2468
rect 9493 2459 9551 2465
rect 9766 2456 9772 2468
rect 9824 2456 9830 2508
rect 12360 2496 12388 2592
rect 13164 2567 13222 2573
rect 13164 2533 13176 2567
rect 13210 2564 13222 2567
rect 13722 2564 13728 2576
rect 13210 2536 13728 2564
rect 13210 2533 13222 2536
rect 13164 2527 13222 2533
rect 13722 2524 13728 2536
rect 13780 2524 13786 2576
rect 14844 2564 14872 2595
rect 16666 2592 16672 2644
rect 16724 2632 16730 2644
rect 16853 2635 16911 2641
rect 16853 2632 16865 2635
rect 16724 2604 16865 2632
rect 16724 2592 16730 2604
rect 16853 2601 16865 2604
rect 16899 2601 16911 2635
rect 17402 2632 17408 2644
rect 17363 2604 17408 2632
rect 16853 2595 16911 2601
rect 17402 2592 17408 2604
rect 17460 2592 17466 2644
rect 19981 2635 20039 2641
rect 19981 2601 19993 2635
rect 20027 2632 20039 2635
rect 20622 2632 20628 2644
rect 20027 2604 20628 2632
rect 20027 2601 20039 2604
rect 19981 2595 20039 2601
rect 20622 2592 20628 2604
rect 20680 2592 20686 2644
rect 22186 2592 22192 2644
rect 22244 2632 22250 2644
rect 22649 2635 22707 2641
rect 22649 2632 22661 2635
rect 22244 2604 22661 2632
rect 22244 2592 22250 2604
rect 22649 2601 22661 2604
rect 22695 2601 22707 2635
rect 22649 2595 22707 2601
rect 23845 2635 23903 2641
rect 23845 2601 23857 2635
rect 23891 2632 23903 2635
rect 24026 2632 24032 2644
rect 23891 2604 24032 2632
rect 23891 2601 23903 2604
rect 23845 2595 23903 2601
rect 24026 2592 24032 2604
rect 24084 2592 24090 2644
rect 24486 2632 24492 2644
rect 24447 2604 24492 2632
rect 24486 2592 24492 2604
rect 24544 2632 24550 2644
rect 25041 2635 25099 2641
rect 25041 2632 25053 2635
rect 24544 2604 25053 2632
rect 24544 2592 24550 2604
rect 25041 2601 25053 2604
rect 25087 2601 25099 2635
rect 25958 2632 25964 2644
rect 25919 2604 25964 2632
rect 25041 2595 25099 2601
rect 25958 2592 25964 2604
rect 26016 2592 26022 2644
rect 26510 2592 26516 2644
rect 26568 2632 26574 2644
rect 26605 2635 26663 2641
rect 26605 2632 26617 2635
rect 26568 2604 26617 2632
rect 26568 2592 26574 2604
rect 26605 2601 26617 2604
rect 26651 2601 26663 2635
rect 26605 2595 26663 2601
rect 15718 2567 15776 2573
rect 15718 2564 15730 2567
rect 14844 2536 15730 2564
rect 15718 2533 15730 2536
rect 15764 2533 15776 2567
rect 15718 2527 15776 2533
rect 18868 2567 18926 2573
rect 18868 2533 18880 2567
rect 18914 2564 18926 2567
rect 19242 2564 19248 2576
rect 18914 2536 19248 2564
rect 18914 2533 18926 2536
rect 18868 2527 18926 2533
rect 19242 2524 19248 2536
rect 19300 2524 19306 2576
rect 21536 2567 21594 2573
rect 21536 2533 21548 2567
rect 21582 2564 21594 2567
rect 22002 2564 22008 2576
rect 21582 2536 22008 2564
rect 21582 2533 21594 2536
rect 21536 2527 21594 2533
rect 22002 2524 22008 2536
rect 22060 2524 22066 2576
rect 24044 2564 24072 2592
rect 24397 2567 24455 2573
rect 24397 2564 24409 2567
rect 24044 2536 24409 2564
rect 24397 2533 24409 2536
rect 24443 2533 24455 2567
rect 24397 2527 24455 2533
rect 25593 2567 25651 2573
rect 25593 2533 25605 2567
rect 25639 2564 25651 2567
rect 26050 2564 26056 2576
rect 25639 2536 26056 2564
rect 25639 2533 25651 2536
rect 25593 2527 25651 2533
rect 26050 2524 26056 2536
rect 26108 2524 26114 2576
rect 12897 2499 12955 2505
rect 12897 2496 12909 2499
rect 12360 2468 12909 2496
rect 12897 2465 12909 2468
rect 12943 2496 12955 2499
rect 15197 2499 15255 2505
rect 15197 2496 15209 2499
rect 12943 2468 15209 2496
rect 12943 2465 12955 2468
rect 12897 2459 12955 2465
rect 15197 2465 15209 2468
rect 15243 2496 15255 2499
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 15243 2468 15485 2496
rect 15243 2465 15255 2468
rect 15197 2459 15255 2465
rect 15473 2465 15485 2468
rect 15519 2465 15531 2499
rect 15473 2459 15531 2465
rect 18046 2456 18052 2508
rect 18104 2496 18110 2508
rect 18141 2499 18199 2505
rect 18141 2496 18153 2499
rect 18104 2468 18153 2496
rect 18104 2456 18110 2468
rect 18141 2465 18153 2468
rect 18187 2496 18199 2499
rect 18601 2499 18659 2505
rect 18601 2496 18613 2499
rect 18187 2468 18613 2496
rect 18187 2465 18199 2468
rect 18141 2459 18199 2465
rect 18601 2465 18613 2468
rect 18647 2465 18659 2499
rect 20622 2496 20628 2508
rect 20583 2468 20628 2496
rect 18601 2459 18659 2465
rect 20622 2456 20628 2468
rect 20680 2456 20686 2508
rect 20990 2496 20996 2508
rect 20903 2468 20996 2496
rect 20990 2456 20996 2468
rect 21048 2496 21054 2508
rect 21269 2499 21327 2505
rect 21269 2496 21281 2499
rect 21048 2468 21281 2496
rect 21048 2456 21054 2468
rect 21269 2465 21281 2468
rect 21315 2465 21327 2499
rect 25774 2496 25780 2508
rect 25735 2468 25780 2496
rect 21269 2459 21327 2465
rect 25774 2456 25780 2468
rect 25832 2456 25838 2508
rect 26620 2496 26648 2595
rect 28166 2592 28172 2644
rect 28224 2632 28230 2644
rect 28261 2635 28319 2641
rect 28261 2632 28273 2635
rect 28224 2604 28273 2632
rect 28224 2592 28230 2604
rect 28261 2601 28273 2604
rect 28307 2601 28319 2635
rect 28261 2595 28319 2601
rect 29178 2592 29184 2644
rect 29236 2632 29242 2644
rect 29457 2635 29515 2641
rect 29457 2632 29469 2635
rect 29236 2604 29469 2632
rect 29236 2592 29242 2604
rect 29457 2601 29469 2604
rect 29503 2601 29515 2635
rect 31938 2632 31944 2644
rect 31899 2604 31944 2632
rect 29457 2595 29515 2601
rect 27154 2573 27160 2576
rect 27148 2564 27160 2573
rect 27115 2536 27160 2564
rect 27148 2527 27160 2536
rect 27154 2524 27160 2527
rect 27212 2524 27218 2576
rect 26881 2499 26939 2505
rect 26881 2496 26893 2499
rect 26620 2468 26893 2496
rect 26881 2465 26893 2468
rect 26927 2465 26939 2499
rect 29472 2496 29500 2595
rect 31938 2592 31944 2604
rect 31996 2592 32002 2644
rect 32122 2592 32128 2644
rect 32180 2632 32186 2644
rect 32309 2635 32367 2641
rect 32309 2632 32321 2635
rect 32180 2604 32321 2632
rect 32180 2592 32186 2604
rect 32309 2601 32321 2604
rect 32355 2601 32367 2635
rect 34238 2632 34244 2644
rect 34199 2604 34244 2632
rect 32309 2595 32367 2601
rect 29914 2524 29920 2576
rect 29972 2564 29978 2576
rect 30070 2567 30128 2573
rect 30070 2564 30082 2567
rect 29972 2536 30082 2564
rect 29972 2524 29978 2536
rect 30070 2533 30082 2536
rect 30116 2533 30128 2567
rect 30070 2527 30128 2533
rect 29825 2499 29883 2505
rect 29825 2496 29837 2499
rect 29472 2468 29837 2496
rect 26881 2459 26939 2465
rect 29825 2465 29837 2468
rect 29871 2465 29883 2499
rect 32324 2496 32352 2595
rect 34238 2592 34244 2604
rect 34296 2632 34302 2644
rect 34296 2604 35848 2632
rect 34296 2592 34302 2604
rect 33128 2567 33186 2573
rect 33128 2533 33140 2567
rect 33174 2564 33186 2567
rect 33686 2564 33692 2576
rect 33174 2536 33692 2564
rect 33174 2533 33186 2536
rect 33128 2527 33186 2533
rect 33686 2524 33692 2536
rect 33744 2564 33750 2576
rect 34793 2567 34851 2573
rect 34793 2564 34805 2567
rect 33744 2536 34805 2564
rect 33744 2524 33750 2536
rect 34793 2533 34805 2536
rect 34839 2533 34851 2567
rect 34793 2527 34851 2533
rect 35704 2567 35762 2573
rect 35704 2533 35716 2567
rect 35750 2564 35762 2567
rect 35820 2564 35848 2604
rect 36538 2592 36544 2644
rect 36596 2632 36602 2644
rect 36817 2635 36875 2641
rect 36817 2632 36829 2635
rect 36596 2604 36829 2632
rect 36596 2592 36602 2604
rect 36817 2601 36829 2604
rect 36863 2601 36875 2635
rect 36817 2595 36875 2601
rect 37369 2567 37427 2573
rect 37369 2564 37381 2567
rect 35750 2536 37381 2564
rect 35750 2533 35762 2536
rect 35704 2527 35762 2533
rect 37369 2533 37381 2536
rect 37415 2533 37427 2567
rect 37369 2527 37427 2533
rect 32861 2499 32919 2505
rect 32861 2496 32873 2499
rect 32324 2468 32873 2496
rect 29825 2459 29883 2465
rect 32861 2465 32873 2468
rect 32907 2496 32919 2499
rect 35161 2499 35219 2505
rect 35161 2496 35173 2499
rect 32907 2468 35173 2496
rect 32907 2465 32919 2468
rect 32861 2459 32919 2465
rect 35161 2465 35173 2468
rect 35207 2496 35219 2499
rect 35250 2496 35256 2508
rect 35207 2468 35256 2496
rect 35207 2465 35219 2468
rect 35161 2459 35219 2465
rect 35250 2456 35256 2468
rect 35308 2496 35314 2508
rect 35437 2499 35495 2505
rect 35437 2496 35449 2499
rect 35308 2468 35449 2496
rect 35308 2456 35314 2468
rect 35437 2465 35449 2468
rect 35483 2465 35495 2499
rect 35437 2459 35495 2465
rect 5810 2428 5816 2440
rect 3559 2400 5672 2428
rect 5771 2400 5816 2428
rect 3559 2397 3571 2400
rect 3513 2391 3571 2397
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 23382 2388 23388 2440
rect 23440 2428 23446 2440
rect 23477 2431 23535 2437
rect 23477 2428 23489 2431
rect 23440 2400 23489 2428
rect 23440 2388 23446 2400
rect 23477 2397 23489 2400
rect 23523 2428 23535 2431
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 23523 2400 24593 2428
rect 23523 2397 23535 2400
rect 23477 2391 23535 2397
rect 24581 2397 24593 2400
rect 24627 2397 24639 2431
rect 24581 2391 24639 2397
rect 25501 2431 25559 2437
rect 25501 2397 25513 2431
rect 25547 2428 25559 2431
rect 25792 2428 25820 2456
rect 25547 2400 25820 2428
rect 25547 2397 25559 2400
rect 25501 2391 25559 2397
rect 4341 2363 4399 2369
rect 4341 2329 4353 2363
rect 4387 2360 4399 2363
rect 4982 2360 4988 2372
rect 4387 2332 4988 2360
rect 4387 2329 4399 2332
rect 4341 2323 4399 2329
rect 4982 2320 4988 2332
rect 5040 2320 5046 2372
rect 29181 2363 29239 2369
rect 29181 2329 29193 2363
rect 29227 2360 29239 2363
rect 29227 2332 29868 2360
rect 29227 2329 29239 2332
rect 29181 2323 29239 2329
rect 566 2252 572 2304
rect 624 2292 630 2304
rect 1581 2295 1639 2301
rect 1581 2292 1593 2295
rect 624 2264 1593 2292
rect 624 2252 630 2264
rect 1581 2261 1593 2264
rect 1627 2261 1639 2295
rect 1581 2255 1639 2261
rect 2685 2295 2743 2301
rect 2685 2261 2697 2295
rect 2731 2292 2743 2295
rect 2774 2292 2780 2304
rect 2731 2264 2780 2292
rect 2731 2261 2743 2264
rect 2685 2255 2743 2261
rect 2774 2252 2780 2264
rect 2832 2252 2838 2304
rect 4798 2292 4804 2304
rect 4759 2264 4804 2292
rect 4798 2252 4804 2264
rect 4856 2252 4862 2304
rect 24026 2292 24032 2304
rect 23987 2264 24032 2292
rect 24026 2252 24032 2264
rect 24084 2252 24090 2304
rect 26050 2252 26056 2304
rect 26108 2292 26114 2304
rect 26237 2295 26295 2301
rect 26237 2292 26249 2295
rect 26108 2264 26249 2292
rect 26108 2252 26114 2264
rect 26237 2261 26249 2264
rect 26283 2261 26295 2295
rect 29840 2292 29868 2332
rect 30006 2292 30012 2304
rect 29840 2264 30012 2292
rect 26237 2255 26295 2261
rect 30006 2252 30012 2264
rect 30064 2292 30070 2304
rect 31205 2295 31263 2301
rect 31205 2292 31217 2295
rect 30064 2264 31217 2292
rect 30064 2252 30070 2264
rect 31205 2261 31217 2264
rect 31251 2261 31263 2295
rect 31205 2255 31263 2261
rect 1104 2202 38824 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 35624 36363 35676 36372
rect 35624 36329 35633 36363
rect 35633 36329 35667 36363
rect 35667 36329 35676 36363
rect 35624 36320 35676 36329
rect 35808 36184 35860 36236
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 35716 35776 35768 35828
rect 33048 35479 33100 35488
rect 33048 35445 33057 35479
rect 33057 35445 33091 35479
rect 33091 35445 33100 35479
rect 33048 35436 33100 35445
rect 33416 35479 33468 35488
rect 33416 35445 33425 35479
rect 33425 35445 33459 35479
rect 33459 35445 33468 35479
rect 33416 35436 33468 35445
rect 34796 35436 34848 35488
rect 35900 35436 35952 35488
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 33416 35232 33468 35284
rect 33048 35164 33100 35216
rect 34520 35096 34572 35148
rect 32128 35071 32180 35080
rect 32128 35037 32137 35071
rect 32137 35037 32171 35071
rect 32171 35037 32180 35071
rect 32128 35028 32180 35037
rect 34612 35071 34664 35080
rect 34612 35037 34621 35071
rect 34621 35037 34655 35071
rect 34655 35037 34664 35071
rect 34612 35028 34664 35037
rect 34520 34935 34572 34944
rect 34520 34901 34529 34935
rect 34529 34901 34563 34935
rect 34563 34901 34572 34935
rect 34520 34892 34572 34901
rect 35900 34892 35952 34944
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 34520 34688 34572 34740
rect 37556 34731 37608 34740
rect 37556 34697 37565 34731
rect 37565 34697 37599 34731
rect 37599 34697 37608 34731
rect 37556 34688 37608 34697
rect 30012 34348 30064 34400
rect 32128 34484 32180 34536
rect 34612 34663 34664 34672
rect 34612 34629 34621 34663
rect 34621 34629 34655 34663
rect 34655 34629 34664 34663
rect 34612 34620 34664 34629
rect 33232 34552 33284 34604
rect 33048 34484 33100 34536
rect 30564 34416 30616 34468
rect 33324 34459 33376 34468
rect 33324 34425 33333 34459
rect 33333 34425 33367 34459
rect 33367 34425 33376 34459
rect 33324 34416 33376 34425
rect 31852 34391 31904 34400
rect 31852 34357 31861 34391
rect 31861 34357 31895 34391
rect 31895 34357 31904 34391
rect 31852 34348 31904 34357
rect 32956 34391 33008 34400
rect 32956 34357 32965 34391
rect 32965 34357 32999 34391
rect 32999 34357 33008 34391
rect 32956 34348 33008 34357
rect 37832 34484 37884 34536
rect 34428 34416 34480 34468
rect 33508 34348 33560 34400
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 30564 34187 30616 34196
rect 30564 34153 30573 34187
rect 30573 34153 30607 34187
rect 30607 34153 30616 34187
rect 30564 34144 30616 34153
rect 33508 34187 33560 34196
rect 33508 34153 33517 34187
rect 33517 34153 33551 34187
rect 33551 34153 33560 34187
rect 33508 34144 33560 34153
rect 31852 34076 31904 34128
rect 32864 34076 32916 34128
rect 33324 34076 33376 34128
rect 34428 34119 34480 34128
rect 34428 34085 34437 34119
rect 34437 34085 34471 34119
rect 34471 34085 34480 34119
rect 34428 34076 34480 34085
rect 34520 34076 34572 34128
rect 35808 34076 35860 34128
rect 32128 33983 32180 33992
rect 32128 33949 32137 33983
rect 32137 33949 32171 33983
rect 32171 33949 32180 33983
rect 32128 33940 32180 33949
rect 34612 33983 34664 33992
rect 34612 33949 34621 33983
rect 34621 33949 34655 33983
rect 34655 33949 34664 33983
rect 34612 33940 34664 33949
rect 30104 33847 30156 33856
rect 30104 33813 30113 33847
rect 30113 33813 30147 33847
rect 30147 33813 30156 33847
rect 30104 33804 30156 33813
rect 33232 33804 33284 33856
rect 35992 33847 36044 33856
rect 35992 33813 36001 33847
rect 36001 33813 36035 33847
rect 36035 33813 36044 33847
rect 35992 33804 36044 33813
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 30656 33600 30708 33652
rect 32496 33600 32548 33652
rect 33876 33600 33928 33652
rect 34520 33600 34572 33652
rect 32128 33575 32180 33584
rect 32128 33541 32137 33575
rect 32137 33541 32171 33575
rect 32171 33541 32180 33575
rect 32128 33532 32180 33541
rect 32496 33464 32548 33516
rect 33232 33464 33284 33516
rect 30012 33439 30064 33448
rect 29460 33260 29512 33312
rect 30012 33405 30021 33439
rect 30021 33405 30055 33439
rect 30055 33405 30064 33439
rect 30012 33396 30064 33405
rect 30104 33396 30156 33448
rect 30288 33439 30340 33448
rect 30288 33405 30311 33439
rect 30311 33405 30340 33439
rect 32864 33439 32916 33448
rect 30288 33396 30340 33405
rect 32864 33405 32873 33439
rect 32873 33405 32907 33439
rect 32907 33405 32916 33439
rect 32864 33396 32916 33405
rect 32312 33260 32364 33312
rect 34612 33303 34664 33312
rect 34612 33269 34621 33303
rect 34621 33269 34655 33303
rect 34655 33269 34664 33303
rect 35348 33396 35400 33448
rect 35992 33396 36044 33448
rect 34612 33260 34664 33269
rect 36636 33303 36688 33312
rect 36636 33269 36645 33303
rect 36645 33269 36679 33303
rect 36679 33269 36688 33303
rect 36636 33260 36688 33269
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 30380 33056 30432 33108
rect 30748 33056 30800 33108
rect 32496 33099 32548 33108
rect 32496 33065 32505 33099
rect 32505 33065 32539 33099
rect 32539 33065 32548 33099
rect 32496 33056 32548 33065
rect 32864 33099 32916 33108
rect 32864 33065 32873 33099
rect 32873 33065 32907 33099
rect 32907 33065 32916 33099
rect 32864 33056 32916 33065
rect 33876 33099 33928 33108
rect 33876 33065 33885 33099
rect 33885 33065 33919 33099
rect 33919 33065 33928 33099
rect 33876 33056 33928 33065
rect 35348 33056 35400 33108
rect 29736 32963 29788 32972
rect 29736 32929 29770 32963
rect 29770 32929 29788 32963
rect 29736 32920 29788 32929
rect 29460 32895 29512 32904
rect 29460 32861 29469 32895
rect 29469 32861 29503 32895
rect 29503 32861 29512 32895
rect 29460 32852 29512 32861
rect 33600 32852 33652 32904
rect 34336 32920 34388 32972
rect 35440 32963 35492 32972
rect 35440 32929 35474 32963
rect 35474 32929 35492 32963
rect 35440 32920 35492 32929
rect 36636 32920 36688 32972
rect 34612 32852 34664 32904
rect 30932 32716 30984 32768
rect 33232 32759 33284 32768
rect 33232 32725 33241 32759
rect 33241 32725 33275 32759
rect 33275 32725 33284 32759
rect 33232 32716 33284 32725
rect 33508 32759 33560 32768
rect 33508 32725 33517 32759
rect 33517 32725 33551 32759
rect 33551 32725 33560 32759
rect 33508 32716 33560 32725
rect 35808 32716 35860 32768
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 29736 32512 29788 32564
rect 33876 32512 33928 32564
rect 34612 32555 34664 32564
rect 34612 32521 34621 32555
rect 34621 32521 34655 32555
rect 34655 32521 34664 32555
rect 34612 32512 34664 32521
rect 36636 32512 36688 32564
rect 36820 32555 36872 32564
rect 36820 32521 36829 32555
rect 36829 32521 36863 32555
rect 36863 32521 36872 32555
rect 36820 32512 36872 32521
rect 33600 32487 33652 32496
rect 30932 32419 30984 32428
rect 30932 32385 30941 32419
rect 30941 32385 30975 32419
rect 30975 32385 30984 32419
rect 30932 32376 30984 32385
rect 33600 32453 33609 32487
rect 33609 32453 33643 32487
rect 33643 32453 33652 32487
rect 33600 32444 33652 32453
rect 32588 32419 32640 32428
rect 32588 32385 32597 32419
rect 32597 32385 32631 32419
rect 32631 32385 32640 32419
rect 32588 32376 32640 32385
rect 35992 32444 36044 32496
rect 35624 32419 35676 32428
rect 35624 32385 35633 32419
rect 35633 32385 35667 32419
rect 35667 32385 35676 32419
rect 35624 32376 35676 32385
rect 30748 32351 30800 32360
rect 30748 32317 30757 32351
rect 30757 32317 30791 32351
rect 30791 32317 30800 32351
rect 30748 32308 30800 32317
rect 32312 32351 32364 32360
rect 32312 32317 32321 32351
rect 32321 32317 32355 32351
rect 32355 32317 32364 32351
rect 32312 32308 32364 32317
rect 28448 32172 28500 32224
rect 29460 32215 29512 32224
rect 29460 32181 29469 32215
rect 29469 32181 29503 32215
rect 29503 32181 29512 32215
rect 29460 32172 29512 32181
rect 31944 32215 31996 32224
rect 31944 32181 31953 32215
rect 31953 32181 31987 32215
rect 31987 32181 31996 32215
rect 31944 32172 31996 32181
rect 33968 32172 34020 32224
rect 34336 32215 34388 32224
rect 34336 32181 34345 32215
rect 34345 32181 34379 32215
rect 34379 32181 34388 32215
rect 34336 32172 34388 32181
rect 34704 32172 34756 32224
rect 35440 32215 35492 32224
rect 35440 32181 35449 32215
rect 35449 32181 35483 32215
rect 35483 32181 35492 32215
rect 35440 32172 35492 32181
rect 37096 32172 37148 32224
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 29736 31968 29788 32020
rect 30748 31968 30800 32020
rect 30932 31968 30984 32020
rect 31668 31968 31720 32020
rect 28540 31875 28592 31884
rect 28540 31841 28574 31875
rect 28574 31841 28592 31875
rect 28540 31832 28592 31841
rect 31024 31832 31076 31884
rect 32956 31968 33008 32020
rect 33232 31968 33284 32020
rect 34612 32011 34664 32020
rect 34612 31977 34621 32011
rect 34621 31977 34655 32011
rect 34655 31977 34664 32011
rect 34612 31968 34664 31977
rect 35440 31968 35492 32020
rect 35900 31968 35952 32020
rect 32772 31900 32824 31952
rect 33508 31900 33560 31952
rect 34520 31832 34572 31884
rect 35808 31832 35860 31884
rect 28448 31628 28500 31680
rect 31852 31671 31904 31680
rect 31852 31637 31861 31671
rect 31861 31637 31895 31671
rect 31895 31637 31904 31671
rect 32588 31764 32640 31816
rect 31852 31628 31904 31637
rect 34060 31671 34112 31680
rect 34060 31637 34069 31671
rect 34069 31637 34103 31671
rect 34103 31637 34112 31671
rect 34060 31628 34112 31637
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 31024 31467 31076 31476
rect 31024 31433 31033 31467
rect 31033 31433 31067 31467
rect 31067 31433 31076 31467
rect 31024 31424 31076 31433
rect 32772 31424 32824 31476
rect 31760 31288 31812 31340
rect 35348 31356 35400 31408
rect 35624 31356 35676 31408
rect 31944 31220 31996 31272
rect 34060 31288 34112 31340
rect 34428 31288 34480 31340
rect 34612 31288 34664 31340
rect 35716 31331 35768 31340
rect 35716 31297 35725 31331
rect 35725 31297 35759 31331
rect 35759 31297 35768 31331
rect 35716 31288 35768 31297
rect 36084 31288 36136 31340
rect 35808 31220 35860 31272
rect 24860 31127 24912 31136
rect 24860 31093 24869 31127
rect 24869 31093 24903 31127
rect 24903 31093 24912 31127
rect 24860 31084 24912 31093
rect 27528 31127 27580 31136
rect 27528 31093 27537 31127
rect 27537 31093 27571 31127
rect 27571 31093 27580 31127
rect 27528 31084 27580 31093
rect 28448 31084 28500 31136
rect 28540 31084 28592 31136
rect 33324 31084 33376 31136
rect 35256 31084 35308 31136
rect 35440 31127 35492 31136
rect 35440 31093 35449 31127
rect 35449 31093 35483 31127
rect 35483 31093 35492 31127
rect 35440 31084 35492 31093
rect 35900 31084 35952 31136
rect 36084 31127 36136 31136
rect 36084 31093 36093 31127
rect 36093 31093 36127 31127
rect 36127 31093 36136 31127
rect 36084 31084 36136 31093
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 24860 30880 24912 30932
rect 25228 30923 25280 30932
rect 25228 30889 25237 30923
rect 25237 30889 25271 30923
rect 25271 30889 25280 30923
rect 25228 30880 25280 30889
rect 32956 30880 33008 30932
rect 33232 30880 33284 30932
rect 35992 30880 36044 30932
rect 27620 30744 27672 30796
rect 32128 30787 32180 30796
rect 32128 30753 32137 30787
rect 32137 30753 32171 30787
rect 32171 30753 32180 30787
rect 32128 30744 32180 30753
rect 33140 30744 33192 30796
rect 35440 30744 35492 30796
rect 35808 30744 35860 30796
rect 24860 30676 24912 30728
rect 26884 30719 26936 30728
rect 24952 30608 25004 30660
rect 26884 30685 26893 30719
rect 26893 30685 26927 30719
rect 26927 30685 26936 30719
rect 26884 30676 26936 30685
rect 26240 30540 26292 30592
rect 29276 30583 29328 30592
rect 29276 30549 29285 30583
rect 29285 30549 29319 30583
rect 29319 30549 29328 30583
rect 29276 30540 29328 30549
rect 29644 30583 29696 30592
rect 29644 30549 29653 30583
rect 29653 30549 29687 30583
rect 29687 30549 29696 30583
rect 29644 30540 29696 30549
rect 32312 30583 32364 30592
rect 32312 30549 32321 30583
rect 32321 30549 32355 30583
rect 32355 30549 32364 30583
rect 32312 30540 32364 30549
rect 33140 30540 33192 30592
rect 34152 30540 34204 30592
rect 34612 30583 34664 30592
rect 34612 30549 34621 30583
rect 34621 30549 34655 30583
rect 34655 30549 34664 30583
rect 34612 30540 34664 30549
rect 35992 30540 36044 30592
rect 37188 30540 37240 30592
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 27896 30336 27948 30388
rect 28540 30336 28592 30388
rect 33140 30336 33192 30388
rect 24216 30268 24268 30320
rect 24860 30268 24912 30320
rect 26884 30268 26936 30320
rect 28448 30268 28500 30320
rect 34612 30336 34664 30388
rect 34704 30311 34756 30320
rect 34704 30277 34713 30311
rect 34713 30277 34747 30311
rect 34747 30277 34756 30311
rect 34704 30268 34756 30277
rect 35164 30268 35216 30320
rect 35992 30336 36044 30388
rect 27528 30200 27580 30252
rect 23940 29996 23992 30048
rect 25228 30175 25280 30184
rect 25228 30141 25262 30175
rect 25262 30141 25280 30175
rect 25228 30132 25280 30141
rect 27620 30132 27672 30184
rect 29276 30200 29328 30252
rect 29644 30175 29696 30184
rect 29644 30141 29653 30175
rect 29653 30141 29687 30175
rect 29687 30141 29696 30175
rect 29644 30132 29696 30141
rect 26332 30039 26384 30048
rect 26332 30005 26341 30039
rect 26341 30005 26375 30039
rect 26375 30005 26384 30039
rect 26332 29996 26384 30005
rect 27436 30039 27488 30048
rect 27436 30005 27445 30039
rect 27445 30005 27479 30039
rect 27479 30005 27488 30039
rect 27436 29996 27488 30005
rect 29000 29996 29052 30048
rect 29460 29996 29512 30048
rect 33048 30200 33100 30252
rect 33232 30200 33284 30252
rect 33784 30200 33836 30252
rect 34336 30200 34388 30252
rect 36728 30268 36780 30320
rect 32128 30132 32180 30184
rect 35256 30175 35308 30184
rect 33416 29996 33468 30048
rect 33600 30039 33652 30048
rect 33600 30005 33609 30039
rect 33609 30005 33643 30039
rect 33643 30005 33652 30039
rect 33600 29996 33652 30005
rect 34244 30039 34296 30048
rect 34244 30005 34253 30039
rect 34253 30005 34287 30039
rect 34287 30005 34296 30039
rect 34244 29996 34296 30005
rect 35256 30141 35265 30175
rect 35265 30141 35299 30175
rect 35299 30141 35308 30175
rect 35256 30132 35308 30141
rect 35164 30064 35216 30116
rect 36176 30064 36228 30116
rect 35900 30039 35952 30048
rect 35900 30005 35909 30039
rect 35909 30005 35943 30039
rect 35943 30005 35952 30039
rect 35900 29996 35952 30005
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 25228 29792 25280 29844
rect 27620 29792 27672 29844
rect 29644 29792 29696 29844
rect 34520 29792 34572 29844
rect 35348 29792 35400 29844
rect 24216 29767 24268 29776
rect 24216 29733 24250 29767
rect 24250 29733 24268 29767
rect 24216 29724 24268 29733
rect 26332 29724 26384 29776
rect 26884 29724 26936 29776
rect 29276 29767 29328 29776
rect 29276 29733 29310 29767
rect 29310 29733 29328 29767
rect 29276 29724 29328 29733
rect 32956 29724 33008 29776
rect 33600 29724 33652 29776
rect 26516 29699 26568 29708
rect 26516 29665 26525 29699
rect 26525 29665 26559 29699
rect 26559 29665 26568 29699
rect 26516 29656 26568 29665
rect 28448 29656 28500 29708
rect 29092 29656 29144 29708
rect 34520 29656 34572 29708
rect 35716 29699 35768 29708
rect 23940 29631 23992 29640
rect 23940 29597 23949 29631
rect 23949 29597 23983 29631
rect 23983 29597 23992 29631
rect 23940 29588 23992 29597
rect 32864 29631 32916 29640
rect 32864 29597 32873 29631
rect 32873 29597 32907 29631
rect 32907 29597 32916 29631
rect 32864 29588 32916 29597
rect 34612 29588 34664 29640
rect 35716 29665 35725 29699
rect 35725 29665 35759 29699
rect 35759 29665 35768 29699
rect 35716 29656 35768 29665
rect 24216 29452 24268 29504
rect 27528 29452 27580 29504
rect 33600 29452 33652 29504
rect 34244 29495 34296 29504
rect 34244 29461 34253 29495
rect 34253 29461 34287 29495
rect 34287 29461 34296 29495
rect 34244 29452 34296 29461
rect 35256 29452 35308 29504
rect 35992 29588 36044 29640
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 24860 29248 24912 29300
rect 26332 29248 26384 29300
rect 27620 29248 27672 29300
rect 32312 29291 32364 29300
rect 32312 29257 32321 29291
rect 32321 29257 32355 29291
rect 32355 29257 32364 29291
rect 32312 29248 32364 29257
rect 32864 29248 32916 29300
rect 33048 29248 33100 29300
rect 35808 29248 35860 29300
rect 37188 29248 37240 29300
rect 26240 29112 26292 29164
rect 28448 29180 28500 29232
rect 30288 29180 30340 29232
rect 36268 29223 36320 29232
rect 36268 29189 36277 29223
rect 36277 29189 36311 29223
rect 36311 29189 36320 29223
rect 36268 29180 36320 29189
rect 27528 29112 27580 29164
rect 23940 29087 23992 29096
rect 23940 29053 23949 29087
rect 23949 29053 23983 29087
rect 23983 29053 23992 29087
rect 23940 29044 23992 29053
rect 24216 29087 24268 29096
rect 24216 29053 24250 29087
rect 24250 29053 24268 29087
rect 24216 29044 24268 29053
rect 26332 29044 26384 29096
rect 27436 29044 27488 29096
rect 26516 28976 26568 29028
rect 32864 29112 32916 29164
rect 33784 29155 33836 29164
rect 33784 29121 33793 29155
rect 33793 29121 33827 29155
rect 33827 29121 33836 29155
rect 33784 29112 33836 29121
rect 34152 29112 34204 29164
rect 33600 29087 33652 29096
rect 29644 28976 29696 29028
rect 33600 29053 33609 29087
rect 33609 29053 33643 29087
rect 33643 29053 33652 29087
rect 33600 29044 33652 29053
rect 34980 29044 35032 29096
rect 33048 28976 33100 29028
rect 34520 28976 34572 29028
rect 35256 28976 35308 29028
rect 38016 29019 38068 29028
rect 38016 28985 38025 29019
rect 38025 28985 38059 29019
rect 38059 28985 38068 29019
rect 38016 28976 38068 28985
rect 23572 28908 23624 28960
rect 27804 28951 27856 28960
rect 27804 28917 27813 28951
rect 27813 28917 27847 28951
rect 27847 28917 27856 28951
rect 27804 28908 27856 28917
rect 28448 28908 28500 28960
rect 28540 28908 28592 28960
rect 29092 28951 29144 28960
rect 29092 28917 29101 28951
rect 29101 28917 29135 28951
rect 29135 28917 29144 28951
rect 29092 28908 29144 28917
rect 33232 28951 33284 28960
rect 33232 28917 33241 28951
rect 33241 28917 33275 28951
rect 33275 28917 33284 28951
rect 33232 28908 33284 28917
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 24216 28704 24268 28756
rect 26332 28747 26384 28756
rect 26332 28713 26341 28747
rect 26341 28713 26375 28747
rect 26375 28713 26384 28747
rect 26332 28704 26384 28713
rect 29276 28704 29328 28756
rect 32956 28747 33008 28756
rect 32956 28713 32965 28747
rect 32965 28713 32999 28747
rect 32999 28713 33008 28747
rect 32956 28704 33008 28713
rect 34520 28704 34572 28756
rect 35348 28747 35400 28756
rect 35348 28713 35357 28747
rect 35357 28713 35391 28747
rect 35391 28713 35400 28747
rect 35348 28704 35400 28713
rect 35992 28704 36044 28756
rect 27068 28636 27120 28688
rect 29552 28636 29604 28688
rect 30288 28636 30340 28688
rect 23480 28568 23532 28620
rect 27620 28568 27672 28620
rect 28080 28611 28132 28620
rect 28080 28577 28089 28611
rect 28089 28577 28123 28611
rect 28123 28577 28132 28611
rect 28080 28568 28132 28577
rect 32864 28568 32916 28620
rect 33048 28568 33100 28620
rect 34244 28568 34296 28620
rect 35992 28568 36044 28620
rect 26976 28543 27028 28552
rect 26976 28509 26985 28543
rect 26985 28509 27019 28543
rect 27019 28509 27028 28543
rect 26976 28500 27028 28509
rect 27160 28543 27212 28552
rect 27160 28509 27169 28543
rect 27169 28509 27203 28543
rect 27203 28509 27212 28543
rect 27160 28500 27212 28509
rect 29092 28500 29144 28552
rect 23572 28364 23624 28416
rect 26332 28364 26384 28416
rect 27620 28407 27672 28416
rect 27620 28373 27629 28407
rect 27629 28373 27663 28407
rect 27663 28373 27672 28407
rect 27620 28364 27672 28373
rect 28264 28407 28316 28416
rect 28264 28373 28273 28407
rect 28273 28373 28307 28407
rect 28307 28373 28316 28407
rect 28264 28364 28316 28373
rect 30288 28364 30340 28416
rect 36084 28364 36136 28416
rect 36728 28364 36780 28416
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 23480 28160 23532 28212
rect 26976 28160 27028 28212
rect 27068 28203 27120 28212
rect 27068 28169 27077 28203
rect 27077 28169 27111 28203
rect 27111 28169 27120 28203
rect 27068 28160 27120 28169
rect 27804 28160 27856 28212
rect 32588 28203 32640 28212
rect 32588 28169 32597 28203
rect 32597 28169 32631 28203
rect 32631 28169 32640 28203
rect 32588 28160 32640 28169
rect 33140 28160 33192 28212
rect 34244 28203 34296 28212
rect 34244 28169 34253 28203
rect 34253 28169 34287 28203
rect 34287 28169 34296 28203
rect 34244 28160 34296 28169
rect 35532 28160 35584 28212
rect 36728 28203 36780 28212
rect 36728 28169 36737 28203
rect 36737 28169 36771 28203
rect 36771 28169 36780 28203
rect 36728 28160 36780 28169
rect 24860 28092 24912 28144
rect 27160 28092 27212 28144
rect 27620 28024 27672 28076
rect 33140 28067 33192 28076
rect 33140 28033 33149 28067
rect 33149 28033 33183 28067
rect 33183 28033 33192 28067
rect 33140 28024 33192 28033
rect 33416 28024 33468 28076
rect 23572 27956 23624 28008
rect 23480 27888 23532 27940
rect 24216 27888 24268 27940
rect 28908 27956 28960 28008
rect 32588 27956 32640 28008
rect 33232 27956 33284 28008
rect 29276 27888 29328 27940
rect 31852 27931 31904 27940
rect 31852 27897 31861 27931
rect 31861 27897 31895 27931
rect 31895 27897 31904 27931
rect 34336 28024 34388 28076
rect 31852 27888 31904 27897
rect 23572 27820 23624 27872
rect 26148 27820 26200 27872
rect 26608 27820 26660 27872
rect 27988 27863 28040 27872
rect 27988 27829 27997 27863
rect 27997 27829 28031 27863
rect 28031 27829 28040 27863
rect 27988 27820 28040 27829
rect 29092 27863 29144 27872
rect 29092 27829 29101 27863
rect 29101 27829 29135 27863
rect 29135 27829 29144 27863
rect 29092 27820 29144 27829
rect 30656 27820 30708 27872
rect 32128 27863 32180 27872
rect 32128 27829 32137 27863
rect 32137 27829 32171 27863
rect 32171 27829 32180 27863
rect 32128 27820 32180 27829
rect 34612 27820 34664 27872
rect 35992 27863 36044 27872
rect 35992 27829 36001 27863
rect 36001 27829 36035 27863
rect 36035 27829 36044 27863
rect 35992 27820 36044 27829
rect 37188 27863 37240 27872
rect 37188 27829 37197 27863
rect 37197 27829 37231 27863
rect 37231 27829 37240 27863
rect 37188 27820 37240 27829
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 24216 27659 24268 27668
rect 24216 27625 24225 27659
rect 24225 27625 24259 27659
rect 24259 27625 24268 27659
rect 24216 27616 24268 27625
rect 27988 27616 28040 27668
rect 24860 27548 24912 27600
rect 28080 27591 28132 27600
rect 28080 27557 28089 27591
rect 28089 27557 28123 27591
rect 28123 27557 28132 27591
rect 28080 27548 28132 27557
rect 28724 27548 28776 27600
rect 29552 27616 29604 27668
rect 33232 27616 33284 27668
rect 33600 27548 33652 27600
rect 35532 27548 35584 27600
rect 24308 27455 24360 27464
rect 24308 27421 24317 27455
rect 24317 27421 24351 27455
rect 24351 27421 24360 27455
rect 24308 27412 24360 27421
rect 26332 27480 26384 27532
rect 29276 27523 29328 27532
rect 29276 27489 29285 27523
rect 29285 27489 29319 27523
rect 29319 27489 29328 27523
rect 30288 27523 30340 27532
rect 29276 27480 29328 27489
rect 30288 27489 30297 27523
rect 30297 27489 30331 27523
rect 30331 27489 30340 27523
rect 30288 27480 30340 27489
rect 30472 27523 30524 27532
rect 30472 27489 30481 27523
rect 30481 27489 30515 27523
rect 30515 27489 30524 27523
rect 30472 27480 30524 27489
rect 30656 27523 30708 27532
rect 30656 27489 30665 27523
rect 30665 27489 30699 27523
rect 30699 27489 30708 27523
rect 30656 27480 30708 27489
rect 31944 27480 31996 27532
rect 33140 27480 33192 27532
rect 26424 27412 26476 27464
rect 27160 27455 27212 27464
rect 27160 27421 27169 27455
rect 27169 27421 27203 27455
rect 27203 27421 27212 27455
rect 27160 27412 27212 27421
rect 27528 27412 27580 27464
rect 29460 27455 29512 27464
rect 29460 27421 29469 27455
rect 29469 27421 29503 27455
rect 29503 27421 29512 27455
rect 29460 27412 29512 27421
rect 32772 27412 32824 27464
rect 35256 27480 35308 27532
rect 33232 27387 33284 27396
rect 33232 27353 33241 27387
rect 33241 27353 33275 27387
rect 33275 27353 33284 27387
rect 33232 27344 33284 27353
rect 34704 27412 34756 27464
rect 23572 27276 23624 27328
rect 23848 27319 23900 27328
rect 23848 27285 23857 27319
rect 23857 27285 23891 27319
rect 23891 27285 23900 27319
rect 23848 27276 23900 27285
rect 26516 27319 26568 27328
rect 26516 27285 26525 27319
rect 26525 27285 26559 27319
rect 26559 27285 26568 27319
rect 26516 27276 26568 27285
rect 32312 27319 32364 27328
rect 32312 27285 32321 27319
rect 32321 27285 32355 27319
rect 32355 27285 32364 27319
rect 32312 27276 32364 27285
rect 33324 27319 33376 27328
rect 33324 27285 33333 27319
rect 33333 27285 33367 27319
rect 33367 27285 33376 27319
rect 33324 27276 33376 27285
rect 34428 27319 34480 27328
rect 34428 27285 34437 27319
rect 34437 27285 34471 27319
rect 34471 27285 34480 27319
rect 34428 27276 34480 27285
rect 36544 27319 36596 27328
rect 36544 27285 36553 27319
rect 36553 27285 36587 27319
rect 36587 27285 36596 27319
rect 36544 27276 36596 27285
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 22376 27115 22428 27124
rect 22376 27081 22385 27115
rect 22385 27081 22419 27115
rect 22419 27081 22428 27115
rect 22376 27072 22428 27081
rect 23480 27072 23532 27124
rect 26424 27072 26476 27124
rect 26608 27072 26660 27124
rect 29276 27072 29328 27124
rect 30656 27072 30708 27124
rect 33140 27115 33192 27124
rect 33140 27081 33149 27115
rect 33149 27081 33183 27115
rect 33183 27081 33192 27115
rect 33140 27072 33192 27081
rect 33600 27072 33652 27124
rect 35716 27072 35768 27124
rect 36452 27072 36504 27124
rect 28724 27047 28776 27056
rect 28724 27013 28733 27047
rect 28733 27013 28767 27047
rect 28767 27013 28776 27047
rect 28724 27004 28776 27013
rect 32772 27047 32824 27056
rect 32772 27013 32781 27047
rect 32781 27013 32815 27047
rect 32815 27013 32824 27047
rect 32772 27004 32824 27013
rect 34520 27004 34572 27056
rect 36820 27047 36872 27056
rect 36820 27013 36829 27047
rect 36829 27013 36863 27047
rect 36863 27013 36872 27047
rect 36820 27004 36872 27013
rect 27804 26979 27856 26988
rect 27804 26945 27813 26979
rect 27813 26945 27847 26979
rect 27847 26945 27856 26979
rect 27804 26936 27856 26945
rect 33876 26979 33928 26988
rect 33876 26945 33885 26979
rect 33885 26945 33919 26979
rect 33919 26945 33928 26979
rect 33876 26936 33928 26945
rect 22376 26868 22428 26920
rect 23572 26868 23624 26920
rect 24308 26800 24360 26852
rect 30656 26868 30708 26920
rect 33232 26868 33284 26920
rect 35532 26868 35584 26920
rect 35716 26911 35768 26920
rect 32864 26800 32916 26852
rect 34336 26800 34388 26852
rect 35716 26877 35750 26911
rect 35750 26877 35768 26911
rect 35716 26868 35768 26877
rect 36544 26868 36596 26920
rect 22652 26775 22704 26784
rect 22652 26741 22661 26775
rect 22661 26741 22695 26775
rect 22695 26741 22704 26775
rect 22652 26732 22704 26741
rect 23572 26732 23624 26784
rect 26608 26775 26660 26784
rect 26608 26741 26617 26775
rect 26617 26741 26651 26775
rect 26651 26741 26660 26775
rect 26608 26732 26660 26741
rect 27712 26732 27764 26784
rect 29092 26775 29144 26784
rect 29092 26741 29101 26775
rect 29101 26741 29135 26775
rect 29135 26741 29144 26775
rect 29092 26732 29144 26741
rect 29276 26732 29328 26784
rect 30840 26732 30892 26784
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 23480 26571 23532 26580
rect 23480 26537 23489 26571
rect 23489 26537 23523 26571
rect 23523 26537 23532 26571
rect 23480 26528 23532 26537
rect 24308 26528 24360 26580
rect 26240 26528 26292 26580
rect 23756 26460 23808 26512
rect 26332 26503 26384 26512
rect 26332 26469 26341 26503
rect 26341 26469 26375 26503
rect 26375 26469 26384 26503
rect 26332 26460 26384 26469
rect 26884 26435 26936 26444
rect 26884 26401 26893 26435
rect 26893 26401 26927 26435
rect 26927 26401 26936 26435
rect 26884 26392 26936 26401
rect 27528 26392 27580 26444
rect 28264 26528 28316 26580
rect 28816 26528 28868 26580
rect 30472 26528 30524 26580
rect 31944 26571 31996 26580
rect 31944 26537 31953 26571
rect 31953 26537 31987 26571
rect 31987 26537 31996 26571
rect 31944 26528 31996 26537
rect 33876 26528 33928 26580
rect 35532 26528 35584 26580
rect 28448 26503 28500 26512
rect 28448 26469 28457 26503
rect 28457 26469 28491 26503
rect 28491 26469 28500 26503
rect 28448 26460 28500 26469
rect 29460 26460 29512 26512
rect 30380 26460 30432 26512
rect 32864 26503 32916 26512
rect 32864 26469 32873 26503
rect 32873 26469 32907 26503
rect 32907 26469 32916 26503
rect 32864 26460 32916 26469
rect 34428 26460 34480 26512
rect 35716 26460 35768 26512
rect 35992 26460 36044 26512
rect 30196 26392 30248 26444
rect 33048 26392 33100 26444
rect 35532 26392 35584 26444
rect 23572 26367 23624 26376
rect 23572 26333 23581 26367
rect 23581 26333 23615 26367
rect 23615 26333 23624 26367
rect 23572 26324 23624 26333
rect 27160 26367 27212 26376
rect 27160 26333 27169 26367
rect 27169 26333 27203 26367
rect 27203 26333 27212 26367
rect 27160 26324 27212 26333
rect 27804 26324 27856 26376
rect 28724 26367 28776 26376
rect 28724 26333 28733 26367
rect 28733 26333 28767 26367
rect 28767 26333 28776 26367
rect 28724 26324 28776 26333
rect 29828 26324 29880 26376
rect 30288 26367 30340 26376
rect 30288 26333 30297 26367
rect 30297 26333 30331 26367
rect 30331 26333 30340 26367
rect 30288 26324 30340 26333
rect 27068 26256 27120 26308
rect 35900 26256 35952 26308
rect 34336 26231 34388 26240
rect 34336 26197 34345 26231
rect 34345 26197 34379 26231
rect 34379 26197 34388 26231
rect 34336 26188 34388 26197
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 26332 25984 26384 26036
rect 26884 25984 26936 26036
rect 28264 25984 28316 26036
rect 32956 25984 33008 26036
rect 34428 25984 34480 26036
rect 34520 25984 34572 26036
rect 26792 25916 26844 25968
rect 28448 25916 28500 25968
rect 33048 25916 33100 25968
rect 27068 25891 27120 25900
rect 27068 25857 27077 25891
rect 27077 25857 27111 25891
rect 27111 25857 27120 25891
rect 27068 25848 27120 25857
rect 33508 25891 33560 25900
rect 33508 25857 33517 25891
rect 33517 25857 33551 25891
rect 33551 25857 33560 25891
rect 33508 25848 33560 25857
rect 34336 25848 34388 25900
rect 23572 25780 23624 25832
rect 23940 25780 23992 25832
rect 27712 25780 27764 25832
rect 28448 25780 28500 25832
rect 29828 25780 29880 25832
rect 33324 25823 33376 25832
rect 23756 25712 23808 25764
rect 24308 25755 24360 25764
rect 23940 25687 23992 25696
rect 23940 25653 23949 25687
rect 23949 25653 23983 25687
rect 23983 25653 23992 25687
rect 23940 25644 23992 25653
rect 24308 25721 24342 25755
rect 24342 25721 24360 25755
rect 24308 25712 24360 25721
rect 33324 25789 33333 25823
rect 33333 25789 33367 25823
rect 33367 25789 33376 25823
rect 33324 25780 33376 25789
rect 34704 25984 34756 26036
rect 35992 25984 36044 26036
rect 36176 26027 36228 26036
rect 36176 25993 36185 26027
rect 36185 25993 36219 26027
rect 36219 25993 36228 26027
rect 36176 25984 36228 25993
rect 35900 25780 35952 25832
rect 26884 25687 26936 25696
rect 26884 25653 26893 25687
rect 26893 25653 26927 25687
rect 26927 25653 26936 25687
rect 26884 25644 26936 25653
rect 27620 25687 27672 25696
rect 27620 25653 27629 25687
rect 27629 25653 27663 25687
rect 27663 25653 27672 25687
rect 27620 25644 27672 25653
rect 28264 25687 28316 25696
rect 28264 25653 28273 25687
rect 28273 25653 28307 25687
rect 28307 25653 28316 25687
rect 28264 25644 28316 25653
rect 29276 25644 29328 25696
rect 30012 25712 30064 25764
rect 30840 25712 30892 25764
rect 31300 25687 31352 25696
rect 31300 25653 31309 25687
rect 31309 25653 31343 25687
rect 31343 25653 31352 25687
rect 31300 25644 31352 25653
rect 32956 25644 33008 25696
rect 35532 25687 35584 25696
rect 35532 25653 35541 25687
rect 35541 25653 35575 25687
rect 35575 25653 35584 25687
rect 35532 25644 35584 25653
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 26332 25483 26384 25492
rect 26332 25449 26341 25483
rect 26341 25449 26375 25483
rect 26375 25449 26384 25483
rect 26332 25440 26384 25449
rect 26884 25440 26936 25492
rect 28264 25440 28316 25492
rect 30104 25440 30156 25492
rect 30196 25440 30248 25492
rect 30840 25483 30892 25492
rect 30840 25449 30849 25483
rect 30849 25449 30883 25483
rect 30883 25449 30892 25483
rect 30840 25440 30892 25449
rect 32956 25483 33008 25492
rect 26792 25415 26844 25424
rect 26792 25381 26826 25415
rect 26826 25381 26844 25415
rect 26792 25372 26844 25381
rect 28448 25415 28500 25424
rect 28448 25381 28457 25415
rect 28457 25381 28491 25415
rect 28491 25381 28500 25415
rect 28448 25372 28500 25381
rect 28724 25372 28776 25424
rect 30380 25372 30432 25424
rect 32956 25449 32965 25483
rect 32965 25449 32999 25483
rect 32999 25449 33008 25483
rect 32956 25440 33008 25449
rect 33508 25372 33560 25424
rect 24216 25347 24268 25356
rect 24216 25313 24250 25347
rect 24250 25313 24268 25347
rect 24216 25304 24268 25313
rect 25228 25304 25280 25356
rect 27068 25304 27120 25356
rect 30932 25347 30984 25356
rect 30932 25313 30941 25347
rect 30941 25313 30975 25347
rect 30975 25313 30984 25347
rect 30932 25304 30984 25313
rect 33140 25347 33192 25356
rect 33140 25313 33149 25347
rect 33149 25313 33183 25347
rect 33183 25313 33192 25347
rect 33140 25304 33192 25313
rect 23940 25279 23992 25288
rect 23940 25245 23949 25279
rect 23949 25245 23983 25279
rect 23983 25245 23992 25279
rect 23940 25236 23992 25245
rect 26516 25279 26568 25288
rect 26516 25245 26525 25279
rect 26525 25245 26559 25279
rect 26559 25245 26568 25279
rect 26516 25236 26568 25245
rect 24308 25100 24360 25152
rect 24952 25100 25004 25152
rect 29000 25100 29052 25152
rect 30012 25279 30064 25288
rect 30012 25245 30021 25279
rect 30021 25245 30055 25279
rect 30055 25245 30064 25279
rect 30012 25236 30064 25245
rect 31760 25143 31812 25152
rect 31760 25109 31769 25143
rect 31769 25109 31803 25143
rect 31803 25109 31812 25143
rect 34520 25143 34572 25152
rect 31760 25100 31812 25109
rect 34520 25109 34529 25143
rect 34529 25109 34563 25143
rect 34563 25109 34572 25143
rect 34520 25100 34572 25109
rect 35440 25100 35492 25152
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 26516 24939 26568 24948
rect 26516 24905 26525 24939
rect 26525 24905 26559 24939
rect 26559 24905 26568 24939
rect 26516 24896 26568 24905
rect 26792 24896 26844 24948
rect 30932 24896 30984 24948
rect 33140 24939 33192 24948
rect 33140 24905 33149 24939
rect 33149 24905 33183 24939
rect 33183 24905 33192 24939
rect 33140 24896 33192 24905
rect 33508 24939 33560 24948
rect 33508 24905 33517 24939
rect 33517 24905 33551 24939
rect 33551 24905 33560 24939
rect 33508 24896 33560 24905
rect 31300 24828 31352 24880
rect 28816 24760 28868 24812
rect 29276 24803 29328 24812
rect 29276 24769 29285 24803
rect 29285 24769 29319 24803
rect 29319 24769 29328 24803
rect 29276 24760 29328 24769
rect 31760 24760 31812 24812
rect 34244 24803 34296 24812
rect 34244 24769 34253 24803
rect 34253 24769 34287 24803
rect 34287 24769 34296 24803
rect 34244 24760 34296 24769
rect 35440 24803 35492 24812
rect 35440 24769 35449 24803
rect 35449 24769 35483 24803
rect 35483 24769 35492 24803
rect 35440 24760 35492 24769
rect 23940 24599 23992 24608
rect 23940 24565 23949 24599
rect 23949 24565 23983 24599
rect 23983 24565 23992 24599
rect 24676 24624 24728 24676
rect 23940 24556 23992 24565
rect 25044 24556 25096 24608
rect 28908 24624 28960 24676
rect 34428 24692 34480 24744
rect 29552 24667 29604 24676
rect 29552 24633 29586 24667
rect 29586 24633 29604 24667
rect 29552 24624 29604 24633
rect 30380 24624 30432 24676
rect 29920 24556 29972 24608
rect 31760 24599 31812 24608
rect 31760 24565 31769 24599
rect 31769 24565 31803 24599
rect 31803 24565 31812 24599
rect 34336 24624 34388 24676
rect 31760 24556 31812 24565
rect 34612 24599 34664 24608
rect 34612 24565 34621 24599
rect 34621 24565 34655 24599
rect 34655 24565 34664 24599
rect 34612 24556 34664 24565
rect 34888 24599 34940 24608
rect 34888 24565 34897 24599
rect 34897 24565 34931 24599
rect 34931 24565 34940 24599
rect 34888 24556 34940 24565
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 24216 24352 24268 24404
rect 25044 24395 25096 24404
rect 25044 24361 25053 24395
rect 25053 24361 25087 24395
rect 25087 24361 25096 24395
rect 25044 24352 25096 24361
rect 30104 24395 30156 24404
rect 30104 24361 30113 24395
rect 30113 24361 30147 24395
rect 30147 24361 30156 24395
rect 30104 24352 30156 24361
rect 30840 24352 30892 24404
rect 31300 24352 31352 24404
rect 35440 24352 35492 24404
rect 24676 24284 24728 24336
rect 24952 24259 25004 24268
rect 24952 24225 24961 24259
rect 24961 24225 24995 24259
rect 24995 24225 25004 24259
rect 24952 24216 25004 24225
rect 28080 24216 28132 24268
rect 29920 24216 29972 24268
rect 30656 24259 30708 24268
rect 30656 24225 30665 24259
rect 30665 24225 30699 24259
rect 30699 24225 30708 24259
rect 30656 24216 30708 24225
rect 33876 24216 33928 24268
rect 34520 24216 34572 24268
rect 25228 24191 25280 24200
rect 25228 24157 25237 24191
rect 25237 24157 25271 24191
rect 25271 24157 25280 24191
rect 25228 24148 25280 24157
rect 26516 24148 26568 24200
rect 27252 24148 27304 24200
rect 28172 24191 28224 24200
rect 28172 24157 28181 24191
rect 28181 24157 28215 24191
rect 28215 24157 28224 24191
rect 28172 24148 28224 24157
rect 33140 24148 33192 24200
rect 33968 24191 34020 24200
rect 33968 24157 33977 24191
rect 33977 24157 34011 24191
rect 34011 24157 34020 24191
rect 33968 24148 34020 24157
rect 36452 24191 36504 24200
rect 36452 24157 36461 24191
rect 36461 24157 36495 24191
rect 36495 24157 36504 24191
rect 36452 24148 36504 24157
rect 24584 24123 24636 24132
rect 24584 24089 24593 24123
rect 24593 24089 24627 24123
rect 24627 24089 24636 24123
rect 24584 24080 24636 24089
rect 30472 24080 30524 24132
rect 28908 24012 28960 24064
rect 35716 24012 35768 24064
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 25044 23808 25096 23860
rect 25228 23808 25280 23860
rect 28080 23851 28132 23860
rect 28080 23817 28089 23851
rect 28089 23817 28123 23851
rect 28123 23817 28132 23851
rect 28080 23808 28132 23817
rect 28172 23808 28224 23860
rect 24952 23783 25004 23792
rect 24952 23749 24961 23783
rect 24961 23749 24995 23783
rect 24995 23749 25004 23783
rect 24952 23740 25004 23749
rect 30656 23808 30708 23860
rect 33968 23808 34020 23860
rect 36820 23851 36872 23860
rect 29920 23715 29972 23724
rect 29920 23681 29929 23715
rect 29929 23681 29963 23715
rect 29963 23681 29972 23715
rect 29920 23672 29972 23681
rect 34980 23740 35032 23792
rect 29276 23604 29328 23656
rect 30012 23604 30064 23656
rect 29736 23579 29788 23588
rect 29736 23545 29745 23579
rect 29745 23545 29779 23579
rect 29779 23545 29788 23579
rect 29736 23536 29788 23545
rect 34612 23672 34664 23724
rect 36820 23817 36829 23851
rect 36829 23817 36863 23851
rect 36863 23817 36872 23851
rect 36820 23808 36872 23817
rect 31300 23647 31352 23656
rect 31300 23613 31334 23647
rect 31334 23613 31352 23647
rect 31300 23604 31352 23613
rect 35716 23647 35768 23656
rect 35716 23613 35750 23647
rect 35750 23613 35768 23647
rect 35716 23604 35768 23613
rect 33140 23536 33192 23588
rect 33876 23536 33928 23588
rect 28172 23511 28224 23520
rect 28172 23477 28181 23511
rect 28181 23477 28215 23511
rect 28215 23477 28224 23511
rect 28172 23468 28224 23477
rect 29092 23468 29144 23520
rect 31944 23468 31996 23520
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 28172 23264 28224 23316
rect 28540 23264 28592 23316
rect 29092 23264 29144 23316
rect 29736 23264 29788 23316
rect 29920 23307 29972 23316
rect 29920 23273 29929 23307
rect 29929 23273 29963 23307
rect 29963 23273 29972 23307
rect 29920 23264 29972 23273
rect 30288 23264 30340 23316
rect 31300 23264 31352 23316
rect 34428 23264 34480 23316
rect 35716 23264 35768 23316
rect 33140 23196 33192 23248
rect 33692 23239 33744 23248
rect 33692 23205 33701 23239
rect 33701 23205 33735 23239
rect 33735 23205 33744 23239
rect 33692 23196 33744 23205
rect 35440 23196 35492 23248
rect 34520 23128 34572 23180
rect 34980 23171 35032 23180
rect 34980 23137 34989 23171
rect 34989 23137 35023 23171
rect 35023 23137 35032 23171
rect 34980 23128 35032 23137
rect 28080 23060 28132 23112
rect 28908 23060 28960 23112
rect 33784 23103 33836 23112
rect 33784 23069 33793 23103
rect 33793 23069 33827 23103
rect 33827 23069 33836 23103
rect 33784 23060 33836 23069
rect 33876 23103 33928 23112
rect 33876 23069 33885 23103
rect 33885 23069 33919 23103
rect 33919 23069 33928 23103
rect 33876 23060 33928 23069
rect 29736 22992 29788 23044
rect 24032 22967 24084 22976
rect 24032 22933 24041 22967
rect 24041 22933 24075 22967
rect 24075 22933 24084 22967
rect 24032 22924 24084 22933
rect 26792 22967 26844 22976
rect 26792 22933 26801 22967
rect 26801 22933 26835 22967
rect 26835 22933 26844 22967
rect 26792 22924 26844 22933
rect 34704 22924 34756 22976
rect 35348 22924 35400 22976
rect 36912 22967 36964 22976
rect 36912 22933 36921 22967
rect 36921 22933 36955 22967
rect 36955 22933 36964 22967
rect 36912 22924 36964 22933
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 28080 22720 28132 22772
rect 28540 22763 28592 22772
rect 28540 22729 28549 22763
rect 28549 22729 28583 22763
rect 28583 22729 28592 22763
rect 28540 22720 28592 22729
rect 33876 22720 33928 22772
rect 34520 22720 34572 22772
rect 36452 22763 36504 22772
rect 36452 22729 36461 22763
rect 36461 22729 36495 22763
rect 36495 22729 36504 22763
rect 36452 22720 36504 22729
rect 36544 22763 36596 22772
rect 36544 22729 36553 22763
rect 36553 22729 36587 22763
rect 36587 22729 36596 22763
rect 36544 22720 36596 22729
rect 36820 22720 36872 22772
rect 26700 22652 26752 22704
rect 33692 22695 33744 22704
rect 26332 22584 26384 22636
rect 26792 22584 26844 22636
rect 33692 22661 33701 22695
rect 33701 22661 33735 22695
rect 33735 22661 33744 22695
rect 33692 22652 33744 22661
rect 36912 22652 36964 22704
rect 29736 22627 29788 22636
rect 29736 22593 29745 22627
rect 29745 22593 29779 22627
rect 29779 22593 29788 22627
rect 29736 22584 29788 22593
rect 35716 22584 35768 22636
rect 23940 22559 23992 22568
rect 23940 22525 23949 22559
rect 23949 22525 23983 22559
rect 23983 22525 23992 22559
rect 23940 22516 23992 22525
rect 24032 22516 24084 22568
rect 29184 22516 29236 22568
rect 30012 22559 30064 22568
rect 30012 22525 30021 22559
rect 30021 22525 30055 22559
rect 30055 22525 30064 22559
rect 30012 22516 30064 22525
rect 36452 22516 36504 22568
rect 33140 22448 33192 22500
rect 25320 22423 25372 22432
rect 25320 22389 25329 22423
rect 25329 22389 25363 22423
rect 25363 22389 25372 22423
rect 25320 22380 25372 22389
rect 26240 22423 26292 22432
rect 26240 22389 26249 22423
rect 26249 22389 26283 22423
rect 26283 22389 26292 22423
rect 26240 22380 26292 22389
rect 26424 22423 26476 22432
rect 26424 22389 26433 22423
rect 26433 22389 26467 22423
rect 26467 22389 26476 22423
rect 26424 22380 26476 22389
rect 30380 22380 30432 22432
rect 33784 22380 33836 22432
rect 34152 22380 34204 22432
rect 34520 22448 34572 22500
rect 34888 22448 34940 22500
rect 35900 22448 35952 22500
rect 35440 22423 35492 22432
rect 35440 22389 35449 22423
rect 35449 22389 35483 22423
rect 35483 22389 35492 22423
rect 35440 22380 35492 22389
rect 35532 22380 35584 22432
rect 36544 22380 36596 22432
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 28908 22176 28960 22228
rect 29736 22219 29788 22228
rect 29736 22185 29745 22219
rect 29745 22185 29779 22219
rect 29779 22185 29788 22219
rect 29736 22176 29788 22185
rect 31760 22176 31812 22228
rect 32404 22176 32456 22228
rect 34152 22219 34204 22228
rect 34152 22185 34161 22219
rect 34161 22185 34195 22219
rect 34195 22185 34204 22219
rect 34152 22176 34204 22185
rect 35440 22176 35492 22228
rect 36820 22219 36872 22228
rect 21916 22040 21968 22092
rect 23940 22083 23992 22092
rect 23940 22049 23949 22083
rect 23949 22049 23983 22083
rect 23983 22049 23992 22083
rect 23940 22040 23992 22049
rect 24676 22083 24728 22092
rect 24676 22049 24685 22083
rect 24685 22049 24719 22083
rect 24719 22049 24728 22083
rect 24676 22040 24728 22049
rect 21824 22015 21876 22024
rect 21824 21981 21833 22015
rect 21833 21981 21867 22015
rect 21867 21981 21876 22015
rect 21824 21972 21876 21981
rect 23756 21972 23808 22024
rect 26792 22083 26844 22092
rect 26792 22049 26826 22083
rect 26826 22049 26844 22083
rect 26792 22040 26844 22049
rect 29276 22083 29328 22092
rect 29276 22049 29285 22083
rect 29285 22049 29319 22083
rect 29319 22049 29328 22083
rect 29276 22040 29328 22049
rect 30196 22040 30248 22092
rect 36820 22185 36829 22219
rect 36829 22185 36863 22219
rect 36863 22185 36872 22219
rect 36820 22176 36872 22185
rect 26516 22015 26568 22024
rect 24032 21904 24084 21956
rect 26516 21981 26525 22015
rect 26525 21981 26559 22015
rect 26559 21981 26568 22015
rect 26516 21972 26568 21981
rect 32588 22015 32640 22024
rect 32588 21981 32597 22015
rect 32597 21981 32631 22015
rect 32631 21981 32640 22015
rect 32588 21972 32640 21981
rect 32680 22015 32732 22024
rect 32680 21981 32689 22015
rect 32689 21981 32723 22015
rect 32723 21981 32732 22015
rect 34336 22015 34388 22024
rect 32680 21972 32732 21981
rect 34336 21981 34345 22015
rect 34345 21981 34379 22015
rect 34379 21981 34388 22015
rect 34336 21972 34388 21981
rect 34520 21972 34572 22024
rect 34888 21972 34940 22024
rect 23204 21879 23256 21888
rect 23204 21845 23213 21879
rect 23213 21845 23247 21879
rect 23247 21845 23256 21879
rect 23204 21836 23256 21845
rect 24308 21879 24360 21888
rect 24308 21845 24317 21879
rect 24317 21845 24351 21879
rect 24351 21845 24360 21879
rect 24308 21836 24360 21845
rect 24768 21836 24820 21888
rect 25596 21836 25648 21888
rect 26240 21836 26292 21888
rect 29184 21904 29236 21956
rect 31944 21947 31996 21956
rect 31944 21913 31953 21947
rect 31953 21913 31987 21947
rect 31987 21913 31996 21947
rect 31944 21904 31996 21913
rect 27896 21879 27948 21888
rect 27896 21845 27905 21879
rect 27905 21845 27939 21879
rect 27939 21845 27948 21879
rect 27896 21836 27948 21845
rect 30196 21879 30248 21888
rect 30196 21845 30205 21879
rect 30205 21845 30239 21879
rect 30239 21845 30248 21879
rect 30196 21836 30248 21845
rect 30656 21879 30708 21888
rect 30656 21845 30665 21879
rect 30665 21845 30699 21879
rect 30699 21845 30708 21879
rect 30656 21836 30708 21845
rect 30748 21836 30800 21888
rect 31668 21836 31720 21888
rect 32128 21879 32180 21888
rect 32128 21845 32137 21879
rect 32137 21845 32171 21879
rect 32171 21845 32180 21879
rect 32128 21836 32180 21845
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 21824 21632 21876 21684
rect 24032 21632 24084 21684
rect 21916 21539 21968 21548
rect 21916 21505 21925 21539
rect 21925 21505 21959 21539
rect 21959 21505 21968 21539
rect 21916 21496 21968 21505
rect 24676 21632 24728 21684
rect 26056 21632 26108 21684
rect 26700 21675 26752 21684
rect 26700 21641 26709 21675
rect 26709 21641 26743 21675
rect 26743 21641 26752 21675
rect 26700 21632 26752 21641
rect 30104 21675 30156 21684
rect 30104 21641 30113 21675
rect 30113 21641 30147 21675
rect 30147 21641 30156 21675
rect 30104 21632 30156 21641
rect 30380 21675 30432 21684
rect 30380 21641 30389 21675
rect 30389 21641 30423 21675
rect 30423 21641 30432 21675
rect 30380 21632 30432 21641
rect 35900 21675 35952 21684
rect 35900 21641 35909 21675
rect 35909 21641 35943 21675
rect 35943 21641 35952 21675
rect 35900 21632 35952 21641
rect 25044 21496 25096 21548
rect 20904 21471 20956 21480
rect 20904 21437 20913 21471
rect 20913 21437 20947 21471
rect 20947 21437 20956 21471
rect 20904 21428 20956 21437
rect 26240 21496 26292 21548
rect 30748 21496 30800 21548
rect 31024 21539 31076 21548
rect 31024 21505 31033 21539
rect 31033 21505 31067 21539
rect 31067 21505 31076 21539
rect 31024 21496 31076 21505
rect 35348 21539 35400 21548
rect 35348 21505 35357 21539
rect 35357 21505 35391 21539
rect 35391 21505 35400 21539
rect 35348 21496 35400 21505
rect 35440 21496 35492 21548
rect 25596 21471 25648 21480
rect 25596 21437 25605 21471
rect 25605 21437 25639 21471
rect 25639 21437 25648 21471
rect 25596 21428 25648 21437
rect 26792 21428 26844 21480
rect 30656 21428 30708 21480
rect 31300 21471 31352 21480
rect 31300 21437 31309 21471
rect 31309 21437 31343 21471
rect 31343 21437 31352 21471
rect 31300 21428 31352 21437
rect 26516 21360 26568 21412
rect 27252 21403 27304 21412
rect 27252 21369 27261 21403
rect 27261 21369 27295 21403
rect 27295 21369 27304 21403
rect 27252 21360 27304 21369
rect 21364 21335 21416 21344
rect 21364 21301 21373 21335
rect 21373 21301 21407 21335
rect 21407 21301 21416 21335
rect 21364 21292 21416 21301
rect 26976 21292 27028 21344
rect 27436 21292 27488 21344
rect 30380 21292 30432 21344
rect 31576 21292 31628 21344
rect 34520 21428 34572 21480
rect 32588 21292 32640 21344
rect 33324 21335 33376 21344
rect 33324 21301 33333 21335
rect 33333 21301 33367 21335
rect 33367 21301 33376 21335
rect 33324 21292 33376 21301
rect 34796 21292 34848 21344
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 21916 21088 21968 21140
rect 24768 21131 24820 21140
rect 24768 21097 24777 21131
rect 24777 21097 24811 21131
rect 24811 21097 24820 21131
rect 24768 21088 24820 21097
rect 25320 21088 25372 21140
rect 26240 21131 26292 21140
rect 26240 21097 26249 21131
rect 26249 21097 26283 21131
rect 26283 21097 26292 21131
rect 26240 21088 26292 21097
rect 28448 21131 28500 21140
rect 28448 21097 28457 21131
rect 28457 21097 28491 21131
rect 28491 21097 28500 21131
rect 28448 21088 28500 21097
rect 31024 21088 31076 21140
rect 31300 21088 31352 21140
rect 33048 21088 33100 21140
rect 34336 21088 34388 21140
rect 21824 21020 21876 21072
rect 23204 21020 23256 21072
rect 23480 21020 23532 21072
rect 21548 20952 21600 21004
rect 23940 20952 23992 21004
rect 32588 21020 32640 21072
rect 34612 21020 34664 21072
rect 35440 21020 35492 21072
rect 26976 20952 27028 21004
rect 30288 20995 30340 21004
rect 30288 20961 30297 20995
rect 30297 20961 30331 20995
rect 30331 20961 30340 20995
rect 30288 20952 30340 20961
rect 32404 20952 32456 21004
rect 27068 20927 27120 20936
rect 27068 20893 27077 20927
rect 27077 20893 27111 20927
rect 27111 20893 27120 20927
rect 27068 20884 27120 20893
rect 27344 20927 27396 20936
rect 27344 20893 27353 20927
rect 27353 20893 27387 20927
rect 27387 20893 27396 20927
rect 27344 20884 27396 20893
rect 29828 20884 29880 20936
rect 30748 20884 30800 20936
rect 31668 20884 31720 20936
rect 33324 20952 33376 21004
rect 32772 20927 32824 20936
rect 32772 20893 32781 20927
rect 32781 20893 32815 20927
rect 32815 20893 32824 20927
rect 32772 20884 32824 20893
rect 20076 20791 20128 20800
rect 20076 20757 20085 20791
rect 20085 20757 20119 20791
rect 20119 20757 20128 20791
rect 20076 20748 20128 20757
rect 25044 20748 25096 20800
rect 30380 20748 30432 20800
rect 32772 20748 32824 20800
rect 34336 20748 34388 20800
rect 35348 20791 35400 20800
rect 35348 20757 35357 20791
rect 35357 20757 35391 20791
rect 35391 20757 35400 20791
rect 35348 20748 35400 20757
rect 36176 20748 36228 20800
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 18328 20408 18380 20460
rect 21548 20544 21600 20596
rect 23940 20544 23992 20596
rect 20996 20476 21048 20528
rect 21824 20476 21876 20528
rect 25412 20544 25464 20596
rect 26792 20544 26844 20596
rect 30748 20587 30800 20596
rect 30748 20553 30757 20587
rect 30757 20553 30791 20587
rect 30791 20553 30800 20587
rect 30748 20544 30800 20553
rect 31300 20587 31352 20596
rect 31300 20553 31309 20587
rect 31309 20553 31343 20587
rect 31343 20553 31352 20587
rect 31300 20544 31352 20553
rect 31576 20544 31628 20596
rect 34612 20587 34664 20596
rect 34612 20553 34621 20587
rect 34621 20553 34655 20587
rect 34655 20553 34664 20587
rect 34612 20544 34664 20553
rect 26516 20476 26568 20528
rect 27896 20408 27948 20460
rect 31852 20476 31904 20528
rect 36636 20519 36688 20528
rect 36636 20485 36645 20519
rect 36645 20485 36679 20519
rect 36679 20485 36688 20519
rect 36636 20476 36688 20485
rect 32588 20451 32640 20460
rect 32588 20417 32597 20451
rect 32597 20417 32631 20451
rect 32631 20417 32640 20451
rect 32588 20408 32640 20417
rect 20076 20340 20128 20392
rect 22468 20383 22520 20392
rect 22468 20349 22477 20383
rect 22477 20349 22511 20383
rect 22511 20349 22520 20383
rect 22468 20340 22520 20349
rect 23664 20383 23716 20392
rect 23664 20349 23673 20383
rect 23673 20349 23707 20383
rect 23707 20349 23716 20383
rect 23664 20340 23716 20349
rect 25320 20383 25372 20392
rect 25320 20349 25354 20383
rect 25354 20349 25372 20383
rect 25320 20340 25372 20349
rect 26976 20340 27028 20392
rect 27528 20340 27580 20392
rect 31760 20340 31812 20392
rect 27344 20272 27396 20324
rect 28080 20272 28132 20324
rect 29460 20272 29512 20324
rect 30380 20272 30432 20324
rect 31576 20272 31628 20324
rect 21548 20204 21600 20256
rect 22652 20247 22704 20256
rect 22652 20213 22661 20247
rect 22661 20213 22695 20247
rect 22695 20213 22704 20247
rect 22652 20204 22704 20213
rect 23848 20247 23900 20256
rect 23848 20213 23857 20247
rect 23857 20213 23891 20247
rect 23891 20213 23900 20247
rect 23848 20204 23900 20213
rect 27528 20247 27580 20256
rect 27528 20213 27537 20247
rect 27537 20213 27571 20247
rect 27571 20213 27580 20247
rect 27528 20204 27580 20213
rect 27988 20247 28040 20256
rect 27988 20213 27997 20247
rect 27997 20213 28031 20247
rect 28031 20213 28040 20247
rect 27988 20204 28040 20213
rect 33692 20247 33744 20256
rect 33692 20213 33701 20247
rect 33701 20213 33735 20247
rect 33735 20213 33744 20247
rect 33692 20204 33744 20213
rect 34336 20247 34388 20256
rect 34336 20213 34345 20247
rect 34345 20213 34379 20247
rect 34379 20213 34388 20247
rect 36176 20272 36228 20324
rect 34336 20204 34388 20213
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 20076 20000 20128 20052
rect 20904 20043 20956 20052
rect 20904 20009 20913 20043
rect 20913 20009 20947 20043
rect 20947 20009 20956 20043
rect 20904 20000 20956 20009
rect 21272 20043 21324 20052
rect 21272 20009 21281 20043
rect 21281 20009 21315 20043
rect 21315 20009 21324 20043
rect 21272 20000 21324 20009
rect 17960 19864 18012 19916
rect 18052 19796 18104 19848
rect 18328 19839 18380 19848
rect 18328 19805 18337 19839
rect 18337 19805 18371 19839
rect 18371 19805 18380 19839
rect 18328 19796 18380 19805
rect 21088 19796 21140 19848
rect 22652 20000 22704 20052
rect 23480 20043 23532 20052
rect 23480 20009 23489 20043
rect 23489 20009 23523 20043
rect 23523 20009 23532 20043
rect 23480 20000 23532 20009
rect 23756 20043 23808 20052
rect 23756 20009 23765 20043
rect 23765 20009 23799 20043
rect 23799 20009 23808 20043
rect 23756 20000 23808 20009
rect 24124 20043 24176 20052
rect 24124 20009 24133 20043
rect 24133 20009 24167 20043
rect 24167 20009 24176 20043
rect 24124 20000 24176 20009
rect 24216 20043 24268 20052
rect 24216 20009 24225 20043
rect 24225 20009 24259 20043
rect 24259 20009 24268 20043
rect 24216 20000 24268 20009
rect 25320 20000 25372 20052
rect 26148 20000 26200 20052
rect 26700 20000 26752 20052
rect 27068 20000 27120 20052
rect 27804 20000 27856 20052
rect 29460 20043 29512 20052
rect 29460 20009 29469 20043
rect 29469 20009 29503 20043
rect 29503 20009 29512 20043
rect 29460 20000 29512 20009
rect 29828 20043 29880 20052
rect 29828 20009 29837 20043
rect 29837 20009 29871 20043
rect 29871 20009 29880 20043
rect 29828 20000 29880 20009
rect 30288 20000 30340 20052
rect 30748 20043 30800 20052
rect 30748 20009 30757 20043
rect 30757 20009 30791 20043
rect 30791 20009 30800 20043
rect 30748 20000 30800 20009
rect 31668 20000 31720 20052
rect 31852 20043 31904 20052
rect 31852 20009 31861 20043
rect 31861 20009 31895 20043
rect 31895 20009 31904 20043
rect 31852 20000 31904 20009
rect 33232 20000 33284 20052
rect 34612 20000 34664 20052
rect 22468 19907 22520 19916
rect 22468 19873 22477 19907
rect 22477 19873 22511 19907
rect 22511 19873 22520 19907
rect 22468 19864 22520 19873
rect 27896 19932 27948 19984
rect 35348 19932 35400 19984
rect 21548 19839 21600 19848
rect 21548 19805 21557 19839
rect 21557 19805 21591 19839
rect 21591 19805 21600 19839
rect 21548 19796 21600 19805
rect 21916 19796 21968 19848
rect 28080 19864 28132 19916
rect 32588 19907 32640 19916
rect 32588 19873 32622 19907
rect 32622 19873 32640 19907
rect 32588 19864 32640 19873
rect 26516 19796 26568 19848
rect 27068 19839 27120 19848
rect 27068 19805 27077 19839
rect 27077 19805 27111 19839
rect 27111 19805 27120 19839
rect 27068 19796 27120 19805
rect 32312 19839 32364 19848
rect 32312 19805 32321 19839
rect 32321 19805 32355 19839
rect 32355 19805 32364 19839
rect 32312 19796 32364 19805
rect 34336 19796 34388 19848
rect 34612 19796 34664 19848
rect 16580 19660 16632 19712
rect 16948 19660 17000 19712
rect 18328 19660 18380 19712
rect 19340 19660 19392 19712
rect 20628 19703 20680 19712
rect 20628 19669 20637 19703
rect 20637 19669 20671 19703
rect 20671 19669 20680 19703
rect 20628 19660 20680 19669
rect 21180 19660 21232 19712
rect 36176 19703 36228 19712
rect 36176 19669 36185 19703
rect 36185 19669 36219 19703
rect 36219 19669 36228 19703
rect 36176 19660 36228 19669
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 21088 19456 21140 19508
rect 21272 19456 21324 19508
rect 21916 19499 21968 19508
rect 21916 19465 21925 19499
rect 21925 19465 21959 19499
rect 21959 19465 21968 19499
rect 21916 19456 21968 19465
rect 24124 19456 24176 19508
rect 26332 19456 26384 19508
rect 26700 19499 26752 19508
rect 26700 19465 26709 19499
rect 26709 19465 26743 19499
rect 26743 19465 26752 19499
rect 26700 19456 26752 19465
rect 27068 19456 27120 19508
rect 27896 19456 27948 19508
rect 31760 19456 31812 19508
rect 32588 19456 32640 19508
rect 34612 19499 34664 19508
rect 34612 19465 34621 19499
rect 34621 19465 34655 19499
rect 34655 19465 34664 19499
rect 34612 19456 34664 19465
rect 35348 19456 35400 19508
rect 16672 19320 16724 19372
rect 18052 19363 18104 19372
rect 18052 19329 18061 19363
rect 18061 19329 18095 19363
rect 18095 19329 18104 19363
rect 18052 19320 18104 19329
rect 21180 19363 21232 19372
rect 16580 19252 16632 19304
rect 17960 19252 18012 19304
rect 21180 19329 21189 19363
rect 21189 19329 21223 19363
rect 21223 19329 21232 19363
rect 21180 19320 21232 19329
rect 24216 19320 24268 19372
rect 25320 19320 25372 19372
rect 27804 19320 27856 19372
rect 33876 19363 33928 19372
rect 33876 19329 33885 19363
rect 33885 19329 33919 19363
rect 33919 19329 33928 19363
rect 33876 19320 33928 19329
rect 20720 19252 20772 19304
rect 25044 19252 25096 19304
rect 25504 19295 25556 19304
rect 25504 19261 25513 19295
rect 25513 19261 25547 19295
rect 25547 19261 25556 19295
rect 25504 19252 25556 19261
rect 26056 19252 26108 19304
rect 27528 19252 27580 19304
rect 33140 19295 33192 19304
rect 33140 19261 33149 19295
rect 33149 19261 33183 19295
rect 33183 19261 33192 19295
rect 33692 19295 33744 19304
rect 33140 19252 33192 19261
rect 33692 19261 33701 19295
rect 33701 19261 33735 19295
rect 33735 19261 33744 19295
rect 33692 19252 33744 19261
rect 36176 19320 36228 19372
rect 18328 19227 18380 19236
rect 18328 19193 18362 19227
rect 18362 19193 18380 19227
rect 18328 19184 18380 19193
rect 20996 19227 21048 19236
rect 20996 19193 21005 19227
rect 21005 19193 21039 19227
rect 21039 19193 21048 19227
rect 20996 19184 21048 19193
rect 27436 19184 27488 19236
rect 15844 19159 15896 19168
rect 15844 19125 15853 19159
rect 15853 19125 15887 19159
rect 15887 19125 15896 19159
rect 15844 19116 15896 19125
rect 16396 19159 16448 19168
rect 16396 19125 16405 19159
rect 16405 19125 16439 19159
rect 16439 19125 16448 19159
rect 16396 19116 16448 19125
rect 19432 19159 19484 19168
rect 19432 19125 19441 19159
rect 19441 19125 19475 19159
rect 19475 19125 19484 19159
rect 19432 19116 19484 19125
rect 20536 19159 20588 19168
rect 20536 19125 20545 19159
rect 20545 19125 20579 19159
rect 20579 19125 20588 19159
rect 20536 19116 20588 19125
rect 22376 19159 22428 19168
rect 22376 19125 22385 19159
rect 22385 19125 22419 19159
rect 22419 19125 22428 19159
rect 22376 19116 22428 19125
rect 23112 19159 23164 19168
rect 23112 19125 23121 19159
rect 23121 19125 23155 19159
rect 23155 19125 23164 19159
rect 23112 19116 23164 19125
rect 25504 19116 25556 19168
rect 31944 19116 31996 19168
rect 32312 19159 32364 19168
rect 32312 19125 32321 19159
rect 32321 19125 32355 19159
rect 32355 19125 32364 19159
rect 35716 19184 35768 19236
rect 32312 19116 32364 19125
rect 33324 19116 33376 19168
rect 34704 19116 34756 19168
rect 35256 19116 35308 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 16396 18912 16448 18964
rect 17960 18912 18012 18964
rect 19432 18912 19484 18964
rect 20996 18912 21048 18964
rect 22468 18912 22520 18964
rect 23112 18912 23164 18964
rect 23480 18912 23532 18964
rect 25044 18955 25096 18964
rect 25044 18921 25053 18955
rect 25053 18921 25087 18955
rect 25087 18921 25096 18955
rect 25044 18912 25096 18921
rect 27528 18955 27580 18964
rect 27528 18921 27537 18955
rect 27537 18921 27571 18955
rect 27571 18921 27580 18955
rect 27528 18912 27580 18921
rect 33232 18955 33284 18964
rect 33232 18921 33241 18955
rect 33241 18921 33275 18955
rect 33275 18921 33284 18955
rect 33232 18912 33284 18921
rect 33876 18912 33928 18964
rect 35256 18955 35308 18964
rect 35256 18921 35265 18955
rect 35265 18921 35299 18955
rect 35299 18921 35308 18955
rect 35256 18912 35308 18921
rect 35716 18955 35768 18964
rect 35716 18921 35725 18955
rect 35725 18921 35759 18955
rect 35759 18921 35768 18955
rect 35716 18912 35768 18921
rect 9956 18887 10008 18896
rect 9956 18853 9990 18887
rect 9990 18853 10008 18887
rect 9956 18844 10008 18853
rect 18052 18844 18104 18896
rect 20904 18887 20956 18896
rect 20904 18853 20913 18887
rect 20913 18853 20947 18887
rect 20947 18853 20956 18887
rect 20904 18844 20956 18853
rect 27896 18844 27948 18896
rect 16212 18776 16264 18828
rect 19432 18776 19484 18828
rect 20076 18776 20128 18828
rect 22836 18776 22888 18828
rect 9680 18751 9732 18760
rect 9680 18717 9689 18751
rect 9689 18717 9723 18751
rect 9723 18717 9732 18751
rect 9680 18708 9732 18717
rect 19708 18751 19760 18760
rect 11060 18615 11112 18624
rect 11060 18581 11069 18615
rect 11069 18581 11103 18615
rect 11103 18581 11112 18615
rect 11060 18572 11112 18581
rect 14924 18615 14976 18624
rect 14924 18581 14933 18615
rect 14933 18581 14967 18615
rect 14967 18581 14976 18615
rect 14924 18572 14976 18581
rect 15936 18615 15988 18624
rect 15936 18581 15945 18615
rect 15945 18581 15979 18615
rect 15979 18581 15988 18615
rect 15936 18572 15988 18581
rect 19708 18717 19717 18751
rect 19717 18717 19751 18751
rect 19751 18717 19760 18751
rect 19708 18708 19760 18717
rect 19984 18708 20036 18760
rect 32036 18708 32088 18760
rect 19340 18640 19392 18692
rect 21824 18640 21876 18692
rect 16304 18572 16356 18624
rect 17500 18615 17552 18624
rect 17500 18581 17509 18615
rect 17509 18581 17543 18615
rect 17543 18581 17552 18615
rect 17500 18572 17552 18581
rect 22008 18615 22060 18624
rect 22008 18581 22017 18615
rect 22017 18581 22051 18615
rect 22051 18581 22060 18615
rect 22008 18572 22060 18581
rect 27160 18572 27212 18624
rect 31116 18572 31168 18624
rect 32680 18615 32732 18624
rect 32680 18581 32689 18615
rect 32689 18581 32723 18615
rect 32723 18581 32732 18615
rect 32680 18572 32732 18581
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 7380 18411 7432 18420
rect 7380 18377 7389 18411
rect 7389 18377 7423 18411
rect 7423 18377 7432 18411
rect 7380 18368 7432 18377
rect 9956 18368 10008 18420
rect 15936 18368 15988 18420
rect 16856 18368 16908 18420
rect 18052 18368 18104 18420
rect 18328 18368 18380 18420
rect 20076 18368 20128 18420
rect 20904 18411 20956 18420
rect 20904 18377 20913 18411
rect 20913 18377 20947 18411
rect 20947 18377 20956 18411
rect 20904 18368 20956 18377
rect 20996 18368 21048 18420
rect 26516 18411 26568 18420
rect 26516 18377 26525 18411
rect 26525 18377 26559 18411
rect 26559 18377 26568 18411
rect 26516 18368 26568 18377
rect 32036 18411 32088 18420
rect 32036 18377 32045 18411
rect 32045 18377 32079 18411
rect 32079 18377 32088 18411
rect 32036 18368 32088 18377
rect 7564 18207 7616 18216
rect 7564 18173 7573 18207
rect 7573 18173 7607 18207
rect 7607 18173 7616 18207
rect 7564 18164 7616 18173
rect 14924 18232 14976 18284
rect 15844 18232 15896 18284
rect 16488 18232 16540 18284
rect 16948 18275 17000 18284
rect 16948 18241 16957 18275
rect 16957 18241 16991 18275
rect 16991 18241 17000 18275
rect 16948 18232 17000 18241
rect 17868 18232 17920 18284
rect 27436 18300 27488 18352
rect 30564 18343 30616 18352
rect 30564 18309 30573 18343
rect 30573 18309 30607 18343
rect 30607 18309 30616 18343
rect 30564 18300 30616 18309
rect 21824 18275 21876 18284
rect 21824 18241 21833 18275
rect 21833 18241 21867 18275
rect 21867 18241 21876 18275
rect 21824 18232 21876 18241
rect 22008 18275 22060 18284
rect 22008 18241 22017 18275
rect 22017 18241 22051 18275
rect 22051 18241 22060 18275
rect 22008 18232 22060 18241
rect 27344 18232 27396 18284
rect 31116 18275 31168 18284
rect 31116 18241 31125 18275
rect 31125 18241 31159 18275
rect 31159 18241 31168 18275
rect 31116 18232 31168 18241
rect 16212 18164 16264 18216
rect 16396 18164 16448 18216
rect 16856 18207 16908 18216
rect 16856 18173 16865 18207
rect 16865 18173 16899 18207
rect 16899 18173 16908 18207
rect 27160 18207 27212 18216
rect 16856 18164 16908 18173
rect 27160 18173 27169 18207
rect 27169 18173 27203 18207
rect 27203 18173 27212 18207
rect 27160 18164 27212 18173
rect 17500 18096 17552 18148
rect 19340 18096 19392 18148
rect 19708 18096 19760 18148
rect 26516 18096 26568 18148
rect 30932 18139 30984 18148
rect 30932 18105 30941 18139
rect 30941 18105 30975 18139
rect 30975 18105 30984 18139
rect 30932 18096 30984 18105
rect 32956 18232 33008 18284
rect 8944 18071 8996 18080
rect 8944 18037 8953 18071
rect 8953 18037 8987 18071
rect 8987 18037 8996 18071
rect 8944 18028 8996 18037
rect 9680 18071 9732 18080
rect 9680 18037 9689 18071
rect 9689 18037 9723 18071
rect 9723 18037 9732 18071
rect 9680 18028 9732 18037
rect 15200 18071 15252 18080
rect 15200 18037 15209 18071
rect 15209 18037 15243 18071
rect 15243 18037 15252 18071
rect 15200 18028 15252 18037
rect 16304 18028 16356 18080
rect 16488 18028 16540 18080
rect 22468 18071 22520 18080
rect 22468 18037 22477 18071
rect 22477 18037 22511 18071
rect 22511 18037 22520 18071
rect 22468 18028 22520 18037
rect 22836 18071 22888 18080
rect 22836 18037 22845 18071
rect 22845 18037 22879 18071
rect 22879 18037 22888 18071
rect 22836 18028 22888 18037
rect 23388 18028 23440 18080
rect 24676 18028 24728 18080
rect 30012 18071 30064 18080
rect 30012 18037 30021 18071
rect 30021 18037 30055 18071
rect 30055 18037 30064 18071
rect 30012 18028 30064 18037
rect 31484 18028 31536 18080
rect 32220 18028 32272 18080
rect 32680 18028 32732 18080
rect 33048 18028 33100 18080
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 15108 17824 15160 17876
rect 15752 17824 15804 17876
rect 17960 17824 18012 17876
rect 18696 17824 18748 17876
rect 19340 17824 19392 17876
rect 19432 17824 19484 17876
rect 22468 17824 22520 17876
rect 30932 17867 30984 17876
rect 30932 17833 30941 17867
rect 30941 17833 30975 17867
rect 30975 17833 30984 17867
rect 30932 17824 30984 17833
rect 32956 17824 33008 17876
rect 21548 17756 21600 17808
rect 32312 17756 32364 17808
rect 16764 17731 16816 17740
rect 16764 17697 16798 17731
rect 16798 17697 16816 17731
rect 16764 17688 16816 17697
rect 18972 17731 19024 17740
rect 18972 17697 18981 17731
rect 18981 17697 19015 17731
rect 19015 17697 19024 17731
rect 18972 17688 19024 17697
rect 20720 17688 20772 17740
rect 22836 17731 22888 17740
rect 22836 17697 22845 17731
rect 22845 17697 22879 17731
rect 22879 17697 22888 17731
rect 22836 17688 22888 17697
rect 24124 17688 24176 17740
rect 27620 17688 27672 17740
rect 28080 17688 28132 17740
rect 28540 17688 28592 17740
rect 35440 17731 35492 17740
rect 35440 17697 35449 17731
rect 35449 17697 35483 17731
rect 35483 17697 35492 17731
rect 35440 17688 35492 17697
rect 16304 17620 16356 17672
rect 19984 17663 20036 17672
rect 19984 17629 19993 17663
rect 19993 17629 20027 17663
rect 20027 17629 20036 17663
rect 19984 17620 20036 17629
rect 21732 17663 21784 17672
rect 21732 17629 21741 17663
rect 21741 17629 21775 17663
rect 21775 17629 21784 17663
rect 21732 17620 21784 17629
rect 21916 17663 21968 17672
rect 21916 17629 21925 17663
rect 21925 17629 21959 17663
rect 21959 17629 21968 17663
rect 21916 17620 21968 17629
rect 24768 17663 24820 17672
rect 24768 17629 24777 17663
rect 24777 17629 24811 17663
rect 24811 17629 24820 17663
rect 24768 17620 24820 17629
rect 26608 17663 26660 17672
rect 7564 17552 7616 17604
rect 8484 17552 8536 17604
rect 24032 17552 24084 17604
rect 24676 17552 24728 17604
rect 26608 17629 26617 17663
rect 26617 17629 26651 17663
rect 26651 17629 26660 17663
rect 26608 17620 26660 17629
rect 27712 17620 27764 17672
rect 28448 17663 28500 17672
rect 28448 17629 28457 17663
rect 28457 17629 28491 17663
rect 28491 17629 28500 17663
rect 28448 17620 28500 17629
rect 32036 17620 32088 17672
rect 30288 17552 30340 17604
rect 31668 17552 31720 17604
rect 35624 17595 35676 17604
rect 35624 17561 35633 17595
rect 35633 17561 35667 17595
rect 35667 17561 35676 17595
rect 35624 17552 35676 17561
rect 8300 17484 8352 17536
rect 16212 17527 16264 17536
rect 16212 17493 16221 17527
rect 16221 17493 16255 17527
rect 16255 17493 16264 17527
rect 16212 17484 16264 17493
rect 18420 17527 18472 17536
rect 18420 17493 18429 17527
rect 18429 17493 18463 17527
rect 18463 17493 18472 17527
rect 18420 17484 18472 17493
rect 21456 17484 21508 17536
rect 24124 17527 24176 17536
rect 24124 17493 24133 17527
rect 24133 17493 24167 17527
rect 24167 17493 24176 17527
rect 24124 17484 24176 17493
rect 29828 17527 29880 17536
rect 29828 17493 29837 17527
rect 29837 17493 29871 17527
rect 29871 17493 29880 17527
rect 29828 17484 29880 17493
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 16212 17280 16264 17332
rect 19432 17280 19484 17332
rect 21732 17280 21784 17332
rect 22192 17280 22244 17332
rect 23480 17280 23532 17332
rect 24768 17280 24820 17332
rect 25136 17280 25188 17332
rect 28540 17280 28592 17332
rect 32128 17323 32180 17332
rect 32128 17289 32137 17323
rect 32137 17289 32171 17323
rect 32171 17289 32180 17323
rect 32128 17280 32180 17289
rect 18972 17212 19024 17264
rect 25412 17255 25464 17264
rect 25412 17221 25421 17255
rect 25421 17221 25455 17255
rect 25455 17221 25464 17255
rect 25412 17212 25464 17221
rect 18696 17187 18748 17196
rect 18696 17153 18705 17187
rect 18705 17153 18739 17187
rect 18739 17153 18748 17187
rect 18696 17144 18748 17153
rect 21456 17187 21508 17196
rect 21456 17153 21465 17187
rect 21465 17153 21499 17187
rect 21499 17153 21508 17187
rect 21456 17144 21508 17153
rect 21548 17187 21600 17196
rect 21548 17153 21557 17187
rect 21557 17153 21591 17187
rect 21591 17153 21600 17187
rect 21548 17144 21600 17153
rect 24032 17144 24084 17196
rect 27988 17212 28040 17264
rect 33140 17280 33192 17332
rect 35440 17323 35492 17332
rect 35440 17289 35449 17323
rect 35449 17289 35483 17323
rect 35483 17289 35492 17323
rect 35440 17280 35492 17289
rect 8484 17076 8536 17128
rect 15476 17119 15528 17128
rect 15476 17085 15485 17119
rect 15485 17085 15519 17119
rect 15519 17085 15528 17119
rect 15476 17076 15528 17085
rect 15752 17119 15804 17128
rect 15752 17085 15786 17119
rect 15786 17085 15804 17119
rect 15752 17076 15804 17085
rect 19892 17076 19944 17128
rect 23480 17076 23532 17128
rect 33416 17144 33468 17196
rect 35256 17212 35308 17264
rect 35624 17212 35676 17264
rect 29736 17076 29788 17128
rect 30288 17119 30340 17128
rect 30288 17085 30297 17119
rect 30297 17085 30331 17119
rect 30331 17085 30340 17119
rect 30288 17076 30340 17085
rect 8300 17008 8352 17060
rect 16304 17008 16356 17060
rect 16580 17008 16632 17060
rect 23664 17008 23716 17060
rect 25688 17008 25740 17060
rect 27620 17008 27672 17060
rect 28448 17008 28500 17060
rect 29828 17008 29880 17060
rect 31668 17076 31720 17128
rect 32220 17076 32272 17128
rect 33876 17187 33928 17196
rect 33876 17153 33885 17187
rect 33885 17153 33919 17187
rect 33919 17153 33928 17187
rect 33876 17144 33928 17153
rect 8392 16940 8444 16992
rect 15384 16940 15436 16992
rect 16764 16940 16816 16992
rect 18236 16940 18288 16992
rect 18420 16983 18472 16992
rect 18420 16949 18429 16983
rect 18429 16949 18463 16983
rect 18463 16949 18472 16983
rect 18420 16940 18472 16949
rect 20720 16940 20772 16992
rect 20996 16983 21048 16992
rect 20996 16949 21005 16983
rect 21005 16949 21039 16983
rect 21039 16949 21048 16983
rect 20996 16940 21048 16949
rect 21272 16940 21324 16992
rect 27712 16983 27764 16992
rect 27712 16949 27721 16983
rect 27721 16949 27755 16983
rect 27755 16949 27764 16983
rect 27712 16940 27764 16949
rect 27988 16983 28040 16992
rect 27988 16949 27997 16983
rect 27997 16949 28031 16983
rect 28031 16949 28040 16983
rect 27988 16940 28040 16949
rect 32128 16940 32180 16992
rect 33048 16940 33100 16992
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 5448 16779 5500 16788
rect 5448 16745 5457 16779
rect 5457 16745 5491 16779
rect 5491 16745 5500 16779
rect 5448 16736 5500 16745
rect 8116 16736 8168 16788
rect 8392 16779 8444 16788
rect 6000 16668 6052 16720
rect 7932 16711 7984 16720
rect 7932 16677 7941 16711
rect 7941 16677 7975 16711
rect 7975 16677 7984 16711
rect 8392 16745 8401 16779
rect 8401 16745 8435 16779
rect 8435 16745 8444 16779
rect 8392 16736 8444 16745
rect 11060 16779 11112 16788
rect 11060 16745 11069 16779
rect 11069 16745 11103 16779
rect 11103 16745 11112 16779
rect 11060 16736 11112 16745
rect 15292 16779 15344 16788
rect 15292 16745 15301 16779
rect 15301 16745 15335 16779
rect 15335 16745 15344 16779
rect 15292 16736 15344 16745
rect 15752 16736 15804 16788
rect 16304 16736 16356 16788
rect 16856 16736 16908 16788
rect 18236 16779 18288 16788
rect 18236 16745 18245 16779
rect 18245 16745 18279 16779
rect 18279 16745 18288 16779
rect 18236 16736 18288 16745
rect 20996 16736 21048 16788
rect 22836 16736 22888 16788
rect 23480 16779 23532 16788
rect 23480 16745 23489 16779
rect 23489 16745 23523 16779
rect 23523 16745 23532 16779
rect 23480 16736 23532 16745
rect 25688 16779 25740 16788
rect 25688 16745 25697 16779
rect 25697 16745 25731 16779
rect 25731 16745 25740 16779
rect 25688 16736 25740 16745
rect 27344 16736 27396 16788
rect 29368 16779 29420 16788
rect 29368 16745 29377 16779
rect 29377 16745 29411 16779
rect 29411 16745 29420 16779
rect 29368 16736 29420 16745
rect 7932 16668 7984 16677
rect 8300 16668 8352 16720
rect 9588 16668 9640 16720
rect 20720 16668 20772 16720
rect 6276 16600 6328 16652
rect 9772 16600 9824 16652
rect 10968 16600 11020 16652
rect 16764 16600 16816 16652
rect 20812 16600 20864 16652
rect 21916 16600 21968 16652
rect 24400 16668 24452 16720
rect 25412 16668 25464 16720
rect 29920 16668 29972 16720
rect 30288 16668 30340 16720
rect 31116 16736 31168 16788
rect 32312 16736 32364 16788
rect 33876 16736 33928 16788
rect 24124 16600 24176 16652
rect 5264 16532 5316 16584
rect 9680 16575 9732 16584
rect 9680 16541 9689 16575
rect 9689 16541 9723 16575
rect 9723 16541 9732 16575
rect 9680 16532 9732 16541
rect 15384 16532 15436 16584
rect 16120 16532 16172 16584
rect 16672 16532 16724 16584
rect 8484 16464 8536 16516
rect 5356 16439 5408 16448
rect 5356 16405 5365 16439
rect 5365 16405 5399 16439
rect 5399 16405 5408 16439
rect 5356 16396 5408 16405
rect 7196 16439 7248 16448
rect 7196 16405 7205 16439
rect 7205 16405 7239 16439
rect 7239 16405 7248 16439
rect 7196 16396 7248 16405
rect 7472 16439 7524 16448
rect 7472 16405 7481 16439
rect 7481 16405 7515 16439
rect 7515 16405 7524 16439
rect 7472 16396 7524 16405
rect 16856 16575 16908 16584
rect 16856 16541 16865 16575
rect 16865 16541 16899 16575
rect 16899 16541 16908 16575
rect 21088 16575 21140 16584
rect 16856 16532 16908 16541
rect 21088 16541 21097 16575
rect 21097 16541 21131 16575
rect 21131 16541 21140 16575
rect 21088 16532 21140 16541
rect 26332 16600 26384 16652
rect 27252 16600 27304 16652
rect 29552 16643 29604 16652
rect 29552 16609 29561 16643
rect 29561 16609 29595 16643
rect 29595 16609 29604 16643
rect 29552 16600 29604 16609
rect 30380 16600 30432 16652
rect 32128 16643 32180 16652
rect 26516 16575 26568 16584
rect 26516 16541 26525 16575
rect 26525 16541 26559 16575
rect 26559 16541 26568 16575
rect 26516 16532 26568 16541
rect 30932 16532 30984 16584
rect 32128 16609 32137 16643
rect 32137 16609 32171 16643
rect 32171 16609 32180 16643
rect 32128 16600 32180 16609
rect 33232 16532 33284 16584
rect 17040 16396 17092 16448
rect 18788 16439 18840 16448
rect 18788 16405 18797 16439
rect 18797 16405 18831 16439
rect 18831 16405 18840 16439
rect 18788 16396 18840 16405
rect 22100 16396 22152 16448
rect 24768 16396 24820 16448
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 5448 16192 5500 16244
rect 8484 16235 8536 16244
rect 8484 16201 8493 16235
rect 8493 16201 8527 16235
rect 8527 16201 8536 16235
rect 8484 16192 8536 16201
rect 9680 16192 9732 16244
rect 10968 16192 11020 16244
rect 15384 16235 15436 16244
rect 15384 16201 15393 16235
rect 15393 16201 15427 16235
rect 15427 16201 15436 16235
rect 15384 16192 15436 16201
rect 15752 16235 15804 16244
rect 15752 16201 15761 16235
rect 15761 16201 15795 16235
rect 15795 16201 15804 16235
rect 15752 16192 15804 16201
rect 16488 16192 16540 16244
rect 18052 16192 18104 16244
rect 21088 16192 21140 16244
rect 22192 16192 22244 16244
rect 23480 16192 23532 16244
rect 24400 16235 24452 16244
rect 24400 16201 24409 16235
rect 24409 16201 24443 16235
rect 24443 16201 24452 16235
rect 24400 16192 24452 16201
rect 26240 16235 26292 16244
rect 7472 16124 7524 16176
rect 5356 16056 5408 16108
rect 6644 16056 6696 16108
rect 7564 16099 7616 16108
rect 7564 16065 7573 16099
rect 7573 16065 7607 16099
rect 7607 16065 7616 16099
rect 7564 16056 7616 16065
rect 16120 16124 16172 16176
rect 17040 16099 17092 16108
rect 7196 15988 7248 16040
rect 8484 15988 8536 16040
rect 17040 16065 17049 16099
rect 17049 16065 17083 16099
rect 17083 16065 17092 16099
rect 17040 16056 17092 16065
rect 26240 16201 26249 16235
rect 26249 16201 26283 16235
rect 26283 16201 26292 16235
rect 26240 16192 26292 16201
rect 26608 16192 26660 16244
rect 26516 16124 26568 16176
rect 27528 16124 27580 16176
rect 9220 15988 9272 16040
rect 18788 15988 18840 16040
rect 23756 16031 23808 16040
rect 23756 15997 23765 16031
rect 23765 15997 23799 16031
rect 23799 15997 23808 16031
rect 23756 15988 23808 15997
rect 25136 16031 25188 16040
rect 25136 15997 25170 16031
rect 25170 15997 25188 16031
rect 25136 15988 25188 15997
rect 30012 16192 30064 16244
rect 30380 16235 30432 16244
rect 30380 16201 30389 16235
rect 30389 16201 30423 16235
rect 30423 16201 30432 16235
rect 30380 16192 30432 16201
rect 32312 16235 32364 16244
rect 32312 16201 32321 16235
rect 32321 16201 32355 16235
rect 32355 16201 32364 16235
rect 32312 16192 32364 16201
rect 33232 16235 33284 16244
rect 33232 16201 33241 16235
rect 33241 16201 33275 16235
rect 33275 16201 33284 16235
rect 33232 16192 33284 16201
rect 27896 16099 27948 16108
rect 27896 16065 27905 16099
rect 27905 16065 27939 16099
rect 27939 16065 27948 16099
rect 27896 16056 27948 16065
rect 29828 16099 29880 16108
rect 29828 16065 29837 16099
rect 29837 16065 29871 16099
rect 29871 16065 29880 16099
rect 29828 16056 29880 16065
rect 30288 16056 30340 16108
rect 30932 16099 30984 16108
rect 30932 16065 30941 16099
rect 30941 16065 30975 16099
rect 30975 16065 30984 16099
rect 30932 16056 30984 16065
rect 29368 15988 29420 16040
rect 30196 15988 30248 16040
rect 17500 15920 17552 15972
rect 22284 15920 22336 15972
rect 27620 15920 27672 15972
rect 31116 15920 31168 15972
rect 4804 15895 4856 15904
rect 4804 15861 4813 15895
rect 4813 15861 4847 15895
rect 4847 15861 4856 15895
rect 4804 15852 4856 15861
rect 5264 15895 5316 15904
rect 5264 15861 5273 15895
rect 5273 15861 5307 15895
rect 5307 15861 5316 15895
rect 5264 15852 5316 15861
rect 6000 15895 6052 15904
rect 6000 15861 6009 15895
rect 6009 15861 6043 15895
rect 6043 15861 6052 15895
rect 6000 15852 6052 15861
rect 6276 15895 6328 15904
rect 6276 15861 6285 15895
rect 6285 15861 6319 15895
rect 6319 15861 6328 15895
rect 6276 15852 6328 15861
rect 7104 15895 7156 15904
rect 7104 15861 7113 15895
rect 7113 15861 7147 15895
rect 7147 15861 7156 15895
rect 7104 15852 7156 15861
rect 16764 15895 16816 15904
rect 16764 15861 16773 15895
rect 16773 15861 16807 15895
rect 16807 15861 16816 15895
rect 16764 15852 16816 15861
rect 17224 15852 17276 15904
rect 19432 15895 19484 15904
rect 19432 15861 19441 15895
rect 19441 15861 19475 15895
rect 19475 15861 19484 15895
rect 19432 15852 19484 15861
rect 33048 15852 33100 15904
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 7104 15648 7156 15700
rect 8024 15648 8076 15700
rect 9772 15648 9824 15700
rect 16120 15691 16172 15700
rect 16120 15657 16129 15691
rect 16129 15657 16163 15691
rect 16163 15657 16172 15691
rect 16120 15648 16172 15657
rect 16764 15648 16816 15700
rect 20720 15691 20772 15700
rect 20720 15657 20729 15691
rect 20729 15657 20763 15691
rect 20763 15657 20772 15691
rect 20720 15648 20772 15657
rect 26332 15691 26384 15700
rect 26332 15657 26341 15691
rect 26341 15657 26375 15691
rect 26375 15657 26384 15691
rect 26332 15648 26384 15657
rect 27896 15691 27948 15700
rect 27896 15657 27905 15691
rect 27905 15657 27939 15691
rect 27939 15657 27948 15691
rect 27896 15648 27948 15657
rect 30288 15648 30340 15700
rect 33416 15691 33468 15700
rect 33416 15657 33425 15691
rect 33425 15657 33459 15691
rect 33459 15657 33468 15691
rect 33416 15648 33468 15657
rect 36544 15691 36596 15700
rect 36544 15657 36553 15691
rect 36553 15657 36587 15691
rect 36587 15657 36596 15691
rect 36544 15648 36596 15657
rect 7564 15580 7616 15632
rect 8208 15580 8260 15632
rect 17500 15623 17552 15632
rect 17500 15589 17534 15623
rect 17534 15589 17552 15623
rect 17500 15580 17552 15589
rect 6000 15512 6052 15564
rect 8300 15512 8352 15564
rect 20720 15512 20772 15564
rect 22192 15512 22244 15564
rect 24400 15580 24452 15632
rect 26976 15580 27028 15632
rect 27344 15580 27396 15632
rect 24032 15512 24084 15564
rect 26516 15555 26568 15564
rect 26516 15521 26525 15555
rect 26525 15521 26559 15555
rect 26559 15521 26568 15555
rect 26516 15512 26568 15521
rect 30564 15555 30616 15564
rect 30564 15521 30573 15555
rect 30573 15521 30607 15555
rect 30607 15521 30616 15555
rect 30564 15512 30616 15521
rect 31668 15555 31720 15564
rect 31668 15521 31677 15555
rect 31677 15521 31711 15555
rect 31711 15521 31720 15555
rect 31668 15512 31720 15521
rect 32128 15555 32180 15564
rect 32128 15521 32137 15555
rect 32137 15521 32171 15555
rect 32171 15521 32180 15555
rect 32128 15512 32180 15521
rect 33232 15555 33284 15564
rect 33232 15521 33241 15555
rect 33241 15521 33275 15555
rect 33275 15521 33284 15555
rect 33232 15512 33284 15521
rect 35256 15512 35308 15564
rect 35900 15512 35952 15564
rect 4988 15487 5040 15496
rect 4988 15453 4997 15487
rect 4997 15453 5031 15487
rect 5031 15453 5040 15487
rect 4988 15444 5040 15453
rect 8668 15487 8720 15496
rect 8668 15453 8677 15487
rect 8677 15453 8711 15487
rect 8711 15453 8720 15487
rect 8668 15444 8720 15453
rect 17224 15487 17276 15496
rect 17224 15453 17233 15487
rect 17233 15453 17267 15487
rect 17267 15453 17276 15487
rect 17224 15444 17276 15453
rect 21088 15487 21140 15496
rect 21088 15453 21097 15487
rect 21097 15453 21131 15487
rect 21131 15453 21140 15487
rect 21088 15444 21140 15453
rect 30656 15487 30708 15496
rect 30656 15453 30665 15487
rect 30665 15453 30699 15487
rect 30699 15453 30708 15487
rect 30656 15444 30708 15453
rect 29920 15376 29972 15428
rect 31392 15444 31444 15496
rect 4620 15308 4672 15360
rect 6276 15308 6328 15360
rect 6644 15308 6696 15360
rect 8300 15308 8352 15360
rect 14556 15308 14608 15360
rect 24124 15308 24176 15360
rect 30196 15351 30248 15360
rect 30196 15317 30205 15351
rect 30205 15317 30239 15351
rect 30239 15317 30248 15351
rect 30196 15308 30248 15317
rect 31760 15308 31812 15360
rect 33692 15308 33744 15360
rect 35348 15308 35400 15360
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 8116 15104 8168 15156
rect 17500 15104 17552 15156
rect 20628 15147 20680 15156
rect 20628 15113 20637 15147
rect 20637 15113 20671 15147
rect 20671 15113 20680 15147
rect 20628 15104 20680 15113
rect 21088 15104 21140 15156
rect 23664 15147 23716 15156
rect 23664 15113 23673 15147
rect 23673 15113 23707 15147
rect 23707 15113 23716 15147
rect 23664 15104 23716 15113
rect 24400 15104 24452 15156
rect 26056 15147 26108 15156
rect 26056 15113 26065 15147
rect 26065 15113 26099 15147
rect 26099 15113 26108 15147
rect 26056 15104 26108 15113
rect 26516 15147 26568 15156
rect 26516 15113 26525 15147
rect 26525 15113 26559 15147
rect 26559 15113 26568 15147
rect 26516 15104 26568 15113
rect 26976 15147 27028 15156
rect 26976 15113 26985 15147
rect 26985 15113 27019 15147
rect 27019 15113 27028 15147
rect 26976 15104 27028 15113
rect 27436 15147 27488 15156
rect 27436 15113 27445 15147
rect 27445 15113 27479 15147
rect 27479 15113 27488 15147
rect 27436 15104 27488 15113
rect 29920 15147 29972 15156
rect 29920 15113 29929 15147
rect 29929 15113 29963 15147
rect 29963 15113 29972 15147
rect 29920 15104 29972 15113
rect 30564 15147 30616 15156
rect 30564 15113 30573 15147
rect 30573 15113 30607 15147
rect 30607 15113 30616 15147
rect 30564 15104 30616 15113
rect 30932 15147 30984 15156
rect 30932 15113 30941 15147
rect 30941 15113 30975 15147
rect 30975 15113 30984 15147
rect 30932 15104 30984 15113
rect 31392 15104 31444 15156
rect 14556 15011 14608 15020
rect 14556 14977 14565 15011
rect 14565 14977 14599 15011
rect 14599 14977 14608 15011
rect 14556 14968 14608 14977
rect 22376 15036 22428 15088
rect 24124 15011 24176 15020
rect 24124 14977 24133 15011
rect 24133 14977 24167 15011
rect 24167 14977 24176 15011
rect 24124 14968 24176 14977
rect 24676 15036 24728 15088
rect 24308 14968 24360 15020
rect 4252 14943 4304 14952
rect 4252 14909 4261 14943
rect 4261 14909 4295 14943
rect 4295 14909 4304 14943
rect 4252 14900 4304 14909
rect 4988 14900 5040 14952
rect 8484 14900 8536 14952
rect 4620 14832 4672 14884
rect 6000 14832 6052 14884
rect 5632 14807 5684 14816
rect 5632 14773 5641 14807
rect 5641 14773 5675 14807
rect 5675 14773 5684 14807
rect 5632 14764 5684 14773
rect 7932 14832 7984 14884
rect 14096 14832 14148 14884
rect 13912 14807 13964 14816
rect 13912 14773 13921 14807
rect 13921 14773 13955 14807
rect 13955 14773 13964 14807
rect 13912 14764 13964 14773
rect 22284 14900 22336 14952
rect 24768 14900 24820 14952
rect 26056 14900 26108 14952
rect 31668 14900 31720 14952
rect 33692 14943 33744 14952
rect 33692 14909 33701 14943
rect 33701 14909 33735 14943
rect 33735 14909 33744 14943
rect 33692 14900 33744 14909
rect 35348 15104 35400 15156
rect 21732 14832 21784 14884
rect 30656 14832 30708 14884
rect 33048 14832 33100 14884
rect 15108 14764 15160 14816
rect 15476 14764 15528 14816
rect 17224 14807 17276 14816
rect 17224 14773 17233 14807
rect 17233 14773 17267 14807
rect 17267 14773 17276 14807
rect 17224 14764 17276 14773
rect 21640 14764 21692 14816
rect 32496 14764 32548 14816
rect 33232 14807 33284 14816
rect 33232 14773 33241 14807
rect 33241 14773 33275 14807
rect 33275 14773 33284 14807
rect 33232 14764 33284 14773
rect 33876 14807 33928 14816
rect 33876 14773 33885 14807
rect 33885 14773 33919 14807
rect 33919 14773 33928 14807
rect 33876 14764 33928 14773
rect 34152 14764 34204 14816
rect 35256 14832 35308 14884
rect 35900 14764 35952 14816
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 7012 14560 7064 14612
rect 7380 14560 7432 14612
rect 7932 14560 7984 14612
rect 8024 14560 8076 14612
rect 8668 14560 8720 14612
rect 13912 14560 13964 14612
rect 14924 14560 14976 14612
rect 21088 14603 21140 14612
rect 21088 14569 21097 14603
rect 21097 14569 21131 14603
rect 21131 14569 21140 14603
rect 21088 14560 21140 14569
rect 21272 14603 21324 14612
rect 21272 14569 21281 14603
rect 21281 14569 21315 14603
rect 21315 14569 21324 14603
rect 21272 14560 21324 14569
rect 21732 14603 21784 14612
rect 21732 14569 21741 14603
rect 21741 14569 21775 14603
rect 21775 14569 21784 14603
rect 21732 14560 21784 14569
rect 22008 14560 22060 14612
rect 24032 14603 24084 14612
rect 24032 14569 24041 14603
rect 24041 14569 24075 14603
rect 24075 14569 24084 14603
rect 24032 14560 24084 14569
rect 24308 14603 24360 14612
rect 24308 14569 24317 14603
rect 24317 14569 24351 14603
rect 24351 14569 24360 14603
rect 24308 14560 24360 14569
rect 30472 14560 30524 14612
rect 30564 14560 30616 14612
rect 32128 14603 32180 14612
rect 21640 14535 21692 14544
rect 21640 14501 21649 14535
rect 21649 14501 21683 14535
rect 21683 14501 21692 14535
rect 21640 14492 21692 14501
rect 32128 14569 32137 14603
rect 32137 14569 32171 14603
rect 32171 14569 32180 14603
rect 32128 14560 32180 14569
rect 32496 14603 32548 14612
rect 32496 14569 32505 14603
rect 32505 14569 32539 14603
rect 32539 14569 32548 14603
rect 32496 14560 32548 14569
rect 35900 14603 35952 14612
rect 35900 14569 35909 14603
rect 35909 14569 35943 14603
rect 35943 14569 35952 14603
rect 35900 14560 35952 14569
rect 36820 14603 36872 14612
rect 36820 14569 36829 14603
rect 36829 14569 36863 14603
rect 36863 14569 36872 14603
rect 36820 14560 36872 14569
rect 33416 14492 33468 14544
rect 3516 14424 3568 14476
rect 4804 14424 4856 14476
rect 5632 14424 5684 14476
rect 7104 14467 7156 14476
rect 7104 14433 7113 14467
rect 7113 14433 7147 14467
rect 7147 14433 7156 14467
rect 7104 14424 7156 14433
rect 8300 14467 8352 14476
rect 8300 14433 8309 14467
rect 8309 14433 8343 14467
rect 8343 14433 8352 14467
rect 8300 14424 8352 14433
rect 9864 14467 9916 14476
rect 9864 14433 9873 14467
rect 9873 14433 9907 14467
rect 9907 14433 9916 14467
rect 9864 14424 9916 14433
rect 11244 14424 11296 14476
rect 12532 14467 12584 14476
rect 12532 14433 12541 14467
rect 12541 14433 12575 14467
rect 12575 14433 12584 14467
rect 12532 14424 12584 14433
rect 12624 14424 12676 14476
rect 3884 14356 3936 14408
rect 4252 14399 4304 14408
rect 4252 14365 4261 14399
rect 4261 14365 4295 14399
rect 4295 14365 4304 14399
rect 4252 14356 4304 14365
rect 6276 14356 6328 14408
rect 8668 14356 8720 14408
rect 11152 14356 11204 14408
rect 22376 14424 22428 14476
rect 29092 14424 29144 14476
rect 30840 14467 30892 14476
rect 5264 14220 5316 14272
rect 5632 14263 5684 14272
rect 5632 14229 5641 14263
rect 5641 14229 5675 14263
rect 5675 14229 5684 14263
rect 5632 14220 5684 14229
rect 6736 14263 6788 14272
rect 6736 14229 6745 14263
rect 6745 14229 6779 14263
rect 6779 14229 6788 14263
rect 6736 14220 6788 14229
rect 8484 14263 8536 14272
rect 8484 14229 8493 14263
rect 8493 14229 8527 14263
rect 8527 14229 8536 14263
rect 8484 14220 8536 14229
rect 10048 14263 10100 14272
rect 10048 14229 10057 14263
rect 10057 14229 10091 14263
rect 10091 14229 10100 14263
rect 10048 14220 10100 14229
rect 10784 14263 10836 14272
rect 10784 14229 10793 14263
rect 10793 14229 10827 14263
rect 10827 14229 10836 14263
rect 10784 14220 10836 14229
rect 13452 14220 13504 14272
rect 19340 14220 19392 14272
rect 26976 14263 27028 14272
rect 26976 14229 26985 14263
rect 26985 14229 27019 14263
rect 27019 14229 27028 14263
rect 26976 14220 27028 14229
rect 29552 14263 29604 14272
rect 29552 14229 29561 14263
rect 29561 14229 29595 14263
rect 29595 14229 29604 14263
rect 29552 14220 29604 14229
rect 30840 14433 30849 14467
rect 30849 14433 30883 14467
rect 30883 14433 30892 14467
rect 30840 14424 30892 14433
rect 32588 14467 32640 14476
rect 32588 14433 32597 14467
rect 32597 14433 32631 14467
rect 32631 14433 32640 14467
rect 32588 14424 32640 14433
rect 33784 14424 33836 14476
rect 34520 14424 34572 14476
rect 35256 14467 35308 14476
rect 35256 14433 35265 14467
rect 35265 14433 35299 14467
rect 35299 14433 35308 14467
rect 35256 14424 35308 14433
rect 37096 14492 37148 14544
rect 36544 14424 36596 14476
rect 30564 14356 30616 14408
rect 33876 14356 33928 14408
rect 35348 14399 35400 14408
rect 35348 14365 35357 14399
rect 35357 14365 35391 14399
rect 35391 14365 35400 14399
rect 35348 14356 35400 14365
rect 34520 14288 34572 14340
rect 31300 14220 31352 14272
rect 33324 14263 33376 14272
rect 33324 14229 33333 14263
rect 33333 14229 33367 14263
rect 33367 14229 33376 14263
rect 33324 14220 33376 14229
rect 33416 14220 33468 14272
rect 34060 14220 34112 14272
rect 35440 14220 35492 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 3516 14059 3568 14068
rect 3516 14025 3525 14059
rect 3525 14025 3559 14059
rect 3559 14025 3568 14059
rect 3516 14016 3568 14025
rect 3884 14059 3936 14068
rect 3884 14025 3893 14059
rect 3893 14025 3927 14059
rect 3927 14025 3936 14059
rect 3884 14016 3936 14025
rect 5540 14016 5592 14068
rect 7104 14016 7156 14068
rect 7380 14059 7432 14068
rect 7380 14025 7389 14059
rect 7389 14025 7423 14059
rect 7423 14025 7432 14059
rect 7380 14016 7432 14025
rect 6276 13991 6328 14000
rect 6276 13957 6285 13991
rect 6285 13957 6319 13991
rect 6319 13957 6328 13991
rect 6276 13948 6328 13957
rect 3884 13812 3936 13864
rect 5632 13812 5684 13864
rect 6736 13812 6788 13864
rect 6920 13812 6972 13864
rect 8484 14016 8536 14068
rect 11152 14016 11204 14068
rect 12532 14016 12584 14068
rect 8668 13812 8720 13864
rect 9496 13812 9548 13864
rect 9864 13855 9916 13864
rect 9864 13821 9873 13855
rect 9873 13821 9907 13855
rect 9907 13821 9916 13855
rect 9864 13812 9916 13821
rect 10876 13880 10928 13932
rect 14372 14016 14424 14068
rect 21732 14016 21784 14068
rect 22376 14016 22428 14068
rect 26700 14059 26752 14068
rect 26700 14025 26709 14059
rect 26709 14025 26743 14059
rect 26743 14025 26752 14059
rect 26700 14016 26752 14025
rect 29092 14059 29144 14068
rect 29092 14025 29101 14059
rect 29101 14025 29135 14059
rect 29135 14025 29144 14059
rect 29092 14016 29144 14025
rect 30564 14059 30616 14068
rect 30564 14025 30573 14059
rect 30573 14025 30607 14059
rect 30607 14025 30616 14059
rect 30564 14016 30616 14025
rect 30656 14016 30708 14068
rect 31300 14016 31352 14068
rect 32588 14016 32640 14068
rect 35256 14016 35308 14068
rect 37096 14059 37148 14068
rect 37096 14025 37105 14059
rect 37105 14025 37139 14059
rect 37139 14025 37148 14059
rect 37096 14016 37148 14025
rect 21640 13991 21692 14000
rect 21640 13957 21649 13991
rect 21649 13957 21683 13991
rect 21683 13957 21692 13991
rect 21640 13948 21692 13957
rect 25596 13991 25648 14000
rect 25596 13957 25605 13991
rect 25605 13957 25639 13991
rect 25639 13957 25648 13991
rect 25596 13948 25648 13957
rect 29552 13948 29604 14000
rect 13452 13923 13504 13932
rect 11152 13855 11204 13864
rect 11152 13821 11161 13855
rect 11161 13821 11195 13855
rect 11195 13821 11204 13855
rect 11152 13812 11204 13821
rect 13452 13889 13461 13923
rect 13461 13889 13495 13923
rect 13495 13889 13504 13923
rect 13452 13880 13504 13889
rect 12532 13812 12584 13864
rect 14648 13812 14700 13864
rect 14924 13880 14976 13932
rect 27436 13923 27488 13932
rect 27436 13889 27445 13923
rect 27445 13889 27479 13923
rect 27479 13889 27488 13923
rect 27436 13880 27488 13889
rect 18604 13855 18656 13864
rect 12440 13744 12492 13796
rect 18604 13821 18613 13855
rect 18613 13821 18647 13855
rect 18647 13821 18656 13855
rect 18604 13812 18656 13821
rect 19432 13812 19484 13864
rect 16120 13744 16172 13796
rect 19340 13744 19392 13796
rect 25688 13744 25740 13796
rect 26976 13812 27028 13864
rect 29000 13812 29052 13864
rect 30840 13812 30892 13864
rect 31576 13948 31628 14000
rect 33876 13991 33928 14000
rect 31668 13923 31720 13932
rect 31668 13889 31677 13923
rect 31677 13889 31711 13923
rect 31711 13889 31720 13923
rect 31668 13880 31720 13889
rect 33876 13957 33885 13991
rect 33885 13957 33919 13991
rect 33919 13957 33928 13991
rect 33876 13948 33928 13957
rect 33416 13923 33468 13932
rect 33416 13889 33425 13923
rect 33425 13889 33459 13923
rect 33459 13889 33468 13923
rect 33416 13880 33468 13889
rect 34152 13812 34204 13864
rect 35348 13855 35400 13864
rect 35348 13821 35382 13855
rect 35382 13821 35400 13855
rect 26700 13744 26752 13796
rect 32404 13744 32456 13796
rect 5080 13676 5132 13728
rect 9956 13676 10008 13728
rect 10784 13676 10836 13728
rect 12808 13719 12860 13728
rect 12808 13685 12817 13719
rect 12817 13685 12851 13719
rect 12851 13685 12860 13719
rect 12808 13676 12860 13685
rect 13268 13676 13320 13728
rect 13912 13676 13964 13728
rect 19156 13719 19208 13728
rect 19156 13685 19165 13719
rect 19165 13685 19199 13719
rect 19199 13685 19208 13719
rect 19156 13676 19208 13685
rect 26884 13719 26936 13728
rect 26884 13685 26893 13719
rect 26893 13685 26927 13719
rect 26927 13685 26936 13719
rect 26884 13676 26936 13685
rect 31944 13676 31996 13728
rect 32496 13676 32548 13728
rect 33140 13719 33192 13728
rect 33140 13685 33149 13719
rect 33149 13685 33183 13719
rect 33183 13685 33192 13719
rect 33140 13676 33192 13685
rect 35348 13812 35400 13821
rect 35900 13744 35952 13796
rect 35256 13676 35308 13728
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 3884 13472 3936 13524
rect 5080 13515 5132 13524
rect 5080 13481 5089 13515
rect 5089 13481 5123 13515
rect 5123 13481 5132 13515
rect 5080 13472 5132 13481
rect 6920 13515 6972 13524
rect 6920 13481 6929 13515
rect 6929 13481 6963 13515
rect 6963 13481 6972 13515
rect 6920 13472 6972 13481
rect 8300 13515 8352 13524
rect 8300 13481 8309 13515
rect 8309 13481 8343 13515
rect 8343 13481 8352 13515
rect 8300 13472 8352 13481
rect 9864 13472 9916 13524
rect 10048 13515 10100 13524
rect 10048 13481 10057 13515
rect 10057 13481 10091 13515
rect 10091 13481 10100 13515
rect 10048 13472 10100 13481
rect 10876 13515 10928 13524
rect 10876 13481 10885 13515
rect 10885 13481 10919 13515
rect 10919 13481 10928 13515
rect 10876 13472 10928 13481
rect 12624 13515 12676 13524
rect 12624 13481 12633 13515
rect 12633 13481 12667 13515
rect 12667 13481 12676 13515
rect 12624 13472 12676 13481
rect 13452 13472 13504 13524
rect 14096 13515 14148 13524
rect 14096 13481 14105 13515
rect 14105 13481 14139 13515
rect 14139 13481 14148 13515
rect 14096 13472 14148 13481
rect 16672 13515 16724 13524
rect 16672 13481 16681 13515
rect 16681 13481 16715 13515
rect 16715 13481 16724 13515
rect 16672 13472 16724 13481
rect 19156 13472 19208 13524
rect 26976 13472 27028 13524
rect 29000 13515 29052 13524
rect 29000 13481 29009 13515
rect 29009 13481 29043 13515
rect 29043 13481 29052 13515
rect 29000 13472 29052 13481
rect 29460 13515 29512 13524
rect 29460 13481 29469 13515
rect 29469 13481 29503 13515
rect 29503 13481 29512 13515
rect 29460 13472 29512 13481
rect 30840 13472 30892 13524
rect 31668 13472 31720 13524
rect 31944 13515 31996 13524
rect 31944 13481 31953 13515
rect 31953 13481 31987 13515
rect 31987 13481 31996 13515
rect 31944 13472 31996 13481
rect 32404 13515 32456 13524
rect 32404 13481 32413 13515
rect 32413 13481 32447 13515
rect 32447 13481 32456 13515
rect 32404 13472 32456 13481
rect 32864 13515 32916 13524
rect 32864 13481 32873 13515
rect 32873 13481 32907 13515
rect 32907 13481 32916 13515
rect 32864 13472 32916 13481
rect 33140 13472 33192 13524
rect 33416 13472 33468 13524
rect 36544 13515 36596 13524
rect 36544 13481 36553 13515
rect 36553 13481 36587 13515
rect 36587 13481 36596 13515
rect 36544 13472 36596 13481
rect 26700 13404 26752 13456
rect 34428 13404 34480 13456
rect 4988 13379 5040 13388
rect 4988 13345 4997 13379
rect 4997 13345 5031 13379
rect 5031 13345 5040 13379
rect 4988 13336 5040 13345
rect 8484 13379 8536 13388
rect 8484 13345 8493 13379
rect 8493 13345 8527 13379
rect 8527 13345 8536 13379
rect 8484 13336 8536 13345
rect 5356 13268 5408 13320
rect 9404 13268 9456 13320
rect 15200 13336 15252 13388
rect 16304 13336 16356 13388
rect 21088 13336 21140 13388
rect 22192 13379 22244 13388
rect 22192 13345 22226 13379
rect 22226 13345 22244 13379
rect 22192 13336 22244 13345
rect 26516 13379 26568 13388
rect 26516 13345 26525 13379
rect 26525 13345 26559 13379
rect 26559 13345 26568 13379
rect 26516 13336 26568 13345
rect 29368 13379 29420 13388
rect 29368 13345 29377 13379
rect 29377 13345 29411 13379
rect 29411 13345 29420 13379
rect 29368 13336 29420 13345
rect 11060 13268 11112 13320
rect 11244 13311 11296 13320
rect 11244 13277 11260 13311
rect 11260 13277 11294 13311
rect 11294 13277 11296 13311
rect 11244 13268 11296 13277
rect 15200 13200 15252 13252
rect 17960 13268 18012 13320
rect 19064 13311 19116 13320
rect 19064 13277 19073 13311
rect 19073 13277 19107 13311
rect 19107 13277 19116 13311
rect 19064 13268 19116 13277
rect 19156 13311 19208 13320
rect 19156 13277 19165 13311
rect 19165 13277 19199 13311
rect 19199 13277 19208 13311
rect 19156 13268 19208 13277
rect 5448 13132 5500 13184
rect 7380 13175 7432 13184
rect 7380 13141 7389 13175
rect 7389 13141 7423 13175
rect 7423 13141 7432 13175
rect 7380 13132 7432 13141
rect 12440 13132 12492 13184
rect 13268 13175 13320 13184
rect 13268 13141 13277 13175
rect 13277 13141 13311 13175
rect 13311 13141 13320 13175
rect 13268 13132 13320 13141
rect 14648 13175 14700 13184
rect 14648 13141 14657 13175
rect 14657 13141 14691 13175
rect 14691 13141 14700 13175
rect 14648 13132 14700 13141
rect 30380 13200 30432 13252
rect 32220 13379 32272 13388
rect 32220 13345 32229 13379
rect 32229 13345 32263 13379
rect 32263 13345 32272 13379
rect 32220 13336 32272 13345
rect 34336 13379 34388 13388
rect 34336 13345 34345 13379
rect 34345 13345 34379 13379
rect 34379 13345 34388 13379
rect 34336 13336 34388 13345
rect 35992 13336 36044 13388
rect 34428 13268 34480 13320
rect 35348 13311 35400 13320
rect 35348 13277 35357 13311
rect 35357 13277 35391 13311
rect 35391 13277 35400 13311
rect 35348 13268 35400 13277
rect 35440 13311 35492 13320
rect 35440 13277 35449 13311
rect 35449 13277 35483 13311
rect 35483 13277 35492 13311
rect 35440 13268 35492 13277
rect 33048 13200 33100 13252
rect 15476 13132 15528 13184
rect 19248 13132 19300 13184
rect 21916 13132 21968 13184
rect 23296 13175 23348 13184
rect 23296 13141 23305 13175
rect 23305 13141 23339 13175
rect 23339 13141 23348 13175
rect 23296 13132 23348 13141
rect 30472 13175 30524 13184
rect 30472 13141 30481 13175
rect 30481 13141 30515 13175
rect 30515 13141 30524 13175
rect 30472 13132 30524 13141
rect 35992 13175 36044 13184
rect 35992 13141 36001 13175
rect 36001 13141 36035 13175
rect 36035 13141 36044 13175
rect 35992 13132 36044 13141
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 3884 12928 3936 12980
rect 4988 12928 5040 12980
rect 6276 12928 6328 12980
rect 10048 12928 10100 12980
rect 11060 12928 11112 12980
rect 15292 12928 15344 12980
rect 19432 12971 19484 12980
rect 19432 12937 19441 12971
rect 19441 12937 19475 12971
rect 19475 12937 19484 12971
rect 19432 12928 19484 12937
rect 25688 12971 25740 12980
rect 25688 12937 25697 12971
rect 25697 12937 25731 12971
rect 25731 12937 25740 12971
rect 25688 12928 25740 12937
rect 26516 12971 26568 12980
rect 26516 12937 26525 12971
rect 26525 12937 26559 12971
rect 26559 12937 26568 12971
rect 26516 12928 26568 12937
rect 30472 12928 30524 12980
rect 32220 12971 32272 12980
rect 32220 12937 32229 12971
rect 32229 12937 32263 12971
rect 32263 12937 32272 12971
rect 32220 12928 32272 12937
rect 35900 12928 35952 12980
rect 9772 12903 9824 12912
rect 9772 12869 9781 12903
rect 9781 12869 9815 12903
rect 9815 12869 9824 12903
rect 9772 12860 9824 12869
rect 19064 12860 19116 12912
rect 3884 12767 3936 12776
rect 3884 12733 3893 12767
rect 3893 12733 3927 12767
rect 3927 12733 3936 12767
rect 3884 12724 3936 12733
rect 16304 12835 16356 12844
rect 5080 12724 5132 12776
rect 7380 12724 7432 12776
rect 7932 12724 7984 12776
rect 8484 12724 8536 12776
rect 9588 12724 9640 12776
rect 16304 12801 16313 12835
rect 16313 12801 16347 12835
rect 16347 12801 16356 12835
rect 16304 12792 16356 12801
rect 17776 12792 17828 12844
rect 29368 12860 29420 12912
rect 26608 12835 26660 12844
rect 26608 12801 26617 12835
rect 26617 12801 26651 12835
rect 26651 12801 26660 12835
rect 26608 12792 26660 12801
rect 29828 12835 29880 12844
rect 29828 12801 29837 12835
rect 29837 12801 29871 12835
rect 29871 12801 29880 12835
rect 29828 12792 29880 12801
rect 30380 12792 30432 12844
rect 31944 12792 31996 12844
rect 33324 12792 33376 12844
rect 34428 12792 34480 12844
rect 11244 12724 11296 12776
rect 15200 12724 15252 12776
rect 16120 12767 16172 12776
rect 16120 12733 16129 12767
rect 16129 12733 16163 12767
rect 16163 12733 16172 12767
rect 16120 12724 16172 12733
rect 21088 12724 21140 12776
rect 22468 12767 22520 12776
rect 22468 12733 22477 12767
rect 22477 12733 22511 12767
rect 22511 12733 22520 12767
rect 22468 12724 22520 12733
rect 6828 12656 6880 12708
rect 10416 12656 10468 12708
rect 13452 12656 13504 12708
rect 18236 12656 18288 12708
rect 19340 12656 19392 12708
rect 20628 12656 20680 12708
rect 21272 12656 21324 12708
rect 5356 12588 5408 12640
rect 6644 12588 6696 12640
rect 7104 12588 7156 12640
rect 7288 12631 7340 12640
rect 7288 12597 7297 12631
rect 7297 12597 7331 12631
rect 7331 12597 7340 12631
rect 7288 12588 7340 12597
rect 13820 12588 13872 12640
rect 16212 12631 16264 12640
rect 16212 12597 16221 12631
rect 16221 12597 16255 12631
rect 16255 12597 16264 12631
rect 16212 12588 16264 12597
rect 17776 12631 17828 12640
rect 17776 12597 17785 12631
rect 17785 12597 17819 12631
rect 17819 12597 17828 12631
rect 17776 12588 17828 12597
rect 22192 12656 22244 12708
rect 24400 12699 24452 12708
rect 24400 12665 24409 12699
rect 24409 12665 24443 12699
rect 24443 12665 24452 12699
rect 24400 12656 24452 12665
rect 26976 12656 27028 12708
rect 28724 12699 28776 12708
rect 28724 12665 28733 12699
rect 28733 12665 28767 12699
rect 28767 12665 28776 12699
rect 28724 12656 28776 12665
rect 30288 12656 30340 12708
rect 33600 12699 33652 12708
rect 33600 12665 33609 12699
rect 33609 12665 33643 12699
rect 33643 12665 33652 12699
rect 33600 12656 33652 12665
rect 35256 12724 35308 12776
rect 35992 12724 36044 12776
rect 35716 12656 35768 12708
rect 27620 12588 27672 12640
rect 31208 12631 31260 12640
rect 31208 12597 31217 12631
rect 31217 12597 31251 12631
rect 31251 12597 31260 12631
rect 31208 12588 31260 12597
rect 32312 12588 32364 12640
rect 34520 12588 34572 12640
rect 34888 12588 34940 12640
rect 35256 12588 35308 12640
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 5080 12384 5132 12436
rect 5448 12384 5500 12436
rect 9404 12427 9456 12436
rect 9404 12393 9413 12427
rect 9413 12393 9447 12427
rect 9447 12393 9456 12427
rect 9404 12384 9456 12393
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 12808 12384 12860 12436
rect 16212 12427 16264 12436
rect 16212 12393 16221 12427
rect 16221 12393 16255 12427
rect 16255 12393 16264 12427
rect 16212 12384 16264 12393
rect 17868 12384 17920 12436
rect 20628 12427 20680 12436
rect 20628 12393 20637 12427
rect 20637 12393 20671 12427
rect 20671 12393 20680 12427
rect 20628 12384 20680 12393
rect 26608 12384 26660 12436
rect 26976 12384 27028 12436
rect 29460 12384 29512 12436
rect 29828 12384 29880 12436
rect 4988 12359 5040 12368
rect 4988 12325 4997 12359
rect 4997 12325 5031 12359
rect 5031 12325 5040 12359
rect 4988 12316 5040 12325
rect 10416 12316 10468 12368
rect 16120 12316 16172 12368
rect 17132 12316 17184 12368
rect 18236 12316 18288 12368
rect 4712 12248 4764 12300
rect 6276 12180 6328 12232
rect 8300 12248 8352 12300
rect 8484 12223 8536 12232
rect 8484 12189 8493 12223
rect 8493 12189 8527 12223
rect 8527 12189 8536 12223
rect 8484 12180 8536 12189
rect 8668 12223 8720 12232
rect 8668 12189 8677 12223
rect 8677 12189 8711 12223
rect 8711 12189 8720 12223
rect 8668 12180 8720 12189
rect 6920 12087 6972 12096
rect 6920 12053 6929 12087
rect 6929 12053 6963 12087
rect 6963 12053 6972 12087
rect 6920 12044 6972 12053
rect 7104 12044 7156 12096
rect 7472 12044 7524 12096
rect 11060 12248 11112 12300
rect 11244 12291 11296 12300
rect 11244 12257 11253 12291
rect 11253 12257 11287 12291
rect 11287 12257 11296 12291
rect 11244 12248 11296 12257
rect 12716 12248 12768 12300
rect 18696 12316 18748 12368
rect 22652 12316 22704 12368
rect 23296 12316 23348 12368
rect 26700 12316 26752 12368
rect 28080 12316 28132 12368
rect 28724 12316 28776 12368
rect 30288 12384 30340 12436
rect 31944 12384 31996 12436
rect 32864 12384 32916 12436
rect 33048 12427 33100 12436
rect 33048 12393 33057 12427
rect 33057 12393 33091 12427
rect 33091 12393 33100 12427
rect 33048 12384 33100 12393
rect 33416 12427 33468 12436
rect 33416 12393 33425 12427
rect 33425 12393 33459 12427
rect 33459 12393 33468 12427
rect 33416 12384 33468 12393
rect 33600 12384 33652 12436
rect 34060 12384 34112 12436
rect 34336 12384 34388 12436
rect 35348 12384 35400 12436
rect 9496 12180 9548 12232
rect 13728 12223 13780 12232
rect 13728 12189 13737 12223
rect 13737 12189 13771 12223
rect 13771 12189 13780 12223
rect 13728 12180 13780 12189
rect 16764 12180 16816 12232
rect 22468 12248 22520 12300
rect 30472 12291 30524 12300
rect 17500 12180 17552 12232
rect 17776 12180 17828 12232
rect 21272 12180 21324 12232
rect 30472 12257 30481 12291
rect 30481 12257 30515 12291
rect 30515 12257 30524 12291
rect 30472 12248 30524 12257
rect 26608 12180 26660 12232
rect 27620 12223 27672 12232
rect 27620 12189 27629 12223
rect 27629 12189 27663 12223
rect 27663 12189 27672 12223
rect 27620 12180 27672 12189
rect 30196 12180 30248 12232
rect 34520 12316 34572 12368
rect 35992 12384 36044 12436
rect 33876 12291 33928 12300
rect 33876 12257 33885 12291
rect 33885 12257 33919 12291
rect 33919 12257 33928 12291
rect 33876 12248 33928 12257
rect 36268 12248 36320 12300
rect 30840 12180 30892 12232
rect 33968 12223 34020 12232
rect 33968 12189 33977 12223
rect 33977 12189 34011 12223
rect 34011 12189 34020 12223
rect 33968 12180 34020 12189
rect 34336 12180 34388 12232
rect 34612 12180 34664 12232
rect 34888 12180 34940 12232
rect 10968 12044 11020 12096
rect 11060 12044 11112 12096
rect 13176 12087 13228 12096
rect 13176 12053 13185 12087
rect 13185 12053 13219 12087
rect 13219 12053 13228 12087
rect 13176 12044 13228 12053
rect 15016 12087 15068 12096
rect 15016 12053 15025 12087
rect 15025 12053 15059 12087
rect 15059 12053 15068 12087
rect 15016 12044 15068 12053
rect 18236 12044 18288 12096
rect 21088 12087 21140 12096
rect 21088 12053 21097 12087
rect 21097 12053 21131 12087
rect 21131 12053 21140 12087
rect 21088 12044 21140 12053
rect 22192 12087 22244 12096
rect 22192 12053 22201 12087
rect 22201 12053 22235 12087
rect 22235 12053 22244 12087
rect 22192 12044 22244 12053
rect 22560 12087 22612 12096
rect 22560 12053 22569 12087
rect 22569 12053 22603 12087
rect 22603 12053 22612 12087
rect 22560 12044 22612 12053
rect 23940 12044 23992 12096
rect 30380 12044 30432 12096
rect 31208 12044 31260 12096
rect 34428 12044 34480 12096
rect 34612 12044 34664 12096
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 3884 11883 3936 11892
rect 3884 11849 3893 11883
rect 3893 11849 3927 11883
rect 3927 11849 3936 11883
rect 3884 11840 3936 11849
rect 6828 11883 6880 11892
rect 6828 11849 6837 11883
rect 6837 11849 6871 11883
rect 6871 11849 6880 11883
rect 6828 11840 6880 11849
rect 6920 11840 6972 11892
rect 8484 11840 8536 11892
rect 9036 11840 9088 11892
rect 9772 11840 9824 11892
rect 10416 11883 10468 11892
rect 10416 11849 10425 11883
rect 10425 11849 10459 11883
rect 10459 11849 10468 11883
rect 10416 11840 10468 11849
rect 12716 11883 12768 11892
rect 12716 11849 12725 11883
rect 12725 11849 12759 11883
rect 12759 11849 12768 11883
rect 12716 11840 12768 11849
rect 16764 11883 16816 11892
rect 16764 11849 16773 11883
rect 16773 11849 16807 11883
rect 16807 11849 16816 11883
rect 16764 11840 16816 11849
rect 17132 11883 17184 11892
rect 17132 11849 17141 11883
rect 17141 11849 17175 11883
rect 17175 11849 17184 11883
rect 17132 11840 17184 11849
rect 20628 11883 20680 11892
rect 20628 11849 20637 11883
rect 20637 11849 20671 11883
rect 20671 11849 20680 11883
rect 20628 11840 20680 11849
rect 21272 11883 21324 11892
rect 21272 11849 21281 11883
rect 21281 11849 21315 11883
rect 21315 11849 21324 11883
rect 21272 11840 21324 11849
rect 21732 11883 21784 11892
rect 21732 11849 21741 11883
rect 21741 11849 21775 11883
rect 21775 11849 21784 11883
rect 21732 11840 21784 11849
rect 22468 11840 22520 11892
rect 26608 11883 26660 11892
rect 7472 11747 7524 11756
rect 3884 11636 3936 11688
rect 7472 11713 7481 11747
rect 7481 11713 7515 11747
rect 7515 11713 7524 11747
rect 7472 11704 7524 11713
rect 22560 11747 22612 11756
rect 4988 11636 5040 11688
rect 8116 11636 8168 11688
rect 9036 11679 9088 11688
rect 9036 11645 9045 11679
rect 9045 11645 9079 11679
rect 9079 11645 9088 11679
rect 9036 11636 9088 11645
rect 22560 11713 22569 11747
rect 22569 11713 22603 11747
rect 22603 11713 22612 11747
rect 22560 11704 22612 11713
rect 26608 11849 26617 11883
rect 26617 11849 26651 11883
rect 26651 11849 26660 11883
rect 26608 11840 26660 11849
rect 28080 11883 28132 11892
rect 28080 11849 28089 11883
rect 28089 11849 28123 11883
rect 28123 11849 28132 11883
rect 28080 11840 28132 11849
rect 30840 11840 30892 11892
rect 32312 11883 32364 11892
rect 32312 11849 32321 11883
rect 32321 11849 32355 11883
rect 32355 11849 32364 11883
rect 32312 11840 32364 11849
rect 33968 11840 34020 11892
rect 34336 11840 34388 11892
rect 36268 11883 36320 11892
rect 36268 11849 36277 11883
rect 36277 11849 36311 11883
rect 36311 11849 36320 11883
rect 36268 11840 36320 11849
rect 33876 11704 33928 11756
rect 6644 11611 6696 11620
rect 6644 11577 6653 11611
rect 6653 11577 6687 11611
rect 6687 11577 6696 11611
rect 6644 11568 6696 11577
rect 9312 11611 9364 11620
rect 9312 11577 9346 11611
rect 9346 11577 9364 11611
rect 9312 11568 9364 11577
rect 12716 11568 12768 11620
rect 13728 11636 13780 11688
rect 21916 11679 21968 11688
rect 5172 11500 5224 11552
rect 7656 11500 7708 11552
rect 8300 11500 8352 11552
rect 11244 11500 11296 11552
rect 12900 11500 12952 11552
rect 13820 11500 13872 11552
rect 17500 11543 17552 11552
rect 17500 11509 17509 11543
rect 17509 11509 17543 11543
rect 17543 11509 17552 11543
rect 17500 11500 17552 11509
rect 17776 11500 17828 11552
rect 21916 11645 21925 11679
rect 21925 11645 21959 11679
rect 21959 11645 21968 11679
rect 21916 11636 21968 11645
rect 23940 11679 23992 11688
rect 19432 11568 19484 11620
rect 23940 11645 23974 11679
rect 23974 11645 23992 11679
rect 23940 11636 23992 11645
rect 26792 11568 26844 11620
rect 27528 11568 27580 11620
rect 29552 11611 29604 11620
rect 29552 11577 29586 11611
rect 29586 11577 29604 11611
rect 29552 11568 29604 11577
rect 32404 11568 32456 11620
rect 35992 11568 36044 11620
rect 18696 11543 18748 11552
rect 18696 11509 18705 11543
rect 18705 11509 18739 11543
rect 18739 11509 18748 11543
rect 18696 11500 18748 11509
rect 22008 11543 22060 11552
rect 22008 11509 22017 11543
rect 22017 11509 22051 11543
rect 22051 11509 22060 11543
rect 22008 11500 22060 11509
rect 22192 11500 22244 11552
rect 22744 11500 22796 11552
rect 25044 11543 25096 11552
rect 25044 11509 25053 11543
rect 25053 11509 25087 11543
rect 25087 11509 25096 11543
rect 25044 11500 25096 11509
rect 28172 11500 28224 11552
rect 30380 11500 30432 11552
rect 33508 11500 33560 11552
rect 34612 11543 34664 11552
rect 34612 11509 34621 11543
rect 34621 11509 34655 11543
rect 34655 11509 34664 11543
rect 34612 11500 34664 11509
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 4712 11339 4764 11348
rect 4712 11305 4721 11339
rect 4721 11305 4755 11339
rect 4755 11305 4764 11339
rect 4712 11296 4764 11305
rect 5172 11339 5224 11348
rect 5172 11305 5181 11339
rect 5181 11305 5215 11339
rect 5215 11305 5224 11339
rect 5172 11296 5224 11305
rect 5448 11296 5500 11348
rect 6276 11296 6328 11348
rect 8392 11296 8444 11348
rect 9496 11339 9548 11348
rect 9496 11305 9505 11339
rect 9505 11305 9539 11339
rect 9539 11305 9548 11339
rect 9496 11296 9548 11305
rect 6644 11228 6696 11280
rect 8484 11228 8536 11280
rect 15016 11296 15068 11348
rect 18696 11296 18748 11348
rect 19432 11296 19484 11348
rect 21088 11296 21140 11348
rect 22652 11339 22704 11348
rect 22652 11305 22661 11339
rect 22661 11305 22695 11339
rect 22695 11305 22704 11339
rect 22652 11296 22704 11305
rect 23940 11296 23992 11348
rect 26792 11339 26844 11348
rect 26792 11305 26801 11339
rect 26801 11305 26835 11339
rect 26835 11305 26844 11339
rect 26792 11296 26844 11305
rect 27620 11339 27672 11348
rect 27620 11305 27629 11339
rect 27629 11305 27663 11339
rect 27663 11305 27672 11339
rect 27620 11296 27672 11305
rect 28080 11339 28132 11348
rect 28080 11305 28089 11339
rect 28089 11305 28123 11339
rect 28123 11305 28132 11339
rect 28080 11296 28132 11305
rect 29552 11339 29604 11348
rect 29552 11305 29561 11339
rect 29561 11305 29595 11339
rect 29595 11305 29604 11339
rect 30472 11339 30524 11348
rect 29552 11296 29604 11305
rect 30472 11305 30481 11339
rect 30481 11305 30515 11339
rect 30515 11305 30524 11339
rect 30472 11296 30524 11305
rect 30840 11339 30892 11348
rect 30840 11305 30849 11339
rect 30849 11305 30883 11339
rect 30883 11305 30892 11339
rect 30840 11296 30892 11305
rect 33508 11339 33560 11348
rect 33508 11305 33517 11339
rect 33517 11305 33551 11339
rect 33551 11305 33560 11339
rect 33508 11296 33560 11305
rect 35992 11339 36044 11348
rect 35992 11305 36001 11339
rect 36001 11305 36035 11339
rect 36035 11305 36044 11339
rect 35992 11296 36044 11305
rect 20996 11228 21048 11280
rect 22008 11228 22060 11280
rect 5448 11160 5500 11212
rect 5356 11092 5408 11144
rect 6276 11135 6328 11144
rect 6276 11101 6285 11135
rect 6285 11101 6319 11135
rect 6319 11101 6328 11135
rect 6276 11092 6328 11101
rect 7656 11067 7708 11076
rect 3792 10956 3844 11008
rect 7656 11033 7665 11067
rect 7665 11033 7699 11067
rect 7699 11033 7708 11067
rect 10508 11160 10560 11212
rect 12440 11160 12492 11212
rect 17776 11160 17828 11212
rect 17960 11160 18012 11212
rect 19156 11160 19208 11212
rect 22744 11228 22796 11280
rect 23204 11228 23256 11280
rect 25044 11228 25096 11280
rect 28632 11228 28684 11280
rect 30196 11271 30248 11280
rect 30196 11237 30205 11271
rect 30205 11237 30239 11271
rect 30239 11237 30248 11271
rect 30196 11228 30248 11237
rect 32404 11271 32456 11280
rect 32404 11237 32438 11271
rect 32438 11237 32456 11271
rect 32404 11228 32456 11237
rect 33968 11228 34020 11280
rect 34796 11228 34848 11280
rect 28172 11203 28224 11212
rect 28172 11169 28181 11203
rect 28181 11169 28215 11203
rect 28215 11169 28224 11203
rect 28172 11160 28224 11169
rect 9036 11092 9088 11144
rect 12716 11135 12768 11144
rect 12716 11101 12725 11135
rect 12725 11101 12759 11135
rect 12759 11101 12768 11135
rect 12716 11092 12768 11101
rect 20720 11092 20772 11144
rect 23480 11135 23532 11144
rect 23480 11101 23489 11135
rect 23489 11101 23523 11135
rect 23523 11101 23532 11135
rect 23480 11092 23532 11101
rect 32128 11135 32180 11144
rect 32128 11101 32137 11135
rect 32137 11101 32171 11135
rect 32171 11101 32180 11135
rect 32128 11092 32180 11101
rect 34612 11135 34664 11144
rect 34612 11101 34621 11135
rect 34621 11101 34655 11135
rect 34655 11101 34664 11135
rect 34612 11092 34664 11101
rect 8668 11067 8720 11076
rect 7656 11024 7708 11033
rect 8668 11033 8677 11067
rect 8677 11033 8711 11067
rect 8711 11033 8720 11067
rect 8668 11024 8720 11033
rect 9588 11024 9640 11076
rect 20812 11024 20864 11076
rect 22560 11024 22612 11076
rect 24860 11067 24912 11076
rect 24860 11033 24869 11067
rect 24869 11033 24903 11067
rect 24903 11033 24912 11067
rect 24860 11024 24912 11033
rect 34336 11024 34388 11076
rect 8300 10956 8352 11008
rect 9312 10956 9364 11008
rect 9496 10956 9548 11008
rect 21272 10999 21324 11008
rect 21272 10965 21281 10999
rect 21281 10965 21315 10999
rect 21315 10965 21324 10999
rect 21272 10956 21324 10965
rect 23020 10999 23072 11008
rect 23020 10965 23029 10999
rect 23029 10965 23063 10999
rect 23063 10965 23072 10999
rect 23020 10956 23072 10965
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 3792 10795 3844 10804
rect 3792 10761 3801 10795
rect 3801 10761 3835 10795
rect 3835 10761 3844 10795
rect 3792 10752 3844 10761
rect 3884 10752 3936 10804
rect 5448 10752 5500 10804
rect 8208 10752 8260 10804
rect 9496 10752 9548 10804
rect 9772 10752 9824 10804
rect 10508 10795 10560 10804
rect 6276 10684 6328 10736
rect 7012 10684 7064 10736
rect 8116 10727 8168 10736
rect 8116 10693 8125 10727
rect 8125 10693 8159 10727
rect 8159 10693 8168 10727
rect 8116 10684 8168 10693
rect 4252 10659 4304 10668
rect 4252 10625 4261 10659
rect 4261 10625 4295 10659
rect 4295 10625 4304 10659
rect 4252 10616 4304 10625
rect 10508 10761 10517 10795
rect 10517 10761 10551 10795
rect 10551 10761 10560 10795
rect 10508 10752 10560 10761
rect 17868 10752 17920 10804
rect 19156 10752 19208 10804
rect 20996 10795 21048 10804
rect 20996 10761 21005 10795
rect 21005 10761 21039 10795
rect 21039 10761 21048 10795
rect 20996 10752 21048 10761
rect 21088 10752 21140 10804
rect 22468 10752 22520 10804
rect 23480 10752 23532 10804
rect 28172 10795 28224 10804
rect 28172 10761 28181 10795
rect 28181 10761 28215 10795
rect 28215 10761 28224 10795
rect 28172 10752 28224 10761
rect 28632 10795 28684 10804
rect 28632 10761 28641 10795
rect 28641 10761 28675 10795
rect 28675 10761 28684 10795
rect 28632 10752 28684 10761
rect 32128 10752 32180 10804
rect 32404 10752 32456 10804
rect 34612 10795 34664 10804
rect 34612 10761 34621 10795
rect 34621 10761 34655 10795
rect 34655 10761 34664 10795
rect 34612 10752 34664 10761
rect 34796 10752 34848 10804
rect 10600 10616 10652 10668
rect 12716 10659 12768 10668
rect 12716 10625 12725 10659
rect 12725 10625 12759 10659
rect 12759 10625 12768 10659
rect 12716 10616 12768 10625
rect 13452 10616 13504 10668
rect 7288 10548 7340 10600
rect 8484 10591 8536 10600
rect 8484 10557 8518 10591
rect 8518 10557 8536 10591
rect 8484 10548 8536 10557
rect 11152 10591 11204 10600
rect 11152 10557 11161 10591
rect 11161 10557 11195 10591
rect 11195 10557 11204 10591
rect 11152 10548 11204 10557
rect 14648 10616 14700 10668
rect 22560 10659 22612 10668
rect 22560 10625 22569 10659
rect 22569 10625 22603 10659
rect 22603 10625 22612 10659
rect 22560 10616 22612 10625
rect 23020 10616 23072 10668
rect 14464 10591 14516 10600
rect 14464 10557 14473 10591
rect 14473 10557 14507 10591
rect 14507 10557 14516 10591
rect 17776 10591 17828 10600
rect 14464 10548 14516 10557
rect 4804 10480 4856 10532
rect 5172 10480 5224 10532
rect 16856 10480 16908 10532
rect 17776 10557 17785 10591
rect 17785 10557 17819 10591
rect 17819 10557 17828 10591
rect 17776 10548 17828 10557
rect 23480 10548 23532 10600
rect 24768 10548 24820 10600
rect 18236 10480 18288 10532
rect 30288 10548 30340 10600
rect 34520 10684 34572 10736
rect 12256 10455 12308 10464
rect 12256 10421 12265 10455
rect 12265 10421 12299 10455
rect 12299 10421 12308 10455
rect 12256 10412 12308 10421
rect 13820 10412 13872 10464
rect 15568 10455 15620 10464
rect 15568 10421 15577 10455
rect 15577 10421 15611 10455
rect 15611 10421 15620 10455
rect 15568 10412 15620 10421
rect 20628 10455 20680 10464
rect 20628 10421 20637 10455
rect 20637 10421 20671 10455
rect 20671 10421 20680 10455
rect 20628 10412 20680 10421
rect 21916 10412 21968 10464
rect 22376 10455 22428 10464
rect 22376 10421 22385 10455
rect 22385 10421 22419 10455
rect 22419 10421 22428 10455
rect 22376 10412 22428 10421
rect 25044 10455 25096 10464
rect 25044 10421 25053 10455
rect 25053 10421 25087 10455
rect 25087 10421 25096 10455
rect 25044 10412 25096 10421
rect 30012 10412 30064 10464
rect 31024 10455 31076 10464
rect 31024 10421 31033 10455
rect 31033 10421 31067 10455
rect 31067 10421 31076 10455
rect 31024 10412 31076 10421
rect 35624 10548 35676 10600
rect 32404 10523 32456 10532
rect 32404 10489 32438 10523
rect 32438 10489 32456 10523
rect 32404 10480 32456 10489
rect 32956 10412 33008 10464
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 4804 10251 4856 10260
rect 4804 10217 4813 10251
rect 4813 10217 4847 10251
rect 4847 10217 4856 10251
rect 4804 10208 4856 10217
rect 6644 10208 6696 10260
rect 7932 10251 7984 10260
rect 7932 10217 7941 10251
rect 7941 10217 7975 10251
rect 7975 10217 7984 10251
rect 7932 10208 7984 10217
rect 8484 10208 8536 10260
rect 9588 10208 9640 10260
rect 10968 10251 11020 10260
rect 10968 10217 10977 10251
rect 10977 10217 11011 10251
rect 11011 10217 11020 10251
rect 10968 10208 11020 10217
rect 23204 10251 23256 10260
rect 23204 10217 23213 10251
rect 23213 10217 23247 10251
rect 23247 10217 23256 10251
rect 23204 10208 23256 10217
rect 5448 10140 5500 10192
rect 13728 10140 13780 10192
rect 22376 10140 22428 10192
rect 23020 10140 23072 10192
rect 25044 10140 25096 10192
rect 30288 10208 30340 10260
rect 31024 10208 31076 10260
rect 32404 10251 32456 10260
rect 32404 10217 32413 10251
rect 32413 10217 32447 10251
rect 32447 10217 32456 10251
rect 32404 10208 32456 10217
rect 32496 10208 32548 10260
rect 34796 10208 34848 10260
rect 30196 10140 30248 10192
rect 33508 10140 33560 10192
rect 4252 10072 4304 10124
rect 5080 10115 5132 10124
rect 5080 10081 5089 10115
rect 5089 10081 5123 10115
rect 5123 10081 5132 10115
rect 5080 10072 5132 10081
rect 8300 10115 8352 10124
rect 8300 10081 8309 10115
rect 8309 10081 8343 10115
rect 8343 10081 8352 10115
rect 8300 10072 8352 10081
rect 9680 10115 9732 10124
rect 9680 10081 9689 10115
rect 9689 10081 9723 10115
rect 9723 10081 9732 10115
rect 9680 10072 9732 10081
rect 10968 10072 11020 10124
rect 12716 10115 12768 10124
rect 12716 10081 12725 10115
rect 12725 10081 12759 10115
rect 12759 10081 12768 10115
rect 12716 10072 12768 10081
rect 16672 10072 16724 10124
rect 19340 10115 19392 10124
rect 19340 10081 19349 10115
rect 19349 10081 19383 10115
rect 19383 10081 19392 10115
rect 19340 10072 19392 10081
rect 21272 10072 21324 10124
rect 22008 10072 22060 10124
rect 27988 10072 28040 10124
rect 30012 10115 30064 10124
rect 30012 10081 30021 10115
rect 30021 10081 30055 10115
rect 30055 10081 30064 10115
rect 30012 10072 30064 10081
rect 35440 10115 35492 10124
rect 35440 10081 35449 10115
rect 35449 10081 35483 10115
rect 35483 10081 35492 10115
rect 35440 10072 35492 10081
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 16304 10004 16356 10056
rect 16856 10047 16908 10056
rect 16856 10013 16865 10047
rect 16865 10013 16899 10047
rect 16899 10013 16908 10047
rect 16856 10004 16908 10013
rect 23296 10047 23348 10056
rect 23296 10013 23305 10047
rect 23305 10013 23339 10047
rect 23339 10013 23348 10047
rect 23296 10004 23348 10013
rect 30196 10047 30248 10056
rect 30196 10013 30205 10047
rect 30205 10013 30239 10047
rect 30239 10013 30248 10047
rect 30196 10004 30248 10013
rect 32956 10047 33008 10056
rect 32956 10013 32965 10047
rect 32965 10013 32999 10047
rect 32999 10013 33008 10047
rect 32956 10004 33008 10013
rect 34520 9936 34572 9988
rect 13820 9868 13872 9920
rect 14648 9911 14700 9920
rect 14648 9877 14657 9911
rect 14657 9877 14691 9911
rect 14691 9877 14700 9911
rect 14648 9868 14700 9877
rect 16488 9911 16540 9920
rect 16488 9877 16497 9911
rect 16497 9877 16531 9911
rect 16531 9877 16540 9911
rect 16488 9868 16540 9877
rect 18236 9911 18288 9920
rect 18236 9877 18245 9911
rect 18245 9877 18279 9911
rect 18279 9877 18288 9911
rect 18236 9868 18288 9877
rect 19340 9868 19392 9920
rect 21088 9911 21140 9920
rect 21088 9877 21097 9911
rect 21097 9877 21131 9911
rect 21131 9877 21140 9911
rect 21088 9868 21140 9877
rect 21548 9911 21600 9920
rect 21548 9877 21557 9911
rect 21557 9877 21591 9911
rect 21591 9877 21600 9911
rect 21548 9868 21600 9877
rect 22560 9868 22612 9920
rect 23204 9868 23256 9920
rect 24676 9911 24728 9920
rect 24676 9877 24685 9911
rect 24685 9877 24719 9911
rect 24719 9877 24728 9911
rect 24676 9868 24728 9877
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 5080 9707 5132 9716
rect 5080 9673 5089 9707
rect 5089 9673 5123 9707
rect 5123 9673 5132 9707
rect 5080 9664 5132 9673
rect 5448 9707 5500 9716
rect 5448 9673 5457 9707
rect 5457 9673 5491 9707
rect 5491 9673 5500 9707
rect 5448 9664 5500 9673
rect 8116 9596 8168 9648
rect 8484 9664 8536 9716
rect 8576 9664 8628 9716
rect 10968 9664 11020 9716
rect 12716 9707 12768 9716
rect 12716 9673 12725 9707
rect 12725 9673 12759 9707
rect 12759 9673 12768 9707
rect 12716 9664 12768 9673
rect 14464 9664 14516 9716
rect 16856 9664 16908 9716
rect 19432 9707 19484 9716
rect 19432 9673 19441 9707
rect 19441 9673 19475 9707
rect 19475 9673 19484 9707
rect 19432 9664 19484 9673
rect 21272 9664 21324 9716
rect 23020 9707 23072 9716
rect 23020 9673 23029 9707
rect 23029 9673 23063 9707
rect 23063 9673 23072 9707
rect 23020 9664 23072 9673
rect 24676 9707 24728 9716
rect 12256 9596 12308 9648
rect 16672 9596 16724 9648
rect 23664 9639 23716 9648
rect 7840 9460 7892 9512
rect 13728 9528 13780 9580
rect 17040 9571 17092 9580
rect 17040 9537 17049 9571
rect 17049 9537 17083 9571
rect 17083 9537 17092 9571
rect 17040 9528 17092 9537
rect 18236 9528 18288 9580
rect 18696 9571 18748 9580
rect 18696 9537 18705 9571
rect 18705 9537 18739 9571
rect 18739 9537 18748 9571
rect 18696 9528 18748 9537
rect 21916 9571 21968 9580
rect 21916 9537 21925 9571
rect 21925 9537 21959 9571
rect 21959 9537 21968 9571
rect 21916 9528 21968 9537
rect 23664 9605 23673 9639
rect 23673 9605 23707 9639
rect 23707 9605 23716 9639
rect 23664 9596 23716 9605
rect 24676 9673 24685 9707
rect 24685 9673 24719 9707
rect 24719 9673 24728 9707
rect 24676 9664 24728 9673
rect 30012 9707 30064 9716
rect 30012 9673 30021 9707
rect 30021 9673 30055 9707
rect 30055 9673 30064 9707
rect 30012 9664 30064 9673
rect 30196 9664 30248 9716
rect 32956 9707 33008 9716
rect 30288 9596 30340 9648
rect 32956 9673 32965 9707
rect 32965 9673 32999 9707
rect 32999 9673 33008 9707
rect 32956 9664 33008 9673
rect 33508 9664 33560 9716
rect 35440 9707 35492 9716
rect 35440 9673 35449 9707
rect 35449 9673 35483 9707
rect 35483 9673 35492 9707
rect 35440 9664 35492 9673
rect 30840 9596 30892 9648
rect 24124 9571 24176 9580
rect 24124 9537 24133 9571
rect 24133 9537 24167 9571
rect 24167 9537 24176 9571
rect 24124 9528 24176 9537
rect 7472 9392 7524 9444
rect 8576 9392 8628 9444
rect 12992 9460 13044 9512
rect 7840 9367 7892 9376
rect 7840 9333 7849 9367
rect 7849 9333 7883 9367
rect 7883 9333 7892 9367
rect 7840 9324 7892 9333
rect 8392 9324 8444 9376
rect 8944 9367 8996 9376
rect 8944 9333 8953 9367
rect 8953 9333 8987 9367
rect 8987 9333 8996 9367
rect 8944 9324 8996 9333
rect 9680 9324 9732 9376
rect 11612 9324 11664 9376
rect 12808 9324 12860 9376
rect 13084 9392 13136 9444
rect 16764 9460 16816 9512
rect 18420 9503 18472 9512
rect 18420 9469 18429 9503
rect 18429 9469 18463 9503
rect 18463 9469 18472 9503
rect 18420 9460 18472 9469
rect 19156 9460 19208 9512
rect 20628 9503 20680 9512
rect 20628 9469 20637 9503
rect 20637 9469 20671 9503
rect 20671 9469 20680 9503
rect 20628 9460 20680 9469
rect 20812 9460 20864 9512
rect 21548 9460 21600 9512
rect 23204 9460 23256 9512
rect 13636 9324 13688 9376
rect 16396 9367 16448 9376
rect 16396 9333 16405 9367
rect 16405 9333 16439 9367
rect 16439 9333 16448 9367
rect 16396 9324 16448 9333
rect 16488 9324 16540 9376
rect 16580 9324 16632 9376
rect 16764 9367 16816 9376
rect 16764 9333 16773 9367
rect 16773 9333 16807 9367
rect 16807 9333 16816 9367
rect 16764 9324 16816 9333
rect 20628 9324 20680 9376
rect 22652 9324 22704 9376
rect 23296 9367 23348 9376
rect 23296 9333 23305 9367
rect 23305 9333 23339 9367
rect 23339 9333 23348 9367
rect 23296 9324 23348 9333
rect 24032 9367 24084 9376
rect 24032 9333 24041 9367
rect 24041 9333 24075 9367
rect 24075 9333 24084 9367
rect 24032 9324 24084 9333
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 13084 9163 13136 9172
rect 13084 9129 13093 9163
rect 13093 9129 13127 9163
rect 13127 9129 13136 9163
rect 13084 9120 13136 9129
rect 13452 9163 13504 9172
rect 13452 9129 13461 9163
rect 13461 9129 13495 9163
rect 13495 9129 13504 9163
rect 13452 9120 13504 9129
rect 13544 9163 13596 9172
rect 13544 9129 13553 9163
rect 13553 9129 13587 9163
rect 13587 9129 13596 9163
rect 13544 9120 13596 9129
rect 16764 9120 16816 9172
rect 17408 9120 17460 9172
rect 18420 9120 18472 9172
rect 18696 9120 18748 9172
rect 19340 9120 19392 9172
rect 21088 9120 21140 9172
rect 24032 9163 24084 9172
rect 24032 9129 24041 9163
rect 24041 9129 24075 9163
rect 24075 9129 24084 9163
rect 24032 9120 24084 9129
rect 12992 9095 13044 9104
rect 12992 9061 13001 9095
rect 13001 9061 13035 9095
rect 13035 9061 13044 9095
rect 12992 9052 13044 9061
rect 16672 9052 16724 9104
rect 23112 9052 23164 9104
rect 24124 9052 24176 9104
rect 7288 9027 7340 9036
rect 7288 8993 7322 9027
rect 7322 8993 7340 9027
rect 7288 8984 7340 8993
rect 10876 9027 10928 9036
rect 10876 8993 10910 9027
rect 10910 8993 10928 9027
rect 10876 8984 10928 8993
rect 12716 8984 12768 9036
rect 16304 8984 16356 9036
rect 21364 8984 21416 9036
rect 26608 8984 26660 9036
rect 28172 9120 28224 9172
rect 28080 8984 28132 9036
rect 6828 8916 6880 8968
rect 7012 8959 7064 8968
rect 7012 8925 7021 8959
rect 7021 8925 7055 8959
rect 7055 8925 7064 8959
rect 7012 8916 7064 8925
rect 10600 8959 10652 8968
rect 10600 8925 10609 8959
rect 10609 8925 10643 8959
rect 10643 8925 10652 8959
rect 10600 8916 10652 8925
rect 13636 8959 13688 8968
rect 13636 8925 13645 8959
rect 13645 8925 13679 8959
rect 13679 8925 13688 8959
rect 13636 8916 13688 8925
rect 18972 8916 19024 8968
rect 19524 8959 19576 8968
rect 19524 8925 19533 8959
rect 19533 8925 19567 8959
rect 19567 8925 19576 8959
rect 19524 8916 19576 8925
rect 21456 8959 21508 8968
rect 21456 8925 21465 8959
rect 21465 8925 21499 8959
rect 21499 8925 21508 8959
rect 21456 8916 21508 8925
rect 22652 8959 22704 8968
rect 22652 8925 22661 8959
rect 22661 8925 22695 8959
rect 22695 8925 22704 8959
rect 22652 8916 22704 8925
rect 6920 8823 6972 8832
rect 6920 8789 6929 8823
rect 6929 8789 6963 8823
rect 6963 8789 6972 8823
rect 6920 8780 6972 8789
rect 8392 8823 8444 8832
rect 8392 8789 8401 8823
rect 8401 8789 8435 8823
rect 8435 8789 8444 8823
rect 8392 8780 8444 8789
rect 10784 8780 10836 8832
rect 18880 8823 18932 8832
rect 18880 8789 18889 8823
rect 18889 8789 18923 8823
rect 18923 8789 18932 8823
rect 18880 8780 18932 8789
rect 20536 8780 20588 8832
rect 20720 8780 20772 8832
rect 25504 8780 25556 8832
rect 29368 8823 29420 8832
rect 29368 8789 29377 8823
rect 29377 8789 29411 8823
rect 29411 8789 29420 8823
rect 29368 8780 29420 8789
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 10600 8576 10652 8628
rect 7840 8508 7892 8560
rect 10324 8508 10376 8560
rect 10876 8483 10928 8492
rect 10876 8449 10885 8483
rect 10885 8449 10919 8483
rect 10919 8449 10928 8483
rect 10876 8440 10928 8449
rect 13636 8576 13688 8628
rect 16580 8576 16632 8628
rect 17408 8619 17460 8628
rect 17408 8585 17417 8619
rect 17417 8585 17451 8619
rect 17451 8585 17460 8619
rect 17408 8576 17460 8585
rect 18972 8619 19024 8628
rect 18972 8585 18981 8619
rect 18981 8585 19015 8619
rect 19015 8585 19024 8619
rect 18972 8576 19024 8585
rect 19340 8619 19392 8628
rect 19340 8585 19349 8619
rect 19349 8585 19383 8619
rect 19383 8585 19392 8619
rect 19340 8576 19392 8585
rect 20628 8619 20680 8628
rect 20628 8585 20637 8619
rect 20637 8585 20671 8619
rect 20671 8585 20680 8619
rect 20628 8576 20680 8585
rect 21088 8576 21140 8628
rect 23112 8619 23164 8628
rect 23112 8585 23121 8619
rect 23121 8585 23155 8619
rect 23155 8585 23164 8619
rect 23112 8576 23164 8585
rect 26608 8619 26660 8628
rect 26608 8585 26617 8619
rect 26617 8585 26651 8619
rect 26651 8585 26660 8619
rect 26608 8576 26660 8585
rect 28080 8619 28132 8628
rect 28080 8585 28089 8619
rect 28089 8585 28123 8619
rect 28123 8585 28132 8619
rect 28080 8576 28132 8585
rect 28172 8576 28224 8628
rect 28724 8576 28776 8628
rect 13820 8551 13872 8560
rect 13820 8517 13829 8551
rect 13829 8517 13863 8551
rect 13863 8517 13872 8551
rect 13820 8508 13872 8517
rect 19892 8508 19944 8560
rect 21364 8508 21416 8560
rect 6828 8415 6880 8424
rect 6184 8279 6236 8288
rect 6184 8245 6193 8279
rect 6193 8245 6227 8279
rect 6227 8245 6236 8279
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 10600 8372 10652 8424
rect 10784 8415 10836 8424
rect 10784 8381 10793 8415
rect 10793 8381 10827 8415
rect 10827 8381 10836 8415
rect 10784 8372 10836 8381
rect 6920 8304 6972 8356
rect 8208 8304 8260 8356
rect 17316 8440 17368 8492
rect 18696 8440 18748 8492
rect 25596 8440 25648 8492
rect 6184 8236 6236 8245
rect 8760 8236 8812 8288
rect 12532 8304 12584 8356
rect 14004 8372 14056 8424
rect 16396 8372 16448 8424
rect 20536 8372 20588 8424
rect 20628 8372 20680 8424
rect 25504 8415 25556 8424
rect 25504 8381 25513 8415
rect 25513 8381 25547 8415
rect 25547 8381 25556 8415
rect 25504 8372 25556 8381
rect 26240 8372 26292 8424
rect 13268 8304 13320 8356
rect 16672 8304 16724 8356
rect 19524 8304 19576 8356
rect 20168 8304 20220 8356
rect 21456 8304 21508 8356
rect 26148 8304 26200 8356
rect 26792 8304 26844 8356
rect 11244 8236 11296 8288
rect 16304 8279 16356 8288
rect 16304 8245 16313 8279
rect 16313 8245 16347 8279
rect 16347 8245 16356 8279
rect 16304 8236 16356 8245
rect 16764 8279 16816 8288
rect 16764 8245 16773 8279
rect 16773 8245 16807 8279
rect 16807 8245 16816 8279
rect 16764 8236 16816 8245
rect 22652 8236 22704 8288
rect 22928 8236 22980 8288
rect 25136 8279 25188 8288
rect 25136 8245 25145 8279
rect 25145 8245 25179 8279
rect 25179 8245 25188 8279
rect 25136 8236 25188 8245
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 8392 8032 8444 8084
rect 12532 8075 12584 8084
rect 12532 8041 12541 8075
rect 12541 8041 12575 8075
rect 12575 8041 12584 8075
rect 12532 8032 12584 8041
rect 13452 8032 13504 8084
rect 16672 8075 16724 8084
rect 16672 8041 16681 8075
rect 16681 8041 16715 8075
rect 16715 8041 16724 8075
rect 16672 8032 16724 8041
rect 17316 8075 17368 8084
rect 17316 8041 17325 8075
rect 17325 8041 17359 8075
rect 17359 8041 17368 8075
rect 17316 8032 17368 8041
rect 19984 8032 20036 8084
rect 20628 8032 20680 8084
rect 21456 8032 21508 8084
rect 26240 8032 26292 8084
rect 27620 8032 27672 8084
rect 28080 8075 28132 8084
rect 28080 8041 28089 8075
rect 28089 8041 28123 8075
rect 28123 8041 28132 8075
rect 28080 8032 28132 8041
rect 5540 7964 5592 8016
rect 7840 7964 7892 8016
rect 13728 7964 13780 8016
rect 6184 7896 6236 7948
rect 10508 7896 10560 7948
rect 13544 7896 13596 7948
rect 16304 7964 16356 8016
rect 21732 8007 21784 8016
rect 21732 7973 21766 8007
rect 21766 7973 21784 8007
rect 21732 7964 21784 7973
rect 25320 7964 25372 8016
rect 26792 8007 26844 8016
rect 26792 7973 26801 8007
rect 26801 7973 26835 8007
rect 26835 7973 26844 8007
rect 26792 7964 26844 7973
rect 27804 7964 27856 8016
rect 28816 7964 28868 8016
rect 29368 7964 29420 8016
rect 7288 7828 7340 7880
rect 8392 7871 8444 7880
rect 8392 7837 8401 7871
rect 8401 7837 8435 7871
rect 8435 7837 8444 7871
rect 8392 7828 8444 7837
rect 8760 7828 8812 7880
rect 9956 7871 10008 7880
rect 9956 7837 9965 7871
rect 9965 7837 9999 7871
rect 9999 7837 10008 7871
rect 9956 7828 10008 7837
rect 14004 7828 14056 7880
rect 15200 7828 15252 7880
rect 17776 7939 17828 7948
rect 17776 7905 17785 7939
rect 17785 7905 17819 7939
rect 17819 7905 17828 7939
rect 17776 7896 17828 7905
rect 28724 7939 28776 7948
rect 28724 7905 28733 7939
rect 28733 7905 28767 7939
rect 28767 7905 28776 7939
rect 28724 7896 28776 7905
rect 18144 7828 18196 7880
rect 18880 7828 18932 7880
rect 19892 7871 19944 7880
rect 19892 7837 19901 7871
rect 19901 7837 19935 7871
rect 19935 7837 19944 7871
rect 19892 7828 19944 7837
rect 21456 7871 21508 7880
rect 21456 7837 21465 7871
rect 21465 7837 21499 7871
rect 21499 7837 21508 7871
rect 21456 7828 21508 7837
rect 23940 7871 23992 7880
rect 23940 7837 23949 7871
rect 23949 7837 23983 7871
rect 23983 7837 23992 7871
rect 23940 7828 23992 7837
rect 26700 7828 26752 7880
rect 19156 7760 19208 7812
rect 6828 7735 6880 7744
rect 6828 7701 6837 7735
rect 6837 7701 6871 7735
rect 6871 7701 6880 7735
rect 6828 7692 6880 7701
rect 7932 7735 7984 7744
rect 7932 7701 7941 7735
rect 7941 7701 7975 7735
rect 7975 7701 7984 7735
rect 7932 7692 7984 7701
rect 11336 7735 11388 7744
rect 11336 7701 11345 7735
rect 11345 7701 11379 7735
rect 11379 7701 11388 7735
rect 11336 7692 11388 7701
rect 19248 7735 19300 7744
rect 19248 7701 19257 7735
rect 19257 7701 19291 7735
rect 19291 7701 19300 7735
rect 19248 7692 19300 7701
rect 21088 7692 21140 7744
rect 25964 7692 26016 7744
rect 30104 7735 30156 7744
rect 30104 7701 30113 7735
rect 30113 7701 30147 7735
rect 30147 7701 30156 7735
rect 30104 7692 30156 7701
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 8392 7488 8444 7540
rect 9956 7488 10008 7540
rect 10508 7531 10560 7540
rect 10508 7497 10517 7531
rect 10517 7497 10551 7531
rect 10551 7497 10560 7531
rect 10508 7488 10560 7497
rect 5816 7395 5868 7404
rect 5540 7327 5592 7336
rect 5540 7293 5549 7327
rect 5549 7293 5583 7327
rect 5583 7293 5592 7327
rect 5540 7284 5592 7293
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 6736 7284 6788 7336
rect 11244 7395 11296 7404
rect 11244 7361 11253 7395
rect 11253 7361 11287 7395
rect 11287 7361 11296 7395
rect 11244 7352 11296 7361
rect 11704 7327 11756 7336
rect 11704 7293 11713 7327
rect 11713 7293 11747 7327
rect 11747 7293 11756 7327
rect 11704 7284 11756 7293
rect 12532 7284 12584 7336
rect 5816 7216 5868 7268
rect 11336 7216 11388 7268
rect 13360 7216 13412 7268
rect 19248 7488 19300 7540
rect 19892 7488 19944 7540
rect 21732 7488 21784 7540
rect 25320 7531 25372 7540
rect 25320 7497 25329 7531
rect 25329 7497 25363 7531
rect 25363 7497 25372 7531
rect 25320 7488 25372 7497
rect 25964 7531 26016 7540
rect 25964 7497 25973 7531
rect 25973 7497 26007 7531
rect 26007 7497 26016 7531
rect 25964 7488 26016 7497
rect 26424 7488 26476 7540
rect 26608 7488 26660 7540
rect 27804 7531 27856 7540
rect 27804 7497 27813 7531
rect 27813 7497 27847 7531
rect 27847 7497 27856 7531
rect 27804 7488 27856 7497
rect 28724 7531 28776 7540
rect 28724 7497 28733 7531
rect 28733 7497 28767 7531
rect 28767 7497 28776 7531
rect 28724 7488 28776 7497
rect 35256 7488 35308 7540
rect 35532 7488 35584 7540
rect 29276 7395 29328 7404
rect 29276 7361 29285 7395
rect 29285 7361 29319 7395
rect 29319 7361 29328 7395
rect 29276 7352 29328 7361
rect 18052 7284 18104 7336
rect 19156 7327 19208 7336
rect 19156 7293 19190 7327
rect 19190 7293 19208 7327
rect 19156 7284 19208 7293
rect 21456 7284 21508 7336
rect 22928 7284 22980 7336
rect 23940 7327 23992 7336
rect 23940 7293 23949 7327
rect 23949 7293 23983 7327
rect 23983 7293 23992 7327
rect 26424 7327 26476 7336
rect 23940 7284 23992 7293
rect 26424 7293 26433 7327
rect 26433 7293 26467 7327
rect 26467 7293 26476 7327
rect 26424 7284 26476 7293
rect 26516 7284 26568 7336
rect 29368 7284 29420 7336
rect 30104 7284 30156 7336
rect 16304 7216 16356 7268
rect 18144 7216 18196 7268
rect 24216 7259 24268 7268
rect 24216 7225 24250 7259
rect 24250 7225 24268 7259
rect 24216 7216 24268 7225
rect 5172 7191 5224 7200
rect 5172 7157 5181 7191
rect 5181 7157 5215 7191
rect 5215 7157 5224 7191
rect 5172 7148 5224 7157
rect 6184 7191 6236 7200
rect 6184 7157 6193 7191
rect 6193 7157 6227 7191
rect 6227 7157 6236 7191
rect 6184 7148 6236 7157
rect 10692 7191 10744 7200
rect 10692 7157 10701 7191
rect 10701 7157 10735 7191
rect 10735 7157 10744 7191
rect 10692 7148 10744 7157
rect 12900 7148 12952 7200
rect 15200 7148 15252 7200
rect 17040 7191 17092 7200
rect 17040 7157 17049 7191
rect 17049 7157 17083 7191
rect 17083 7157 17092 7191
rect 17040 7148 17092 7157
rect 17776 7148 17828 7200
rect 18236 7148 18288 7200
rect 20260 7191 20312 7200
rect 20260 7157 20269 7191
rect 20269 7157 20303 7191
rect 20303 7157 20312 7191
rect 20260 7148 20312 7157
rect 30380 7148 30432 7200
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 7748 6987 7800 6996
rect 7748 6953 7757 6987
rect 7757 6953 7791 6987
rect 7791 6953 7800 6987
rect 7748 6944 7800 6953
rect 7932 6944 7984 6996
rect 8484 6987 8536 6996
rect 8484 6953 8493 6987
rect 8493 6953 8527 6987
rect 8527 6953 8536 6987
rect 8484 6944 8536 6953
rect 11704 6987 11756 6996
rect 11704 6953 11713 6987
rect 11713 6953 11747 6987
rect 11747 6953 11756 6987
rect 11704 6944 11756 6953
rect 13452 6944 13504 6996
rect 14004 6987 14056 6996
rect 14004 6953 14013 6987
rect 14013 6953 14047 6987
rect 14047 6953 14056 6987
rect 14004 6944 14056 6953
rect 19984 6987 20036 6996
rect 19984 6953 19993 6987
rect 19993 6953 20027 6987
rect 20027 6953 20036 6987
rect 19984 6944 20036 6953
rect 27804 6944 27856 6996
rect 5448 6808 5500 6860
rect 6828 6808 6880 6860
rect 9956 6808 10008 6860
rect 10600 6851 10652 6860
rect 10600 6817 10634 6851
rect 10634 6817 10652 6851
rect 10600 6808 10652 6817
rect 16856 6808 16908 6860
rect 18144 6876 18196 6928
rect 20260 6808 20312 6860
rect 20904 6851 20956 6860
rect 20904 6817 20913 6851
rect 20913 6817 20947 6851
rect 20947 6817 20956 6851
rect 20904 6808 20956 6817
rect 21088 6851 21140 6860
rect 21088 6817 21097 6851
rect 21097 6817 21131 6851
rect 21131 6817 21140 6851
rect 21088 6808 21140 6817
rect 24216 6876 24268 6928
rect 24768 6876 24820 6928
rect 27620 6919 27672 6928
rect 27620 6885 27629 6919
rect 27629 6885 27663 6919
rect 27663 6885 27672 6919
rect 27620 6876 27672 6885
rect 29368 6944 29420 6996
rect 4896 6783 4948 6792
rect 4896 6749 4905 6783
rect 4905 6749 4939 6783
rect 4939 6749 4948 6783
rect 4896 6740 4948 6749
rect 8024 6783 8076 6792
rect 8024 6749 8033 6783
rect 8033 6749 8067 6783
rect 8067 6749 8076 6783
rect 8024 6740 8076 6749
rect 13636 6740 13688 6792
rect 14188 6783 14240 6792
rect 14188 6749 14197 6783
rect 14197 6749 14231 6783
rect 14231 6749 14240 6783
rect 14188 6740 14240 6749
rect 15200 6740 15252 6792
rect 17408 6740 17460 6792
rect 18052 6783 18104 6792
rect 18052 6749 18061 6783
rect 18061 6749 18095 6783
rect 18095 6749 18104 6783
rect 18052 6740 18104 6749
rect 20720 6740 20772 6792
rect 24400 6808 24452 6860
rect 25136 6808 25188 6860
rect 25412 6808 25464 6860
rect 27252 6808 27304 6860
rect 28080 6851 28132 6860
rect 28080 6817 28089 6851
rect 28089 6817 28123 6851
rect 28123 6817 28132 6851
rect 28816 6851 28868 6860
rect 28080 6808 28132 6817
rect 28816 6817 28825 6851
rect 28825 6817 28859 6851
rect 28859 6817 28868 6851
rect 28816 6808 28868 6817
rect 29276 6851 29328 6860
rect 29276 6817 29285 6851
rect 29285 6817 29319 6851
rect 29319 6817 29328 6851
rect 29276 6808 29328 6817
rect 30380 6808 30432 6860
rect 13912 6672 13964 6724
rect 22100 6672 22152 6724
rect 25872 6672 25924 6724
rect 26700 6672 26752 6724
rect 28448 6740 28500 6792
rect 28356 6672 28408 6724
rect 6276 6647 6328 6656
rect 6276 6613 6285 6647
rect 6285 6613 6319 6647
rect 6319 6613 6328 6647
rect 6276 6604 6328 6613
rect 7380 6647 7432 6656
rect 7380 6613 7389 6647
rect 7389 6613 7423 6647
rect 7423 6613 7432 6647
rect 7380 6604 7432 6613
rect 8760 6647 8812 6656
rect 8760 6613 8769 6647
rect 8769 6613 8803 6647
rect 8803 6613 8812 6647
rect 8760 6604 8812 6613
rect 14372 6604 14424 6656
rect 14648 6604 14700 6656
rect 14832 6604 14884 6656
rect 17132 6647 17184 6656
rect 17132 6613 17141 6647
rect 17141 6613 17175 6647
rect 17175 6613 17184 6647
rect 17132 6604 17184 6613
rect 17592 6647 17644 6656
rect 17592 6613 17601 6647
rect 17601 6613 17635 6647
rect 17635 6613 17644 6647
rect 17592 6604 17644 6613
rect 19156 6604 19208 6656
rect 23664 6647 23716 6656
rect 23664 6613 23673 6647
rect 23673 6613 23707 6647
rect 23707 6613 23716 6647
rect 23664 6604 23716 6613
rect 24768 6647 24820 6656
rect 24768 6613 24777 6647
rect 24777 6613 24811 6647
rect 24811 6613 24820 6647
rect 24768 6604 24820 6613
rect 25504 6647 25556 6656
rect 25504 6613 25513 6647
rect 25513 6613 25547 6647
rect 25547 6613 25556 6647
rect 25504 6604 25556 6613
rect 27344 6604 27396 6656
rect 27712 6647 27764 6656
rect 27712 6613 27721 6647
rect 27721 6613 27755 6647
rect 27755 6613 27764 6647
rect 27712 6604 27764 6613
rect 30656 6647 30708 6656
rect 30656 6613 30665 6647
rect 30665 6613 30699 6647
rect 30699 6613 30708 6647
rect 30656 6604 30708 6613
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 4896 6443 4948 6452
rect 4896 6409 4905 6443
rect 4905 6409 4939 6443
rect 4939 6409 4948 6443
rect 4896 6400 4948 6409
rect 5448 6400 5500 6452
rect 8208 6443 8260 6452
rect 8208 6409 8217 6443
rect 8217 6409 8251 6443
rect 8251 6409 8260 6443
rect 8208 6400 8260 6409
rect 9956 6400 10008 6452
rect 11060 6400 11112 6452
rect 13452 6443 13504 6452
rect 13452 6409 13461 6443
rect 13461 6409 13495 6443
rect 13495 6409 13504 6443
rect 13452 6400 13504 6409
rect 16856 6443 16908 6452
rect 16856 6409 16865 6443
rect 16865 6409 16899 6443
rect 16899 6409 16908 6443
rect 16856 6400 16908 6409
rect 17408 6443 17460 6452
rect 17408 6409 17417 6443
rect 17417 6409 17451 6443
rect 17451 6409 17460 6443
rect 17408 6400 17460 6409
rect 19156 6443 19208 6452
rect 19156 6409 19165 6443
rect 19165 6409 19199 6443
rect 19199 6409 19208 6443
rect 19156 6400 19208 6409
rect 19432 6443 19484 6452
rect 19432 6409 19441 6443
rect 19441 6409 19475 6443
rect 19475 6409 19484 6443
rect 19432 6400 19484 6409
rect 21088 6400 21140 6452
rect 24768 6400 24820 6452
rect 25412 6400 25464 6452
rect 26148 6443 26200 6452
rect 26148 6409 26157 6443
rect 26157 6409 26191 6443
rect 26191 6409 26200 6443
rect 26148 6400 26200 6409
rect 28080 6400 28132 6452
rect 28356 6443 28408 6452
rect 28356 6409 28365 6443
rect 28365 6409 28399 6443
rect 28399 6409 28408 6443
rect 28356 6400 28408 6409
rect 30380 6443 30432 6452
rect 6184 6332 6236 6384
rect 13544 6332 13596 6384
rect 10324 6307 10376 6316
rect 10324 6273 10333 6307
rect 10333 6273 10367 6307
rect 10367 6273 10376 6307
rect 10324 6264 10376 6273
rect 10508 6307 10560 6316
rect 10508 6273 10517 6307
rect 10517 6273 10551 6307
rect 10551 6273 10560 6307
rect 10508 6264 10560 6273
rect 14372 6307 14424 6316
rect 6920 6196 6972 6248
rect 8484 6196 8536 6248
rect 9956 6196 10008 6248
rect 10692 6196 10744 6248
rect 13912 6239 13964 6248
rect 8024 6128 8076 6180
rect 10508 6128 10560 6180
rect 13912 6205 13921 6239
rect 13921 6205 13955 6239
rect 13955 6205 13964 6239
rect 13912 6196 13964 6205
rect 14372 6273 14381 6307
rect 14381 6273 14415 6307
rect 14415 6273 14424 6307
rect 14372 6264 14424 6273
rect 17868 6264 17920 6316
rect 19984 6332 20036 6384
rect 18696 6307 18748 6316
rect 18696 6273 18705 6307
rect 18705 6273 18739 6307
rect 18739 6273 18748 6307
rect 18696 6264 18748 6273
rect 19156 6264 19208 6316
rect 20076 6307 20128 6316
rect 20076 6273 20085 6307
rect 20085 6273 20119 6307
rect 20119 6273 20128 6307
rect 20076 6264 20128 6273
rect 20260 6307 20312 6316
rect 20260 6273 20269 6307
rect 20269 6273 20303 6307
rect 20303 6273 20312 6307
rect 20260 6264 20312 6273
rect 17408 6196 17460 6248
rect 19432 6196 19484 6248
rect 25320 6332 25372 6384
rect 29276 6332 29328 6384
rect 26700 6264 26752 6316
rect 28448 6264 28500 6316
rect 30380 6409 30389 6443
rect 30389 6409 30423 6443
rect 30423 6409 30432 6443
rect 30380 6400 30432 6409
rect 30656 6443 30708 6452
rect 30656 6409 30665 6443
rect 30665 6409 30699 6443
rect 30699 6409 30708 6443
rect 30656 6400 30708 6409
rect 29920 6307 29972 6316
rect 29920 6273 29929 6307
rect 29929 6273 29963 6307
rect 29963 6273 29972 6307
rect 29920 6264 29972 6273
rect 21364 6196 21416 6248
rect 23296 6196 23348 6248
rect 23572 6196 23624 6248
rect 26516 6239 26568 6248
rect 26516 6205 26525 6239
rect 26525 6205 26559 6239
rect 26559 6205 26568 6239
rect 26516 6196 26568 6205
rect 28356 6196 28408 6248
rect 29644 6239 29696 6248
rect 29644 6205 29653 6239
rect 29653 6205 29687 6239
rect 29687 6205 29696 6239
rect 29644 6196 29696 6205
rect 30656 6196 30708 6248
rect 20904 6128 20956 6180
rect 21640 6128 21692 6180
rect 24400 6128 24452 6180
rect 12624 6103 12676 6112
rect 12624 6069 12633 6103
rect 12633 6069 12667 6103
rect 12667 6069 12676 6103
rect 12624 6060 12676 6069
rect 13820 6103 13872 6112
rect 13820 6069 13829 6103
rect 13829 6069 13863 6103
rect 13863 6069 13872 6103
rect 13820 6060 13872 6069
rect 14648 6060 14700 6112
rect 15568 6060 15620 6112
rect 16948 6103 17000 6112
rect 16948 6069 16957 6103
rect 16957 6069 16991 6103
rect 16991 6069 17000 6103
rect 16948 6060 17000 6069
rect 17960 6060 18012 6112
rect 18512 6060 18564 6112
rect 21456 6060 21508 6112
rect 22652 6103 22704 6112
rect 22652 6069 22661 6103
rect 22661 6069 22695 6103
rect 22695 6069 22704 6103
rect 22652 6060 22704 6069
rect 22928 6060 22980 6112
rect 23572 6060 23624 6112
rect 27252 6103 27304 6112
rect 27252 6069 27261 6103
rect 27261 6069 27295 6103
rect 27295 6069 27304 6103
rect 27252 6060 27304 6069
rect 27528 6060 27580 6112
rect 29276 6103 29328 6112
rect 29276 6069 29285 6103
rect 29285 6069 29319 6103
rect 29319 6069 29328 6103
rect 29276 6060 29328 6069
rect 31392 6060 31444 6112
rect 33324 6103 33376 6112
rect 33324 6069 33333 6103
rect 33333 6069 33367 6103
rect 33367 6069 33376 6103
rect 33324 6060 33376 6069
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 4620 5856 4672 5908
rect 6276 5856 6328 5908
rect 6920 5899 6972 5908
rect 6920 5865 6929 5899
rect 6929 5865 6963 5899
rect 6963 5865 6972 5899
rect 6920 5856 6972 5865
rect 7932 5856 7984 5908
rect 9956 5899 10008 5908
rect 9956 5865 9965 5899
rect 9965 5865 9999 5899
rect 9999 5865 10008 5899
rect 9956 5856 10008 5865
rect 10600 5856 10652 5908
rect 11244 5856 11296 5908
rect 13636 5899 13688 5908
rect 13636 5865 13645 5899
rect 13645 5865 13679 5899
rect 13679 5865 13688 5899
rect 13636 5856 13688 5865
rect 14372 5856 14424 5908
rect 15568 5856 15620 5908
rect 5448 5788 5500 5840
rect 6184 5788 6236 5840
rect 14188 5788 14240 5840
rect 7380 5720 7432 5772
rect 8300 5720 8352 5772
rect 10600 5720 10652 5772
rect 11704 5720 11756 5772
rect 13636 5720 13688 5772
rect 16212 5720 16264 5772
rect 17592 5856 17644 5908
rect 17868 5899 17920 5908
rect 17868 5865 17877 5899
rect 17877 5865 17911 5899
rect 17911 5865 17920 5899
rect 17868 5856 17920 5865
rect 20076 5856 20128 5908
rect 20260 5899 20312 5908
rect 20260 5865 20269 5899
rect 20269 5865 20303 5899
rect 20303 5865 20312 5899
rect 20260 5856 20312 5865
rect 21364 5899 21416 5908
rect 21364 5865 21373 5899
rect 21373 5865 21407 5899
rect 21407 5865 21416 5899
rect 21364 5856 21416 5865
rect 22100 5899 22152 5908
rect 22100 5865 22109 5899
rect 22109 5865 22143 5899
rect 22143 5865 22152 5899
rect 22100 5856 22152 5865
rect 24400 5899 24452 5908
rect 24400 5865 24409 5899
rect 24409 5865 24443 5899
rect 24443 5865 24452 5899
rect 24400 5856 24452 5865
rect 26516 5856 26568 5908
rect 27712 5856 27764 5908
rect 28356 5899 28408 5908
rect 28356 5865 28365 5899
rect 28365 5865 28399 5899
rect 28399 5865 28408 5899
rect 28356 5856 28408 5865
rect 28448 5856 28500 5908
rect 29920 5856 29972 5908
rect 18696 5788 18748 5840
rect 23020 5788 23072 5840
rect 29644 5788 29696 5840
rect 5816 5652 5868 5704
rect 7196 5695 7248 5704
rect 7196 5661 7205 5695
rect 7205 5661 7239 5695
rect 7239 5661 7248 5695
rect 7196 5652 7248 5661
rect 7748 5652 7800 5704
rect 14096 5695 14148 5704
rect 14096 5661 14105 5695
rect 14105 5661 14139 5695
rect 14139 5661 14148 5695
rect 14096 5652 14148 5661
rect 9036 5584 9088 5636
rect 13360 5584 13412 5636
rect 15108 5652 15160 5704
rect 15844 5695 15896 5704
rect 15844 5661 15853 5695
rect 15853 5661 15887 5695
rect 15887 5661 15896 5695
rect 15844 5652 15896 5661
rect 14832 5584 14884 5636
rect 18052 5720 18104 5772
rect 21916 5763 21968 5772
rect 21916 5729 21925 5763
rect 21925 5729 21959 5763
rect 21959 5729 21968 5763
rect 21916 5720 21968 5729
rect 29276 5720 29328 5772
rect 34336 5763 34388 5772
rect 34336 5729 34345 5763
rect 34345 5729 34379 5763
rect 34379 5729 34388 5763
rect 34336 5720 34388 5729
rect 17868 5652 17920 5704
rect 20904 5695 20956 5704
rect 20904 5661 20913 5695
rect 20913 5661 20947 5695
rect 20947 5661 20956 5695
rect 20904 5652 20956 5661
rect 22928 5652 22980 5704
rect 26792 5652 26844 5704
rect 29184 5695 29236 5704
rect 29184 5661 29193 5695
rect 29193 5661 29227 5695
rect 29227 5661 29236 5695
rect 29184 5652 29236 5661
rect 32680 5695 32732 5704
rect 32680 5661 32689 5695
rect 32689 5661 32723 5695
rect 32723 5661 32732 5695
rect 32680 5652 32732 5661
rect 33968 5652 34020 5704
rect 5632 5559 5684 5568
rect 5632 5525 5641 5559
rect 5641 5525 5675 5559
rect 5675 5525 5684 5559
rect 5632 5516 5684 5525
rect 9312 5516 9364 5568
rect 10692 5559 10744 5568
rect 10692 5525 10701 5559
rect 10701 5525 10735 5559
rect 10735 5525 10744 5559
rect 10692 5516 10744 5525
rect 10968 5516 11020 5568
rect 13820 5516 13872 5568
rect 15016 5559 15068 5568
rect 15016 5525 15025 5559
rect 15025 5525 15059 5559
rect 15059 5525 15068 5559
rect 15016 5516 15068 5525
rect 15108 5516 15160 5568
rect 17684 5516 17736 5568
rect 28356 5584 28408 5636
rect 31944 5627 31996 5636
rect 31944 5593 31953 5627
rect 31953 5593 31987 5627
rect 31987 5593 31996 5627
rect 31944 5584 31996 5593
rect 32496 5584 32548 5636
rect 34244 5584 34296 5636
rect 17960 5516 18012 5568
rect 19340 5559 19392 5568
rect 19340 5525 19349 5559
rect 19349 5525 19383 5559
rect 19383 5525 19392 5559
rect 19340 5516 19392 5525
rect 22468 5559 22520 5568
rect 22468 5525 22477 5559
rect 22477 5525 22511 5559
rect 22511 5525 22520 5559
rect 22468 5516 22520 5525
rect 23020 5516 23072 5568
rect 24952 5559 25004 5568
rect 24952 5525 24961 5559
rect 24961 5525 24995 5559
rect 24995 5525 25004 5559
rect 24952 5516 25004 5525
rect 30564 5559 30616 5568
rect 30564 5525 30573 5559
rect 30573 5525 30607 5559
rect 30607 5525 30616 5559
rect 30564 5516 30616 5525
rect 31208 5559 31260 5568
rect 31208 5525 31217 5559
rect 31217 5525 31251 5559
rect 31251 5525 31260 5559
rect 31208 5516 31260 5525
rect 32312 5559 32364 5568
rect 32312 5525 32321 5559
rect 32321 5525 32355 5559
rect 32355 5525 32364 5559
rect 32312 5516 32364 5525
rect 33140 5559 33192 5568
rect 33140 5525 33149 5559
rect 33149 5525 33183 5559
rect 33183 5525 33192 5559
rect 33140 5516 33192 5525
rect 34520 5516 34572 5568
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 4068 5176 4120 5228
rect 4896 5312 4948 5364
rect 6184 5355 6236 5364
rect 6184 5321 6193 5355
rect 6193 5321 6227 5355
rect 6227 5321 6236 5355
rect 6184 5312 6236 5321
rect 8024 5312 8076 5364
rect 8300 5312 8352 5364
rect 10600 5355 10652 5364
rect 10600 5321 10609 5355
rect 10609 5321 10643 5355
rect 10643 5321 10652 5355
rect 10600 5312 10652 5321
rect 12440 5312 12492 5364
rect 13544 5312 13596 5364
rect 15200 5312 15252 5364
rect 16212 5355 16264 5364
rect 16212 5321 16221 5355
rect 16221 5321 16255 5355
rect 16255 5321 16264 5355
rect 16212 5312 16264 5321
rect 17960 5312 18012 5364
rect 18696 5312 18748 5364
rect 19340 5312 19392 5364
rect 20168 5312 20220 5364
rect 20628 5355 20680 5364
rect 20628 5321 20637 5355
rect 20637 5321 20671 5355
rect 20671 5321 20680 5355
rect 20628 5312 20680 5321
rect 20812 5312 20864 5364
rect 20996 5312 21048 5364
rect 22928 5312 22980 5364
rect 25596 5355 25648 5364
rect 22100 5244 22152 5296
rect 9864 5219 9916 5228
rect 9864 5185 9873 5219
rect 9873 5185 9907 5219
rect 9907 5185 9916 5219
rect 9864 5176 9916 5185
rect 10692 5176 10744 5228
rect 13820 5176 13872 5228
rect 7932 5151 7984 5160
rect 4620 5040 4672 5092
rect 7932 5117 7941 5151
rect 7941 5117 7975 5151
rect 7975 5117 7984 5151
rect 7932 5108 7984 5117
rect 10968 5151 11020 5160
rect 10968 5117 10977 5151
rect 10977 5117 11011 5151
rect 11011 5117 11020 5151
rect 10968 5108 11020 5117
rect 13084 5108 13136 5160
rect 17684 5176 17736 5228
rect 18880 5176 18932 5228
rect 22468 5219 22520 5228
rect 22468 5185 22477 5219
rect 22477 5185 22511 5219
rect 22511 5185 22520 5219
rect 22468 5176 22520 5185
rect 25596 5321 25605 5355
rect 25605 5321 25639 5355
rect 25639 5321 25648 5355
rect 25596 5312 25648 5321
rect 26240 5312 26292 5364
rect 26792 5312 26844 5364
rect 29184 5312 29236 5364
rect 30656 5312 30708 5364
rect 32680 5312 32732 5364
rect 33968 5355 34020 5364
rect 33968 5321 33977 5355
rect 33977 5321 34011 5355
rect 34011 5321 34020 5355
rect 33968 5312 34020 5321
rect 34336 5355 34388 5364
rect 34336 5321 34345 5355
rect 34345 5321 34379 5355
rect 34379 5321 34388 5355
rect 34336 5312 34388 5321
rect 33232 5244 33284 5296
rect 28264 5219 28316 5228
rect 16396 5151 16448 5160
rect 7472 5083 7524 5092
rect 7472 5049 7481 5083
rect 7481 5049 7515 5083
rect 7515 5049 7524 5083
rect 7472 5040 7524 5049
rect 9312 5040 9364 5092
rect 11060 5040 11112 5092
rect 16396 5117 16405 5151
rect 16405 5117 16439 5151
rect 16439 5117 16448 5151
rect 16396 5108 16448 5117
rect 20536 5108 20588 5160
rect 20720 5151 20772 5160
rect 20720 5117 20729 5151
rect 20729 5117 20763 5151
rect 20763 5117 20772 5151
rect 20720 5108 20772 5117
rect 23020 5108 23072 5160
rect 28264 5185 28273 5219
rect 28273 5185 28307 5219
rect 28307 5185 28316 5219
rect 28264 5176 28316 5185
rect 29920 5219 29972 5228
rect 29920 5185 29929 5219
rect 29929 5185 29963 5219
rect 29963 5185 29972 5219
rect 29920 5176 29972 5185
rect 31392 5219 31444 5228
rect 31392 5185 31401 5219
rect 31401 5185 31435 5219
rect 31435 5185 31444 5219
rect 31392 5176 31444 5185
rect 33048 5176 33100 5228
rect 24768 5108 24820 5160
rect 24860 5108 24912 5160
rect 27160 5151 27212 5160
rect 27160 5117 27169 5151
rect 27169 5117 27203 5151
rect 27203 5117 27212 5151
rect 27160 5108 27212 5117
rect 27988 5108 28040 5160
rect 32680 5108 32732 5160
rect 14004 5040 14056 5092
rect 18052 5040 18104 5092
rect 21916 5083 21968 5092
rect 21916 5049 21925 5083
rect 21925 5049 21959 5083
rect 21959 5049 21968 5083
rect 21916 5040 21968 5049
rect 22744 5040 22796 5092
rect 23940 5083 23992 5092
rect 23940 5049 23974 5083
rect 23974 5049 23992 5083
rect 23940 5040 23992 5049
rect 29460 5040 29512 5092
rect 31760 5040 31812 5092
rect 33140 5040 33192 5092
rect 34244 5040 34296 5092
rect 4988 4972 5040 5024
rect 5816 4972 5868 5024
rect 7196 4972 7248 5024
rect 8392 4972 8444 5024
rect 10508 4972 10560 5024
rect 11152 5015 11204 5024
rect 11152 4981 11161 5015
rect 11161 4981 11195 5015
rect 11195 4981 11204 5015
rect 11152 4972 11204 4981
rect 11704 5015 11756 5024
rect 11704 4981 11713 5015
rect 11713 4981 11747 5015
rect 11747 4981 11756 5015
rect 11704 4972 11756 4981
rect 12256 5015 12308 5024
rect 12256 4981 12265 5015
rect 12265 4981 12299 5015
rect 12299 4981 12308 5015
rect 12256 4972 12308 4981
rect 13084 5015 13136 5024
rect 13084 4981 13093 5015
rect 13093 4981 13127 5015
rect 13127 4981 13136 5015
rect 13084 4972 13136 4981
rect 15568 4972 15620 5024
rect 16580 5015 16632 5024
rect 16580 4981 16589 5015
rect 16589 4981 16623 5015
rect 16623 4981 16632 5015
rect 17500 5015 17552 5024
rect 16580 4972 16632 4981
rect 17500 4981 17509 5015
rect 17509 4981 17543 5015
rect 17543 4981 17552 5015
rect 17500 4972 17552 4981
rect 18144 4972 18196 5024
rect 18512 5015 18564 5024
rect 18512 4981 18521 5015
rect 18521 4981 18555 5015
rect 18555 4981 18564 5015
rect 18512 4972 18564 4981
rect 18696 4972 18748 5024
rect 22008 5015 22060 5024
rect 22008 4981 22017 5015
rect 22017 4981 22051 5015
rect 22051 4981 22060 5015
rect 22008 4972 22060 4981
rect 25044 5015 25096 5024
rect 25044 4981 25053 5015
rect 25053 4981 25087 5015
rect 25087 4981 25096 5015
rect 25044 4972 25096 4981
rect 26332 5015 26384 5024
rect 26332 4981 26341 5015
rect 26341 4981 26375 5015
rect 26375 4981 26384 5015
rect 26332 4972 26384 4981
rect 27436 5015 27488 5024
rect 27436 4981 27445 5015
rect 27445 4981 27479 5015
rect 27479 4981 27488 5015
rect 27436 4972 27488 4981
rect 27620 5015 27672 5024
rect 27620 4981 27629 5015
rect 27629 4981 27663 5015
rect 27663 4981 27672 5015
rect 27620 4972 27672 4981
rect 27988 5015 28040 5024
rect 27988 4981 27997 5015
rect 27997 4981 28031 5015
rect 28031 4981 28040 5015
rect 27988 4972 28040 4981
rect 29276 5015 29328 5024
rect 29276 4981 29285 5015
rect 29285 4981 29319 5015
rect 29319 4981 29328 5015
rect 29276 4972 29328 4981
rect 29736 5015 29788 5024
rect 29736 4981 29745 5015
rect 29745 4981 29779 5015
rect 29779 4981 29788 5015
rect 30656 5015 30708 5024
rect 29736 4972 29788 4981
rect 30656 4981 30665 5015
rect 30665 4981 30699 5015
rect 30699 4981 30708 5015
rect 30656 4972 30708 4981
rect 30840 5015 30892 5024
rect 30840 4981 30849 5015
rect 30849 4981 30883 5015
rect 30883 4981 30892 5015
rect 30840 4972 30892 4981
rect 31208 5015 31260 5024
rect 31208 4981 31217 5015
rect 31217 4981 31251 5015
rect 31251 4981 31260 5015
rect 31208 4972 31260 4981
rect 32680 4972 32732 5024
rect 34704 4972 34756 5024
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 4988 4811 5040 4820
rect 4988 4777 4997 4811
rect 4997 4777 5031 4811
rect 5031 4777 5040 4811
rect 4988 4768 5040 4777
rect 5632 4768 5684 4820
rect 6184 4768 6236 4820
rect 8392 4811 8444 4820
rect 8392 4777 8401 4811
rect 8401 4777 8435 4811
rect 8435 4777 8444 4811
rect 8392 4768 8444 4777
rect 9312 4768 9364 4820
rect 10968 4768 11020 4820
rect 13820 4811 13872 4820
rect 13820 4777 13829 4811
rect 13829 4777 13863 4811
rect 13863 4777 13872 4811
rect 13820 4768 13872 4777
rect 6460 4743 6512 4752
rect 6460 4709 6469 4743
rect 6469 4709 6503 4743
rect 6503 4709 6512 4743
rect 6460 4700 6512 4709
rect 8024 4700 8076 4752
rect 10508 4743 10560 4752
rect 10508 4709 10517 4743
rect 10517 4709 10551 4743
rect 10551 4709 10560 4743
rect 10508 4700 10560 4709
rect 10784 4743 10836 4752
rect 10784 4709 10793 4743
rect 10793 4709 10827 4743
rect 10827 4709 10836 4743
rect 10784 4700 10836 4709
rect 12256 4700 12308 4752
rect 15108 4768 15160 4820
rect 17040 4768 17092 4820
rect 17500 4768 17552 4820
rect 17960 4768 18012 4820
rect 19432 4768 19484 4820
rect 19984 4768 20036 4820
rect 22468 4768 22520 4820
rect 23940 4811 23992 4820
rect 23940 4777 23949 4811
rect 23949 4777 23983 4811
rect 23983 4777 23992 4811
rect 23940 4768 23992 4777
rect 24308 4811 24360 4820
rect 24308 4777 24317 4811
rect 24317 4777 24351 4811
rect 24351 4777 24360 4811
rect 24308 4768 24360 4777
rect 25504 4768 25556 4820
rect 25872 4811 25924 4820
rect 25872 4777 25881 4811
rect 25881 4777 25915 4811
rect 25915 4777 25924 4811
rect 25872 4768 25924 4777
rect 26240 4811 26292 4820
rect 26240 4777 26249 4811
rect 26249 4777 26283 4811
rect 26283 4777 26292 4811
rect 26240 4768 26292 4777
rect 28264 4768 28316 4820
rect 29736 4768 29788 4820
rect 29920 4811 29972 4820
rect 29920 4777 29929 4811
rect 29929 4777 29963 4811
rect 29963 4777 29972 4811
rect 29920 4768 29972 4777
rect 31392 4811 31444 4820
rect 31392 4777 31401 4811
rect 31401 4777 31435 4811
rect 31435 4777 31444 4811
rect 31392 4768 31444 4777
rect 31760 4811 31812 4820
rect 31760 4777 31769 4811
rect 31769 4777 31803 4811
rect 31803 4777 31812 4811
rect 31760 4768 31812 4777
rect 32312 4768 32364 4820
rect 33324 4768 33376 4820
rect 34520 4811 34572 4820
rect 34520 4777 34529 4811
rect 34529 4777 34563 4811
rect 34563 4777 34572 4811
rect 34520 4768 34572 4777
rect 16396 4700 16448 4752
rect 16764 4743 16816 4752
rect 16764 4709 16773 4743
rect 16773 4709 16807 4743
rect 16807 4709 16816 4743
rect 16764 4700 16816 4709
rect 23112 4743 23164 4752
rect 23112 4709 23121 4743
rect 23121 4709 23155 4743
rect 23155 4709 23164 4743
rect 23112 4700 23164 4709
rect 24584 4700 24636 4752
rect 27712 4700 27764 4752
rect 29276 4700 29328 4752
rect 31484 4700 31536 4752
rect 4896 4675 4948 4684
rect 4896 4641 4905 4675
rect 4905 4641 4939 4675
rect 4939 4641 4948 4675
rect 4896 4632 4948 4641
rect 6276 4632 6328 4684
rect 7840 4632 7892 4684
rect 9772 4675 9824 4684
rect 9772 4641 9781 4675
rect 9781 4641 9815 4675
rect 9815 4641 9824 4675
rect 9772 4632 9824 4641
rect 9864 4632 9916 4684
rect 11060 4632 11112 4684
rect 11244 4675 11296 4684
rect 11244 4641 11278 4675
rect 11278 4641 11296 4675
rect 15660 4675 15712 4684
rect 11244 4632 11296 4641
rect 15660 4641 15669 4675
rect 15669 4641 15703 4675
rect 15703 4641 15712 4675
rect 15660 4632 15712 4641
rect 17960 4632 18012 4684
rect 20996 4632 21048 4684
rect 21180 4675 21232 4684
rect 21180 4641 21214 4675
rect 21214 4641 21232 4675
rect 21180 4632 21232 4641
rect 23848 4632 23900 4684
rect 27620 4632 27672 4684
rect 28632 4632 28684 4684
rect 30380 4632 30432 4684
rect 34704 4632 34756 4684
rect 4988 4564 5040 4616
rect 4620 4496 4672 4548
rect 8024 4564 8076 4616
rect 14280 4564 14332 4616
rect 15200 4564 15252 4616
rect 16488 4564 16540 4616
rect 18420 4564 18472 4616
rect 18696 4607 18748 4616
rect 18696 4573 18705 4607
rect 18705 4573 18739 4607
rect 18739 4573 18748 4607
rect 18696 4564 18748 4573
rect 19708 4607 19760 4616
rect 19708 4573 19717 4607
rect 19717 4573 19751 4607
rect 19751 4573 19760 4607
rect 19708 4564 19760 4573
rect 5816 4496 5868 4548
rect 14188 4496 14240 4548
rect 15752 4496 15804 4548
rect 16304 4539 16356 4548
rect 16304 4505 16313 4539
rect 16313 4505 16347 4539
rect 16347 4505 16356 4539
rect 16304 4496 16356 4505
rect 17868 4496 17920 4548
rect 19340 4496 19392 4548
rect 24676 4564 24728 4616
rect 26516 4607 26568 4616
rect 24952 4496 25004 4548
rect 26516 4573 26525 4607
rect 26525 4573 26559 4607
rect 26559 4573 26568 4607
rect 26516 4564 26568 4573
rect 30840 4607 30892 4616
rect 30840 4573 30849 4607
rect 30849 4573 30883 4607
rect 30883 4573 30892 4607
rect 30840 4564 30892 4573
rect 33784 4607 33836 4616
rect 26148 4496 26200 4548
rect 27896 4539 27948 4548
rect 27896 4505 27905 4539
rect 27905 4505 27939 4539
rect 27939 4505 27948 4539
rect 27896 4496 27948 4505
rect 33048 4496 33100 4548
rect 6092 4471 6144 4480
rect 6092 4437 6101 4471
rect 6101 4437 6135 4471
rect 6135 4437 6144 4471
rect 6092 4428 6144 4437
rect 7288 4428 7340 4480
rect 7472 4471 7524 4480
rect 7472 4437 7481 4471
rect 7481 4437 7515 4471
rect 7515 4437 7524 4471
rect 7472 4428 7524 4437
rect 8300 4428 8352 4480
rect 12348 4471 12400 4480
rect 12348 4437 12357 4471
rect 12357 4437 12391 4471
rect 12391 4437 12400 4471
rect 12348 4428 12400 4437
rect 12900 4471 12952 4480
rect 12900 4437 12909 4471
rect 12909 4437 12943 4471
rect 12943 4437 12952 4471
rect 12900 4428 12952 4437
rect 13360 4428 13412 4480
rect 13820 4428 13872 4480
rect 14096 4428 14148 4480
rect 15292 4471 15344 4480
rect 15292 4437 15301 4471
rect 15301 4437 15335 4471
rect 15335 4437 15344 4471
rect 15292 4428 15344 4437
rect 19248 4471 19300 4480
rect 19248 4437 19257 4471
rect 19257 4437 19291 4471
rect 19291 4437 19300 4471
rect 19248 4428 19300 4437
rect 20352 4471 20404 4480
rect 20352 4437 20361 4471
rect 20361 4437 20395 4471
rect 20395 4437 20404 4471
rect 20352 4428 20404 4437
rect 23572 4471 23624 4480
rect 23572 4437 23581 4471
rect 23581 4437 23615 4471
rect 23615 4437 23624 4471
rect 23572 4428 23624 4437
rect 27436 4428 27488 4480
rect 29000 4428 29052 4480
rect 30288 4471 30340 4480
rect 30288 4437 30297 4471
rect 30297 4437 30331 4471
rect 30331 4437 30340 4471
rect 30288 4428 30340 4437
rect 33784 4573 33793 4607
rect 33793 4573 33827 4607
rect 33827 4573 33836 4607
rect 33784 4564 33836 4573
rect 35440 4564 35492 4616
rect 34796 4496 34848 4548
rect 36084 4496 36136 4548
rect 34428 4428 34480 4480
rect 35716 4471 35768 4480
rect 35716 4437 35725 4471
rect 35725 4437 35759 4471
rect 35759 4437 35768 4471
rect 35716 4428 35768 4437
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 4068 4267 4120 4276
rect 4068 4233 4077 4267
rect 4077 4233 4111 4267
rect 4111 4233 4120 4267
rect 4068 4224 4120 4233
rect 6184 4267 6236 4276
rect 6184 4233 6193 4267
rect 6193 4233 6227 4267
rect 6227 4233 6236 4267
rect 6184 4224 6236 4233
rect 6460 4224 6512 4276
rect 7932 4224 7984 4276
rect 11060 4267 11112 4276
rect 11060 4233 11069 4267
rect 11069 4233 11103 4267
rect 11103 4233 11112 4267
rect 11060 4224 11112 4233
rect 11152 4224 11204 4276
rect 14004 4224 14056 4276
rect 3056 4131 3108 4140
rect 3056 4097 3065 4131
rect 3065 4097 3099 4131
rect 3099 4097 3108 4131
rect 8024 4156 8076 4208
rect 3056 4088 3108 4097
rect 4068 4020 4120 4072
rect 7932 4131 7984 4140
rect 7932 4097 7941 4131
rect 7941 4097 7975 4131
rect 7975 4097 7984 4131
rect 7932 4088 7984 4097
rect 9036 4131 9088 4140
rect 9036 4097 9045 4131
rect 9045 4097 9079 4131
rect 9079 4097 9088 4131
rect 9036 4088 9088 4097
rect 10508 4088 10560 4140
rect 11888 4088 11940 4140
rect 12348 4088 12400 4140
rect 13728 4088 13780 4140
rect 15660 4224 15712 4276
rect 18420 4224 18472 4276
rect 21180 4224 21232 4276
rect 26516 4224 26568 4276
rect 28264 4267 28316 4276
rect 28264 4233 28273 4267
rect 28273 4233 28307 4267
rect 28307 4233 28316 4267
rect 28264 4224 28316 4233
rect 28632 4267 28684 4276
rect 28632 4233 28641 4267
rect 28641 4233 28675 4267
rect 28675 4233 28684 4267
rect 28632 4224 28684 4233
rect 29460 4267 29512 4276
rect 29460 4233 29469 4267
rect 29469 4233 29503 4267
rect 29503 4233 29512 4267
rect 29460 4224 29512 4233
rect 30380 4267 30432 4276
rect 30380 4233 30389 4267
rect 30389 4233 30423 4267
rect 30423 4233 30432 4267
rect 30380 4224 30432 4233
rect 34704 4267 34756 4276
rect 34704 4233 34713 4267
rect 34713 4233 34747 4267
rect 34747 4233 34756 4267
rect 34704 4224 34756 4233
rect 17776 4131 17828 4140
rect 17776 4097 17785 4131
rect 17785 4097 17819 4131
rect 17819 4097 17828 4131
rect 17776 4088 17828 4097
rect 4988 4020 5040 4072
rect 7472 4020 7524 4072
rect 8392 4020 8444 4072
rect 8484 3952 8536 4004
rect 3332 3927 3384 3936
rect 3332 3893 3341 3927
rect 3341 3893 3375 3927
rect 3375 3893 3384 3927
rect 3332 3884 3384 3893
rect 4896 3884 4948 3936
rect 7288 3927 7340 3936
rect 7288 3893 7297 3927
rect 7297 3893 7331 3927
rect 7331 3893 7340 3927
rect 7288 3884 7340 3893
rect 10784 4020 10836 4072
rect 12164 4063 12216 4072
rect 12164 4029 12173 4063
rect 12173 4029 12207 4063
rect 12207 4029 12216 4063
rect 12164 4020 12216 4029
rect 15016 4020 15068 4072
rect 16764 4063 16816 4072
rect 16764 4029 16773 4063
rect 16773 4029 16807 4063
rect 16807 4029 16816 4063
rect 16764 4020 16816 4029
rect 9864 3952 9916 4004
rect 9772 3927 9824 3936
rect 9772 3893 9781 3927
rect 9781 3893 9815 3927
rect 9815 3893 9824 3927
rect 9772 3884 9824 3893
rect 9956 3927 10008 3936
rect 9956 3893 9965 3927
rect 9965 3893 9999 3927
rect 9999 3893 10008 3927
rect 9956 3884 10008 3893
rect 11888 3927 11940 3936
rect 11888 3893 11897 3927
rect 11897 3893 11931 3927
rect 11931 3893 11940 3927
rect 11888 3884 11940 3893
rect 13728 3952 13780 4004
rect 12900 3927 12952 3936
rect 12900 3893 12909 3927
rect 12909 3893 12943 3927
rect 12943 3893 12952 3927
rect 12900 3884 12952 3893
rect 15660 3927 15712 3936
rect 15660 3893 15669 3927
rect 15669 3893 15703 3927
rect 15703 3893 15712 3927
rect 15660 3884 15712 3893
rect 16672 3927 16724 3936
rect 16672 3893 16681 3927
rect 16681 3893 16715 3927
rect 16715 3893 16724 3927
rect 16672 3884 16724 3893
rect 16948 3927 17000 3936
rect 16948 3893 16957 3927
rect 16957 3893 16991 3927
rect 16991 3893 17000 3927
rect 16948 3884 17000 3893
rect 18052 3884 18104 3936
rect 18880 4063 18932 4072
rect 18880 4029 18914 4063
rect 18914 4029 18932 4063
rect 20352 4156 20404 4208
rect 23572 4156 23624 4208
rect 21548 4088 21600 4140
rect 22836 4131 22888 4140
rect 22836 4097 22845 4131
rect 22845 4097 22879 4131
rect 22879 4097 22888 4131
rect 22836 4088 22888 4097
rect 25596 4156 25648 4208
rect 24676 4131 24728 4140
rect 24676 4097 24685 4131
rect 24685 4097 24719 4131
rect 24719 4097 24728 4131
rect 24676 4088 24728 4097
rect 20996 4063 21048 4072
rect 18880 4020 18932 4029
rect 20996 4029 21005 4063
rect 21005 4029 21039 4063
rect 21039 4029 21048 4063
rect 20996 4020 21048 4029
rect 21456 4063 21508 4072
rect 21456 4029 21465 4063
rect 21465 4029 21499 4063
rect 21499 4029 21508 4063
rect 21456 4020 21508 4029
rect 23664 4020 23716 4072
rect 24308 4020 24360 4072
rect 24768 4020 24820 4072
rect 25504 4020 25556 4072
rect 27712 4088 27764 4140
rect 29000 4131 29052 4140
rect 29000 4097 29009 4131
rect 29009 4097 29043 4131
rect 29043 4097 29052 4131
rect 30012 4131 30064 4140
rect 29000 4088 29052 4097
rect 30012 4097 30021 4131
rect 30021 4097 30055 4131
rect 30055 4097 30064 4131
rect 30840 4156 30892 4208
rect 30012 4088 30064 4097
rect 30748 4088 30800 4140
rect 31760 4088 31812 4140
rect 25872 4063 25924 4072
rect 25872 4029 25906 4063
rect 25906 4029 25924 4063
rect 21088 3927 21140 3936
rect 21088 3893 21097 3927
rect 21097 3893 21131 3927
rect 21131 3893 21140 3927
rect 21088 3884 21140 3893
rect 23848 3952 23900 4004
rect 25872 4020 25924 4029
rect 28264 4020 28316 4072
rect 30380 4020 30432 4072
rect 26516 3952 26568 4004
rect 22376 3884 22428 3936
rect 23296 3884 23348 3936
rect 26976 3927 27028 3936
rect 26976 3893 26985 3927
rect 26985 3893 27019 3927
rect 27019 3893 27028 3927
rect 26976 3884 27028 3893
rect 31668 3952 31720 4004
rect 35164 4020 35216 4072
rect 35716 4063 35768 4072
rect 35716 4029 35750 4063
rect 35750 4029 35768 4063
rect 35716 4020 35768 4029
rect 35256 3952 35308 4004
rect 35532 3952 35584 4004
rect 31208 3927 31260 3936
rect 31208 3893 31217 3927
rect 31217 3893 31251 3927
rect 31251 3893 31260 3927
rect 31852 3927 31904 3936
rect 31208 3884 31260 3893
rect 31852 3893 31861 3927
rect 31861 3893 31895 3927
rect 31895 3893 31904 3927
rect 31852 3884 31904 3893
rect 32128 3927 32180 3936
rect 32128 3893 32137 3927
rect 32137 3893 32171 3927
rect 32171 3893 32180 3927
rect 32128 3884 32180 3893
rect 32956 3884 33008 3936
rect 33692 3927 33744 3936
rect 33692 3893 33701 3927
rect 33701 3893 33735 3927
rect 33735 3893 33744 3927
rect 33692 3884 33744 3893
rect 33784 3884 33836 3936
rect 35900 3884 35952 3936
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 4068 3680 4120 3732
rect 4712 3544 4764 3596
rect 4896 3680 4948 3732
rect 7472 3680 7524 3732
rect 9036 3680 9088 3732
rect 10508 3723 10560 3732
rect 10508 3689 10517 3723
rect 10517 3689 10551 3723
rect 10551 3689 10560 3723
rect 10508 3680 10560 3689
rect 10876 3723 10928 3732
rect 10876 3689 10885 3723
rect 10885 3689 10919 3723
rect 10919 3689 10928 3723
rect 10876 3680 10928 3689
rect 13912 3680 13964 3732
rect 15660 3680 15712 3732
rect 15844 3723 15896 3732
rect 15844 3689 15853 3723
rect 15853 3689 15887 3723
rect 15887 3689 15896 3723
rect 15844 3680 15896 3689
rect 16304 3680 16356 3732
rect 16856 3723 16908 3732
rect 16856 3689 16865 3723
rect 16865 3689 16899 3723
rect 16899 3689 16908 3723
rect 16856 3680 16908 3689
rect 17500 3680 17552 3732
rect 19984 3680 20036 3732
rect 23296 3723 23348 3732
rect 23296 3689 23305 3723
rect 23305 3689 23339 3723
rect 23339 3689 23348 3723
rect 23296 3680 23348 3689
rect 23664 3723 23716 3732
rect 23664 3689 23673 3723
rect 23673 3689 23707 3723
rect 23707 3689 23716 3723
rect 23664 3680 23716 3689
rect 24860 3723 24912 3732
rect 5540 3612 5592 3664
rect 11888 3612 11940 3664
rect 14464 3612 14516 3664
rect 15108 3612 15160 3664
rect 19432 3612 19484 3664
rect 20628 3612 20680 3664
rect 24860 3689 24869 3723
rect 24869 3689 24903 3723
rect 24903 3689 24912 3723
rect 24860 3680 24912 3689
rect 25320 3723 25372 3732
rect 25320 3689 25329 3723
rect 25329 3689 25363 3723
rect 25363 3689 25372 3723
rect 25320 3680 25372 3689
rect 26332 3680 26384 3732
rect 27068 3680 27120 3732
rect 27528 3680 27580 3732
rect 29920 3680 29972 3732
rect 31484 3723 31536 3732
rect 31484 3689 31493 3723
rect 31493 3689 31527 3723
rect 31527 3689 31536 3723
rect 31484 3680 31536 3689
rect 34520 3680 34572 3732
rect 24952 3612 25004 3664
rect 6184 3544 6236 3596
rect 8208 3587 8260 3596
rect 8208 3553 8217 3587
rect 8217 3553 8251 3587
rect 8251 3553 8260 3587
rect 8208 3544 8260 3553
rect 10968 3587 11020 3596
rect 10968 3553 10977 3587
rect 10977 3553 11011 3587
rect 11011 3553 11020 3587
rect 10968 3544 11020 3553
rect 8116 3476 8168 3528
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 8760 3476 8812 3528
rect 11244 3476 11296 3528
rect 12348 3519 12400 3528
rect 12348 3485 12357 3519
rect 12357 3485 12391 3519
rect 12391 3485 12400 3519
rect 12348 3476 12400 3485
rect 16396 3519 16448 3528
rect 16396 3485 16405 3519
rect 16405 3485 16439 3519
rect 16439 3485 16448 3519
rect 16396 3476 16448 3485
rect 17592 3476 17644 3528
rect 17868 3519 17920 3528
rect 17868 3485 17877 3519
rect 17877 3485 17911 3519
rect 17911 3485 17920 3519
rect 17868 3476 17920 3485
rect 18144 3519 18196 3528
rect 18144 3485 18153 3519
rect 18153 3485 18187 3519
rect 18187 3485 18196 3519
rect 18144 3476 18196 3485
rect 20812 3544 20864 3596
rect 21548 3544 21600 3596
rect 23756 3587 23808 3596
rect 23756 3553 23765 3587
rect 23765 3553 23799 3587
rect 23799 3553 23808 3587
rect 23756 3544 23808 3553
rect 25228 3587 25280 3596
rect 25228 3553 25237 3587
rect 25237 3553 25271 3587
rect 25271 3553 25280 3587
rect 34612 3612 34664 3664
rect 25228 3544 25280 3553
rect 27068 3544 27120 3596
rect 28172 3544 28224 3596
rect 31300 3544 31352 3596
rect 32312 3544 32364 3596
rect 33232 3587 33284 3596
rect 33232 3553 33241 3587
rect 33241 3553 33275 3587
rect 33275 3553 33284 3587
rect 33232 3544 33284 3553
rect 34796 3544 34848 3596
rect 19984 3476 20036 3528
rect 20996 3519 21048 3528
rect 20996 3485 21005 3519
rect 21005 3485 21039 3519
rect 21039 3485 21048 3519
rect 20996 3476 21048 3485
rect 25596 3476 25648 3528
rect 26148 3476 26200 3528
rect 28448 3519 28500 3528
rect 28448 3485 28457 3519
rect 28457 3485 28491 3519
rect 28491 3485 28500 3519
rect 28448 3476 28500 3485
rect 32496 3519 32548 3528
rect 32496 3485 32505 3519
rect 32505 3485 32539 3519
rect 32539 3485 32548 3519
rect 32496 3476 32548 3485
rect 32680 3476 32732 3528
rect 33048 3476 33100 3528
rect 36820 3519 36872 3528
rect 2780 3340 2832 3392
rect 4620 3340 4672 3392
rect 19340 3408 19392 3460
rect 31208 3408 31260 3460
rect 32404 3408 32456 3460
rect 35440 3408 35492 3460
rect 6092 3340 6144 3392
rect 6736 3383 6788 3392
rect 6736 3349 6745 3383
rect 6745 3349 6779 3383
rect 6779 3349 6788 3383
rect 6736 3340 6788 3349
rect 9956 3383 10008 3392
rect 9956 3349 9965 3383
rect 9965 3349 9999 3383
rect 9999 3349 10008 3383
rect 9956 3340 10008 3349
rect 13728 3383 13780 3392
rect 13728 3349 13737 3383
rect 13737 3349 13771 3383
rect 13771 3349 13780 3383
rect 13728 3340 13780 3349
rect 14188 3340 14240 3392
rect 15752 3340 15804 3392
rect 22100 3340 22152 3392
rect 23388 3340 23440 3392
rect 24400 3383 24452 3392
rect 24400 3349 24409 3383
rect 24409 3349 24443 3383
rect 24443 3349 24452 3383
rect 24400 3340 24452 3349
rect 24768 3383 24820 3392
rect 24768 3349 24777 3383
rect 24777 3349 24811 3383
rect 24811 3349 24820 3383
rect 24768 3340 24820 3349
rect 27160 3340 27212 3392
rect 28264 3383 28316 3392
rect 28264 3349 28273 3383
rect 28273 3349 28307 3383
rect 28307 3349 28316 3383
rect 28264 3340 28316 3349
rect 31852 3340 31904 3392
rect 32312 3383 32364 3392
rect 32312 3349 32321 3383
rect 32321 3349 32355 3383
rect 32355 3349 32364 3383
rect 32312 3340 32364 3349
rect 34336 3383 34388 3392
rect 34336 3349 34345 3383
rect 34345 3349 34379 3383
rect 34379 3349 34388 3383
rect 34336 3340 34388 3349
rect 35716 3408 35768 3460
rect 36820 3485 36829 3519
rect 36829 3485 36863 3519
rect 36863 3485 36872 3519
rect 36820 3476 36872 3485
rect 36544 3383 36596 3392
rect 36544 3349 36553 3383
rect 36553 3349 36587 3383
rect 36587 3349 36596 3383
rect 36544 3340 36596 3349
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 2044 3179 2096 3188
rect 2044 3145 2053 3179
rect 2053 3145 2087 3179
rect 2087 3145 2096 3179
rect 2044 3136 2096 3145
rect 3792 3179 3844 3188
rect 3792 3145 3801 3179
rect 3801 3145 3835 3179
rect 3835 3145 3844 3179
rect 3792 3136 3844 3145
rect 6184 3179 6236 3188
rect 6184 3145 6193 3179
rect 6193 3145 6227 3179
rect 6227 3145 6236 3179
rect 6184 3136 6236 3145
rect 3884 3068 3936 3120
rect 4160 3111 4212 3120
rect 4160 3077 4169 3111
rect 4169 3077 4203 3111
rect 4203 3077 4212 3111
rect 4160 3068 4212 3077
rect 4068 3000 4120 3052
rect 8116 3136 8168 3188
rect 8392 3136 8444 3188
rect 8852 3136 8904 3188
rect 10968 3136 11020 3188
rect 11244 3179 11296 3188
rect 11244 3145 11253 3179
rect 11253 3145 11287 3179
rect 11287 3145 11296 3179
rect 11244 3136 11296 3145
rect 11888 3179 11940 3188
rect 11888 3145 11897 3179
rect 11897 3145 11931 3179
rect 11931 3145 11940 3179
rect 11888 3136 11940 3145
rect 15752 3136 15804 3188
rect 17040 3179 17092 3188
rect 17040 3145 17049 3179
rect 17049 3145 17083 3179
rect 17083 3145 17092 3179
rect 17040 3136 17092 3145
rect 17500 3179 17552 3188
rect 17500 3145 17509 3179
rect 17509 3145 17543 3179
rect 17543 3145 17552 3179
rect 17500 3136 17552 3145
rect 19984 3179 20036 3188
rect 19984 3145 19993 3179
rect 19993 3145 20027 3179
rect 20027 3145 20036 3179
rect 19984 3136 20036 3145
rect 22836 3136 22888 3188
rect 25228 3136 25280 3188
rect 25504 3136 25556 3188
rect 27160 3179 27212 3188
rect 6644 3000 6696 3052
rect 11060 3000 11112 3052
rect 12348 3000 12400 3052
rect 13452 3043 13504 3052
rect 13452 3009 13461 3043
rect 13461 3009 13495 3043
rect 13495 3009 13504 3043
rect 13452 3000 13504 3009
rect 13912 3000 13964 3052
rect 2044 2932 2096 2984
rect 3792 2932 3844 2984
rect 4896 2932 4948 2984
rect 9772 2975 9824 2984
rect 9772 2941 9781 2975
rect 9781 2941 9815 2975
rect 9815 2941 9824 2975
rect 9772 2932 9824 2941
rect 13268 2932 13320 2984
rect 14832 2932 14884 2984
rect 15108 3000 15160 3052
rect 24584 3068 24636 3120
rect 15568 2932 15620 2984
rect 18052 2975 18104 2984
rect 18052 2941 18061 2975
rect 18061 2941 18095 2975
rect 18095 2941 18104 2975
rect 18052 2932 18104 2941
rect 20444 2932 20496 2984
rect 20720 3000 20772 3052
rect 21456 3000 21508 3052
rect 24400 3000 24452 3052
rect 27160 3145 27169 3179
rect 27169 3145 27203 3179
rect 27203 3145 27212 3179
rect 27160 3136 27212 3145
rect 28448 3136 28500 3188
rect 29184 3136 29236 3188
rect 30748 3179 30800 3188
rect 30748 3145 30757 3179
rect 30757 3145 30791 3179
rect 30791 3145 30800 3179
rect 30748 3136 30800 3145
rect 31300 3179 31352 3188
rect 31300 3145 31309 3179
rect 31309 3145 31343 3179
rect 31343 3145 31352 3179
rect 31300 3136 31352 3145
rect 32496 3136 32548 3188
rect 33232 3136 33284 3188
rect 34796 3136 34848 3188
rect 35256 3179 35308 3188
rect 35256 3145 35265 3179
rect 35265 3145 35299 3179
rect 35299 3145 35308 3179
rect 35256 3136 35308 3145
rect 36820 3179 36872 3188
rect 36820 3145 36829 3179
rect 36829 3145 36863 3179
rect 36863 3145 36872 3179
rect 36820 3136 36872 3145
rect 37372 3179 37424 3188
rect 37372 3145 37381 3179
rect 37381 3145 37415 3179
rect 37415 3145 37424 3179
rect 37372 3136 37424 3145
rect 33968 3068 34020 3120
rect 5908 2864 5960 2916
rect 6736 2864 6788 2916
rect 9956 2864 10008 2916
rect 10968 2864 11020 2916
rect 18236 2864 18288 2916
rect 23756 2864 23808 2916
rect 1676 2796 1728 2848
rect 5540 2796 5592 2848
rect 12992 2839 13044 2848
rect 12992 2805 13001 2839
rect 13001 2805 13035 2839
rect 13035 2805 13044 2839
rect 12992 2796 13044 2805
rect 14648 2796 14700 2848
rect 17500 2796 17552 2848
rect 19340 2796 19392 2848
rect 20076 2796 20128 2848
rect 21916 2796 21968 2848
rect 22376 2839 22428 2848
rect 22376 2805 22385 2839
rect 22385 2805 22419 2839
rect 22419 2805 22428 2839
rect 22376 2796 22428 2805
rect 23388 2796 23440 2848
rect 24768 2864 24820 2916
rect 26976 2932 27028 2984
rect 30012 2932 30064 2984
rect 31944 2932 31996 2984
rect 32404 3000 32456 3052
rect 34336 3000 34388 3052
rect 33048 2932 33100 2984
rect 36544 2932 36596 2984
rect 24952 2796 25004 2848
rect 28172 2839 28224 2848
rect 28172 2805 28181 2839
rect 28181 2805 28215 2839
rect 28215 2805 28224 2839
rect 28172 2796 28224 2805
rect 32680 2796 32732 2848
rect 34428 2796 34480 2848
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 2688 2592 2740 2644
rect 3148 2635 3200 2644
rect 3148 2601 3157 2635
rect 3157 2601 3191 2635
rect 3191 2601 3200 2635
rect 3148 2592 3200 2601
rect 4896 2592 4948 2644
rect 5264 2635 5316 2644
rect 5264 2601 5273 2635
rect 5273 2601 5307 2635
rect 5307 2601 5316 2635
rect 5264 2592 5316 2601
rect 6644 2635 6696 2644
rect 6644 2601 6653 2635
rect 6653 2601 6687 2635
rect 6687 2601 6696 2635
rect 6644 2592 6696 2601
rect 8208 2592 8260 2644
rect 2044 2499 2096 2508
rect 2044 2465 2053 2499
rect 2053 2465 2087 2499
rect 2087 2465 2096 2499
rect 2044 2456 2096 2465
rect 5540 2524 5592 2576
rect 4804 2456 4856 2508
rect 5908 2456 5960 2508
rect 8392 2524 8444 2576
rect 8852 2592 8904 2644
rect 11060 2592 11112 2644
rect 12348 2635 12400 2644
rect 12348 2601 12357 2635
rect 12357 2601 12391 2635
rect 12391 2601 12400 2635
rect 12348 2592 12400 2601
rect 14280 2635 14332 2644
rect 14280 2601 14289 2635
rect 14289 2601 14323 2635
rect 14323 2601 14332 2635
rect 14280 2592 14332 2601
rect 9772 2499 9824 2508
rect 9772 2465 9781 2499
rect 9781 2465 9815 2499
rect 9815 2465 9824 2499
rect 9772 2456 9824 2465
rect 13728 2524 13780 2576
rect 16672 2592 16724 2644
rect 17408 2635 17460 2644
rect 17408 2601 17417 2635
rect 17417 2601 17451 2635
rect 17451 2601 17460 2635
rect 17408 2592 17460 2601
rect 20628 2592 20680 2644
rect 22192 2592 22244 2644
rect 24032 2592 24084 2644
rect 24492 2635 24544 2644
rect 24492 2601 24501 2635
rect 24501 2601 24535 2635
rect 24535 2601 24544 2635
rect 24492 2592 24544 2601
rect 25964 2635 26016 2644
rect 25964 2601 25973 2635
rect 25973 2601 26007 2635
rect 26007 2601 26016 2635
rect 25964 2592 26016 2601
rect 26516 2592 26568 2644
rect 19248 2524 19300 2576
rect 22008 2524 22060 2576
rect 26056 2524 26108 2576
rect 18052 2456 18104 2508
rect 20628 2499 20680 2508
rect 20628 2465 20637 2499
rect 20637 2465 20671 2499
rect 20671 2465 20680 2499
rect 20628 2456 20680 2465
rect 20996 2499 21048 2508
rect 20996 2465 21005 2499
rect 21005 2465 21039 2499
rect 21039 2465 21048 2499
rect 20996 2456 21048 2465
rect 25780 2499 25832 2508
rect 25780 2465 25789 2499
rect 25789 2465 25823 2499
rect 25823 2465 25832 2499
rect 25780 2456 25832 2465
rect 28172 2592 28224 2644
rect 29184 2592 29236 2644
rect 31944 2635 31996 2644
rect 27160 2567 27212 2576
rect 27160 2533 27194 2567
rect 27194 2533 27212 2567
rect 27160 2524 27212 2533
rect 31944 2601 31953 2635
rect 31953 2601 31987 2635
rect 31987 2601 31996 2635
rect 31944 2592 31996 2601
rect 32128 2592 32180 2644
rect 34244 2635 34296 2644
rect 29920 2524 29972 2576
rect 34244 2601 34253 2635
rect 34253 2601 34287 2635
rect 34287 2601 34296 2635
rect 34244 2592 34296 2601
rect 33692 2524 33744 2576
rect 36544 2592 36596 2644
rect 35256 2456 35308 2508
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 23388 2388 23440 2440
rect 4988 2320 5040 2372
rect 572 2252 624 2304
rect 2780 2252 2832 2304
rect 4804 2295 4856 2304
rect 4804 2261 4813 2295
rect 4813 2261 4847 2295
rect 4847 2261 4856 2295
rect 4804 2252 4856 2261
rect 24032 2295 24084 2304
rect 24032 2261 24041 2295
rect 24041 2261 24075 2295
rect 24075 2261 24084 2295
rect 24032 2252 24084 2261
rect 26056 2252 26108 2304
rect 30012 2252 30064 2304
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
<< metal2 >>
rect 9954 39520 10010 40000
rect 29918 39520 29974 40000
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 9968 35193 9996 39520
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 9954 35184 10010 35193
rect 9954 35119 10010 35128
rect 22742 35184 22798 35193
rect 22742 35119 22798 35128
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 22374 27296 22430 27305
rect 4220 27228 4516 27248
rect 22374 27231 22430 27240
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 22388 27130 22416 27231
rect 22376 27124 22428 27130
rect 22376 27066 22428 27072
rect 22388 26926 22416 27066
rect 22376 26920 22428 26926
rect 22376 26862 22428 26868
rect 22652 26784 22704 26790
rect 22650 26752 22652 26761
rect 22704 26752 22706 26761
rect 19580 26684 19876 26704
rect 22650 26687 22706 26696
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 21916 22092 21968 22098
rect 21916 22034 21968 22040
rect 21824 22024 21876 22030
rect 21824 21966 21876 21972
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 21836 21690 21864 21966
rect 21824 21684 21876 21690
rect 21824 21626 21876 21632
rect 20904 21480 20956 21486
rect 20904 21422 20956 21428
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 20076 20800 20128 20806
rect 20076 20742 20128 20748
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 9954 20632 10010 20641
rect 9954 20567 10010 20576
rect 7378 20088 7434 20097
rect 7378 20023 7434 20032
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 7392 18426 7420 20023
rect 9968 18902 9996 20567
rect 18328 20460 18380 20466
rect 18328 20402 18380 20408
rect 17960 19916 18012 19922
rect 17960 19858 18012 19864
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 16948 19712 17000 19718
rect 16948 19654 17000 19660
rect 16592 19310 16620 19654
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 16396 19168 16448 19174
rect 16396 19110 16448 19116
rect 9956 18896 10008 18902
rect 9956 18838 10008 18844
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 7380 18420 7432 18426
rect 7380 18362 7432 18368
rect 7564 18216 7616 18222
rect 7564 18158 7616 18164
rect 7576 17610 7604 18158
rect 9692 18086 9720 18702
rect 9968 18426 9996 18838
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 14924 18624 14976 18630
rect 14924 18566 14976 18572
rect 9956 18420 10008 18426
rect 9956 18362 10008 18368
rect 8944 18080 8996 18086
rect 8944 18022 8996 18028
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 7564 17604 7616 17610
rect 7564 17546 7616 17552
rect 8484 17604 8536 17610
rect 8484 17546 8536 17552
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 8312 17066 8340 17478
rect 8496 17134 8524 17546
rect 8484 17128 8536 17134
rect 8484 17070 8536 17076
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 7562 16824 7618 16833
rect 5448 16788 5500 16794
rect 7562 16759 7618 16768
rect 8116 16788 8168 16794
rect 5448 16730 5500 16736
rect 5460 16697 5488 16730
rect 6000 16720 6052 16726
rect 5446 16688 5502 16697
rect 6000 16662 6052 16668
rect 7010 16688 7066 16697
rect 5446 16623 5502 16632
rect 5264 16584 5316 16590
rect 5264 16526 5316 16532
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 5276 15910 5304 16526
rect 5356 16448 5408 16454
rect 5356 16390 5408 16396
rect 5368 16114 5396 16390
rect 5448 16244 5500 16250
rect 5448 16186 5500 16192
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 4620 15360 4672 15366
rect 4620 15302 4672 15308
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4252 14952 4304 14958
rect 4252 14894 4304 14900
rect 3516 14476 3568 14482
rect 3516 14418 3568 14424
rect 3528 14074 3556 14418
rect 4264 14414 4292 14894
rect 4632 14890 4660 15302
rect 4620 14884 4672 14890
rect 4620 14826 4672 14832
rect 4816 14482 4844 15846
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 5000 14958 5028 15438
rect 4988 14952 5040 14958
rect 4988 14894 5040 14900
rect 4804 14476 4856 14482
rect 4804 14418 4856 14424
rect 3884 14408 3936 14414
rect 3884 14350 3936 14356
rect 4252 14408 4304 14414
rect 4252 14350 4304 14356
rect 3896 14074 3924 14350
rect 5276 14278 5304 15846
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 5460 14090 5488 16186
rect 6012 15910 6040 16662
rect 6276 16652 6328 16658
rect 7010 16623 7066 16632
rect 6276 16594 6328 16600
rect 6288 15910 6316 16594
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 6276 15904 6328 15910
rect 6276 15846 6328 15852
rect 6012 15570 6040 15846
rect 6000 15564 6052 15570
rect 6000 15506 6052 15512
rect 6012 14890 6040 15506
rect 6288 15366 6316 15846
rect 6656 15366 6684 16050
rect 6276 15360 6328 15366
rect 6276 15302 6328 15308
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6000 14884 6052 14890
rect 6000 14826 6052 14832
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5644 14482 5672 14758
rect 5632 14476 5684 14482
rect 5632 14418 5684 14424
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5460 14074 5580 14090
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3884 14068 3936 14074
rect 5460 14068 5592 14074
rect 5460 14062 5540 14068
rect 3884 14010 3936 14016
rect 5540 14010 5592 14016
rect 3896 13870 3924 14010
rect 5644 13870 5672 14214
rect 6288 14006 6316 14350
rect 6276 14000 6328 14006
rect 6276 13942 6328 13948
rect 3884 13864 3936 13870
rect 3884 13806 3936 13812
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 3896 13530 3924 13806
rect 5080 13728 5132 13734
rect 5080 13670 5132 13676
rect 5092 13530 5120 13670
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 5080 13524 5132 13530
rect 5080 13466 5132 13472
rect 3896 12986 3924 13466
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 5000 12986 5028 13330
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 3896 12782 3924 12922
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 3896 11898 3924 12718
rect 5000 12374 5028 12922
rect 5092 12782 5120 13466
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5080 12776 5132 12782
rect 5080 12718 5132 12724
rect 5092 12442 5120 12718
rect 5368 12646 5396 13262
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 4988 12368 5040 12374
rect 4988 12310 5040 12316
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 3896 11694 3924 11834
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3804 10810 3832 10950
rect 3896 10810 3924 11630
rect 4724 11354 4752 12242
rect 5000 11694 5028 12310
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 5184 11354 5212 11494
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 4264 10130 4292 10610
rect 5184 10538 5212 11290
rect 5368 11150 5396 12582
rect 5460 12442 5488 13126
rect 6288 12986 6316 13942
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5460 11354 5488 12378
rect 6288 12238 6316 12922
rect 6656 12646 6684 15302
rect 7024 14618 7052 16623
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7472 16448 7524 16454
rect 7472 16390 7524 16396
rect 7208 16046 7236 16390
rect 7484 16182 7512 16390
rect 7472 16176 7524 16182
rect 7472 16118 7524 16124
rect 7576 16114 7604 16759
rect 8116 16730 8168 16736
rect 7932 16720 7984 16726
rect 7932 16662 7984 16668
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 7116 15706 7144 15846
rect 7104 15700 7156 15706
rect 7104 15642 7156 15648
rect 7576 15638 7604 16050
rect 7564 15632 7616 15638
rect 7564 15574 7616 15580
rect 7944 14890 7972 16662
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 7932 14884 7984 14890
rect 7932 14826 7984 14832
rect 7944 14618 7972 14826
rect 8036 14618 8064 15642
rect 8128 15450 8156 16730
rect 8312 16726 8340 17002
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8404 16794 8432 16934
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 8312 16538 8340 16662
rect 8220 16510 8340 16538
rect 8496 16522 8524 17070
rect 8484 16516 8536 16522
rect 8220 15638 8248 16510
rect 8484 16458 8536 16464
rect 8496 16250 8524 16458
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8496 16046 8524 16186
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8312 15450 8340 15506
rect 8128 15422 8340 15450
rect 8128 15162 8156 15422
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6748 13870 6776 14214
rect 7116 14074 7144 14418
rect 7392 14074 7420 14554
rect 8312 14482 8340 15302
rect 8496 14958 8524 15982
rect 8668 15496 8720 15502
rect 8668 15438 8720 15444
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8680 14618 8708 15438
rect 8956 15065 8984 18022
rect 9588 16720 9640 16726
rect 9218 16688 9274 16697
rect 9588 16662 9640 16668
rect 9218 16623 9274 16632
rect 9232 16046 9260 16623
rect 9600 16266 9628 16662
rect 9692 16590 9720 18022
rect 11072 16946 11100 18566
rect 14936 18290 14964 18566
rect 15856 18290 15884 19110
rect 16408 18970 16436 19110
rect 16396 18964 16448 18970
rect 16396 18906 16448 18912
rect 16212 18828 16264 18834
rect 16212 18770 16264 18776
rect 15936 18624 15988 18630
rect 15936 18566 15988 18572
rect 15948 18426 15976 18566
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 14924 18284 14976 18290
rect 14924 18226 14976 18232
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 16224 18222 16252 18770
rect 16304 18624 16356 18630
rect 16304 18566 16356 18572
rect 16212 18216 16264 18222
rect 16212 18158 16264 18164
rect 15200 18080 15252 18086
rect 15120 18028 15200 18034
rect 15120 18022 15252 18028
rect 15120 18006 15240 18022
rect 15120 17882 15148 18006
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 15764 17134 15792 17818
rect 16224 17542 16252 18158
rect 16316 18086 16344 18566
rect 16408 18222 16436 18906
rect 16684 18306 16712 19314
rect 16856 18420 16908 18426
rect 16856 18362 16908 18368
rect 16500 18290 16712 18306
rect 16488 18284 16712 18290
rect 16540 18278 16712 18284
rect 16488 18226 16540 18232
rect 16396 18216 16448 18222
rect 16396 18158 16448 18164
rect 16486 18184 16542 18193
rect 16486 18119 16542 18128
rect 16500 18086 16528 18119
rect 16304 18080 16356 18086
rect 16304 18022 16356 18028
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 16316 17678 16344 18022
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16212 17536 16264 17542
rect 16212 17478 16264 17484
rect 16224 17338 16252 17478
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15752 17128 15804 17134
rect 15752 17070 15804 17076
rect 15384 16992 15436 16998
rect 10980 16918 11100 16946
rect 15290 16960 15346 16969
rect 9770 16824 9826 16833
rect 9770 16759 9826 16768
rect 9784 16658 9812 16759
rect 10980 16658 11008 16918
rect 15384 16934 15436 16940
rect 15290 16895 15346 16904
rect 15304 16794 15332 16895
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 11072 16697 11100 16730
rect 11058 16688 11114 16697
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 10968 16652 11020 16658
rect 11058 16623 11114 16632
rect 10968 16594 11020 16600
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9692 16402 9720 16526
rect 9692 16374 9812 16402
rect 9600 16250 9720 16266
rect 9600 16244 9732 16250
rect 9600 16238 9680 16244
rect 9680 16186 9732 16192
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 9784 15706 9812 16374
rect 10980 16250 11008 16594
rect 15396 16590 15424 16934
rect 15384 16584 15436 16590
rect 15384 16526 15436 16532
rect 15396 16250 15424 16526
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 8942 15056 8998 15065
rect 8942 14991 8998 15000
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 7380 14068 7432 14074
rect 7380 14010 7432 14016
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6932 13530 6960 13806
rect 8312 13530 8340 14418
rect 8680 14414 8708 14554
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8496 14074 8524 14214
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7392 12782 7420 13126
rect 8496 12782 8524 13330
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7932 12776 7984 12782
rect 7932 12718 7984 12724
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 6828 12708 6880 12714
rect 6828 12650 6880 12656
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 6288 11354 6316 12174
rect 6840 11898 6868 12650
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7116 12102 7144 12582
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 6932 11898 6960 12038
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 6644 11620 6696 11626
rect 6644 11562 6696 11568
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6656 11286 6684 11562
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5356 11144 5408 11150
rect 5356 11086 5408 11092
rect 5460 10810 5488 11154
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 4804 10532 4856 10538
rect 4804 10474 4856 10480
rect 5172 10532 5224 10538
rect 5172 10474 5224 10480
rect 4816 10266 4844 10474
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 5460 10198 5488 10746
rect 6288 10742 6316 11086
rect 6276 10736 6328 10742
rect 6276 10678 6328 10684
rect 6656 10266 6684 11222
rect 7012 10736 7064 10742
rect 7012 10678 7064 10684
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 5092 9722 5120 10066
rect 5460 9722 5488 10134
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 5448 9716 5500 9722
rect 5448 9658 5500 9664
rect 7024 8974 7052 10678
rect 7300 10606 7328 12582
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7484 11762 7512 12038
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7484 9450 7512 11698
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7668 11082 7696 11494
rect 7656 11076 7708 11082
rect 7656 11018 7708 11024
rect 7944 10266 7972 12718
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 8128 10742 8156 11630
rect 8312 11558 8340 12242
rect 8680 12238 8708 13806
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9416 12442 9444 13262
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 9508 12238 9536 13806
rect 9784 12918 9812 15642
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 14568 15026 14596 15302
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14096 14884 14148 14890
rect 14096 14826 14148 14832
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13924 14618 13952 14758
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 9864 14476 9916 14482
rect 9864 14418 9916 14424
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 9876 13870 9904 14418
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 9864 13524 9916 13530
rect 9968 13512 9996 13670
rect 10060 13530 10088 14214
rect 10796 13734 10824 14214
rect 11164 14074 11192 14350
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10784 13728 10836 13734
rect 10784 13670 10836 13676
rect 10888 13530 10916 13874
rect 11164 13870 11192 14010
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 9916 13484 9996 13512
rect 10048 13524 10100 13530
rect 9864 13466 9916 13472
rect 10048 13466 10100 13472
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10060 12986 10088 13466
rect 11256 13326 11284 14418
rect 12544 14074 12572 14418
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12532 13864 12584 13870
rect 12636 13818 12664 14418
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13464 13938 13492 14214
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 12584 13812 12664 13818
rect 12532 13806 12664 13812
rect 12440 13796 12492 13802
rect 12544 13790 12664 13806
rect 12440 13738 12492 13744
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11072 12986 11100 13262
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 9772 12912 9824 12918
rect 9772 12854 9824 12860
rect 9588 12776 9640 12782
rect 9640 12724 9720 12730
rect 9588 12718 9720 12724
rect 9600 12702 9720 12718
rect 9692 12442 9720 12702
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 8496 11898 8524 12174
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8300 11552 8352 11558
rect 8220 11500 8300 11506
rect 8220 11494 8352 11500
rect 8220 11478 8340 11494
rect 8220 10810 8248 11478
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8116 10736 8168 10742
rect 8116 10678 8168 10684
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 8312 10130 8340 10950
rect 8300 10124 8352 10130
rect 8128 10084 8300 10112
rect 8128 9654 8156 10084
rect 8300 10066 8352 10072
rect 8116 9648 8168 9654
rect 8116 9590 8168 9596
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7472 9444 7524 9450
rect 7472 9386 7524 9392
rect 7852 9382 7880 9454
rect 8404 9382 8432 11290
rect 8484 11280 8536 11286
rect 8484 11222 8536 11228
rect 8496 10606 8524 11222
rect 8680 11082 8708 12174
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 9048 11694 9076 11834
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 9048 11150 9076 11630
rect 9312 11620 9364 11626
rect 9312 11562 9364 11568
rect 9036 11144 9088 11150
rect 9036 11086 9088 11092
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 9324 11014 9352 11562
rect 9508 11354 9536 12174
rect 9784 11898 9812 12854
rect 11256 12782 11284 13262
rect 12452 13190 12480 13738
rect 12636 13530 12664 13790
rect 12808 13728 12860 13734
rect 12808 13670 12860 13676
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 10416 12708 10468 12714
rect 10416 12650 10468 12656
rect 10428 12374 10456 12650
rect 12820 12442 12848 13670
rect 13280 13190 13308 13670
rect 13464 13530 13492 13874
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 14002 13696 14058 13705
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13268 13184 13320 13190
rect 13266 13152 13268 13161
rect 13320 13152 13322 13161
rect 13266 13087 13322 13096
rect 13464 12714 13492 13466
rect 13452 12708 13504 12714
rect 13452 12650 13504 12656
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 12808 12436 12860 12442
rect 12808 12378 12860 12384
rect 10416 12368 10468 12374
rect 10416 12310 10468 12316
rect 10428 11898 10456 12310
rect 11060 12300 11112 12306
rect 11244 12300 11296 12306
rect 11112 12260 11192 12288
rect 11060 12242 11112 12248
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 9496 11348 9548 11354
rect 9496 11290 9548 11296
rect 9588 11076 9640 11082
rect 9588 11018 9640 11024
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9508 10810 9536 10950
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 8484 10600 8536 10606
rect 8484 10542 8536 10548
rect 8496 10266 8524 10542
rect 9600 10266 9628 11018
rect 9784 10810 9812 11834
rect 10508 11212 10560 11218
rect 10508 11154 10560 11160
rect 10520 10810 10548 11154
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 8496 9722 8524 10202
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8588 9722 8616 9998
rect 8484 9716 8536 9722
rect 8484 9658 8536 9664
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 8588 9450 8616 9658
rect 8576 9444 8628 9450
rect 8576 9386 8628 9392
rect 9692 9382 9720 10066
rect 7840 9376 7892 9382
rect 7838 9344 7840 9353
rect 8392 9376 8444 9382
rect 7892 9344 7894 9353
rect 8392 9318 8444 9324
rect 8944 9376 8996 9382
rect 9680 9376 9732 9382
rect 8944 9318 8996 9324
rect 9402 9344 9458 9353
rect 7838 9279 7894 9288
rect 8956 9217 8984 9318
rect 9680 9318 9732 9324
rect 9402 9279 9458 9288
rect 8942 9208 8998 9217
rect 8942 9143 8998 9152
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 6840 8430 6868 8910
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6932 8362 6960 8774
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6184 8288 6236 8294
rect 6932 8242 6960 8298
rect 6184 8230 6236 8236
rect 5540 8016 5592 8022
rect 5540 7958 5592 7964
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 5552 7342 5580 7958
rect 6196 7954 6224 8230
rect 6748 8214 6960 8242
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5828 7274 5856 7346
rect 5816 7268 5868 7274
rect 5816 7210 5868 7216
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5184 7041 5212 7142
rect 5170 7032 5226 7041
rect 5170 6967 5226 6976
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 4896 6792 4948 6798
rect 4894 6760 4896 6769
rect 4948 6760 4950 6769
rect 4894 6695 4950 6704
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 4908 6458 4936 6695
rect 5460 6458 5488 6802
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 4080 4282 4108 5170
rect 4632 5098 4660 5850
rect 4908 5370 4936 6394
rect 5460 5846 5488 6394
rect 5448 5840 5500 5846
rect 5448 5782 5500 5788
rect 5828 5710 5856 7210
rect 6196 7206 6224 7890
rect 6748 7342 6776 8214
rect 7300 7886 7328 8978
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 7840 8560 7892 8566
rect 7840 8502 7892 8508
rect 7852 8022 7880 8502
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 7840 8016 7892 8022
rect 7840 7958 7892 7964
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 6196 6390 6224 7142
rect 6840 6866 6868 7686
rect 7746 7032 7802 7041
rect 7944 7002 7972 7686
rect 7746 6967 7748 6976
rect 7800 6967 7802 6976
rect 7932 6996 7984 7002
rect 7748 6938 7800 6944
rect 7932 6938 7984 6944
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 6184 6384 6236 6390
rect 6184 6326 6236 6332
rect 6288 5914 6316 6598
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6932 5914 6960 6190
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6184 5840 6236 5846
rect 6184 5782 6236 5788
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 4620 5092 4672 5098
rect 4620 5034 4672 5040
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 5000 4826 5028 4966
rect 5644 4826 5672 5510
rect 5828 5030 5856 5646
rect 6196 5370 6224 5782
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4620 4548 4672 4554
rect 4620 4490 4672 4496
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 3054 4176 3110 4185
rect 3054 4111 3056 4120
rect 3108 4111 3110 4120
rect 3056 4082 3108 4088
rect 4080 4078 4108 4218
rect 4068 4072 4120 4078
rect 3330 4040 3386 4049
rect 4068 4014 4120 4020
rect 3330 3975 3386 3984
rect 3344 3942 3372 3975
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 2042 3768 2098 3777
rect 2042 3703 2098 3712
rect 3790 3768 3846 3777
rect 4080 3738 4108 4014
rect 3790 3703 3846 3712
rect 4068 3732 4120 3738
rect 2056 3194 2084 3703
rect 2780 3392 2832 3398
rect 2700 3340 2780 3346
rect 2700 3334 2832 3340
rect 2700 3318 2820 3334
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 2056 2990 2084 3130
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 572 2304 624 2310
rect 572 2246 624 2252
rect 584 480 612 2246
rect 1688 480 1716 2790
rect 2700 2650 2728 3318
rect 3804 3194 3832 3703
rect 4068 3674 4120 3680
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3804 2990 3832 3130
rect 3884 3120 3936 3126
rect 3884 3062 3936 3068
rect 3792 2984 3844 2990
rect 3792 2926 3844 2932
rect 3146 2680 3202 2689
rect 2688 2644 2740 2650
rect 3146 2615 3148 2624
rect 2688 2586 2740 2592
rect 3200 2615 3202 2624
rect 3148 2586 3200 2592
rect 2042 2544 2098 2553
rect 2042 2479 2044 2488
rect 2096 2479 2098 2488
rect 2044 2450 2096 2456
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 2792 480 2820 2246
rect 3896 480 3924 3062
rect 4080 3058 4108 3674
rect 4632 3398 4660 4490
rect 4908 3942 4936 4626
rect 5000 4622 5028 4762
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 5000 4078 5028 4558
rect 5828 4554 5856 4966
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 5816 4548 5868 4554
rect 5816 4490 5868 4496
rect 4988 4072 5040 4078
rect 4988 4014 5040 4020
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 5262 3904 5318 3913
rect 4908 3738 4936 3878
rect 5262 3839 5318 3848
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 4160 3120 4212 3126
rect 4158 3088 4160 3097
rect 4724 3097 4752 3538
rect 4212 3088 4214 3097
rect 4068 3052 4120 3058
rect 4158 3023 4214 3032
rect 4710 3088 4766 3097
rect 4710 3023 4766 3032
rect 4068 2994 4120 3000
rect 4908 2990 4936 3674
rect 4896 2984 4948 2990
rect 4896 2926 4948 2932
rect 4908 2650 4936 2926
rect 5276 2650 5304 3839
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 5552 2854 5580 3606
rect 5828 3505 5856 4490
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6104 4185 6132 4422
rect 6196 4282 6224 4762
rect 6288 4690 6316 5850
rect 7392 5778 7420 6598
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 7760 5710 7788 6938
rect 7944 5914 7972 6938
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 8036 6186 8064 6734
rect 8220 6458 8248 8298
rect 8404 8090 8432 8774
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8392 8084 8444 8090
rect 8444 8044 8524 8072
rect 8392 8026 8444 8032
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8404 7546 8432 7822
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8496 7002 8524 8044
rect 8772 7886 8800 8230
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8496 6254 8524 6938
rect 8772 6662 8800 7822
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 7196 5704 7248 5710
rect 7194 5672 7196 5681
rect 7748 5704 7800 5710
rect 7248 5672 7250 5681
rect 7748 5646 7800 5652
rect 7194 5607 7250 5616
rect 8036 5370 8064 6122
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8312 5370 8340 5714
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 7932 5160 7984 5166
rect 7470 5128 7526 5137
rect 7932 5102 7984 5108
rect 7470 5063 7472 5072
rect 7524 5063 7526 5072
rect 7472 5034 7524 5040
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 6460 4752 6512 4758
rect 6460 4694 6512 4700
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 6472 4282 6500 4694
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 6460 4276 6512 4282
rect 6460 4218 6512 4224
rect 6090 4176 6146 4185
rect 6090 4111 6146 4120
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 5814 3496 5870 3505
rect 5814 3431 5870 3440
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 5552 2582 5580 2790
rect 5540 2576 5592 2582
rect 5540 2518 5592 2524
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 4816 2310 4844 2450
rect 5828 2446 5856 3431
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 5908 2916 5960 2922
rect 5908 2858 5960 2864
rect 5920 2514 5948 2858
rect 5908 2508 5960 2514
rect 5908 2450 5960 2456
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 4988 2372 5040 2378
rect 4988 2314 5040 2320
rect 4804 2304 4856 2310
rect 4804 2246 4856 2252
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 4816 2145 4844 2246
rect 4802 2136 4858 2145
rect 4802 2071 4858 2080
rect 5000 480 5028 2314
rect 6104 480 6132 3334
rect 6196 3194 6224 3538
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6656 2650 6684 2994
rect 6748 2922 6776 3334
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 7208 480 7236 4966
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7300 3942 7328 4422
rect 7484 4078 7512 4422
rect 7852 4162 7880 4626
rect 7944 4282 7972 5102
rect 8036 4758 8064 5306
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 8404 4826 8432 4966
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8024 4752 8076 4758
rect 8024 4694 8076 4700
rect 8036 4622 8064 4694
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 7932 4276 7984 4282
rect 7932 4218 7984 4224
rect 8036 4214 8064 4558
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8024 4208 8076 4214
rect 7930 4176 7986 4185
rect 7852 4134 7930 4162
rect 8024 4150 8076 4156
rect 7930 4111 7932 4120
rect 7984 4111 7986 4120
rect 7932 4082 7984 4088
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7288 3936 7340 3942
rect 7286 3904 7288 3913
rect 7340 3904 7342 3913
rect 7286 3839 7342 3848
rect 7484 3738 7512 4014
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8128 3194 8156 3470
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8220 2650 8248 3538
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 8312 480 8340 4422
rect 8404 4078 8432 4762
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8482 4040 8538 4049
rect 8482 3975 8484 3984
rect 8536 3975 8538 3984
rect 8484 3946 8536 3952
rect 8772 3534 8800 6598
rect 9036 5636 9088 5642
rect 9036 5578 9088 5584
rect 9048 4146 9076 5578
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9324 5098 9352 5510
rect 9312 5092 9364 5098
rect 9312 5034 9364 5040
rect 9324 4826 9352 5034
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 9048 3738 9076 4082
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 8392 3528 8444 3534
rect 8390 3496 8392 3505
rect 8760 3528 8812 3534
rect 8444 3496 8446 3505
rect 8760 3470 8812 3476
rect 8390 3431 8446 3440
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 8404 2582 8432 3130
rect 8864 2650 8892 3130
rect 8852 2644 8904 2650
rect 8852 2586 8904 2592
rect 8392 2576 8444 2582
rect 8392 2518 8444 2524
rect 9416 480 9444 9279
rect 10414 9208 10470 9217
rect 10414 9143 10470 9152
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 9968 7546 9996 7822
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 9968 6866 9996 7482
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9968 6458 9996 6802
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 10336 6322 10364 8502
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 9968 5914 9996 6190
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 9862 5264 9918 5273
rect 9862 5199 9864 5208
rect 9916 5199 9918 5208
rect 9864 5170 9916 5176
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 9784 3942 9812 4626
rect 9876 4010 9904 4626
rect 9954 4040 10010 4049
rect 9864 4004 9916 4010
rect 9954 3975 10010 3984
rect 9864 3946 9916 3952
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9784 3505 9812 3878
rect 9876 3754 9904 3946
rect 9968 3942 9996 3975
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9876 3726 9996 3754
rect 9770 3496 9826 3505
rect 9770 3431 9826 3440
rect 9968 3398 9996 3726
rect 10428 3618 10456 9143
rect 10612 8974 10640 10610
rect 10980 10266 11008 12038
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10968 10124 11020 10130
rect 11072 10112 11100 12038
rect 11164 10606 11192 12260
rect 11244 12242 11296 12248
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 11256 11558 11284 12242
rect 12728 11898 12756 12242
rect 13728 12232 13780 12238
rect 13832 12220 13860 12582
rect 13780 12192 13860 12220
rect 13728 12174 13780 12180
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12716 11620 12768 11626
rect 12716 11562 12768 11568
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 12256 10464 12308 10470
rect 12452 10452 12480 11154
rect 12728 11150 12756 11562
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12728 10674 12756 11086
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12308 10424 12480 10452
rect 12256 10406 12308 10412
rect 11020 10084 11100 10112
rect 10968 10066 11020 10072
rect 10980 9722 11008 10066
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 12268 9654 12296 10406
rect 12728 10130 12756 10610
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 12728 9722 12756 10066
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12256 9648 12308 9654
rect 12256 9590 12308 9596
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10612 8634 10640 8910
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10796 8430 10824 8774
rect 10888 8537 10916 8978
rect 10874 8528 10930 8537
rect 10874 8463 10876 8472
rect 10928 8463 10930 8472
rect 10876 8434 10928 8440
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10520 7546 10548 7890
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10612 6866 10640 8366
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11256 7410 11284 8230
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10520 6225 10548 6258
rect 10506 6216 10562 6225
rect 10506 6151 10508 6160
rect 10560 6151 10562 6160
rect 10508 6122 10560 6128
rect 10520 6091 10548 6122
rect 10612 5914 10640 6802
rect 10704 6254 10732 7142
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 10612 5409 10640 5714
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 10598 5400 10654 5409
rect 10598 5335 10600 5344
rect 10652 5335 10654 5344
rect 10600 5306 10652 5312
rect 10704 5234 10732 5510
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10980 5166 11008 5510
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10782 4992 10838 5001
rect 10520 4865 10548 4966
rect 10782 4927 10838 4936
rect 10506 4856 10562 4865
rect 10506 4791 10562 4800
rect 10520 4758 10548 4791
rect 10796 4758 10824 4927
rect 10980 4826 11008 5102
rect 11072 5098 11100 6394
rect 11256 5914 11284 7346
rect 11348 7274 11376 7686
rect 11336 7268 11388 7274
rect 11336 7210 11388 7216
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11060 5092 11112 5098
rect 11060 5034 11112 5040
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 10508 4752 10560 4758
rect 10508 4694 10560 4700
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 10874 4720 10930 4729
rect 10520 4146 10548 4694
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10796 4078 10824 4694
rect 11072 4690 11100 5034
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 10874 4655 10930 4664
rect 11060 4684 11112 4690
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10506 3904 10562 3913
rect 10506 3839 10562 3848
rect 10520 3738 10548 3839
rect 10888 3738 10916 4655
rect 11060 4626 11112 4632
rect 11072 4282 11100 4626
rect 11164 4282 11192 4966
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 10508 3732 10560 3738
rect 10508 3674 10560 3680
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10966 3632 11022 3641
rect 10428 3590 10548 3618
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 9784 2514 9812 2926
rect 9968 2922 9996 3334
rect 9956 2916 10008 2922
rect 9956 2858 10008 2864
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 10520 480 10548 3590
rect 10966 3567 10968 3576
rect 11020 3567 11022 3576
rect 10968 3538 11020 3544
rect 10980 3194 11008 3538
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 11072 3058 11100 4218
rect 11256 3534 11284 4626
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11256 3194 11284 3470
rect 11244 3188 11296 3194
rect 11244 3130 11296 3136
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 10968 2916 11020 2922
rect 11020 2876 11100 2904
rect 10968 2858 11020 2864
rect 11072 2650 11100 2876
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11624 480 11652 9318
rect 12728 9042 12756 9658
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12544 8090 12572 8298
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 11716 7002 11744 7278
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 12438 6216 12494 6225
rect 12438 6151 12494 6160
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11716 5030 11744 5714
rect 12162 5672 12218 5681
rect 12162 5607 12218 5616
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11716 2825 11744 4966
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11900 3942 11928 4082
rect 12176 4078 12204 5607
rect 12452 5370 12480 6151
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12256 5024 12308 5030
rect 12544 5001 12572 7278
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12636 5273 12664 6054
rect 12622 5264 12678 5273
rect 12622 5199 12678 5208
rect 12256 4966 12308 4972
rect 12530 4992 12586 5001
rect 12268 4758 12296 4966
rect 12530 4927 12586 4936
rect 12256 4752 12308 4758
rect 12256 4694 12308 4700
rect 12348 4480 12400 4486
rect 12820 4434 12848 9318
rect 12912 8956 12940 11494
rect 13188 11121 13216 12038
rect 13740 11694 13768 12174
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13174 11112 13230 11121
rect 13174 11047 13230 11056
rect 13452 10668 13504 10674
rect 13452 10610 13504 10616
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 13004 9110 13032 9454
rect 13084 9444 13136 9450
rect 13084 9386 13136 9392
rect 13096 9178 13124 9386
rect 13464 9178 13492 10610
rect 13832 10554 13860 11494
rect 13740 10526 13860 10554
rect 13740 10198 13768 10526
rect 13820 10464 13872 10470
rect 13924 10452 13952 13670
rect 14002 13631 14058 13640
rect 13872 10424 13952 10452
rect 13820 10406 13872 10412
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13740 10010 13768 10134
rect 13648 9982 13768 10010
rect 13542 9752 13598 9761
rect 13542 9687 13598 9696
rect 13556 9178 13584 9687
rect 13648 9382 13676 9982
rect 13820 9920 13872 9926
rect 13740 9868 13820 9874
rect 13740 9862 13872 9868
rect 13740 9846 13860 9862
rect 13740 9586 13768 9846
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 12992 9104 13044 9110
rect 12992 9046 13044 9052
rect 12912 8928 13124 8956
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12912 4593 12940 7142
rect 13096 5250 13124 8928
rect 13268 8356 13320 8362
rect 13268 8298 13320 8304
rect 13004 5222 13124 5250
rect 12898 4584 12954 4593
rect 12898 4519 12954 4528
rect 12348 4422 12400 4428
rect 12360 4146 12388 4422
rect 12636 4406 12848 4434
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12164 4072 12216 4078
rect 12164 4014 12216 4020
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11900 3670 11928 3878
rect 11888 3664 11940 3670
rect 11888 3606 11940 3612
rect 11900 3194 11928 3606
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 12360 3058 12388 3470
rect 12636 3369 12664 4406
rect 12912 3942 12940 4422
rect 12900 3936 12952 3942
rect 12898 3904 12900 3913
rect 12952 3904 12954 3913
rect 12898 3839 12954 3848
rect 13004 3618 13032 5222
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 13096 5030 13124 5102
rect 13084 5024 13136 5030
rect 13082 4992 13084 5001
rect 13136 4992 13138 5001
rect 13082 4927 13138 4936
rect 12728 3590 13032 3618
rect 12622 3360 12678 3369
rect 12622 3295 12678 3304
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 11702 2816 11758 2825
rect 11702 2751 11758 2760
rect 12360 2650 12388 2994
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 12636 2553 12664 3295
rect 12622 2544 12678 2553
rect 12622 2479 12678 2488
rect 12728 480 12756 3590
rect 13280 2990 13308 8298
rect 13464 8090 13492 9114
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13556 7954 13584 9114
rect 13648 8974 13676 9318
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13648 8634 13676 8910
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 13820 8560 13872 8566
rect 13818 8528 13820 8537
rect 13872 8528 13874 8537
rect 13818 8463 13874 8472
rect 13924 8378 13952 10424
rect 14016 8430 14044 13631
rect 14108 13530 14136 14826
rect 14372 14068 14424 14074
rect 14424 14028 14504 14056
rect 14372 14010 14424 14016
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 14476 10606 14504 14028
rect 14568 13705 14596 14962
rect 15488 14822 15516 17070
rect 15764 16794 15792 17070
rect 16316 17066 16344 17614
rect 16304 17060 16356 17066
rect 16304 17002 16356 17008
rect 16580 17060 16632 17066
rect 16580 17002 16632 17008
rect 16316 16794 16344 17002
rect 16592 16946 16620 17002
rect 16500 16918 16620 16946
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 15764 16250 15792 16730
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 16132 16182 16160 16526
rect 16500 16250 16528 16918
rect 16684 16590 16712 18278
rect 16868 18222 16896 18362
rect 16960 18290 16988 19654
rect 17972 19310 18000 19858
rect 18340 19854 18368 20402
rect 20088 20398 20116 20742
rect 20076 20392 20128 20398
rect 20076 20334 20128 20340
rect 20534 20360 20590 20369
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 20088 20058 20116 20334
rect 20534 20295 20590 20304
rect 20076 20052 20128 20058
rect 20076 19994 20128 20000
rect 18052 19848 18104 19854
rect 18052 19790 18104 19796
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 18064 19378 18092 19790
rect 18328 19712 18380 19718
rect 18328 19654 18380 19660
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 18052 19372 18104 19378
rect 18052 19314 18104 19320
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 17972 18970 18000 19246
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 18064 18902 18092 19314
rect 18340 19242 18368 19654
rect 18328 19236 18380 19242
rect 18328 19178 18380 19184
rect 18052 18896 18104 18902
rect 18052 18838 18104 18844
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 16856 18216 16908 18222
rect 16856 18158 16908 18164
rect 17512 18154 17540 18566
rect 18064 18426 18092 18838
rect 18340 18426 18368 19178
rect 19352 18698 19380 19654
rect 19432 19168 19484 19174
rect 19432 19110 19484 19116
rect 19444 18970 19472 19110
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 20088 18834 20116 19994
rect 20548 19174 20576 20295
rect 20916 20058 20944 21422
rect 21364 21344 21416 21350
rect 21364 21286 21416 21292
rect 20996 20528 21048 20534
rect 20996 20470 21048 20476
rect 20904 20052 20956 20058
rect 20904 19994 20956 20000
rect 20902 19952 20958 19961
rect 20902 19887 20958 19896
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20640 19258 20668 19654
rect 20720 19304 20772 19310
rect 20640 19252 20720 19258
rect 20640 19246 20772 19252
rect 20640 19230 20760 19246
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 20916 18902 20944 19887
rect 21008 19394 21036 20470
rect 21376 20233 21404 21286
rect 21836 21078 21864 21626
rect 21928 21554 21956 22034
rect 21916 21548 21968 21554
rect 21916 21490 21968 21496
rect 21928 21146 21956 21490
rect 21916 21140 21968 21146
rect 21916 21082 21968 21088
rect 21824 21072 21876 21078
rect 21824 21014 21876 21020
rect 21548 21004 21600 21010
rect 21548 20946 21600 20952
rect 21560 20602 21588 20946
rect 21548 20596 21600 20602
rect 21548 20538 21600 20544
rect 21560 20262 21588 20538
rect 21836 20534 21864 21014
rect 21824 20528 21876 20534
rect 21824 20470 21876 20476
rect 22468 20392 22520 20398
rect 22466 20360 22468 20369
rect 22520 20360 22522 20369
rect 22466 20295 22522 20304
rect 21548 20256 21600 20262
rect 21362 20224 21418 20233
rect 21548 20198 21600 20204
rect 22652 20256 22704 20262
rect 22652 20198 22704 20204
rect 21362 20159 21418 20168
rect 21270 20088 21326 20097
rect 21270 20023 21272 20032
rect 21324 20023 21326 20032
rect 21272 19994 21324 20000
rect 21088 19848 21140 19854
rect 21088 19790 21140 19796
rect 21100 19514 21128 19790
rect 21180 19712 21232 19718
rect 21180 19654 21232 19660
rect 21088 19508 21140 19514
rect 21088 19450 21140 19456
rect 21008 19366 21128 19394
rect 21192 19378 21220 19654
rect 21284 19514 21312 19994
rect 21560 19854 21588 20198
rect 22664 20058 22692 20198
rect 22652 20052 22704 20058
rect 22652 19994 22704 20000
rect 22468 19916 22520 19922
rect 22468 19858 22520 19864
rect 21548 19848 21600 19854
rect 21548 19790 21600 19796
rect 21916 19848 21968 19854
rect 21916 19790 21968 19796
rect 21928 19514 21956 19790
rect 21272 19508 21324 19514
rect 21272 19450 21324 19456
rect 21916 19508 21968 19514
rect 21916 19450 21968 19456
rect 20994 19272 21050 19281
rect 20994 19207 20996 19216
rect 21048 19207 21050 19216
rect 20996 19178 21048 19184
rect 21008 18970 21036 19178
rect 20996 18964 21048 18970
rect 20996 18906 21048 18912
rect 20904 18896 20956 18902
rect 20904 18838 20956 18844
rect 19432 18828 19484 18834
rect 19432 18770 19484 18776
rect 20076 18828 20128 18834
rect 20076 18770 20128 18776
rect 19340 18692 19392 18698
rect 19340 18634 19392 18640
rect 18052 18420 18104 18426
rect 18052 18362 18104 18368
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 17868 18284 17920 18290
rect 17868 18226 17920 18232
rect 17500 18148 17552 18154
rect 17500 18090 17552 18096
rect 17880 17898 17908 18226
rect 17880 17882 18000 17898
rect 17880 17876 18012 17882
rect 17880 17870 17960 17876
rect 17960 17818 18012 17824
rect 16764 17740 16816 17746
rect 16764 17682 16816 17688
rect 16776 16998 16804 17682
rect 16764 16992 16816 16998
rect 16764 16934 16816 16940
rect 16856 16788 16908 16794
rect 16856 16730 16908 16736
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16488 16244 16540 16250
rect 16488 16186 16540 16192
rect 16120 16176 16172 16182
rect 16120 16118 16172 16124
rect 16132 15706 16160 16118
rect 16776 15910 16804 16594
rect 16868 16590 16896 16730
rect 17038 16688 17094 16697
rect 17038 16623 17094 16632
rect 16856 16584 16908 16590
rect 16856 16526 16908 16532
rect 17052 16454 17080 16623
rect 17040 16448 17092 16454
rect 17040 16390 17092 16396
rect 17052 16114 17080 16390
rect 18064 16250 18092 18362
rect 19340 18148 19392 18154
rect 19340 18090 19392 18096
rect 19352 17882 19380 18090
rect 19444 17882 19472 18770
rect 19708 18760 19760 18766
rect 19708 18702 19760 18708
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 19720 18154 19748 18702
rect 19890 18184 19946 18193
rect 19708 18148 19760 18154
rect 19890 18119 19946 18128
rect 19708 18090 19760 18096
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 18696 17876 18748 17882
rect 18696 17818 18748 17824
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18432 16998 18460 17478
rect 18708 17202 18736 17818
rect 18972 17740 19024 17746
rect 18972 17682 19024 17688
rect 18984 17270 19012 17682
rect 19444 17338 19472 17818
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 18972 17264 19024 17270
rect 18972 17206 19024 17212
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 19904 17134 19932 18119
rect 19996 17678 20024 18702
rect 20088 18426 20116 18770
rect 20916 18426 20944 18838
rect 21008 18426 21036 18906
rect 20076 18420 20128 18426
rect 20076 18362 20128 18368
rect 20904 18420 20956 18426
rect 20904 18362 20956 18368
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 20720 17740 20772 17746
rect 20720 17682 20772 17688
rect 19984 17672 20036 17678
rect 19982 17640 19984 17649
rect 20036 17640 20038 17649
rect 19982 17575 20038 17584
rect 19892 17128 19944 17134
rect 19892 17070 19944 17076
rect 20732 16998 20760 17682
rect 18236 16992 18288 16998
rect 18420 16992 18472 16998
rect 18236 16934 18288 16940
rect 18418 16960 18420 16969
rect 20720 16992 20772 16998
rect 18472 16960 18474 16969
rect 18248 16794 18276 16934
rect 20720 16934 20772 16940
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 18418 16895 18474 16904
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 18236 16788 18288 16794
rect 18236 16730 18288 16736
rect 20732 16726 20760 16934
rect 21008 16794 21036 16934
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 20720 16720 20772 16726
rect 20720 16662 20772 16668
rect 20810 16688 20866 16697
rect 18788 16448 18840 16454
rect 18788 16390 18840 16396
rect 18052 16244 18104 16250
rect 18052 16186 18104 16192
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 18800 16046 18828 16390
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 17500 15972 17552 15978
rect 17500 15914 17552 15920
rect 16764 15904 16816 15910
rect 16764 15846 16816 15852
rect 17224 15904 17276 15910
rect 17224 15846 17276 15852
rect 16776 15706 16804 15846
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 16764 15700 16816 15706
rect 16764 15642 16816 15648
rect 17236 15502 17264 15846
rect 17512 15745 17540 15914
rect 17498 15736 17554 15745
rect 17498 15671 17554 15680
rect 17512 15638 17540 15671
rect 17500 15632 17552 15638
rect 17500 15574 17552 15580
rect 17224 15496 17276 15502
rect 17224 15438 17276 15444
rect 16118 15192 16174 15201
rect 16118 15127 16174 15136
rect 15108 14816 15160 14822
rect 15476 14816 15528 14822
rect 15160 14764 15332 14770
rect 15108 14758 15332 14764
rect 15476 14758 15528 14764
rect 15120 14742 15332 14758
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14936 13938 14964 14554
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14554 13696 14610 13705
rect 14554 13631 14610 13640
rect 14660 13190 14688 13806
rect 15200 13388 15252 13394
rect 15028 13348 15200 13376
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14660 10674 14688 13126
rect 15028 12102 15056 13348
rect 15200 13330 15252 13336
rect 15200 13252 15252 13258
rect 15200 13194 15252 13200
rect 15212 12782 15240 13194
rect 15304 12986 15332 14742
rect 15488 13190 15516 14758
rect 16132 13802 16160 15127
rect 17236 14822 17264 15438
rect 17512 15162 17540 15574
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 18800 14929 18828 15982
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 19444 15745 19472 15846
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19430 15736 19486 15745
rect 19580 15728 19876 15748
rect 20732 15706 20760 16662
rect 20810 16623 20812 16632
rect 20864 16623 20866 16632
rect 20812 16594 20864 16600
rect 21100 16590 21128 19366
rect 21180 19372 21232 19378
rect 21180 19314 21232 19320
rect 22376 19168 22428 19174
rect 22376 19110 22428 19116
rect 22388 19009 22416 19110
rect 22374 19000 22430 19009
rect 22480 18970 22508 19858
rect 22374 18935 22430 18944
rect 22468 18964 22520 18970
rect 22468 18906 22520 18912
rect 21824 18692 21876 18698
rect 21824 18634 21876 18640
rect 21836 18290 21864 18634
rect 22008 18624 22060 18630
rect 22008 18566 22060 18572
rect 22020 18290 22048 18566
rect 22756 18465 22784 35119
rect 29932 34649 29960 39520
rect 35714 39400 35770 39409
rect 35714 39335 35770 39344
rect 35622 38176 35678 38185
rect 35622 38111 35678 38120
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 35636 36378 35664 38111
rect 35624 36372 35676 36378
rect 35624 36314 35676 36320
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 35728 35834 35756 39335
rect 37554 36952 37610 36961
rect 37554 36887 37610 36896
rect 35808 36236 35860 36242
rect 35808 36178 35860 36184
rect 35716 35828 35768 35834
rect 35716 35770 35768 35776
rect 33966 35728 34022 35737
rect 33966 35663 34022 35672
rect 33048 35488 33100 35494
rect 33048 35430 33100 35436
rect 33416 35488 33468 35494
rect 33416 35430 33468 35436
rect 33060 35222 33088 35430
rect 33428 35290 33456 35430
rect 33416 35284 33468 35290
rect 33416 35226 33468 35232
rect 33048 35216 33100 35222
rect 33048 35158 33100 35164
rect 32128 35080 32180 35086
rect 32128 35022 32180 35028
rect 28354 34640 28410 34649
rect 28354 34575 28410 34584
rect 29918 34640 29974 34649
rect 29918 34575 29974 34584
rect 24860 31136 24912 31142
rect 24860 31078 24912 31084
rect 27528 31136 27580 31142
rect 27528 31078 27580 31084
rect 24872 30938 24900 31078
rect 24860 30932 24912 30938
rect 24860 30874 24912 30880
rect 25228 30932 25280 30938
rect 25228 30874 25280 30880
rect 24860 30728 24912 30734
rect 24860 30670 24912 30676
rect 24872 30326 24900 30670
rect 24952 30660 25004 30666
rect 24952 30602 25004 30608
rect 24216 30320 24268 30326
rect 24216 30262 24268 30268
rect 24860 30320 24912 30326
rect 24860 30262 24912 30268
rect 23940 30048 23992 30054
rect 23940 29990 23992 29996
rect 23952 29646 23980 29990
rect 24228 29782 24256 30262
rect 24216 29776 24268 29782
rect 24216 29718 24268 29724
rect 23940 29640 23992 29646
rect 23940 29582 23992 29588
rect 23952 29102 23980 29582
rect 24216 29504 24268 29510
rect 24216 29446 24268 29452
rect 24228 29102 24256 29446
rect 24872 29306 24900 30262
rect 24860 29300 24912 29306
rect 24860 29242 24912 29248
rect 24964 29186 24992 30602
rect 25240 30190 25268 30874
rect 26884 30728 26936 30734
rect 26884 30670 26936 30676
rect 26240 30592 26292 30598
rect 26240 30534 26292 30540
rect 25228 30184 25280 30190
rect 25228 30126 25280 30132
rect 25240 29850 25268 30126
rect 25228 29844 25280 29850
rect 25228 29786 25280 29792
rect 24872 29158 24992 29186
rect 26252 29170 26280 30534
rect 26896 30326 26924 30670
rect 26884 30320 26936 30326
rect 26884 30262 26936 30268
rect 26332 30048 26384 30054
rect 26332 29990 26384 29996
rect 26344 29782 26372 29990
rect 26896 29782 26924 30262
rect 27540 30258 27568 31078
rect 27620 30796 27672 30802
rect 27620 30738 27672 30744
rect 27528 30252 27580 30258
rect 27528 30194 27580 30200
rect 27632 30190 27660 30738
rect 27896 30388 27948 30394
rect 27896 30330 27948 30336
rect 27620 30184 27672 30190
rect 27620 30126 27672 30132
rect 27436 30048 27488 30054
rect 27436 29990 27488 29996
rect 26332 29776 26384 29782
rect 26332 29718 26384 29724
rect 26884 29776 26936 29782
rect 26884 29718 26936 29724
rect 26344 29306 26372 29718
rect 26516 29708 26568 29714
rect 26516 29650 26568 29656
rect 26332 29300 26384 29306
rect 26332 29242 26384 29248
rect 26240 29164 26292 29170
rect 23940 29096 23992 29102
rect 23940 29038 23992 29044
rect 24216 29096 24268 29102
rect 24216 29038 24268 29044
rect 23572 28960 23624 28966
rect 23572 28902 23624 28908
rect 23480 28620 23532 28626
rect 23480 28562 23532 28568
rect 23492 28218 23520 28562
rect 23584 28422 23612 28902
rect 24228 28762 24256 29038
rect 24216 28756 24268 28762
rect 24216 28698 24268 28704
rect 23572 28416 23624 28422
rect 23572 28358 23624 28364
rect 23480 28212 23532 28218
rect 23480 28154 23532 28160
rect 23584 28014 23612 28358
rect 24872 28150 24900 29158
rect 26240 29106 26292 29112
rect 26332 29096 26384 29102
rect 26332 29038 26384 29044
rect 26344 28762 26372 29038
rect 26528 29034 26556 29650
rect 27448 29102 27476 29990
rect 27632 29850 27660 30126
rect 27620 29844 27672 29850
rect 27620 29786 27672 29792
rect 27528 29504 27580 29510
rect 27528 29446 27580 29452
rect 27540 29170 27568 29446
rect 27620 29300 27672 29306
rect 27620 29242 27672 29248
rect 27528 29164 27580 29170
rect 27528 29106 27580 29112
rect 27436 29096 27488 29102
rect 27436 29038 27488 29044
rect 26516 29028 26568 29034
rect 26516 28970 26568 28976
rect 26332 28756 26384 28762
rect 26332 28698 26384 28704
rect 27068 28688 27120 28694
rect 27068 28630 27120 28636
rect 26976 28552 27028 28558
rect 26976 28494 27028 28500
rect 26332 28416 26384 28422
rect 26332 28358 26384 28364
rect 24860 28144 24912 28150
rect 24860 28086 24912 28092
rect 23572 28008 23624 28014
rect 23572 27950 23624 27956
rect 23480 27940 23532 27946
rect 23480 27882 23532 27888
rect 23492 27130 23520 27882
rect 23584 27878 23612 27950
rect 24216 27940 24268 27946
rect 24216 27882 24268 27888
rect 23572 27872 23624 27878
rect 23572 27814 23624 27820
rect 23584 27334 23612 27814
rect 24228 27674 24256 27882
rect 24216 27668 24268 27674
rect 24216 27610 24268 27616
rect 24872 27606 24900 28086
rect 26148 27872 26200 27878
rect 26200 27820 26280 27826
rect 26148 27814 26280 27820
rect 26160 27798 26280 27814
rect 24860 27600 24912 27606
rect 24860 27542 24912 27548
rect 24308 27464 24360 27470
rect 24308 27406 24360 27412
rect 23572 27328 23624 27334
rect 23572 27270 23624 27276
rect 23848 27328 23900 27334
rect 23848 27270 23900 27276
rect 23480 27124 23532 27130
rect 23480 27066 23532 27072
rect 23492 26586 23520 27066
rect 23584 26926 23612 27270
rect 23860 27169 23888 27270
rect 23846 27160 23902 27169
rect 23846 27095 23902 27104
rect 23572 26920 23624 26926
rect 23572 26862 23624 26868
rect 23584 26790 23612 26862
rect 24320 26858 24348 27406
rect 24308 26852 24360 26858
rect 24308 26794 24360 26800
rect 23572 26784 23624 26790
rect 23572 26726 23624 26732
rect 23480 26580 23532 26586
rect 23480 26522 23532 26528
rect 23584 26382 23612 26726
rect 24320 26586 24348 26794
rect 26252 26586 26280 27798
rect 26344 27538 26372 28358
rect 26988 28218 27016 28494
rect 27080 28218 27108 28630
rect 27160 28552 27212 28558
rect 27160 28494 27212 28500
rect 27540 28506 27568 29106
rect 27632 28626 27660 29242
rect 27804 28960 27856 28966
rect 27804 28902 27856 28908
rect 27620 28620 27672 28626
rect 27620 28562 27672 28568
rect 26976 28212 27028 28218
rect 26976 28154 27028 28160
rect 27068 28212 27120 28218
rect 27068 28154 27120 28160
rect 27172 28150 27200 28494
rect 27540 28478 27660 28506
rect 27632 28422 27660 28478
rect 27620 28416 27672 28422
rect 27620 28358 27672 28364
rect 27160 28144 27212 28150
rect 27160 28086 27212 28092
rect 26608 27872 26660 27878
rect 26608 27814 26660 27820
rect 26332 27532 26384 27538
rect 26332 27474 26384 27480
rect 24308 26580 24360 26586
rect 24308 26522 24360 26528
rect 26240 26580 26292 26586
rect 26240 26522 26292 26528
rect 26344 26518 26372 27474
rect 26424 27464 26476 27470
rect 26424 27406 26476 27412
rect 26436 27169 26464 27406
rect 26516 27328 26568 27334
rect 26514 27296 26516 27305
rect 26568 27296 26570 27305
rect 26514 27231 26570 27240
rect 26422 27160 26478 27169
rect 26620 27130 26648 27814
rect 27172 27554 27200 28086
rect 27632 28082 27660 28358
rect 27816 28218 27844 28902
rect 27804 28212 27856 28218
rect 27804 28154 27856 28160
rect 27620 28076 27672 28082
rect 27620 28018 27672 28024
rect 27632 27962 27660 28018
rect 27080 27526 27200 27554
rect 27540 27934 27660 27962
rect 26422 27095 26424 27104
rect 26476 27095 26478 27104
rect 26608 27124 26660 27130
rect 26424 27066 26476 27072
rect 26608 27066 26660 27072
rect 26608 26784 26660 26790
rect 26606 26752 26608 26761
rect 26660 26752 26662 26761
rect 26606 26687 26662 26696
rect 23756 26512 23808 26518
rect 23756 26454 23808 26460
rect 26332 26512 26384 26518
rect 26332 26454 26384 26460
rect 23572 26376 23624 26382
rect 23572 26318 23624 26324
rect 23584 25838 23612 26318
rect 23572 25832 23624 25838
rect 23572 25774 23624 25780
rect 23768 25770 23796 26454
rect 26884 26444 26936 26450
rect 26884 26386 26936 26392
rect 26896 26042 26924 26386
rect 27080 26314 27108 27526
rect 27540 27470 27568 27934
rect 27160 27464 27212 27470
rect 27160 27406 27212 27412
rect 27528 27464 27580 27470
rect 27528 27406 27580 27412
rect 27172 26382 27200 27406
rect 27804 26988 27856 26994
rect 27804 26930 27856 26936
rect 27712 26784 27764 26790
rect 27712 26726 27764 26732
rect 27528 26444 27580 26450
rect 27528 26386 27580 26392
rect 27160 26376 27212 26382
rect 27158 26344 27160 26353
rect 27212 26344 27214 26353
rect 27068 26308 27120 26314
rect 27158 26279 27214 26288
rect 27068 26250 27120 26256
rect 26332 26036 26384 26042
rect 26332 25978 26384 25984
rect 26884 26036 26936 26042
rect 26884 25978 26936 25984
rect 23940 25832 23992 25838
rect 23940 25774 23992 25780
rect 23756 25764 23808 25770
rect 23756 25706 23808 25712
rect 23952 25702 23980 25774
rect 24308 25764 24360 25770
rect 24308 25706 24360 25712
rect 23940 25696 23992 25702
rect 23940 25638 23992 25644
rect 23952 25294 23980 25638
rect 24216 25356 24268 25362
rect 24216 25298 24268 25304
rect 23940 25288 23992 25294
rect 23940 25230 23992 25236
rect 23952 24614 23980 25230
rect 23940 24608 23992 24614
rect 23940 24550 23992 24556
rect 23952 22574 23980 24550
rect 24228 24410 24256 25298
rect 24320 25158 24348 25706
rect 26344 25498 26372 25978
rect 26792 25968 26844 25974
rect 26792 25910 26844 25916
rect 26332 25492 26384 25498
rect 26332 25434 26384 25440
rect 26804 25430 26832 25910
rect 27080 25906 27108 26250
rect 27540 26194 27568 26386
rect 27540 26166 27660 26194
rect 27068 25900 27120 25906
rect 27068 25842 27120 25848
rect 26884 25696 26936 25702
rect 26884 25638 26936 25644
rect 26896 25498 26924 25638
rect 26884 25492 26936 25498
rect 26884 25434 26936 25440
rect 26792 25424 26844 25430
rect 26792 25366 26844 25372
rect 25228 25356 25280 25362
rect 25228 25298 25280 25304
rect 24308 25152 24360 25158
rect 24308 25094 24360 25100
rect 24952 25152 25004 25158
rect 24952 25094 25004 25100
rect 24582 24848 24638 24857
rect 24582 24783 24638 24792
rect 24216 24404 24268 24410
rect 24216 24346 24268 24352
rect 24596 24138 24624 24783
rect 24676 24676 24728 24682
rect 24676 24618 24728 24624
rect 24688 24342 24716 24618
rect 24676 24336 24728 24342
rect 24676 24278 24728 24284
rect 24584 24132 24636 24138
rect 24584 24074 24636 24080
rect 24688 23633 24716 24278
rect 24964 24274 24992 25094
rect 25044 24608 25096 24614
rect 25044 24550 25096 24556
rect 25056 24410 25084 24550
rect 25044 24404 25096 24410
rect 25044 24346 25096 24352
rect 24952 24268 25004 24274
rect 24952 24210 25004 24216
rect 24964 23798 24992 24210
rect 25056 23866 25084 24346
rect 25240 24206 25268 25298
rect 26516 25288 26568 25294
rect 26516 25230 26568 25236
rect 26528 24954 26556 25230
rect 26804 24954 26832 25366
rect 27080 25362 27108 25842
rect 27632 25702 27660 26166
rect 27724 25838 27752 26726
rect 27816 26382 27844 26930
rect 27804 26376 27856 26382
rect 27804 26318 27856 26324
rect 27712 25832 27764 25838
rect 27712 25774 27764 25780
rect 27620 25696 27672 25702
rect 27620 25638 27672 25644
rect 27068 25356 27120 25362
rect 27068 25298 27120 25304
rect 26516 24948 26568 24954
rect 26516 24890 26568 24896
rect 26792 24948 26844 24954
rect 26792 24890 26844 24896
rect 26528 24206 26556 24890
rect 27632 24857 27660 25638
rect 27618 24848 27674 24857
rect 27618 24783 27674 24792
rect 25228 24200 25280 24206
rect 25228 24142 25280 24148
rect 26516 24200 26568 24206
rect 26516 24142 26568 24148
rect 27252 24200 27304 24206
rect 27252 24142 27304 24148
rect 25240 23866 25268 24142
rect 25044 23860 25096 23866
rect 25044 23802 25096 23808
rect 25228 23860 25280 23866
rect 25228 23802 25280 23808
rect 24952 23792 25004 23798
rect 24952 23734 25004 23740
rect 24674 23624 24730 23633
rect 24674 23559 24730 23568
rect 24032 22976 24084 22982
rect 24032 22918 24084 22924
rect 26792 22976 26844 22982
rect 26792 22918 26844 22924
rect 24044 22574 24072 22918
rect 26700 22704 26752 22710
rect 26700 22646 26752 22652
rect 26332 22636 26384 22642
rect 26332 22578 26384 22584
rect 23940 22568 23992 22574
rect 23940 22510 23992 22516
rect 24032 22568 24084 22574
rect 24032 22510 24084 22516
rect 23952 22098 23980 22510
rect 23940 22092 23992 22098
rect 23940 22034 23992 22040
rect 23756 22024 23808 22030
rect 23756 21966 23808 21972
rect 23204 21888 23256 21894
rect 23204 21830 23256 21836
rect 23216 21078 23244 21830
rect 23204 21072 23256 21078
rect 23204 21014 23256 21020
rect 23480 21072 23532 21078
rect 23480 21014 23532 21020
rect 23492 20058 23520 21014
rect 23664 20392 23716 20398
rect 23664 20334 23716 20340
rect 23480 20052 23532 20058
rect 23480 19994 23532 20000
rect 23112 19168 23164 19174
rect 23112 19110 23164 19116
rect 23124 18970 23152 19110
rect 23492 18970 23520 19994
rect 23676 19281 23704 20334
rect 23768 20058 23796 21966
rect 23952 21010 23980 22034
rect 24044 21962 24072 22510
rect 25320 22432 25372 22438
rect 25320 22374 25372 22380
rect 26240 22432 26292 22438
rect 26240 22374 26292 22380
rect 24676 22092 24728 22098
rect 24676 22034 24728 22040
rect 24032 21956 24084 21962
rect 24032 21898 24084 21904
rect 24044 21690 24072 21898
rect 24308 21888 24360 21894
rect 24308 21830 24360 21836
rect 24032 21684 24084 21690
rect 24032 21626 24084 21632
rect 24214 21448 24270 21457
rect 24214 21383 24270 21392
rect 23940 21004 23992 21010
rect 23940 20946 23992 20952
rect 23952 20602 23980 20946
rect 23940 20596 23992 20602
rect 23940 20538 23992 20544
rect 23848 20256 23900 20262
rect 23848 20198 23900 20204
rect 24122 20224 24178 20233
rect 23860 20097 23888 20198
rect 24122 20159 24178 20168
rect 23846 20088 23902 20097
rect 23756 20052 23808 20058
rect 24136 20058 24164 20159
rect 24228 20058 24256 21383
rect 24320 21185 24348 21830
rect 24688 21690 24716 22034
rect 24768 21888 24820 21894
rect 24768 21830 24820 21836
rect 24676 21684 24728 21690
rect 24676 21626 24728 21632
rect 24306 21176 24362 21185
rect 24780 21146 24808 21830
rect 25044 21548 25096 21554
rect 25044 21490 25096 21496
rect 24306 21111 24362 21120
rect 24768 21140 24820 21146
rect 24768 21082 24820 21088
rect 25056 20806 25084 21490
rect 25332 21146 25360 22374
rect 26252 22250 26280 22374
rect 26160 22222 26280 22250
rect 25596 21888 25648 21894
rect 25596 21830 25648 21836
rect 25608 21486 25636 21830
rect 26056 21684 26108 21690
rect 26056 21626 26108 21632
rect 25596 21480 25648 21486
rect 25594 21448 25596 21457
rect 25648 21448 25650 21457
rect 25594 21383 25650 21392
rect 25320 21140 25372 21146
rect 25320 21082 25372 21088
rect 25044 20800 25096 20806
rect 25044 20742 25096 20748
rect 23846 20023 23902 20032
rect 24124 20052 24176 20058
rect 23756 19994 23808 20000
rect 24124 19994 24176 20000
rect 24216 20052 24268 20058
rect 24216 19994 24268 20000
rect 24136 19514 24164 19994
rect 24124 19508 24176 19514
rect 24124 19450 24176 19456
rect 24228 19378 24256 19994
rect 24216 19372 24268 19378
rect 24216 19314 24268 19320
rect 25056 19310 25084 20742
rect 25332 20398 25360 21082
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25320 20392 25372 20398
rect 25320 20334 25372 20340
rect 25332 20058 25360 20334
rect 25320 20052 25372 20058
rect 25320 19994 25372 20000
rect 25332 19378 25360 19994
rect 25320 19372 25372 19378
rect 25320 19314 25372 19320
rect 25044 19304 25096 19310
rect 23662 19272 23718 19281
rect 25044 19246 25096 19252
rect 23662 19207 23718 19216
rect 25056 19009 25084 19246
rect 25042 19000 25098 19009
rect 23112 18964 23164 18970
rect 23112 18906 23164 18912
rect 23480 18964 23532 18970
rect 25042 18935 25044 18944
rect 23480 18906 23532 18912
rect 25096 18935 25098 18944
rect 25044 18906 25096 18912
rect 22836 18828 22888 18834
rect 22836 18770 22888 18776
rect 22742 18456 22798 18465
rect 22742 18391 22798 18400
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 21548 17808 21600 17814
rect 21548 17750 21600 17756
rect 21456 17536 21508 17542
rect 21456 17478 21508 17484
rect 21468 17202 21496 17478
rect 21560 17202 21588 17750
rect 21732 17672 21784 17678
rect 21732 17614 21784 17620
rect 21916 17672 21968 17678
rect 22020 17649 22048 18226
rect 22848 18086 22876 18770
rect 22468 18080 22520 18086
rect 22468 18022 22520 18028
rect 22836 18080 22888 18086
rect 22836 18022 22888 18028
rect 23388 18080 23440 18086
rect 24676 18080 24728 18086
rect 23440 18028 23520 18034
rect 23388 18022 23520 18028
rect 24676 18022 24728 18028
rect 22480 17882 22508 18022
rect 23400 18006 23520 18022
rect 22468 17876 22520 17882
rect 22468 17818 22520 17824
rect 22836 17740 22888 17746
rect 22836 17682 22888 17688
rect 21916 17614 21968 17620
rect 22006 17640 22062 17649
rect 21744 17338 21772 17614
rect 21732 17332 21784 17338
rect 21732 17274 21784 17280
rect 21456 17196 21508 17202
rect 21456 17138 21508 17144
rect 21548 17196 21600 17202
rect 21548 17138 21600 17144
rect 21272 16992 21324 16998
rect 21272 16934 21324 16940
rect 21088 16584 21140 16590
rect 21088 16526 21140 16532
rect 21100 16250 21128 16526
rect 21088 16244 21140 16250
rect 21088 16186 21140 16192
rect 19430 15671 19486 15680
rect 20720 15700 20772 15706
rect 20720 15642 20772 15648
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20732 15450 20760 15506
rect 21100 15502 21128 16186
rect 20640 15422 20760 15450
rect 21088 15496 21140 15502
rect 21088 15438 21140 15444
rect 20640 15162 20668 15422
rect 21100 15162 21128 15438
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 21088 15156 21140 15162
rect 21088 15098 21140 15104
rect 18786 14920 18842 14929
rect 18786 14855 18842 14864
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 21100 14618 21128 15098
rect 21284 14618 21312 16934
rect 21560 16833 21588 17138
rect 21546 16824 21602 16833
rect 21546 16759 21602 16768
rect 21928 16697 21956 17614
rect 22006 17575 22062 17584
rect 22192 17332 22244 17338
rect 22192 17274 22244 17280
rect 21914 16688 21970 16697
rect 21914 16623 21916 16632
rect 21968 16623 21970 16632
rect 21916 16594 21968 16600
rect 21928 16563 21956 16594
rect 22100 16448 22152 16454
rect 22100 16390 22152 16396
rect 21638 14920 21694 14929
rect 21638 14855 21694 14864
rect 21732 14884 21784 14890
rect 21652 14822 21680 14855
rect 21732 14826 21784 14832
rect 21640 14816 21692 14822
rect 21640 14758 21692 14764
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 21272 14612 21324 14618
rect 21272 14554 21324 14560
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 18604 13864 18656 13870
rect 18604 13806 18656 13812
rect 16120 13796 16172 13802
rect 16120 13738 16172 13744
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 16132 12782 16160 13738
rect 16670 13696 16726 13705
rect 16670 13631 16726 13640
rect 16684 13530 16712 13631
rect 16672 13524 16724 13530
rect 16672 13466 16724 13472
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 16210 13152 16266 13161
rect 16210 13087 16266 13096
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16132 12374 16160 12718
rect 16224 12646 16252 13087
rect 16316 12850 16344 13330
rect 17960 13320 18012 13326
rect 17880 13268 17960 13274
rect 17880 13262 18012 13268
rect 17880 13246 18000 13262
rect 16304 12844 16356 12850
rect 16304 12786 16356 12792
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17788 12646 17816 12786
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 17776 12640 17828 12646
rect 17776 12582 17828 12588
rect 16224 12442 16252 12582
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 16120 12368 16172 12374
rect 16120 12310 16172 12316
rect 17132 12368 17184 12374
rect 17132 12310 17184 12316
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 15028 11354 15056 12038
rect 16776 11898 16804 12174
rect 17144 11898 17172 12310
rect 17788 12238 17816 12582
rect 17880 12442 17908 13246
rect 18236 12708 18288 12714
rect 18236 12650 18288 12656
rect 17868 12436 17920 12442
rect 17868 12378 17920 12384
rect 18248 12374 18276 12650
rect 18236 12368 18288 12374
rect 18236 12310 18288 12316
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 17512 11558 17540 12174
rect 17788 11558 17816 12174
rect 18248 12102 18276 12310
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 17512 11121 17540 11494
rect 17788 11218 17816 11494
rect 17776 11212 17828 11218
rect 17776 11154 17828 11160
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17498 11112 17554 11121
rect 17498 11047 17554 11056
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14476 9722 14504 10542
rect 14660 9926 14688 10610
rect 17788 10606 17816 11154
rect 17972 10826 18000 11154
rect 18616 11098 18644 13806
rect 19352 13802 19380 14214
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19340 13796 19392 13802
rect 19340 13738 19392 13744
rect 19156 13728 19208 13734
rect 19156 13670 19208 13676
rect 19168 13530 19196 13670
rect 19156 13524 19208 13530
rect 19156 13466 19208 13472
rect 19064 13320 19116 13326
rect 19064 13262 19116 13268
rect 19156 13320 19208 13326
rect 19156 13262 19208 13268
rect 19076 12918 19104 13262
rect 19064 12912 19116 12918
rect 19064 12854 19116 12860
rect 18696 12368 18748 12374
rect 18696 12310 18748 12316
rect 18708 11558 18736 12310
rect 19168 11801 19196 13262
rect 19248 13184 19300 13190
rect 19248 13126 19300 13132
rect 19154 11792 19210 11801
rect 19154 11727 19210 11736
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18708 11354 18736 11494
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 19156 11212 19208 11218
rect 19156 11154 19208 11160
rect 18694 11112 18750 11121
rect 18616 11070 18694 11098
rect 18694 11047 18750 11056
rect 17880 10810 18000 10826
rect 17868 10804 18000 10810
rect 17920 10798 18000 10804
rect 17868 10746 17920 10752
rect 17776 10600 17828 10606
rect 17776 10542 17828 10548
rect 16856 10532 16908 10538
rect 16856 10474 16908 10480
rect 18236 10532 18288 10538
rect 18236 10474 18288 10480
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 14648 9920 14700 9926
rect 14648 9862 14700 9868
rect 14464 9716 14516 9722
rect 14464 9658 14516 9664
rect 13832 8350 13952 8378
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 13728 8016 13780 8022
rect 13728 7958 13780 7964
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 13360 7268 13412 7274
rect 13360 7210 13412 7216
rect 13372 5642 13400 7210
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13464 6458 13492 6938
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13556 6390 13584 7890
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13544 6384 13596 6390
rect 13544 6326 13596 6332
rect 13556 5794 13584 6326
rect 13648 5914 13676 6734
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 13556 5778 13676 5794
rect 13556 5772 13688 5778
rect 13556 5766 13636 5772
rect 13360 5636 13412 5642
rect 13360 5578 13412 5584
rect 13556 5370 13584 5766
rect 13636 5714 13688 5720
rect 13544 5364 13596 5370
rect 13544 5306 13596 5312
rect 13740 5012 13768 7958
rect 13832 6118 13860 8350
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 14016 7002 14044 7822
rect 14004 6996 14056 7002
rect 14004 6938 14056 6944
rect 14188 6792 14240 6798
rect 14188 6734 14240 6740
rect 13912 6724 13964 6730
rect 13912 6666 13964 6672
rect 13924 6254 13952 6666
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 14200 5846 14228 6734
rect 14660 6662 14688 9862
rect 15580 9761 15608 10406
rect 16672 10124 16724 10130
rect 16672 10066 16724 10072
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 15566 9752 15622 9761
rect 15566 9687 15622 9696
rect 16316 9042 16344 9998
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16500 9382 16528 9862
rect 16684 9654 16712 10066
rect 16868 10062 16896 10474
rect 16856 10056 16908 10062
rect 16856 9998 16908 10004
rect 16868 9722 16896 9998
rect 18248 9926 18276 10474
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 17038 9616 17094 9625
rect 16396 9376 16448 9382
rect 16396 9318 16448 9324
rect 16488 9376 16540 9382
rect 16488 9318 16540 9324
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16316 8294 16344 8978
rect 16408 8430 16436 9318
rect 16592 8634 16620 9318
rect 16684 9194 16712 9590
rect 18248 9586 18276 9862
rect 18708 9586 18736 11047
rect 19168 10810 19196 11154
rect 19260 10826 19288 13126
rect 19352 12714 19380 13738
rect 19444 12986 19472 13806
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 21100 13394 21128 14554
rect 21652 14550 21680 14758
rect 21744 14618 21772 14826
rect 22112 14634 22140 16390
rect 22204 16250 22232 17274
rect 22848 16794 22876 17682
rect 23492 17338 23520 18006
rect 24124 17740 24176 17746
rect 24124 17682 24176 17688
rect 24032 17604 24084 17610
rect 24032 17546 24084 17552
rect 23480 17332 23532 17338
rect 23480 17274 23532 17280
rect 24044 17202 24072 17546
rect 24136 17542 24164 17682
rect 24688 17610 24716 18022
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 24676 17604 24728 17610
rect 24676 17546 24728 17552
rect 24124 17536 24176 17542
rect 24124 17478 24176 17484
rect 24032 17196 24084 17202
rect 24032 17138 24084 17144
rect 23480 17128 23532 17134
rect 23480 17070 23532 17076
rect 23492 16833 23520 17070
rect 23664 17060 23716 17066
rect 23664 17002 23716 17008
rect 23478 16824 23534 16833
rect 22836 16788 22888 16794
rect 23478 16759 23480 16768
rect 22836 16730 22888 16736
rect 23532 16759 23534 16768
rect 23480 16730 23532 16736
rect 22374 16688 22430 16697
rect 22374 16623 22430 16632
rect 22192 16244 22244 16250
rect 22192 16186 22244 16192
rect 22204 15570 22232 16186
rect 22284 15972 22336 15978
rect 22284 15914 22336 15920
rect 22192 15564 22244 15570
rect 22192 15506 22244 15512
rect 22296 14958 22324 15914
rect 22388 15094 22416 16623
rect 23492 16250 23520 16730
rect 23480 16244 23532 16250
rect 23480 16186 23532 16192
rect 23676 15162 23704 17002
rect 24136 16810 24164 17478
rect 24044 16782 24164 16810
rect 24044 16289 24072 16782
rect 24400 16720 24452 16726
rect 24400 16662 24452 16668
rect 24124 16652 24176 16658
rect 24124 16594 24176 16600
rect 24030 16280 24086 16289
rect 24030 16215 24086 16224
rect 23756 16040 23808 16046
rect 23754 16008 23756 16017
rect 23808 16008 23810 16017
rect 23754 15943 23810 15952
rect 24044 15570 24072 16215
rect 24032 15564 24084 15570
rect 24032 15506 24084 15512
rect 23664 15156 23716 15162
rect 23664 15098 23716 15104
rect 22376 15088 22428 15094
rect 22376 15030 22428 15036
rect 22284 14952 22336 14958
rect 22284 14894 22336 14900
rect 22020 14618 22140 14634
rect 21732 14612 21784 14618
rect 21732 14554 21784 14560
rect 22008 14612 22140 14618
rect 22060 14606 22140 14612
rect 22008 14554 22060 14560
rect 21640 14544 21692 14550
rect 21640 14486 21692 14492
rect 21652 14006 21680 14486
rect 21744 14074 21772 14554
rect 22388 14482 22416 15030
rect 24044 14618 24072 15506
rect 24136 15366 24164 16594
rect 24412 16250 24440 16662
rect 24400 16244 24452 16250
rect 24400 16186 24452 16192
rect 24412 15638 24440 16186
rect 24400 15632 24452 15638
rect 24400 15574 24452 15580
rect 24124 15360 24176 15366
rect 24124 15302 24176 15308
rect 24136 15026 24164 15302
rect 24412 15162 24440 15574
rect 24400 15156 24452 15162
rect 24400 15098 24452 15104
rect 24688 15094 24716 17546
rect 24780 17338 24808 17614
rect 24768 17332 24820 17338
rect 24768 17274 24820 17280
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 24768 16448 24820 16454
rect 24768 16390 24820 16396
rect 24676 15088 24728 15094
rect 24676 15030 24728 15036
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 24308 15020 24360 15026
rect 24308 14962 24360 14968
rect 24320 14618 24348 14962
rect 24780 14958 24808 16390
rect 25148 16046 25176 17274
rect 25424 17270 25452 20538
rect 26068 19310 26096 21626
rect 26160 20058 26188 22222
rect 26240 21888 26292 21894
rect 26240 21830 26292 21836
rect 26252 21554 26280 21830
rect 26240 21548 26292 21554
rect 26240 21490 26292 21496
rect 26252 21146 26280 21490
rect 26240 21140 26292 21146
rect 26240 21082 26292 21088
rect 26148 20052 26200 20058
rect 26148 19994 26200 20000
rect 26344 19514 26372 22578
rect 26422 22536 26478 22545
rect 26422 22471 26478 22480
rect 26436 22438 26464 22471
rect 26424 22432 26476 22438
rect 26424 22374 26476 22380
rect 26712 22386 26740 22646
rect 26804 22642 26832 22918
rect 26792 22636 26844 22642
rect 26792 22578 26844 22584
rect 26712 22358 26832 22386
rect 26804 22098 26832 22358
rect 26792 22092 26844 22098
rect 26792 22034 26844 22040
rect 26516 22024 26568 22030
rect 26516 21966 26568 21972
rect 26528 21418 26556 21966
rect 26698 21720 26754 21729
rect 26698 21655 26700 21664
rect 26752 21655 26754 21664
rect 26700 21626 26752 21632
rect 26804 21486 26832 22034
rect 26792 21480 26844 21486
rect 26792 21422 26844 21428
rect 26516 21412 26568 21418
rect 26516 21354 26568 21360
rect 26528 20534 26556 21354
rect 26804 20602 26832 21422
rect 27264 21418 27292 24142
rect 27908 21978 27936 30330
rect 28080 28620 28132 28626
rect 28080 28562 28132 28568
rect 27988 27872 28040 27878
rect 27988 27814 28040 27820
rect 28000 27674 28028 27814
rect 27988 27668 28040 27674
rect 27988 27610 28040 27616
rect 28092 27606 28120 28562
rect 28264 28416 28316 28422
rect 28264 28358 28316 28364
rect 28080 27600 28132 27606
rect 28080 27542 28132 27548
rect 28276 26586 28304 28358
rect 28264 26580 28316 26586
rect 28264 26522 28316 26528
rect 28276 26042 28304 26522
rect 28264 26036 28316 26042
rect 28264 25978 28316 25984
rect 28264 25696 28316 25702
rect 28264 25638 28316 25644
rect 28276 25498 28304 25638
rect 28264 25492 28316 25498
rect 28264 25434 28316 25440
rect 28080 24268 28132 24274
rect 28080 24210 28132 24216
rect 28092 23866 28120 24210
rect 28172 24200 28224 24206
rect 28172 24142 28224 24148
rect 28184 23866 28212 24142
rect 28080 23860 28132 23866
rect 28080 23802 28132 23808
rect 28172 23860 28224 23866
rect 28172 23802 28224 23808
rect 28078 23624 28134 23633
rect 28078 23559 28134 23568
rect 28092 23118 28120 23559
rect 28172 23520 28224 23526
rect 28172 23462 28224 23468
rect 28184 23322 28212 23462
rect 28172 23316 28224 23322
rect 28172 23258 28224 23264
rect 28080 23112 28132 23118
rect 28080 23054 28132 23060
rect 28092 22778 28120 23054
rect 28080 22772 28132 22778
rect 28080 22714 28132 22720
rect 28368 22080 28396 34575
rect 32140 34542 32168 35022
rect 33060 34542 33088 35158
rect 33428 34626 33456 35226
rect 33232 34604 33284 34610
rect 33232 34546 33284 34552
rect 33336 34598 33456 34626
rect 32128 34536 32180 34542
rect 32128 34478 32180 34484
rect 33048 34536 33100 34542
rect 33048 34478 33100 34484
rect 30564 34468 30616 34474
rect 30564 34410 30616 34416
rect 30012 34400 30064 34406
rect 30012 34342 30064 34348
rect 30024 33454 30052 34342
rect 30576 34202 30604 34410
rect 31852 34400 31904 34406
rect 31852 34342 31904 34348
rect 30564 34196 30616 34202
rect 30564 34138 30616 34144
rect 30104 33856 30156 33862
rect 30104 33798 30156 33804
rect 30116 33454 30144 33798
rect 30576 33674 30604 34138
rect 31864 34134 31892 34342
rect 31852 34128 31904 34134
rect 31852 34070 31904 34076
rect 32140 33998 32168 34478
rect 32956 34400 33008 34406
rect 32956 34342 33008 34348
rect 32864 34128 32916 34134
rect 32864 34070 32916 34076
rect 32128 33992 32180 33998
rect 32128 33934 32180 33940
rect 30576 33658 30696 33674
rect 30576 33652 30708 33658
rect 30576 33646 30656 33652
rect 30656 33594 30708 33600
rect 32140 33590 32168 33934
rect 32496 33652 32548 33658
rect 32496 33594 32548 33600
rect 32128 33584 32180 33590
rect 32128 33526 32180 33532
rect 32508 33522 32536 33594
rect 32496 33516 32548 33522
rect 32496 33458 32548 33464
rect 30012 33448 30064 33454
rect 30012 33390 30064 33396
rect 30104 33448 30156 33454
rect 30104 33390 30156 33396
rect 30288 33448 30340 33454
rect 30340 33408 30420 33436
rect 30288 33390 30340 33396
rect 29460 33312 29512 33318
rect 29460 33254 29512 33260
rect 29472 32910 29500 33254
rect 30392 33114 30420 33408
rect 32312 33312 32364 33318
rect 32312 33254 32364 33260
rect 30380 33108 30432 33114
rect 30380 33050 30432 33056
rect 30748 33108 30800 33114
rect 30748 33050 30800 33056
rect 29736 32972 29788 32978
rect 29736 32914 29788 32920
rect 29460 32904 29512 32910
rect 29460 32846 29512 32852
rect 29472 32230 29500 32846
rect 29748 32570 29776 32914
rect 29736 32564 29788 32570
rect 29736 32506 29788 32512
rect 28448 32224 28500 32230
rect 28448 32166 28500 32172
rect 29460 32224 29512 32230
rect 29460 32166 29512 32172
rect 28460 31686 28488 32166
rect 29748 32026 29776 32506
rect 30760 32366 30788 33050
rect 30932 32768 30984 32774
rect 30932 32710 30984 32716
rect 30944 32434 30972 32710
rect 30932 32428 30984 32434
rect 30932 32370 30984 32376
rect 30748 32360 30800 32366
rect 30748 32302 30800 32308
rect 30760 32026 30788 32302
rect 30944 32026 30972 32370
rect 32324 32366 32352 33254
rect 32508 33114 32536 33458
rect 32876 33454 32904 34070
rect 32864 33448 32916 33454
rect 32864 33390 32916 33396
rect 32876 33114 32904 33390
rect 32496 33108 32548 33114
rect 32496 33050 32548 33056
rect 32864 33108 32916 33114
rect 32864 33050 32916 33056
rect 32588 32428 32640 32434
rect 32588 32370 32640 32376
rect 32312 32360 32364 32366
rect 32312 32302 32364 32308
rect 31944 32224 31996 32230
rect 31944 32166 31996 32172
rect 29736 32020 29788 32026
rect 29736 31962 29788 31968
rect 30748 32020 30800 32026
rect 30748 31962 30800 31968
rect 30932 32020 30984 32026
rect 30932 31962 30984 31968
rect 31668 32020 31720 32026
rect 31668 31962 31720 31968
rect 28540 31884 28592 31890
rect 28540 31826 28592 31832
rect 31024 31884 31076 31890
rect 31024 31826 31076 31832
rect 28448 31680 28500 31686
rect 28448 31622 28500 31628
rect 28460 31142 28488 31622
rect 28552 31142 28580 31826
rect 31036 31482 31064 31826
rect 31680 31498 31708 31962
rect 31852 31680 31904 31686
rect 31852 31622 31904 31628
rect 31024 31476 31076 31482
rect 31680 31470 31800 31498
rect 31024 31418 31076 31424
rect 31772 31346 31800 31470
rect 31760 31340 31812 31346
rect 31760 31282 31812 31288
rect 28448 31136 28500 31142
rect 28448 31078 28500 31084
rect 28540 31136 28592 31142
rect 28540 31078 28592 31084
rect 28460 30326 28488 31078
rect 28552 30394 28580 31078
rect 29276 30592 29328 30598
rect 29276 30534 29328 30540
rect 29644 30592 29696 30598
rect 29644 30534 29696 30540
rect 28540 30388 28592 30394
rect 28540 30330 28592 30336
rect 28448 30320 28500 30326
rect 28448 30262 28500 30268
rect 28460 29714 28488 30262
rect 29288 30258 29316 30534
rect 29276 30252 29328 30258
rect 29276 30194 29328 30200
rect 29000 30048 29052 30054
rect 29000 29990 29052 29996
rect 28448 29708 28500 29714
rect 28448 29650 28500 29656
rect 28448 29232 28500 29238
rect 28448 29174 28500 29180
rect 28460 28966 28488 29174
rect 28448 28960 28500 28966
rect 28448 28902 28500 28908
rect 28540 28960 28592 28966
rect 28540 28902 28592 28908
rect 28448 26512 28500 26518
rect 28552 26500 28580 28902
rect 29012 28098 29040 29990
rect 29288 29782 29316 30194
rect 29656 30190 29684 30534
rect 29644 30184 29696 30190
rect 29644 30126 29696 30132
rect 29460 30048 29512 30054
rect 29460 29990 29512 29996
rect 29276 29776 29328 29782
rect 29276 29718 29328 29724
rect 29092 29708 29144 29714
rect 29092 29650 29144 29656
rect 29104 28966 29132 29650
rect 29092 28960 29144 28966
rect 29092 28902 29144 28908
rect 29104 28558 29132 28902
rect 29288 28762 29316 29718
rect 29276 28756 29328 28762
rect 29276 28698 29328 28704
rect 29092 28552 29144 28558
rect 29092 28494 29144 28500
rect 28920 28070 29040 28098
rect 28920 28014 28948 28070
rect 28908 28008 28960 28014
rect 28908 27950 28960 27956
rect 29104 27878 29132 28494
rect 29276 27940 29328 27946
rect 29276 27882 29328 27888
rect 29092 27872 29144 27878
rect 29092 27814 29144 27820
rect 28724 27600 28776 27606
rect 28724 27542 28776 27548
rect 28736 27062 28764 27542
rect 28724 27056 28776 27062
rect 28724 26998 28776 27004
rect 29104 26790 29132 27814
rect 29288 27538 29316 27882
rect 29276 27532 29328 27538
rect 29276 27474 29328 27480
rect 29288 27130 29316 27474
rect 29472 27470 29500 29990
rect 29656 29850 29684 30126
rect 29644 29844 29696 29850
rect 29644 29786 29696 29792
rect 29656 29034 29684 29786
rect 30288 29232 30340 29238
rect 30288 29174 30340 29180
rect 29644 29028 29696 29034
rect 29644 28970 29696 28976
rect 30300 28694 30328 29174
rect 29552 28688 29604 28694
rect 29552 28630 29604 28636
rect 30288 28688 30340 28694
rect 30288 28630 30340 28636
rect 29564 27674 29592 28630
rect 30288 28416 30340 28422
rect 30288 28358 30340 28364
rect 29552 27668 29604 27674
rect 29552 27610 29604 27616
rect 30300 27538 30328 28358
rect 31864 27946 31892 31622
rect 31956 31278 31984 32166
rect 32600 31822 32628 32370
rect 32968 32026 32996 34342
rect 33244 33862 33272 34546
rect 33336 34474 33364 34598
rect 33324 34468 33376 34474
rect 33324 34410 33376 34416
rect 33336 34134 33364 34410
rect 33508 34400 33560 34406
rect 33508 34342 33560 34348
rect 33520 34202 33548 34342
rect 33508 34196 33560 34202
rect 33508 34138 33560 34144
rect 33324 34128 33376 34134
rect 33324 34070 33376 34076
rect 33232 33856 33284 33862
rect 33232 33798 33284 33804
rect 33244 33522 33272 33798
rect 33876 33652 33928 33658
rect 33876 33594 33928 33600
rect 33232 33516 33284 33522
rect 33232 33458 33284 33464
rect 33244 32774 33272 33458
rect 33888 33114 33916 33594
rect 33876 33108 33928 33114
rect 33876 33050 33928 33056
rect 33600 32904 33652 32910
rect 33600 32846 33652 32852
rect 33232 32768 33284 32774
rect 33232 32710 33284 32716
rect 33508 32768 33560 32774
rect 33508 32710 33560 32716
rect 33244 32026 33272 32710
rect 32956 32020 33008 32026
rect 32956 31962 33008 31968
rect 33232 32020 33284 32026
rect 33232 31962 33284 31968
rect 32772 31952 32824 31958
rect 32772 31894 32824 31900
rect 32588 31816 32640 31822
rect 32588 31758 32640 31764
rect 32784 31482 32812 31894
rect 32772 31476 32824 31482
rect 32772 31418 32824 31424
rect 31944 31272 31996 31278
rect 31944 31214 31996 31220
rect 32968 30938 32996 31962
rect 33244 30938 33272 31962
rect 33520 31958 33548 32710
rect 33612 32502 33640 32846
rect 33888 32570 33916 33050
rect 33876 32564 33928 32570
rect 33876 32506 33928 32512
rect 33600 32496 33652 32502
rect 33600 32438 33652 32444
rect 33980 32230 34008 35663
rect 34796 35488 34848 35494
rect 35820 35442 35848 36178
rect 35900 35488 35952 35494
rect 34796 35430 34848 35436
rect 35544 35436 35900 35442
rect 35544 35430 35952 35436
rect 34520 35148 34572 35154
rect 34520 35090 34572 35096
rect 34532 34950 34560 35090
rect 34612 35080 34664 35086
rect 34612 35022 34664 35028
rect 34520 34944 34572 34950
rect 34348 34904 34520 34932
rect 34348 32978 34376 34904
rect 34520 34886 34572 34892
rect 34532 34746 34560 34886
rect 34520 34740 34572 34746
rect 34520 34682 34572 34688
rect 34624 34678 34652 35022
rect 34612 34672 34664 34678
rect 34612 34614 34664 34620
rect 34428 34468 34480 34474
rect 34428 34410 34480 34416
rect 34440 34134 34468 34410
rect 34428 34128 34480 34134
rect 34428 34070 34480 34076
rect 34520 34128 34572 34134
rect 34520 34070 34572 34076
rect 34532 33658 34560 34070
rect 34624 33998 34652 34614
rect 34612 33992 34664 33998
rect 34612 33934 34664 33940
rect 34520 33652 34572 33658
rect 34520 33594 34572 33600
rect 34624 33318 34652 33934
rect 34612 33312 34664 33318
rect 34612 33254 34664 33260
rect 34336 32972 34388 32978
rect 34336 32914 34388 32920
rect 34624 32910 34652 33254
rect 34612 32904 34664 32910
rect 34612 32846 34664 32852
rect 34624 32570 34652 32846
rect 34612 32564 34664 32570
rect 34612 32506 34664 32512
rect 33968 32224 34020 32230
rect 34336 32224 34388 32230
rect 33968 32166 34020 32172
rect 34334 32192 34336 32201
rect 34388 32192 34390 32201
rect 34624 32178 34652 32506
rect 34334 32127 34390 32136
rect 34532 32150 34652 32178
rect 34704 32224 34756 32230
rect 34704 32166 34756 32172
rect 33508 31952 33560 31958
rect 33508 31894 33560 31900
rect 34532 31890 34560 32150
rect 34612 32020 34664 32026
rect 34612 31962 34664 31968
rect 34520 31884 34572 31890
rect 34520 31826 34572 31832
rect 34060 31680 34112 31686
rect 34060 31622 34112 31628
rect 34072 31346 34100 31622
rect 34624 31346 34652 31962
rect 34060 31340 34112 31346
rect 34060 31282 34112 31288
rect 34428 31340 34480 31346
rect 34428 31282 34480 31288
rect 34612 31340 34664 31346
rect 34612 31282 34664 31288
rect 33324 31136 33376 31142
rect 33324 31078 33376 31084
rect 32956 30932 33008 30938
rect 32956 30874 33008 30880
rect 33232 30932 33284 30938
rect 33232 30874 33284 30880
rect 32128 30796 32180 30802
rect 32128 30738 32180 30744
rect 33140 30796 33192 30802
rect 33140 30738 33192 30744
rect 32140 30190 32168 30738
rect 33152 30682 33180 30738
rect 33060 30654 33180 30682
rect 32312 30592 32364 30598
rect 32312 30534 32364 30540
rect 32324 30433 32352 30534
rect 32310 30424 32366 30433
rect 32310 30359 32366 30368
rect 33060 30258 33088 30654
rect 33140 30592 33192 30598
rect 33140 30534 33192 30540
rect 33152 30394 33180 30534
rect 33140 30388 33192 30394
rect 33140 30330 33192 30336
rect 33048 30252 33100 30258
rect 33048 30194 33100 30200
rect 32128 30184 32180 30190
rect 32128 30126 32180 30132
rect 32956 29776 33008 29782
rect 32956 29718 33008 29724
rect 32864 29640 32916 29646
rect 32310 29608 32366 29617
rect 32864 29582 32916 29588
rect 32310 29543 32366 29552
rect 32324 29306 32352 29543
rect 32876 29306 32904 29582
rect 32312 29300 32364 29306
rect 32312 29242 32364 29248
rect 32864 29300 32916 29306
rect 32864 29242 32916 29248
rect 32876 29170 32904 29242
rect 32864 29164 32916 29170
rect 32864 29106 32916 29112
rect 32876 28626 32904 29106
rect 32968 28762 32996 29718
rect 33152 29322 33180 30330
rect 33244 30258 33272 30874
rect 33232 30252 33284 30258
rect 33232 30194 33284 30200
rect 33060 29306 33180 29322
rect 33048 29300 33180 29306
rect 33100 29294 33180 29300
rect 33048 29242 33100 29248
rect 33060 29034 33180 29050
rect 33048 29028 33180 29034
rect 33100 29022 33180 29028
rect 33048 28970 33100 28976
rect 32956 28756 33008 28762
rect 32956 28698 33008 28704
rect 32864 28620 32916 28626
rect 32864 28562 32916 28568
rect 33048 28620 33100 28626
rect 33048 28562 33100 28568
rect 32586 28520 32642 28529
rect 32586 28455 32642 28464
rect 32600 28218 32628 28455
rect 32588 28212 32640 28218
rect 32588 28154 32640 28160
rect 32600 28014 32628 28154
rect 33060 28098 33088 28562
rect 33152 28218 33180 29022
rect 33232 28960 33284 28966
rect 33232 28902 33284 28908
rect 33140 28212 33192 28218
rect 33140 28154 33192 28160
rect 33060 28082 33180 28098
rect 33060 28076 33192 28082
rect 33060 28070 33140 28076
rect 32588 28008 32640 28014
rect 32588 27950 32640 27956
rect 31852 27940 31904 27946
rect 31852 27882 31904 27888
rect 30656 27872 30708 27878
rect 30656 27814 30708 27820
rect 32128 27872 32180 27878
rect 32128 27814 32180 27820
rect 30668 27538 30696 27814
rect 30288 27532 30340 27538
rect 30288 27474 30340 27480
rect 30472 27532 30524 27538
rect 30472 27474 30524 27480
rect 30656 27532 30708 27538
rect 30656 27474 30708 27480
rect 31944 27532 31996 27538
rect 31944 27474 31996 27480
rect 29460 27464 29512 27470
rect 29460 27406 29512 27412
rect 29276 27124 29328 27130
rect 29276 27066 29328 27072
rect 29092 26784 29144 26790
rect 28722 26752 28778 26761
rect 29092 26726 29144 26732
rect 29276 26784 29328 26790
rect 29276 26726 29328 26732
rect 28722 26687 28778 26696
rect 28500 26472 28580 26500
rect 28448 26454 28500 26460
rect 28460 25974 28488 26454
rect 28736 26382 28764 26687
rect 28816 26580 28868 26586
rect 28816 26522 28868 26528
rect 28724 26376 28776 26382
rect 28724 26318 28776 26324
rect 28448 25968 28500 25974
rect 28448 25910 28500 25916
rect 28448 25832 28500 25838
rect 28448 25774 28500 25780
rect 28460 25430 28488 25774
rect 28736 25430 28764 26318
rect 28448 25424 28500 25430
rect 28448 25366 28500 25372
rect 28724 25424 28776 25430
rect 28724 25366 28776 25372
rect 28828 24818 28856 26522
rect 29288 25702 29316 26726
rect 29472 26518 29500 27406
rect 30484 27305 30512 27474
rect 30470 27296 30526 27305
rect 30470 27231 30526 27240
rect 30484 26586 30512 27231
rect 30668 27130 30696 27474
rect 30656 27124 30708 27130
rect 30656 27066 30708 27072
rect 30668 26926 30696 27066
rect 30656 26920 30708 26926
rect 30656 26862 30708 26868
rect 30840 26784 30892 26790
rect 30840 26726 30892 26732
rect 30472 26580 30524 26586
rect 30472 26522 30524 26528
rect 29460 26512 29512 26518
rect 30380 26512 30432 26518
rect 29460 26454 29512 26460
rect 30286 26480 30342 26489
rect 30196 26444 30248 26450
rect 30380 26454 30432 26460
rect 30286 26415 30342 26424
rect 30196 26386 30248 26392
rect 29828 26376 29880 26382
rect 29828 26318 29880 26324
rect 29840 25838 29868 26318
rect 29828 25832 29880 25838
rect 29828 25774 29880 25780
rect 30012 25764 30064 25770
rect 30012 25706 30064 25712
rect 29276 25696 29328 25702
rect 29276 25638 29328 25644
rect 29000 25152 29052 25158
rect 28920 25112 29000 25140
rect 28816 24812 28868 24818
rect 28816 24754 28868 24760
rect 28920 24682 28948 25112
rect 29000 25094 29052 25100
rect 29288 24818 29316 25638
rect 30024 25294 30052 25706
rect 30208 25498 30236 26386
rect 30300 26382 30328 26415
rect 30288 26376 30340 26382
rect 30288 26318 30340 26324
rect 30104 25492 30156 25498
rect 30104 25434 30156 25440
rect 30196 25492 30248 25498
rect 30196 25434 30248 25440
rect 30012 25288 30064 25294
rect 30012 25230 30064 25236
rect 29276 24812 29328 24818
rect 29276 24754 29328 24760
rect 28908 24676 28960 24682
rect 28908 24618 28960 24624
rect 29552 24676 29604 24682
rect 29552 24618 29604 24624
rect 29564 24177 29592 24618
rect 29920 24608 29972 24614
rect 29920 24550 29972 24556
rect 29932 24274 29960 24550
rect 30116 24410 30144 25434
rect 30104 24404 30156 24410
rect 30104 24346 30156 24352
rect 29920 24268 29972 24274
rect 29920 24210 29972 24216
rect 29550 24168 29606 24177
rect 29550 24103 29606 24112
rect 28908 24064 28960 24070
rect 28908 24006 28960 24012
rect 28540 23316 28592 23322
rect 28540 23258 28592 23264
rect 28552 22778 28580 23258
rect 28920 23118 28948 24006
rect 29932 23730 29960 24210
rect 29920 23724 29972 23730
rect 29920 23666 29972 23672
rect 29276 23656 29328 23662
rect 29276 23598 29328 23604
rect 29734 23624 29790 23633
rect 29092 23520 29144 23526
rect 29092 23462 29144 23468
rect 29104 23322 29132 23462
rect 29092 23316 29144 23322
rect 29092 23258 29144 23264
rect 28908 23112 28960 23118
rect 28908 23054 28960 23060
rect 28540 22772 28592 22778
rect 28540 22714 28592 22720
rect 28908 22228 28960 22234
rect 29104 22216 29132 23258
rect 29184 22568 29236 22574
rect 29184 22510 29236 22516
rect 28960 22188 29132 22216
rect 28908 22170 28960 22176
rect 28368 22052 28580 22080
rect 27816 21950 27936 21978
rect 27252 21412 27304 21418
rect 27252 21354 27304 21360
rect 26976 21344 27028 21350
rect 26976 21286 27028 21292
rect 27436 21344 27488 21350
rect 27436 21286 27488 21292
rect 26988 21010 27016 21286
rect 26976 21004 27028 21010
rect 26976 20946 27028 20952
rect 26792 20596 26844 20602
rect 26792 20538 26844 20544
rect 26516 20528 26568 20534
rect 26516 20470 26568 20476
rect 26528 19854 26556 20470
rect 26988 20398 27016 20946
rect 27068 20936 27120 20942
rect 27068 20878 27120 20884
rect 27344 20936 27396 20942
rect 27344 20878 27396 20884
rect 26976 20392 27028 20398
rect 26976 20334 27028 20340
rect 27080 20058 27108 20878
rect 27356 20330 27384 20878
rect 27344 20324 27396 20330
rect 27344 20266 27396 20272
rect 26700 20052 26752 20058
rect 26700 19994 26752 20000
rect 27068 20052 27120 20058
rect 27068 19994 27120 20000
rect 26516 19848 26568 19854
rect 26516 19790 26568 19796
rect 26712 19514 26740 19994
rect 27068 19848 27120 19854
rect 27068 19790 27120 19796
rect 27080 19514 27108 19790
rect 26332 19508 26384 19514
rect 26332 19450 26384 19456
rect 26700 19508 26752 19514
rect 26700 19450 26752 19456
rect 27068 19508 27120 19514
rect 27068 19450 27120 19456
rect 25504 19304 25556 19310
rect 25504 19246 25556 19252
rect 26056 19304 26108 19310
rect 26056 19246 26108 19252
rect 25516 19174 25544 19246
rect 27448 19242 27476 21286
rect 27528 20392 27580 20398
rect 27580 20352 27660 20380
rect 27528 20334 27580 20340
rect 27528 20256 27580 20262
rect 27528 20198 27580 20204
rect 27540 19310 27568 20198
rect 27528 19304 27580 19310
rect 27528 19246 27580 19252
rect 27436 19236 27488 19242
rect 27436 19178 27488 19184
rect 25504 19168 25556 19174
rect 25504 19110 25556 19116
rect 27540 18970 27568 19246
rect 27528 18964 27580 18970
rect 27528 18906 27580 18912
rect 27160 18624 27212 18630
rect 27160 18566 27212 18572
rect 26514 18456 26570 18465
rect 26514 18391 26516 18400
rect 26568 18391 26570 18400
rect 26516 18362 26568 18368
rect 26528 18154 26556 18362
rect 27172 18222 27200 18566
rect 27436 18352 27488 18358
rect 27436 18294 27488 18300
rect 27344 18284 27396 18290
rect 27344 18226 27396 18232
rect 27160 18216 27212 18222
rect 27160 18158 27212 18164
rect 26516 18148 26568 18154
rect 26516 18090 26568 18096
rect 26608 17672 26660 17678
rect 26608 17614 26660 17620
rect 25412 17264 25464 17270
rect 25412 17206 25464 17212
rect 25424 16726 25452 17206
rect 25688 17060 25740 17066
rect 25688 17002 25740 17008
rect 25700 16794 25728 17002
rect 25688 16788 25740 16794
rect 25688 16730 25740 16736
rect 25412 16720 25464 16726
rect 25412 16662 25464 16668
rect 25700 16153 25728 16730
rect 26514 16688 26570 16697
rect 26332 16652 26384 16658
rect 26514 16623 26570 16632
rect 26332 16594 26384 16600
rect 26238 16280 26294 16289
rect 26238 16215 26240 16224
rect 26292 16215 26294 16224
rect 26240 16186 26292 16192
rect 25686 16144 25742 16153
rect 25686 16079 25742 16088
rect 25136 16040 25188 16046
rect 25136 15982 25188 15988
rect 26054 15736 26110 15745
rect 26344 15706 26372 16594
rect 26528 16590 26556 16623
rect 26516 16584 26568 16590
rect 26516 16526 26568 16532
rect 26528 16182 26556 16526
rect 26620 16250 26648 17614
rect 27172 16833 27200 18158
rect 27250 17912 27306 17921
rect 27250 17847 27306 17856
rect 27158 16824 27214 16833
rect 27158 16759 27214 16768
rect 27264 16658 27292 17847
rect 27356 16794 27384 18226
rect 27344 16788 27396 16794
rect 27344 16730 27396 16736
rect 27252 16652 27304 16658
rect 27252 16594 27304 16600
rect 26608 16244 26660 16250
rect 26608 16186 26660 16192
rect 26516 16176 26568 16182
rect 26516 16118 26568 16124
rect 26054 15671 26110 15680
rect 26332 15700 26384 15706
rect 26068 15162 26096 15671
rect 26332 15642 26384 15648
rect 26528 15570 26556 16118
rect 27356 15638 27384 16730
rect 27448 15994 27476 18294
rect 27632 17746 27660 20352
rect 27816 20058 27844 21950
rect 27896 21888 27948 21894
rect 27896 21830 27948 21836
rect 27908 20466 27936 21830
rect 28446 21448 28502 21457
rect 28446 21383 28502 21392
rect 28460 21146 28488 21383
rect 28448 21140 28500 21146
rect 28448 21082 28500 21088
rect 27896 20460 27948 20466
rect 27896 20402 27948 20408
rect 27804 20052 27856 20058
rect 27804 19994 27856 20000
rect 27816 19378 27844 19994
rect 27908 19990 27936 20402
rect 28080 20324 28132 20330
rect 28080 20266 28132 20272
rect 27988 20256 28040 20262
rect 27986 20224 27988 20233
rect 28040 20224 28042 20233
rect 27986 20159 28042 20168
rect 27896 19984 27948 19990
rect 27896 19926 27948 19932
rect 27908 19514 27936 19926
rect 28092 19922 28120 20266
rect 28080 19916 28132 19922
rect 28080 19858 28132 19864
rect 28092 19553 28120 19858
rect 28078 19544 28134 19553
rect 27896 19508 27948 19514
rect 28078 19479 28134 19488
rect 27896 19450 27948 19456
rect 27804 19372 27856 19378
rect 27804 19314 27856 19320
rect 27802 19272 27858 19281
rect 27802 19207 27858 19216
rect 27620 17740 27672 17746
rect 27620 17682 27672 17688
rect 27712 17672 27764 17678
rect 27712 17614 27764 17620
rect 27620 17060 27672 17066
rect 27620 17002 27672 17008
rect 27632 16946 27660 17002
rect 27724 16998 27752 17614
rect 27540 16918 27660 16946
rect 27712 16992 27764 16998
rect 27712 16934 27764 16940
rect 27540 16182 27568 16918
rect 27528 16176 27580 16182
rect 27528 16118 27580 16124
rect 27448 15978 27660 15994
rect 27448 15972 27672 15978
rect 27448 15966 27620 15972
rect 26976 15632 27028 15638
rect 26976 15574 27028 15580
rect 27344 15632 27396 15638
rect 27344 15574 27396 15580
rect 26516 15564 26568 15570
rect 26516 15506 26568 15512
rect 26528 15162 26556 15506
rect 26988 15162 27016 15574
rect 27448 15162 27476 15966
rect 27620 15914 27672 15920
rect 26056 15156 26108 15162
rect 26056 15098 26108 15104
rect 26516 15156 26568 15162
rect 26516 15098 26568 15104
rect 26976 15156 27028 15162
rect 26976 15098 27028 15104
rect 27436 15156 27488 15162
rect 27436 15098 27488 15104
rect 26068 14958 26096 15098
rect 24768 14952 24820 14958
rect 24768 14894 24820 14900
rect 26056 14952 26108 14958
rect 26056 14894 26108 14900
rect 24032 14612 24084 14618
rect 24032 14554 24084 14560
rect 24308 14612 24360 14618
rect 24308 14554 24360 14560
rect 22376 14476 22428 14482
rect 22376 14418 22428 14424
rect 22388 14074 22416 14418
rect 21732 14068 21784 14074
rect 21732 14010 21784 14016
rect 22376 14068 22428 14074
rect 22376 14010 22428 14016
rect 21640 14000 21692 14006
rect 25596 14000 25648 14006
rect 21640 13942 21692 13948
rect 25594 13968 25596 13977
rect 25648 13968 25650 13977
rect 25594 13903 25650 13912
rect 25688 13796 25740 13802
rect 25688 13738 25740 13744
rect 21088 13388 21140 13394
rect 21088 13330 21140 13336
rect 22192 13388 22244 13394
rect 22192 13330 22244 13336
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19340 12708 19392 12714
rect 19340 12650 19392 12656
rect 19444 11626 19472 12922
rect 21100 12782 21128 13330
rect 21916 13184 21968 13190
rect 21916 13126 21968 13132
rect 21928 13025 21956 13126
rect 21914 13016 21970 13025
rect 21914 12951 21970 12960
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 20628 12708 20680 12714
rect 20628 12650 20680 12656
rect 21272 12708 21324 12714
rect 21272 12650 21324 12656
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 20640 12442 20668 12650
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 20640 11898 20668 12378
rect 21284 12238 21312 12650
rect 21730 12336 21786 12345
rect 21730 12271 21786 12280
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21088 12096 21140 12102
rect 21088 12038 21140 12044
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20626 11792 20682 11801
rect 20626 11727 20682 11736
rect 19432 11620 19484 11626
rect 19432 11562 19484 11568
rect 19444 11354 19472 11562
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 20640 11098 20668 11727
rect 21100 11354 21128 12038
rect 21284 11898 21312 12174
rect 21744 11898 21772 12271
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 21732 11892 21784 11898
rect 21732 11834 21784 11840
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 20996 11280 21048 11286
rect 20996 11222 21048 11228
rect 20720 11144 20772 11150
rect 20640 11092 20720 11098
rect 20640 11086 20772 11092
rect 20810 11112 20866 11121
rect 20640 11070 20760 11086
rect 19156 10804 19208 10810
rect 19260 10798 19380 10826
rect 19156 10746 19208 10752
rect 17038 9551 17040 9560
rect 17092 9551 17094 9560
rect 18236 9580 18288 9586
rect 17040 9522 17092 9528
rect 18236 9522 18288 9528
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 18420 9512 18472 9518
rect 18420 9454 18472 9460
rect 16776 9382 16804 9454
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16684 9178 16804 9194
rect 18432 9178 18460 9454
rect 18708 9178 18736 9522
rect 19168 9518 19196 10746
rect 19352 10130 19380 10798
rect 20640 10470 20668 11070
rect 20810 11047 20812 11056
rect 20864 11047 20866 11056
rect 20812 11018 20864 11024
rect 21008 10810 21036 11222
rect 21100 10810 21128 11290
rect 21272 11008 21324 11014
rect 21272 10950 21324 10956
rect 20996 10804 21048 10810
rect 20996 10746 21048 10752
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19352 10010 19380 10066
rect 19352 9982 19472 10010
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19156 9512 19208 9518
rect 19156 9454 19208 9460
rect 19352 9178 19380 9862
rect 19444 9722 19472 9982
rect 19432 9716 19484 9722
rect 19432 9658 19484 9664
rect 20640 9625 20668 10406
rect 21284 10130 21312 10950
rect 21272 10124 21324 10130
rect 21272 10066 21324 10072
rect 21088 9920 21140 9926
rect 21088 9862 21140 9868
rect 20626 9616 20682 9625
rect 20626 9551 20682 9560
rect 20640 9518 20668 9551
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 16684 9172 16816 9178
rect 16684 9166 16764 9172
rect 16764 9114 16816 9120
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 18420 9172 18472 9178
rect 18420 9114 18472 9120
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 16672 9104 16724 9110
rect 16672 9046 16724 9052
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16684 8362 16712 9046
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16316 8022 16344 8230
rect 16684 8090 16712 8298
rect 16776 8294 16804 9114
rect 17420 8634 17448 9114
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 18708 8498 18736 9114
rect 18972 8968 19024 8974
rect 18972 8910 19024 8916
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 17328 8090 17356 8434
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 16304 8016 16356 8022
rect 16304 7958 16356 7964
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15212 7206 15240 7822
rect 16316 7274 16344 7958
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 17038 7304 17094 7313
rect 16304 7268 16356 7274
rect 17038 7239 17094 7248
rect 16304 7210 16356 7216
rect 17052 7206 17080 7239
rect 17788 7206 17816 7890
rect 18892 7886 18920 8774
rect 18984 8634 19012 8910
rect 19352 8634 19380 9114
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19536 8362 19564 8910
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 19892 8560 19944 8566
rect 19892 8502 19944 8508
rect 19524 8356 19576 8362
rect 19524 8298 19576 8304
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 19904 7886 19932 8502
rect 20548 8430 20576 8774
rect 20640 8634 20668 9318
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 20640 8430 20668 8570
rect 20536 8424 20588 8430
rect 20536 8366 20588 8372
rect 20628 8424 20680 8430
rect 20628 8366 20680 8372
rect 20168 8356 20220 8362
rect 20168 8298 20220 8304
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 17040 7200 17092 7206
rect 17040 7142 17092 7148
rect 17776 7200 17828 7206
rect 17776 7142 17828 7148
rect 15212 6798 15240 7142
rect 16856 6860 16908 6866
rect 16856 6802 16908 6808
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14384 6322 14412 6598
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 14384 5914 14412 6258
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14372 5908 14424 5914
rect 14372 5850 14424 5856
rect 14188 5840 14240 5846
rect 14188 5782 14240 5788
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13832 5234 13860 5510
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 13832 5114 13860 5170
rect 13832 5086 13952 5114
rect 13740 4984 13860 5012
rect 13360 4480 13412 4486
rect 13360 4422 13412 4428
rect 13372 3777 13400 4422
rect 13740 4146 13768 4984
rect 13832 4826 13860 4984
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13832 4026 13860 4422
rect 13740 4010 13860 4026
rect 13728 4004 13860 4010
rect 13780 3998 13860 4004
rect 13728 3946 13780 3952
rect 13450 3904 13506 3913
rect 13450 3839 13506 3848
rect 13358 3768 13414 3777
rect 13358 3703 13414 3712
rect 13372 3369 13400 3703
rect 13358 3360 13414 3369
rect 13358 3295 13414 3304
rect 13464 3058 13492 3839
rect 13924 3738 13952 5086
rect 14004 5092 14056 5098
rect 14004 5034 14056 5040
rect 14016 4282 14044 5034
rect 14108 4486 14136 5646
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14462 4584 14518 4593
rect 14188 4548 14240 4554
rect 14188 4490 14240 4496
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 13268 2984 13320 2990
rect 12990 2952 13046 2961
rect 13268 2926 13320 2932
rect 12990 2887 13046 2896
rect 13004 2854 13032 2887
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 13004 2689 13032 2790
rect 12990 2680 13046 2689
rect 12990 2615 13046 2624
rect 13740 2582 13768 3334
rect 13924 3058 13952 3674
rect 14200 3398 14228 4490
rect 14188 3392 14240 3398
rect 14188 3334 14240 3340
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 13910 2816 13966 2825
rect 13910 2751 13966 2760
rect 13728 2576 13780 2582
rect 13728 2518 13780 2524
rect 13924 480 13952 2751
rect 14292 2650 14320 4558
rect 14462 4519 14518 4528
rect 14476 3670 14504 4519
rect 14464 3664 14516 3670
rect 14464 3606 14516 3612
rect 14660 2854 14688 6054
rect 14844 5642 14872 6598
rect 16868 6458 16896 6802
rect 18064 6798 18092 7278
rect 18156 7274 18184 7822
rect 19156 7812 19208 7818
rect 19156 7754 19208 7760
rect 19168 7449 19196 7754
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 19260 7546 19288 7686
rect 19904 7546 19932 7822
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 19892 7540 19944 7546
rect 19892 7482 19944 7488
rect 19154 7440 19210 7449
rect 19154 7375 19210 7384
rect 19168 7342 19196 7375
rect 19156 7336 19208 7342
rect 19156 7278 19208 7284
rect 18144 7268 18196 7274
rect 18144 7210 18196 7216
rect 18156 6934 18184 7210
rect 18236 7200 18288 7206
rect 18236 7142 18288 7148
rect 18144 6928 18196 6934
rect 18144 6870 18196 6876
rect 17408 6792 17460 6798
rect 17408 6734 17460 6740
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 17132 6656 17184 6662
rect 17132 6598 17184 6604
rect 17144 6497 17172 6598
rect 17130 6488 17186 6497
rect 16856 6452 16908 6458
rect 17420 6458 17448 6734
rect 17592 6656 17644 6662
rect 17592 6598 17644 6604
rect 17130 6423 17186 6432
rect 17408 6452 17460 6458
rect 16856 6394 16908 6400
rect 17408 6394 17460 6400
rect 17420 6254 17448 6394
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 15580 5914 15608 6054
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15108 5704 15160 5710
rect 15160 5652 15240 5658
rect 15108 5646 15240 5652
rect 14832 5636 14884 5642
rect 15120 5630 15240 5646
rect 14832 5578 14884 5584
rect 14844 2990 14872 5578
rect 15016 5568 15068 5574
rect 15016 5510 15068 5516
rect 15108 5568 15160 5574
rect 15108 5510 15160 5516
rect 14922 4992 14978 5001
rect 14922 4927 14978 4936
rect 14936 3924 14964 4927
rect 15028 4604 15056 5510
rect 15120 4826 15148 5510
rect 15212 5370 15240 5630
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15580 5030 15608 5850
rect 16212 5772 16264 5778
rect 16212 5714 16264 5720
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 15568 5024 15620 5030
rect 15568 4966 15620 4972
rect 15108 4820 15160 4826
rect 15108 4762 15160 4768
rect 15200 4616 15252 4622
rect 15028 4576 15200 4604
rect 15028 4078 15056 4576
rect 15200 4558 15252 4564
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 14936 3896 15056 3924
rect 15304 3913 15332 4422
rect 14832 2984 14884 2990
rect 14832 2926 14884 2932
rect 14648 2848 14700 2854
rect 14648 2790 14700 2796
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 15028 480 15056 3896
rect 15290 3904 15346 3913
rect 15290 3839 15346 3848
rect 15108 3664 15160 3670
rect 15108 3606 15160 3612
rect 15120 3058 15148 3606
rect 15108 3052 15160 3058
rect 15108 2994 15160 3000
rect 15580 2990 15608 4966
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15672 4593 15700 4626
rect 15658 4584 15714 4593
rect 15856 4570 15884 5646
rect 16118 5400 16174 5409
rect 16224 5370 16252 5714
rect 16960 5681 16988 6054
rect 17604 5914 17632 6598
rect 17868 6316 17920 6322
rect 17868 6258 17920 6264
rect 17880 5914 17908 6258
rect 17960 6112 18012 6118
rect 18064 6100 18092 6734
rect 18012 6072 18092 6100
rect 17960 6054 18012 6060
rect 17592 5908 17644 5914
rect 17592 5850 17644 5856
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 16946 5672 17002 5681
rect 16946 5607 17002 5616
rect 17604 5409 17632 5850
rect 18064 5778 18092 6072
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 17684 5568 17736 5574
rect 17684 5510 17736 5516
rect 17590 5400 17646 5409
rect 16118 5335 16174 5344
rect 16212 5364 16264 5370
rect 15764 4554 15884 4570
rect 15658 4519 15714 4528
rect 15752 4548 15884 4554
rect 15672 4282 15700 4519
rect 15804 4542 15884 4548
rect 15752 4490 15804 4496
rect 15764 4321 15792 4490
rect 15842 4448 15898 4457
rect 15842 4383 15898 4392
rect 15750 4312 15806 4321
rect 15660 4276 15712 4282
rect 15750 4247 15806 4256
rect 15660 4218 15712 4224
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15672 3738 15700 3878
rect 15856 3738 15884 4383
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15844 3732 15896 3738
rect 15844 3674 15896 3680
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 15764 3194 15792 3334
rect 15752 3188 15804 3194
rect 15752 3130 15804 3136
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 16132 480 16160 5335
rect 17590 5335 17646 5344
rect 16212 5306 16264 5312
rect 16396 5160 16448 5166
rect 16396 5102 16448 5108
rect 16408 4865 16436 5102
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 16394 4856 16450 4865
rect 16394 4791 16450 4800
rect 16396 4752 16448 4758
rect 16592 4729 16620 4966
rect 16762 4856 16818 4865
rect 17512 4826 17540 4966
rect 16762 4791 16818 4800
rect 17040 4820 17092 4826
rect 16776 4758 16804 4791
rect 17040 4762 17092 4768
rect 17500 4820 17552 4826
rect 17500 4762 17552 4768
rect 16764 4752 16816 4758
rect 16396 4694 16448 4700
rect 16578 4720 16634 4729
rect 16302 4584 16358 4593
rect 16302 4519 16304 4528
rect 16356 4519 16358 4528
rect 16304 4490 16356 4496
rect 16316 3738 16344 4490
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 16408 3534 16436 4694
rect 16764 4694 16816 4700
rect 16578 4655 16634 4664
rect 16488 4616 16540 4622
rect 16540 4564 16712 4570
rect 16488 4558 16712 4564
rect 16500 4542 16712 4558
rect 16684 3942 16712 4542
rect 16764 4072 16816 4078
rect 16762 4040 16764 4049
rect 16816 4040 16818 4049
rect 16762 3975 16818 3984
rect 16672 3936 16724 3942
rect 16948 3936 17000 3942
rect 16672 3878 16724 3884
rect 16854 3904 16910 3913
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16684 2650 16712 3878
rect 16948 3878 17000 3884
rect 16854 3839 16910 3848
rect 16868 3738 16896 3839
rect 16856 3732 16908 3738
rect 16856 3674 16908 3680
rect 16960 3641 16988 3878
rect 16946 3632 17002 3641
rect 16946 3567 17002 3576
rect 17052 3194 17080 4762
rect 17406 4312 17462 4321
rect 17406 4247 17462 4256
rect 17222 3496 17278 3505
rect 17222 3431 17278 3440
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 17236 480 17264 3431
rect 17420 2650 17448 4247
rect 17500 3732 17552 3738
rect 17500 3674 17552 3680
rect 17512 3233 17540 3674
rect 17604 3534 17632 5335
rect 17696 5234 17724 5510
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17880 4706 17908 5646
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 17972 5370 18000 5510
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17972 4826 18000 5306
rect 18064 5098 18092 5714
rect 18052 5092 18104 5098
rect 18052 5034 18104 5040
rect 17960 4820 18012 4826
rect 17960 4762 18012 4768
rect 17788 4690 18000 4706
rect 17788 4684 18012 4690
rect 17788 4678 17960 4684
rect 17788 4146 17816 4678
rect 17960 4626 18012 4632
rect 17868 4548 17920 4554
rect 17868 4490 17920 4496
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 17880 3534 17908 4490
rect 18064 3942 18092 5034
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 18248 4978 18276 7142
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 19996 7002 20024 8026
rect 20074 7304 20130 7313
rect 20074 7239 20130 7248
rect 19984 6996 20036 7002
rect 19984 6938 20036 6944
rect 19156 6656 19208 6662
rect 19156 6598 19208 6604
rect 19168 6458 19196 6598
rect 19430 6488 19486 6497
rect 19156 6452 19208 6458
rect 19430 6423 19432 6432
rect 19156 6394 19208 6400
rect 19484 6423 19486 6432
rect 19432 6394 19484 6400
rect 19168 6322 19196 6394
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 18512 6112 18564 6118
rect 18512 6054 18564 6060
rect 18524 5030 18552 6054
rect 18708 5846 18736 6258
rect 19444 6254 19472 6394
rect 19996 6390 20024 6938
rect 19984 6384 20036 6390
rect 19984 6326 20036 6332
rect 20088 6322 20116 7239
rect 20076 6316 20128 6322
rect 20076 6258 20128 6264
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 20088 5914 20116 6258
rect 20076 5908 20128 5914
rect 20076 5850 20128 5856
rect 18696 5840 18748 5846
rect 18696 5782 18748 5788
rect 18708 5370 18736 5782
rect 19430 5672 19486 5681
rect 19430 5607 19486 5616
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19352 5370 19380 5510
rect 18696 5364 18748 5370
rect 18696 5306 18748 5312
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 18880 5228 18932 5234
rect 18880 5170 18932 5176
rect 18512 5024 18564 5030
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17498 3224 17554 3233
rect 17498 3159 17500 3168
rect 17552 3159 17554 3168
rect 17500 3130 17552 3136
rect 17512 2854 17540 3130
rect 18064 2990 18092 3878
rect 18156 3534 18184 4966
rect 18248 4950 18368 4978
rect 18512 4966 18564 4972
rect 18696 5024 18748 5030
rect 18696 4966 18748 4972
rect 18234 4856 18290 4865
rect 18234 4791 18290 4800
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 18052 2984 18104 2990
rect 18052 2926 18104 2932
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17408 2644 17460 2650
rect 17408 2586 17460 2592
rect 18064 2514 18092 2926
rect 18248 2922 18276 4791
rect 18236 2916 18288 2922
rect 18236 2858 18288 2864
rect 18052 2508 18104 2514
rect 18052 2450 18104 2456
rect 18340 480 18368 4950
rect 18708 4622 18736 4966
rect 18420 4616 18472 4622
rect 18696 4616 18748 4622
rect 18420 4558 18472 4564
rect 18694 4584 18696 4593
rect 18748 4584 18750 4593
rect 18432 4282 18460 4558
rect 18694 4519 18750 4528
rect 18420 4276 18472 4282
rect 18420 4218 18472 4224
rect 18892 4078 18920 5170
rect 19352 4865 19380 5306
rect 19338 4856 19394 4865
rect 19444 4826 19472 5607
rect 20180 5370 20208 8298
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20272 6866 20300 7142
rect 20260 6860 20312 6866
rect 20260 6802 20312 6808
rect 20272 6322 20300 6802
rect 20548 6746 20576 8366
rect 20628 8084 20680 8090
rect 20732 8072 20760 8774
rect 20680 8044 20760 8072
rect 20628 8026 20680 8032
rect 20720 6792 20772 6798
rect 20548 6740 20720 6746
rect 20548 6734 20772 6740
rect 20548 6718 20760 6734
rect 20260 6316 20312 6322
rect 20260 6258 20312 6264
rect 20272 5914 20300 6258
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 20626 5400 20682 5409
rect 20168 5364 20220 5370
rect 20824 5370 20852 9454
rect 21100 9178 21128 9862
rect 21284 9722 21312 10066
rect 21548 9920 21600 9926
rect 21548 9862 21600 9868
rect 21272 9716 21324 9722
rect 21272 9658 21324 9664
rect 21560 9625 21588 9862
rect 21546 9616 21602 9625
rect 21546 9551 21602 9560
rect 21560 9518 21588 9551
rect 21548 9512 21600 9518
rect 21548 9454 21600 9460
rect 21744 9364 21772 11834
rect 21928 11694 21956 12951
rect 22204 12714 22232 13330
rect 23296 13184 23348 13190
rect 23296 13126 23348 13132
rect 22468 12776 22520 12782
rect 22468 12718 22520 12724
rect 22192 12708 22244 12714
rect 22192 12650 22244 12656
rect 22480 12306 22508 12718
rect 23308 12374 23336 13126
rect 25700 13025 25728 13738
rect 26528 13394 26556 15098
rect 26698 15056 26754 15065
rect 26698 14991 26754 15000
rect 26712 14074 26740 14991
rect 26976 14272 27028 14278
rect 26976 14214 27028 14220
rect 26700 14068 26752 14074
rect 26700 14010 26752 14016
rect 26712 13802 26740 14010
rect 26988 13870 27016 14214
rect 27436 13932 27488 13938
rect 27436 13874 27488 13880
rect 26976 13864 27028 13870
rect 26976 13806 27028 13812
rect 26700 13796 26752 13802
rect 26700 13738 26752 13744
rect 26712 13462 26740 13738
rect 26884 13728 26936 13734
rect 26884 13670 26936 13676
rect 26896 13569 26924 13670
rect 26882 13560 26938 13569
rect 26988 13530 27016 13806
rect 26882 13495 26938 13504
rect 26976 13524 27028 13530
rect 26976 13466 27028 13472
rect 26700 13456 26752 13462
rect 26700 13398 26752 13404
rect 26516 13388 26568 13394
rect 26516 13330 26568 13336
rect 25686 13016 25742 13025
rect 26528 12986 26556 13330
rect 25686 12951 25688 12960
rect 25740 12951 25742 12960
rect 26516 12980 26568 12986
rect 25688 12922 25740 12928
rect 26516 12922 26568 12928
rect 26608 12844 26660 12850
rect 26608 12786 26660 12792
rect 24400 12708 24452 12714
rect 24400 12650 24452 12656
rect 24412 12617 24440 12650
rect 24398 12608 24454 12617
rect 24398 12543 24454 12552
rect 26620 12442 26648 12786
rect 26608 12436 26660 12442
rect 26608 12378 26660 12384
rect 22652 12368 22704 12374
rect 22652 12310 22704 12316
rect 23296 12368 23348 12374
rect 23296 12310 23348 12316
rect 22468 12300 22520 12306
rect 22468 12242 22520 12248
rect 22192 12096 22244 12102
rect 22192 12038 22244 12044
rect 21916 11688 21968 11694
rect 21916 11630 21968 11636
rect 22204 11558 22232 12038
rect 22480 11898 22508 12242
rect 22560 12096 22612 12102
rect 22560 12038 22612 12044
rect 22468 11892 22520 11898
rect 22468 11834 22520 11840
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 22192 11552 22244 11558
rect 22192 11494 22244 11500
rect 22020 11286 22048 11494
rect 22008 11280 22060 11286
rect 22008 11222 22060 11228
rect 22480 10810 22508 11834
rect 22572 11762 22600 12038
rect 22560 11756 22612 11762
rect 22560 11698 22612 11704
rect 22572 11082 22600 11698
rect 22664 11354 22692 12310
rect 26620 12238 26648 12378
rect 26712 12374 26740 13398
rect 26988 12714 27016 13466
rect 27448 12889 27476 13874
rect 27434 12880 27490 12889
rect 27434 12815 27490 12824
rect 26976 12708 27028 12714
rect 26976 12650 27028 12656
rect 26988 12442 27016 12650
rect 27620 12640 27672 12646
rect 27540 12588 27620 12594
rect 27540 12582 27672 12588
rect 27540 12566 27660 12582
rect 26976 12436 27028 12442
rect 26976 12378 27028 12384
rect 26700 12368 26752 12374
rect 26700 12310 26752 12316
rect 26608 12232 26660 12238
rect 26608 12174 26660 12180
rect 23940 12096 23992 12102
rect 23940 12038 23992 12044
rect 23952 11694 23980 12038
rect 26620 11898 26648 12174
rect 26608 11892 26660 11898
rect 26608 11834 26660 11840
rect 23940 11688 23992 11694
rect 23940 11630 23992 11636
rect 22744 11552 22796 11558
rect 22744 11494 22796 11500
rect 22652 11348 22704 11354
rect 22652 11290 22704 11296
rect 22756 11286 22784 11494
rect 23952 11354 23980 11630
rect 27540 11626 27568 12566
rect 27724 12345 27752 16934
rect 27816 15201 27844 19207
rect 27908 18902 27936 19450
rect 27896 18896 27948 18902
rect 27896 18838 27948 18844
rect 28552 17746 28580 22052
rect 29196 21962 29224 22510
rect 29288 22098 29316 23598
rect 29734 23559 29736 23568
rect 29788 23559 29790 23568
rect 29736 23530 29788 23536
rect 29748 23322 29776 23530
rect 29932 23322 29960 23666
rect 30012 23656 30064 23662
rect 30012 23598 30064 23604
rect 29736 23316 29788 23322
rect 29736 23258 29788 23264
rect 29920 23316 29972 23322
rect 29920 23258 29972 23264
rect 29736 23044 29788 23050
rect 29736 22986 29788 22992
rect 29748 22642 29776 22986
rect 29736 22636 29788 22642
rect 29736 22578 29788 22584
rect 29748 22234 29776 22578
rect 30024 22574 30052 23598
rect 30012 22568 30064 22574
rect 30012 22510 30064 22516
rect 29736 22228 29788 22234
rect 29736 22170 29788 22176
rect 30208 22098 30236 25434
rect 30392 25430 30420 26454
rect 30470 26344 30526 26353
rect 30470 26279 30526 26288
rect 30380 25424 30432 25430
rect 30380 25366 30432 25372
rect 30380 24676 30432 24682
rect 30380 24618 30432 24624
rect 30392 24562 30420 24618
rect 30300 24534 30420 24562
rect 30300 23322 30328 24534
rect 30484 24138 30512 26279
rect 30852 25770 30880 26726
rect 31956 26586 31984 27474
rect 32140 26761 32168 27814
rect 32772 27464 32824 27470
rect 32772 27406 32824 27412
rect 32312 27328 32364 27334
rect 32312 27270 32364 27276
rect 32126 26752 32182 26761
rect 32126 26687 32182 26696
rect 31944 26580 31996 26586
rect 31944 26522 31996 26528
rect 32324 26489 32352 27270
rect 32784 27062 32812 27406
rect 32772 27056 32824 27062
rect 32772 26998 32824 27004
rect 32864 26852 32916 26858
rect 32864 26794 32916 26800
rect 32876 26518 32904 26794
rect 32864 26512 32916 26518
rect 32310 26480 32366 26489
rect 32864 26454 32916 26460
rect 33060 26450 33088 28070
rect 33140 28018 33192 28024
rect 33244 28014 33272 28902
rect 33232 28008 33284 28014
rect 33232 27950 33284 27956
rect 33244 27674 33272 27950
rect 33232 27668 33284 27674
rect 33232 27610 33284 27616
rect 33140 27532 33192 27538
rect 33140 27474 33192 27480
rect 33152 27130 33180 27474
rect 33336 27418 33364 31078
rect 34152 30592 34204 30598
rect 34152 30534 34204 30540
rect 33784 30252 33836 30258
rect 33784 30194 33836 30200
rect 33416 30048 33468 30054
rect 33416 29990 33468 29996
rect 33600 30048 33652 30054
rect 33600 29990 33652 29996
rect 33428 28082 33456 29990
rect 33612 29782 33640 29990
rect 33600 29776 33652 29782
rect 33600 29718 33652 29724
rect 33600 29504 33652 29510
rect 33600 29446 33652 29452
rect 33612 29209 33640 29446
rect 33598 29200 33654 29209
rect 33796 29170 33824 30194
rect 34164 29170 34192 30534
rect 34336 30252 34388 30258
rect 34336 30194 34388 30200
rect 34244 30048 34296 30054
rect 34244 29990 34296 29996
rect 34256 29510 34284 29990
rect 34244 29504 34296 29510
rect 34244 29446 34296 29452
rect 33598 29135 33654 29144
rect 33784 29164 33836 29170
rect 33612 29102 33640 29135
rect 33784 29106 33836 29112
rect 34152 29164 34204 29170
rect 34152 29106 34204 29112
rect 33600 29096 33652 29102
rect 33600 29038 33652 29044
rect 33416 28076 33468 28082
rect 33416 28018 33468 28024
rect 33612 27606 33640 29038
rect 34256 28626 34284 29446
rect 34244 28620 34296 28626
rect 34244 28562 34296 28568
rect 34256 28218 34284 28562
rect 34244 28212 34296 28218
rect 34244 28154 34296 28160
rect 34348 28082 34376 30194
rect 34440 29730 34468 31282
rect 34612 30592 34664 30598
rect 34612 30534 34664 30540
rect 34518 30424 34574 30433
rect 34624 30394 34652 30534
rect 34518 30359 34574 30368
rect 34612 30388 34664 30394
rect 34532 29850 34560 30359
rect 34612 30330 34664 30336
rect 34716 30326 34744 32166
rect 34704 30320 34756 30326
rect 34704 30262 34756 30268
rect 34520 29844 34572 29850
rect 34520 29786 34572 29792
rect 34702 29744 34758 29753
rect 34440 29714 34560 29730
rect 34440 29708 34572 29714
rect 34440 29702 34520 29708
rect 34702 29679 34758 29688
rect 34520 29650 34572 29656
rect 34612 29640 34664 29646
rect 34612 29582 34664 29588
rect 34520 29028 34572 29034
rect 34520 28970 34572 28976
rect 34532 28762 34560 28970
rect 34520 28756 34572 28762
rect 34520 28698 34572 28704
rect 34336 28076 34388 28082
rect 34336 28018 34388 28024
rect 34624 27962 34652 29582
rect 34532 27934 34652 27962
rect 34532 27690 34560 27934
rect 34612 27872 34664 27878
rect 34612 27814 34664 27820
rect 34348 27662 34560 27690
rect 33600 27600 33652 27606
rect 33600 27542 33652 27548
rect 33244 27402 33364 27418
rect 33232 27396 33364 27402
rect 33284 27390 33364 27396
rect 33232 27338 33284 27344
rect 33140 27124 33192 27130
rect 33140 27066 33192 27072
rect 33244 26926 33272 27338
rect 33324 27328 33376 27334
rect 33324 27270 33376 27276
rect 33232 26920 33284 26926
rect 33232 26862 33284 26868
rect 32310 26415 32366 26424
rect 33048 26444 33100 26450
rect 33048 26386 33100 26392
rect 33060 26058 33088 26386
rect 32968 26042 33180 26058
rect 32956 26036 33180 26042
rect 33008 26030 33180 26036
rect 32956 25978 33008 25984
rect 33048 25968 33100 25974
rect 30930 25936 30986 25945
rect 33048 25910 33100 25916
rect 30930 25871 30986 25880
rect 30840 25764 30892 25770
rect 30840 25706 30892 25712
rect 30852 25498 30880 25706
rect 30840 25492 30892 25498
rect 30840 25434 30892 25440
rect 30654 24712 30710 24721
rect 30654 24647 30710 24656
rect 30668 24274 30696 24647
rect 30852 24410 30880 25434
rect 30944 25362 30972 25871
rect 31300 25696 31352 25702
rect 31300 25638 31352 25644
rect 32956 25696 33008 25702
rect 32956 25638 33008 25644
rect 30932 25356 30984 25362
rect 30932 25298 30984 25304
rect 30944 24954 30972 25298
rect 30932 24948 30984 24954
rect 30932 24890 30984 24896
rect 31312 24886 31340 25638
rect 32968 25498 32996 25638
rect 32956 25492 33008 25498
rect 32956 25434 33008 25440
rect 31760 25152 31812 25158
rect 31760 25094 31812 25100
rect 31300 24880 31352 24886
rect 31300 24822 31352 24828
rect 31312 24410 31340 24822
rect 31772 24818 31800 25094
rect 31760 24812 31812 24818
rect 31760 24754 31812 24760
rect 31760 24608 31812 24614
rect 31760 24550 31812 24556
rect 30840 24404 30892 24410
rect 30840 24346 30892 24352
rect 31300 24404 31352 24410
rect 31300 24346 31352 24352
rect 30656 24268 30708 24274
rect 30656 24210 30708 24216
rect 30472 24132 30524 24138
rect 30472 24074 30524 24080
rect 30668 23866 30696 24210
rect 30656 23860 30708 23866
rect 30656 23802 30708 23808
rect 31312 23662 31340 24346
rect 31300 23656 31352 23662
rect 31300 23598 31352 23604
rect 31312 23322 31340 23598
rect 30288 23316 30340 23322
rect 30288 23258 30340 23264
rect 31300 23316 31352 23322
rect 31300 23258 31352 23264
rect 30380 22432 30432 22438
rect 30380 22374 30432 22380
rect 29276 22092 29328 22098
rect 30196 22092 30248 22098
rect 29276 22034 29328 22040
rect 30116 22052 30196 22080
rect 29184 21956 29236 21962
rect 29184 21898 29236 21904
rect 29288 21729 29316 22034
rect 29274 21720 29330 21729
rect 30116 21690 30144 22052
rect 30196 22034 30248 22040
rect 30196 21888 30248 21894
rect 30196 21830 30248 21836
rect 29274 21655 29330 21664
rect 30104 21684 30156 21690
rect 30104 21626 30156 21632
rect 29828 20936 29880 20942
rect 29828 20878 29880 20884
rect 29460 20324 29512 20330
rect 29460 20266 29512 20272
rect 29472 20058 29500 20266
rect 29840 20058 29868 20878
rect 30208 20777 30236 21830
rect 30392 21690 30420 22374
rect 31772 22234 31800 24550
rect 33060 23633 33088 25910
rect 33152 25362 33180 26030
rect 33336 25838 33364 27270
rect 33612 27130 33640 27542
rect 33600 27124 33652 27130
rect 33600 27066 33652 27072
rect 33876 26988 33928 26994
rect 33876 26930 33928 26936
rect 33888 26897 33916 26930
rect 33874 26888 33930 26897
rect 34348 26858 34376 27662
rect 34428 27328 34480 27334
rect 34428 27270 34480 27276
rect 34440 27033 34468 27270
rect 34520 27056 34572 27062
rect 34426 27024 34482 27033
rect 34520 26998 34572 27004
rect 34426 26959 34482 26968
rect 33874 26823 33930 26832
rect 34336 26852 34388 26858
rect 33888 26586 33916 26823
rect 34336 26794 34388 26800
rect 33876 26580 33928 26586
rect 33876 26522 33928 26528
rect 34348 26330 34376 26794
rect 34440 26518 34468 26959
rect 34428 26512 34480 26518
rect 34428 26454 34480 26460
rect 34256 26302 34376 26330
rect 33508 25900 33560 25906
rect 33508 25842 33560 25848
rect 33324 25832 33376 25838
rect 33324 25774 33376 25780
rect 33520 25430 33548 25842
rect 33508 25424 33560 25430
rect 33508 25366 33560 25372
rect 33140 25356 33192 25362
rect 33140 25298 33192 25304
rect 33152 24954 33180 25298
rect 33520 24954 33548 25366
rect 33140 24948 33192 24954
rect 33140 24890 33192 24896
rect 33508 24948 33560 24954
rect 33508 24890 33560 24896
rect 33152 24206 33180 24890
rect 34256 24818 34284 26302
rect 34336 26240 34388 26246
rect 34336 26182 34388 26188
rect 34348 25906 34376 26182
rect 34440 26042 34468 26454
rect 34532 26042 34560 26998
rect 34428 26036 34480 26042
rect 34428 25978 34480 25984
rect 34520 26036 34572 26042
rect 34520 25978 34572 25984
rect 34624 25922 34652 27814
rect 34716 27577 34744 29679
rect 34702 27568 34758 27577
rect 34702 27503 34758 27512
rect 34704 27464 34756 27470
rect 34704 27406 34756 27412
rect 34716 26042 34744 27406
rect 34704 26036 34756 26042
rect 34704 25978 34756 25984
rect 34336 25900 34388 25906
rect 34624 25894 34744 25922
rect 34336 25842 34388 25848
rect 34520 25152 34572 25158
rect 34520 25094 34572 25100
rect 34244 24812 34296 24818
rect 34244 24754 34296 24760
rect 34428 24744 34480 24750
rect 34428 24686 34480 24692
rect 34336 24676 34388 24682
rect 34336 24618 34388 24624
rect 33876 24268 33928 24274
rect 33876 24210 33928 24216
rect 33140 24200 33192 24206
rect 33140 24142 33192 24148
rect 33046 23624 33102 23633
rect 33152 23594 33180 24142
rect 33888 23594 33916 24210
rect 33968 24200 34020 24206
rect 33968 24142 34020 24148
rect 33980 23866 34008 24142
rect 33968 23860 34020 23866
rect 33968 23802 34020 23808
rect 33046 23559 33102 23568
rect 33140 23588 33192 23594
rect 31944 23520 31996 23526
rect 31944 23462 31996 23468
rect 33060 23474 33088 23559
rect 33140 23530 33192 23536
rect 33876 23588 33928 23594
rect 33876 23530 33928 23536
rect 31760 22228 31812 22234
rect 31760 22170 31812 22176
rect 31956 21962 31984 23462
rect 33060 23446 33180 23474
rect 33152 23254 33180 23446
rect 33140 23248 33192 23254
rect 33140 23190 33192 23196
rect 33692 23248 33744 23254
rect 33692 23190 33744 23196
rect 33704 22710 33732 23190
rect 33888 23118 33916 23530
rect 33784 23112 33836 23118
rect 33784 23054 33836 23060
rect 33876 23112 33928 23118
rect 33876 23054 33928 23060
rect 33692 22704 33744 22710
rect 33692 22646 33744 22652
rect 33140 22500 33192 22506
rect 33140 22442 33192 22448
rect 32404 22228 32456 22234
rect 32404 22170 32456 22176
rect 31944 21956 31996 21962
rect 31944 21898 31996 21904
rect 30656 21888 30708 21894
rect 30656 21830 30708 21836
rect 30748 21888 30800 21894
rect 30748 21830 30800 21836
rect 31668 21888 31720 21894
rect 32128 21888 32180 21894
rect 31758 21856 31814 21865
rect 31720 21836 31758 21842
rect 31668 21830 31758 21836
rect 30380 21684 30432 21690
rect 30380 21626 30432 21632
rect 30392 21350 30420 21626
rect 30668 21486 30696 21830
rect 30760 21554 30788 21830
rect 31680 21814 31758 21830
rect 32128 21830 32180 21836
rect 31758 21791 31814 21800
rect 30748 21548 30800 21554
rect 30748 21490 30800 21496
rect 31024 21548 31076 21554
rect 31024 21490 31076 21496
rect 30656 21480 30708 21486
rect 30656 21422 30708 21428
rect 30380 21344 30432 21350
rect 30380 21286 30432 21292
rect 31036 21146 31064 21490
rect 31300 21480 31352 21486
rect 31300 21422 31352 21428
rect 31312 21146 31340 21422
rect 31576 21344 31628 21350
rect 31576 21286 31628 21292
rect 31024 21140 31076 21146
rect 31024 21082 31076 21088
rect 31300 21140 31352 21146
rect 31300 21082 31352 21088
rect 30288 21004 30340 21010
rect 30288 20946 30340 20952
rect 30194 20768 30250 20777
rect 30194 20703 30250 20712
rect 30300 20058 30328 20946
rect 30748 20936 30800 20942
rect 30748 20878 30800 20884
rect 30380 20800 30432 20806
rect 30380 20742 30432 20748
rect 30392 20330 30420 20742
rect 30760 20641 30788 20878
rect 30746 20632 30802 20641
rect 31312 20602 31340 21082
rect 31588 20602 31616 21286
rect 31668 20936 31720 20942
rect 31668 20878 31720 20884
rect 30746 20567 30748 20576
rect 30800 20567 30802 20576
rect 31300 20596 31352 20602
rect 30748 20538 30800 20544
rect 31300 20538 31352 20544
rect 31576 20596 31628 20602
rect 31576 20538 31628 20544
rect 30380 20324 30432 20330
rect 30380 20266 30432 20272
rect 30760 20058 30788 20538
rect 31588 20330 31616 20538
rect 31576 20324 31628 20330
rect 31576 20266 31628 20272
rect 29460 20052 29512 20058
rect 29460 19994 29512 20000
rect 29828 20052 29880 20058
rect 29828 19994 29880 20000
rect 30288 20052 30340 20058
rect 30288 19994 30340 20000
rect 30748 20052 30800 20058
rect 30748 19994 30800 20000
rect 31116 18624 31168 18630
rect 31116 18566 31168 18572
rect 30564 18352 30616 18358
rect 30562 18320 30564 18329
rect 30616 18320 30618 18329
rect 31128 18290 31156 18566
rect 30562 18255 30618 18264
rect 31116 18284 31168 18290
rect 31116 18226 31168 18232
rect 30932 18148 30984 18154
rect 30932 18090 30984 18096
rect 30012 18080 30064 18086
rect 30012 18022 30064 18028
rect 28080 17740 28132 17746
rect 28000 17700 28080 17728
rect 28000 17270 28028 17700
rect 28080 17682 28132 17688
rect 28540 17740 28592 17746
rect 28540 17682 28592 17688
rect 28448 17672 28500 17678
rect 28448 17614 28500 17620
rect 27988 17264 28040 17270
rect 27988 17206 28040 17212
rect 28000 16998 28028 17206
rect 28460 17066 28488 17614
rect 28552 17338 28580 17682
rect 29828 17536 29880 17542
rect 29828 17478 29880 17484
rect 28540 17332 28592 17338
rect 28540 17274 28592 17280
rect 29736 17128 29788 17134
rect 29736 17070 29788 17076
rect 28448 17060 28500 17066
rect 28448 17002 28500 17008
rect 27988 16992 28040 16998
rect 27988 16934 28040 16940
rect 27894 16144 27950 16153
rect 27894 16079 27896 16088
rect 27948 16079 27950 16088
rect 27896 16050 27948 16056
rect 27908 15706 27936 16050
rect 27896 15700 27948 15706
rect 27896 15642 27948 15648
rect 27802 15192 27858 15201
rect 27802 15127 27858 15136
rect 27710 12336 27766 12345
rect 27710 12271 27766 12280
rect 27620 12232 27672 12238
rect 27620 12174 27672 12180
rect 26792 11620 26844 11626
rect 26792 11562 26844 11568
rect 27528 11620 27580 11626
rect 27528 11562 27580 11568
rect 25044 11552 25096 11558
rect 25044 11494 25096 11500
rect 23940 11348 23992 11354
rect 23940 11290 23992 11296
rect 25056 11286 25084 11494
rect 26804 11354 26832 11562
rect 27632 11354 27660 12174
rect 26792 11348 26844 11354
rect 26792 11290 26844 11296
rect 27620 11348 27672 11354
rect 27620 11290 27672 11296
rect 22744 11280 22796 11286
rect 22744 11222 22796 11228
rect 23204 11280 23256 11286
rect 23204 11222 23256 11228
rect 25044 11280 25096 11286
rect 25044 11222 25096 11228
rect 22560 11076 22612 11082
rect 22560 11018 22612 11024
rect 22468 10804 22520 10810
rect 22468 10746 22520 10752
rect 22572 10674 22600 11018
rect 23020 11008 23072 11014
rect 23020 10950 23072 10956
rect 23032 10674 23060 10950
rect 22560 10668 22612 10674
rect 22560 10610 22612 10616
rect 23020 10668 23072 10674
rect 23020 10610 23072 10616
rect 21916 10464 21968 10470
rect 21916 10406 21968 10412
rect 22376 10464 22428 10470
rect 22376 10406 22428 10412
rect 21928 9586 21956 10406
rect 22388 10198 22416 10406
rect 22376 10192 22428 10198
rect 22376 10134 22428 10140
rect 22008 10124 22060 10130
rect 22008 10066 22060 10072
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 21560 9336 21772 9364
rect 21088 9172 21140 9178
rect 21088 9114 21140 9120
rect 21100 8634 21128 9114
rect 21364 9036 21416 9042
rect 21364 8978 21416 8984
rect 21088 8628 21140 8634
rect 21088 8570 21140 8576
rect 21376 8566 21404 8978
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21364 8560 21416 8566
rect 21364 8502 21416 8508
rect 21468 8362 21496 8910
rect 21456 8356 21508 8362
rect 21456 8298 21508 8304
rect 21468 8090 21496 8298
rect 21456 8084 21508 8090
rect 21456 8026 21508 8032
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 21088 7744 21140 7750
rect 21088 7686 21140 7692
rect 21100 7449 21128 7686
rect 21086 7440 21142 7449
rect 21086 7375 21142 7384
rect 21100 6866 21128 7375
rect 21468 7342 21496 7822
rect 21456 7336 21508 7342
rect 21456 7278 21508 7284
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 21088 6860 21140 6866
rect 21088 6802 21140 6808
rect 20916 6186 20944 6802
rect 21100 6458 21128 6802
rect 21088 6452 21140 6458
rect 21088 6394 21140 6400
rect 21364 6248 21416 6254
rect 21364 6190 21416 6196
rect 20904 6180 20956 6186
rect 20904 6122 20956 6128
rect 21376 5914 21404 6190
rect 21456 6112 21508 6118
rect 21456 6054 21508 6060
rect 21364 5908 21416 5914
rect 21364 5850 21416 5856
rect 20904 5704 20956 5710
rect 20902 5672 20904 5681
rect 20956 5672 20958 5681
rect 20902 5607 20958 5616
rect 20168 5306 20220 5312
rect 20456 5344 20626 5352
rect 20456 5324 20628 5344
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 19338 4791 19394 4800
rect 19432 4820 19484 4826
rect 19432 4762 19484 4768
rect 19984 4820 20036 4826
rect 19984 4762 20036 4768
rect 19708 4616 19760 4622
rect 19708 4558 19760 4564
rect 19340 4548 19392 4554
rect 19340 4490 19392 4496
rect 19248 4480 19300 4486
rect 19248 4422 19300 4428
rect 18880 4072 18932 4078
rect 18880 4014 18932 4020
rect 19260 3097 19288 4422
rect 19352 3466 19380 4490
rect 19720 4457 19748 4558
rect 19706 4448 19762 4457
rect 19706 4383 19762 4392
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 19996 3738 20024 4762
rect 20352 4480 20404 4486
rect 20350 4448 20352 4457
rect 20404 4448 20406 4457
rect 20350 4383 20406 4392
rect 20364 4214 20392 4383
rect 20352 4208 20404 4214
rect 20352 4150 20404 4156
rect 19984 3732 20036 3738
rect 19984 3674 20036 3680
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 19340 3460 19392 3466
rect 19340 3402 19392 3408
rect 19246 3088 19302 3097
rect 19246 3023 19302 3032
rect 19352 2854 19380 3402
rect 19340 2848 19392 2854
rect 19260 2796 19340 2802
rect 19260 2790 19392 2796
rect 19260 2774 19380 2790
rect 19260 2582 19288 2774
rect 19248 2576 19300 2582
rect 19248 2518 19300 2524
rect 19444 480 19472 3606
rect 19984 3528 20036 3534
rect 19984 3470 20036 3476
rect 19996 3194 20024 3470
rect 20074 3224 20130 3233
rect 19984 3188 20036 3194
rect 20074 3159 20130 3168
rect 19984 3130 20036 3136
rect 20088 2854 20116 3159
rect 20456 2990 20484 5324
rect 20680 5335 20682 5344
rect 20812 5364 20864 5370
rect 20628 5306 20680 5312
rect 20812 5306 20864 5312
rect 20996 5364 21048 5370
rect 20996 5306 21048 5312
rect 20536 5160 20588 5166
rect 20720 5160 20772 5166
rect 20536 5102 20588 5108
rect 20640 5120 20720 5148
rect 20444 2984 20496 2990
rect 20444 2926 20496 2932
rect 20076 2848 20128 2854
rect 20076 2790 20128 2796
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 20548 480 20576 5102
rect 20640 3670 20668 5120
rect 20720 5102 20772 5108
rect 21008 4690 21036 5306
rect 20996 4684 21048 4690
rect 20996 4626 21048 4632
rect 21180 4684 21232 4690
rect 21180 4626 21232 4632
rect 21008 4078 21036 4626
rect 21192 4282 21220 4626
rect 21180 4276 21232 4282
rect 21180 4218 21232 4224
rect 21468 4078 21496 6054
rect 21560 5409 21588 9336
rect 21730 8392 21786 8401
rect 21730 8327 21786 8336
rect 21744 8022 21772 8327
rect 21732 8016 21784 8022
rect 21732 7958 21784 7964
rect 21744 7546 21772 7958
rect 21732 7540 21784 7546
rect 21732 7482 21784 7488
rect 21640 6180 21692 6186
rect 21640 6122 21692 6128
rect 21546 5400 21602 5409
rect 21546 5335 21602 5344
rect 21548 4140 21600 4146
rect 21548 4082 21600 4088
rect 20996 4072 21048 4078
rect 20996 4014 21048 4020
rect 21456 4072 21508 4078
rect 21456 4014 21508 4020
rect 20628 3664 20680 3670
rect 20628 3606 20680 3612
rect 20812 3596 20864 3602
rect 20812 3538 20864 3544
rect 20824 3482 20852 3538
rect 21008 3534 21036 4014
rect 21088 3936 21140 3942
rect 21088 3878 21140 3884
rect 20640 3454 20852 3482
rect 20996 3528 21048 3534
rect 20996 3470 21048 3476
rect 20640 2650 20668 3454
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 20732 2530 20760 2994
rect 20640 2514 20760 2530
rect 21008 2514 21036 3470
rect 21100 2689 21128 3878
rect 21468 3058 21496 4014
rect 21560 3602 21588 4082
rect 21548 3596 21600 3602
rect 21548 3538 21600 3544
rect 21456 3052 21508 3058
rect 21456 2994 21508 3000
rect 21086 2680 21142 2689
rect 21086 2615 21142 2624
rect 20628 2508 20760 2514
rect 20680 2502 20760 2508
rect 20996 2508 21048 2514
rect 20628 2450 20680 2456
rect 20996 2450 21048 2456
rect 21652 480 21680 6122
rect 22020 5896 22048 10066
rect 22572 9926 22600 10610
rect 23216 10266 23244 11222
rect 23480 11144 23532 11150
rect 23480 11086 23532 11092
rect 23492 10810 23520 11086
rect 24860 11076 24912 11082
rect 24860 11018 24912 11024
rect 23480 10804 23532 10810
rect 23480 10746 23532 10752
rect 23492 10606 23520 10746
rect 24872 10690 24900 11018
rect 24780 10662 24900 10690
rect 24780 10606 24808 10662
rect 23480 10600 23532 10606
rect 23480 10542 23532 10548
rect 24768 10600 24820 10606
rect 24768 10542 24820 10548
rect 25044 10464 25096 10470
rect 25044 10406 25096 10412
rect 23204 10260 23256 10266
rect 23204 10202 23256 10208
rect 25056 10198 25084 10406
rect 23020 10192 23072 10198
rect 23020 10134 23072 10140
rect 25044 10192 25096 10198
rect 25044 10134 25096 10140
rect 22560 9920 22612 9926
rect 22560 9862 22612 9868
rect 23032 9722 23060 10134
rect 28000 10130 28028 16934
rect 29366 16824 29422 16833
rect 29366 16759 29368 16768
rect 29420 16759 29422 16768
rect 29368 16730 29420 16736
rect 29380 16046 29408 16730
rect 29550 16688 29606 16697
rect 29550 16623 29552 16632
rect 29604 16623 29606 16632
rect 29552 16594 29604 16600
rect 29368 16040 29420 16046
rect 29368 15982 29420 15988
rect 29092 14476 29144 14482
rect 29092 14418 29144 14424
rect 29104 14074 29132 14418
rect 29552 14272 29604 14278
rect 29552 14214 29604 14220
rect 29092 14068 29144 14074
rect 29092 14010 29144 14016
rect 29564 14006 29592 14214
rect 29552 14000 29604 14006
rect 29748 13977 29776 17070
rect 29840 17066 29868 17478
rect 29828 17060 29880 17066
rect 29828 17002 29880 17008
rect 29840 16114 29868 17002
rect 29920 16720 29972 16726
rect 29920 16662 29972 16668
rect 29828 16108 29880 16114
rect 29828 16050 29880 16056
rect 29932 15434 29960 16662
rect 30024 16250 30052 18022
rect 30944 17882 30972 18090
rect 30932 17876 30984 17882
rect 30932 17818 30984 17824
rect 30288 17604 30340 17610
rect 30288 17546 30340 17552
rect 30300 17134 30328 17546
rect 30288 17128 30340 17134
rect 30288 17070 30340 17076
rect 31128 16794 31156 18226
rect 31484 18080 31536 18086
rect 31484 18022 31536 18028
rect 31496 17921 31524 18022
rect 31482 17912 31538 17921
rect 31482 17847 31538 17856
rect 31588 17490 31616 20266
rect 31680 20058 31708 20878
rect 31772 20398 31800 21791
rect 32140 21593 32168 21830
rect 32126 21584 32182 21593
rect 32126 21519 32182 21528
rect 32416 21010 32444 22170
rect 33152 22114 33180 22442
rect 33796 22438 33824 23054
rect 33888 22778 33916 23054
rect 33876 22772 33928 22778
rect 33876 22714 33928 22720
rect 34348 22658 34376 24618
rect 34440 23322 34468 24686
rect 34532 24274 34560 25094
rect 34612 24608 34664 24614
rect 34612 24550 34664 24556
rect 34520 24268 34572 24274
rect 34520 24210 34572 24216
rect 34624 23730 34652 24550
rect 34612 23724 34664 23730
rect 34612 23666 34664 23672
rect 34716 23610 34744 25894
rect 34624 23582 34744 23610
rect 34428 23316 34480 23322
rect 34428 23258 34480 23264
rect 34520 23180 34572 23186
rect 34520 23122 34572 23128
rect 34532 22778 34560 23122
rect 34520 22772 34572 22778
rect 34520 22714 34572 22720
rect 34348 22630 34560 22658
rect 34532 22506 34560 22630
rect 34520 22500 34572 22506
rect 34520 22442 34572 22448
rect 33784 22432 33836 22438
rect 33784 22374 33836 22380
rect 34152 22432 34204 22438
rect 34152 22374 34204 22380
rect 34164 22234 34192 22374
rect 34152 22228 34204 22234
rect 34152 22170 34204 22176
rect 33060 22086 33180 22114
rect 32588 22024 32640 22030
rect 32588 21966 32640 21972
rect 32680 22024 32732 22030
rect 32680 21966 32732 21972
rect 32600 21350 32628 21966
rect 32588 21344 32640 21350
rect 32588 21286 32640 21292
rect 32600 21078 32628 21286
rect 32588 21072 32640 21078
rect 32588 21014 32640 21020
rect 32404 21004 32456 21010
rect 32404 20946 32456 20952
rect 31850 20768 31906 20777
rect 31850 20703 31906 20712
rect 31864 20534 31892 20703
rect 31852 20528 31904 20534
rect 31852 20470 31904 20476
rect 31760 20392 31812 20398
rect 31760 20334 31812 20340
rect 31668 20052 31720 20058
rect 31668 19994 31720 20000
rect 31772 19514 31800 20334
rect 31864 20058 31892 20470
rect 32600 20466 32628 21014
rect 32588 20460 32640 20466
rect 32588 20402 32640 20408
rect 32692 20346 32720 21966
rect 33060 21146 33088 22086
rect 34336 22024 34388 22030
rect 34336 21966 34388 21972
rect 34520 22024 34572 22030
rect 34520 21966 34572 21972
rect 34348 21865 34376 21966
rect 34334 21856 34390 21865
rect 34334 21791 34390 21800
rect 33324 21344 33376 21350
rect 33324 21286 33376 21292
rect 33048 21140 33100 21146
rect 33048 21082 33100 21088
rect 33336 21010 33364 21286
rect 34348 21146 34376 21791
rect 34532 21486 34560 21966
rect 34520 21480 34572 21486
rect 34520 21422 34572 21428
rect 34624 21162 34652 23582
rect 34704 22976 34756 22982
rect 34704 22918 34756 22924
rect 34336 21140 34388 21146
rect 34336 21082 34388 21088
rect 34532 21134 34652 21162
rect 33324 21004 33376 21010
rect 33324 20946 33376 20952
rect 32772 20936 32824 20942
rect 32772 20878 32824 20884
rect 32784 20806 32812 20878
rect 32772 20800 32824 20806
rect 32772 20742 32824 20748
rect 34336 20800 34388 20806
rect 34336 20742 34388 20748
rect 32784 20505 32812 20742
rect 32770 20496 32826 20505
rect 32770 20431 32826 20440
rect 32600 20318 32720 20346
rect 31852 20052 31904 20058
rect 31852 19994 31904 20000
rect 32600 19922 32628 20318
rect 34348 20262 34376 20742
rect 33692 20256 33744 20262
rect 33692 20198 33744 20204
rect 34336 20256 34388 20262
rect 34336 20198 34388 20204
rect 33232 20052 33284 20058
rect 33232 19994 33284 20000
rect 32588 19916 32640 19922
rect 32588 19858 32640 19864
rect 32312 19848 32364 19854
rect 32312 19790 32364 19796
rect 32126 19544 32182 19553
rect 31760 19508 31812 19514
rect 32126 19479 32182 19488
rect 31760 19450 31812 19456
rect 31772 17898 31800 19450
rect 31944 19168 31996 19174
rect 31944 19110 31996 19116
rect 31680 17870 31800 17898
rect 31956 17898 31984 19110
rect 32036 18760 32088 18766
rect 32036 18702 32088 18708
rect 32048 18426 32076 18702
rect 32036 18420 32088 18426
rect 32036 18362 32088 18368
rect 31956 17870 32076 17898
rect 31680 17610 31708 17870
rect 32048 17678 32076 17870
rect 32036 17672 32088 17678
rect 32036 17614 32088 17620
rect 31668 17604 31720 17610
rect 31668 17546 31720 17552
rect 31588 17462 31708 17490
rect 31680 17134 31708 17462
rect 32048 17218 32076 17614
rect 32140 17338 32168 19479
rect 32324 19174 32352 19790
rect 32600 19514 32628 19858
rect 32588 19508 32640 19514
rect 32588 19450 32640 19456
rect 33140 19304 33192 19310
rect 33138 19272 33140 19281
rect 33192 19272 33194 19281
rect 33138 19207 33194 19216
rect 32312 19168 32364 19174
rect 32312 19110 32364 19116
rect 33244 19122 33272 19994
rect 33704 19310 33732 20198
rect 34348 19854 34376 20198
rect 34336 19848 34388 19854
rect 34336 19790 34388 19796
rect 33876 19372 33928 19378
rect 33876 19314 33928 19320
rect 33692 19304 33744 19310
rect 33692 19246 33744 19252
rect 33324 19168 33376 19174
rect 33244 19116 33324 19122
rect 33244 19110 33376 19116
rect 33244 19094 33364 19110
rect 33244 18970 33272 19094
rect 33888 18970 33916 19314
rect 33232 18964 33284 18970
rect 33232 18906 33284 18912
rect 33876 18964 33928 18970
rect 33876 18906 33928 18912
rect 32680 18624 32732 18630
rect 32680 18566 32732 18572
rect 32692 18086 32720 18566
rect 32956 18284 33008 18290
rect 32956 18226 33008 18232
rect 32220 18080 32272 18086
rect 32218 18048 32220 18057
rect 32680 18080 32732 18086
rect 32272 18048 32274 18057
rect 32680 18022 32732 18028
rect 32218 17983 32274 17992
rect 32968 17882 32996 18226
rect 33048 18080 33100 18086
rect 33100 18040 33180 18068
rect 34532 18057 34560 21134
rect 34612 21072 34664 21078
rect 34612 21014 34664 21020
rect 34624 20602 34652 21014
rect 34612 20596 34664 20602
rect 34612 20538 34664 20544
rect 34624 20058 34652 20538
rect 34612 20052 34664 20058
rect 34612 19994 34664 20000
rect 34612 19848 34664 19854
rect 34612 19790 34664 19796
rect 34624 19514 34652 19790
rect 34612 19508 34664 19514
rect 34612 19450 34664 19456
rect 34716 19174 34744 22918
rect 34808 21350 34836 35430
rect 35544 35414 35940 35430
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 35348 33448 35400 33454
rect 35348 33390 35400 33396
rect 35360 33114 35388 33390
rect 35348 33108 35400 33114
rect 35348 33050 35400 33056
rect 35440 32972 35492 32978
rect 35440 32914 35492 32920
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 35452 32230 35480 32914
rect 35440 32224 35492 32230
rect 35346 32192 35402 32201
rect 35440 32166 35492 32172
rect 35346 32127 35402 32136
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 35360 31414 35388 32127
rect 35452 32026 35480 32166
rect 35440 32020 35492 32026
rect 35440 31962 35492 31968
rect 35348 31408 35400 31414
rect 35348 31350 35400 31356
rect 35544 31226 35572 35414
rect 35900 34944 35952 34950
rect 35900 34886 35952 34892
rect 35912 34218 35940 34886
rect 37568 34746 37596 36887
rect 37556 34740 37608 34746
rect 37556 34682 37608 34688
rect 37832 34536 37884 34542
rect 36818 34504 36874 34513
rect 37832 34478 37884 34484
rect 36818 34439 36874 34448
rect 35820 34190 35940 34218
rect 35820 34134 35848 34190
rect 35808 34128 35860 34134
rect 35808 34070 35860 34076
rect 35992 33856 36044 33862
rect 35992 33798 36044 33804
rect 36004 33454 36032 33798
rect 35992 33448 36044 33454
rect 35992 33390 36044 33396
rect 35808 32768 35860 32774
rect 35808 32710 35860 32716
rect 35624 32428 35676 32434
rect 35624 32370 35676 32376
rect 35636 31634 35664 32370
rect 35820 31890 35848 32710
rect 36004 32502 36032 33390
rect 36636 33312 36688 33318
rect 36636 33254 36688 33260
rect 36726 33280 36782 33289
rect 36648 32978 36676 33254
rect 36726 33215 36782 33224
rect 36636 32972 36688 32978
rect 36636 32914 36688 32920
rect 36648 32570 36676 32914
rect 36636 32564 36688 32570
rect 36636 32506 36688 32512
rect 35992 32496 36044 32502
rect 35992 32438 36044 32444
rect 35990 32056 36046 32065
rect 35900 32020 35952 32026
rect 35990 31991 36046 32000
rect 35900 31962 35952 31968
rect 35808 31884 35860 31890
rect 35808 31826 35860 31832
rect 35636 31606 35756 31634
rect 35624 31408 35676 31414
rect 35624 31350 35676 31356
rect 35360 31198 35572 31226
rect 35256 31136 35308 31142
rect 35256 31078 35308 31084
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 35164 30320 35216 30326
rect 35164 30262 35216 30268
rect 35176 30122 35204 30262
rect 35268 30190 35296 31078
rect 35256 30184 35308 30190
rect 35256 30126 35308 30132
rect 35164 30116 35216 30122
rect 35164 30058 35216 30064
rect 35360 30002 35388 31198
rect 35440 31136 35492 31142
rect 35440 31078 35492 31084
rect 35452 30802 35480 31078
rect 35530 30832 35586 30841
rect 35440 30796 35492 30802
rect 35530 30767 35586 30776
rect 35440 30738 35492 30744
rect 35360 29974 35480 30002
rect 35348 29844 35400 29850
rect 35348 29786 35400 29792
rect 35256 29504 35308 29510
rect 35256 29446 35308 29452
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 34980 29096 35032 29102
rect 34980 29038 35032 29044
rect 34992 28506 35020 29038
rect 35268 29034 35296 29446
rect 35256 29028 35308 29034
rect 35256 28970 35308 28976
rect 35360 28762 35388 29786
rect 35348 28756 35400 28762
rect 35348 28698 35400 28704
rect 34992 28478 35296 28506
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 35268 27538 35296 28478
rect 35256 27532 35308 27538
rect 35256 27474 35308 27480
rect 35346 27296 35402 27305
rect 35268 27254 35346 27282
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 35268 24721 35296 27254
rect 35346 27231 35402 27240
rect 35452 25242 35480 29974
rect 35544 28218 35572 30767
rect 35636 29186 35664 31350
rect 35728 31346 35756 31606
rect 35716 31340 35768 31346
rect 35716 31282 35768 31288
rect 35820 31278 35848 31826
rect 35808 31272 35860 31278
rect 35808 31214 35860 31220
rect 35912 31142 35940 31962
rect 35900 31136 35952 31142
rect 35900 31078 35952 31084
rect 36004 30938 36032 31991
rect 36084 31340 36136 31346
rect 36084 31282 36136 31288
rect 36096 31142 36124 31282
rect 36084 31136 36136 31142
rect 36084 31078 36136 31084
rect 35992 30932 36044 30938
rect 35992 30874 36044 30880
rect 35808 30796 35860 30802
rect 35808 30738 35860 30744
rect 35820 30274 35848 30738
rect 35992 30592 36044 30598
rect 35992 30534 36044 30540
rect 36004 30394 36032 30534
rect 35992 30388 36044 30394
rect 35992 30330 36044 30336
rect 35820 30246 35940 30274
rect 35912 30054 35940 30246
rect 35900 30048 35952 30054
rect 35900 29990 35952 29996
rect 35716 29708 35768 29714
rect 35716 29650 35768 29656
rect 35728 29617 35756 29650
rect 35714 29608 35770 29617
rect 35770 29566 35848 29594
rect 35714 29543 35770 29552
rect 35820 29306 35848 29566
rect 35808 29300 35860 29306
rect 35808 29242 35860 29248
rect 35636 29158 35756 29186
rect 35622 29064 35678 29073
rect 35622 28999 35678 29008
rect 35532 28212 35584 28218
rect 35532 28154 35584 28160
rect 35532 27600 35584 27606
rect 35532 27542 35584 27548
rect 35544 26926 35572 27542
rect 35532 26920 35584 26926
rect 35532 26862 35584 26868
rect 35544 26586 35572 26862
rect 35532 26580 35584 26586
rect 35532 26522 35584 26528
rect 35532 26444 35584 26450
rect 35532 26386 35584 26392
rect 35544 25702 35572 26386
rect 35532 25696 35584 25702
rect 35532 25638 35584 25644
rect 35360 25214 35480 25242
rect 35254 24712 35310 24721
rect 35254 24647 35310 24656
rect 34888 24608 34940 24614
rect 34886 24576 34888 24585
rect 34940 24576 34942 24585
rect 34886 24511 34942 24520
rect 35254 24576 35310 24585
rect 35254 24511 35310 24520
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 34980 23792 35032 23798
rect 34980 23734 35032 23740
rect 34992 23186 35020 23734
rect 34980 23180 35032 23186
rect 34980 23122 35032 23128
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 34888 22500 34940 22506
rect 34888 22442 34940 22448
rect 34900 22030 34928 22442
rect 34888 22024 34940 22030
rect 34888 21966 34940 21972
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 34796 21344 34848 21350
rect 34796 21286 34848 21292
rect 34704 19168 34756 19174
rect 34704 19110 34756 19116
rect 33048 18022 33100 18028
rect 32956 17876 33008 17882
rect 32956 17818 33008 17824
rect 32312 17808 32364 17814
rect 32312 17750 32364 17756
rect 32128 17332 32180 17338
rect 32128 17274 32180 17280
rect 32048 17190 32168 17218
rect 31668 17128 31720 17134
rect 31668 17070 31720 17076
rect 32140 16998 32168 17190
rect 32220 17128 32272 17134
rect 32220 17070 32272 17076
rect 32128 16992 32180 16998
rect 32128 16934 32180 16940
rect 31116 16788 31168 16794
rect 31116 16730 31168 16736
rect 30288 16720 30340 16726
rect 30288 16662 30340 16668
rect 30012 16244 30064 16250
rect 30012 16186 30064 16192
rect 30300 16114 30328 16662
rect 30380 16652 30432 16658
rect 30380 16594 30432 16600
rect 30392 16250 30420 16594
rect 30932 16584 30984 16590
rect 30932 16526 30984 16532
rect 30380 16244 30432 16250
rect 30380 16186 30432 16192
rect 30944 16114 30972 16526
rect 30288 16108 30340 16114
rect 30288 16050 30340 16056
rect 30932 16108 30984 16114
rect 30932 16050 30984 16056
rect 30196 16040 30248 16046
rect 30196 15982 30248 15988
rect 29920 15428 29972 15434
rect 29920 15370 29972 15376
rect 29932 15162 29960 15370
rect 30208 15366 30236 15982
rect 30300 15706 30328 16050
rect 30288 15700 30340 15706
rect 30288 15642 30340 15648
rect 30564 15564 30616 15570
rect 30564 15506 30616 15512
rect 30196 15360 30248 15366
rect 30196 15302 30248 15308
rect 30576 15162 30604 15506
rect 30656 15496 30708 15502
rect 30656 15438 30708 15444
rect 29920 15156 29972 15162
rect 29920 15098 29972 15104
rect 30564 15156 30616 15162
rect 30564 15098 30616 15104
rect 30668 14890 30696 15438
rect 30944 15162 30972 16050
rect 31128 15978 31156 16730
rect 32140 16658 32168 16934
rect 32128 16652 32180 16658
rect 32128 16594 32180 16600
rect 32232 16130 32260 17070
rect 32324 16794 32352 17750
rect 33152 17338 33180 18040
rect 34518 18048 34574 18057
rect 34518 17983 34574 17992
rect 33140 17332 33192 17338
rect 33140 17274 33192 17280
rect 33416 17196 33468 17202
rect 33416 17138 33468 17144
rect 33876 17196 33928 17202
rect 33876 17138 33928 17144
rect 33048 16992 33100 16998
rect 33048 16934 33100 16940
rect 32312 16788 32364 16794
rect 32312 16730 32364 16736
rect 32324 16250 32352 16730
rect 32312 16244 32364 16250
rect 32312 16186 32364 16192
rect 32232 16102 32352 16130
rect 31116 15972 31168 15978
rect 31116 15914 31168 15920
rect 31666 15600 31722 15609
rect 31666 15535 31668 15544
rect 31720 15535 31722 15544
rect 32128 15564 32180 15570
rect 31668 15506 31720 15512
rect 32128 15506 32180 15512
rect 31392 15496 31444 15502
rect 31392 15438 31444 15444
rect 31404 15162 31432 15438
rect 30932 15156 30984 15162
rect 30932 15098 30984 15104
rect 31392 15156 31444 15162
rect 31392 15098 31444 15104
rect 31680 14958 31708 15506
rect 31760 15360 31812 15366
rect 31760 15302 31812 15308
rect 31668 14952 31720 14958
rect 31668 14894 31720 14900
rect 30656 14884 30708 14890
rect 30656 14826 30708 14832
rect 30472 14612 30524 14618
rect 30564 14612 30616 14618
rect 30524 14572 30564 14600
rect 30472 14554 30524 14560
rect 30564 14554 30616 14560
rect 30564 14408 30616 14414
rect 30564 14350 30616 14356
rect 30576 14074 30604 14350
rect 30668 14074 30696 14826
rect 30840 14476 30892 14482
rect 30840 14418 30892 14424
rect 30564 14068 30616 14074
rect 30564 14010 30616 14016
rect 30656 14068 30708 14074
rect 30656 14010 30708 14016
rect 29552 13942 29604 13948
rect 29734 13968 29790 13977
rect 29734 13903 29790 13912
rect 29000 13864 29052 13870
rect 29000 13806 29052 13812
rect 29012 13530 29040 13806
rect 29458 13560 29514 13569
rect 29000 13524 29052 13530
rect 29458 13495 29460 13504
rect 29000 13466 29052 13472
rect 29512 13495 29514 13504
rect 29460 13466 29512 13472
rect 29368 13388 29420 13394
rect 29368 13330 29420 13336
rect 29380 12918 29408 13330
rect 29368 12912 29420 12918
rect 29368 12854 29420 12860
rect 28724 12708 28776 12714
rect 28724 12650 28776 12656
rect 28736 12374 28764 12650
rect 29472 12442 29500 13466
rect 29460 12436 29512 12442
rect 29460 12378 29512 12384
rect 28080 12368 28132 12374
rect 28080 12310 28132 12316
rect 28724 12368 28776 12374
rect 28724 12310 28776 12316
rect 28092 11898 28120 12310
rect 28080 11892 28132 11898
rect 28080 11834 28132 11840
rect 28092 11354 28120 11834
rect 29552 11620 29604 11626
rect 29552 11562 29604 11568
rect 28172 11552 28224 11558
rect 28172 11494 28224 11500
rect 28080 11348 28132 11354
rect 28080 11290 28132 11296
rect 28184 11218 28212 11494
rect 29564 11354 29592 11562
rect 29552 11348 29604 11354
rect 29552 11290 29604 11296
rect 28632 11280 28684 11286
rect 28632 11222 28684 11228
rect 28172 11212 28224 11218
rect 28172 11154 28224 11160
rect 28184 10810 28212 11154
rect 28644 10810 28672 11222
rect 28172 10804 28224 10810
rect 28172 10746 28224 10752
rect 28632 10804 28684 10810
rect 28632 10746 28684 10752
rect 27988 10124 28040 10130
rect 27988 10066 28040 10072
rect 23296 10056 23348 10062
rect 23296 9998 23348 10004
rect 23204 9920 23256 9926
rect 23204 9862 23256 9868
rect 23020 9716 23072 9722
rect 23020 9658 23072 9664
rect 23216 9518 23244 9862
rect 23204 9512 23256 9518
rect 23204 9454 23256 9460
rect 23308 9382 23336 9998
rect 24676 9920 24728 9926
rect 24676 9862 24728 9868
rect 24688 9722 24716 9862
rect 24676 9716 24728 9722
rect 24676 9658 24728 9664
rect 23664 9648 23716 9654
rect 23662 9616 23664 9625
rect 23716 9616 23718 9625
rect 23662 9551 23718 9560
rect 24124 9580 24176 9586
rect 24124 9522 24176 9528
rect 22652 9376 22704 9382
rect 22652 9318 22704 9324
rect 23296 9376 23348 9382
rect 23296 9318 23348 9324
rect 24032 9376 24084 9382
rect 24032 9318 24084 9324
rect 22664 8974 22692 9318
rect 24044 9178 24072 9318
rect 24032 9172 24084 9178
rect 24032 9114 24084 9120
rect 23112 9104 23164 9110
rect 23112 9046 23164 9052
rect 22652 8968 22704 8974
rect 22652 8910 22704 8916
rect 22664 8294 22692 8910
rect 23124 8634 23152 9046
rect 23112 8628 23164 8634
rect 23112 8570 23164 8576
rect 24044 8401 24072 9114
rect 24136 9110 24164 9522
rect 28184 9178 28212 10746
rect 28172 9172 28224 9178
rect 28172 9114 28224 9120
rect 24124 9104 24176 9110
rect 24124 9046 24176 9052
rect 26608 9036 26660 9042
rect 26608 8978 26660 8984
rect 28080 9036 28132 9042
rect 28080 8978 28132 8984
rect 25504 8832 25556 8838
rect 25504 8774 25556 8780
rect 25516 8430 25544 8774
rect 26620 8634 26648 8978
rect 28092 8634 28120 8978
rect 28184 8634 28212 9114
rect 29368 8832 29420 8838
rect 29368 8774 29420 8780
rect 26608 8628 26660 8634
rect 26608 8570 26660 8576
rect 28080 8628 28132 8634
rect 28080 8570 28132 8576
rect 28172 8628 28224 8634
rect 28172 8570 28224 8576
rect 28724 8628 28776 8634
rect 28724 8570 28776 8576
rect 25596 8492 25648 8498
rect 25596 8434 25648 8440
rect 25504 8424 25556 8430
rect 24030 8392 24086 8401
rect 25504 8366 25556 8372
rect 24030 8327 24086 8336
rect 22652 8288 22704 8294
rect 22652 8230 22704 8236
rect 22928 8288 22980 8294
rect 22928 8230 22980 8236
rect 25136 8288 25188 8294
rect 25136 8230 25188 8236
rect 22940 7342 22968 8230
rect 23940 7880 23992 7886
rect 23940 7822 23992 7828
rect 23952 7342 23980 7822
rect 22928 7336 22980 7342
rect 22928 7278 22980 7284
rect 23940 7336 23992 7342
rect 23940 7278 23992 7284
rect 22100 6724 22152 6730
rect 22100 6666 22152 6672
rect 22112 5914 22140 6666
rect 22940 6118 22968 7278
rect 24216 7268 24268 7274
rect 24216 7210 24268 7216
rect 24228 6934 24256 7210
rect 24216 6928 24268 6934
rect 24216 6870 24268 6876
rect 24768 6928 24820 6934
rect 24768 6870 24820 6876
rect 24400 6860 24452 6866
rect 24400 6802 24452 6808
rect 23664 6656 23716 6662
rect 23664 6598 23716 6604
rect 23296 6248 23348 6254
rect 23296 6190 23348 6196
rect 23572 6248 23624 6254
rect 23572 6190 23624 6196
rect 22652 6112 22704 6118
rect 22652 6054 22704 6060
rect 22928 6112 22980 6118
rect 22928 6054 22980 6060
rect 21836 5868 22048 5896
rect 22100 5908 22152 5914
rect 21836 2938 21864 5868
rect 22100 5850 22152 5856
rect 21916 5772 21968 5778
rect 21916 5714 21968 5720
rect 21928 5098 21956 5714
rect 22112 5302 22140 5850
rect 22468 5568 22520 5574
rect 22468 5510 22520 5516
rect 22100 5296 22152 5302
rect 22100 5238 22152 5244
rect 22480 5234 22508 5510
rect 22468 5228 22520 5234
rect 22468 5170 22520 5176
rect 21916 5092 21968 5098
rect 21916 5034 21968 5040
rect 22008 5024 22060 5030
rect 22008 4966 22060 4972
rect 22020 4865 22048 4966
rect 22006 4856 22062 4865
rect 22480 4826 22508 5170
rect 22006 4791 22062 4800
rect 22468 4820 22520 4826
rect 22468 4762 22520 4768
rect 22190 4448 22246 4457
rect 22190 4383 22246 4392
rect 22100 3392 22152 3398
rect 22100 3334 22152 3340
rect 21836 2910 21956 2938
rect 21928 2854 21956 2910
rect 21916 2848 21968 2854
rect 21916 2790 21968 2796
rect 22008 2576 22060 2582
rect 22112 2530 22140 3334
rect 22204 2650 22232 4383
rect 22664 4321 22692 6054
rect 22940 5710 22968 6054
rect 23020 5840 23072 5846
rect 23020 5782 23072 5788
rect 22928 5704 22980 5710
rect 22928 5646 22980 5652
rect 22940 5370 22968 5646
rect 23032 5574 23060 5782
rect 23020 5568 23072 5574
rect 23020 5510 23072 5516
rect 22928 5364 22980 5370
rect 22928 5306 22980 5312
rect 23032 5166 23060 5510
rect 23020 5160 23072 5166
rect 23020 5102 23072 5108
rect 22744 5092 22796 5098
rect 22744 5034 22796 5040
rect 22650 4312 22706 4321
rect 22650 4247 22706 4256
rect 22376 3936 22428 3942
rect 22376 3878 22428 3884
rect 22388 2854 22416 3878
rect 22376 2848 22428 2854
rect 22374 2816 22376 2825
rect 22428 2816 22430 2825
rect 22374 2751 22430 2760
rect 22192 2644 22244 2650
rect 22192 2586 22244 2592
rect 22060 2524 22140 2530
rect 22008 2518 22140 2524
rect 22020 2502 22140 2518
rect 22756 480 22784 5034
rect 23032 4978 23060 5102
rect 23110 4992 23166 5001
rect 23032 4950 23110 4978
rect 23110 4927 23166 4936
rect 23124 4758 23152 4927
rect 23112 4752 23164 4758
rect 23112 4694 23164 4700
rect 22836 4140 22888 4146
rect 22836 4082 22888 4088
rect 22848 3194 22876 4082
rect 23308 3942 23336 6190
rect 23584 6118 23612 6190
rect 23572 6112 23624 6118
rect 23572 6054 23624 6060
rect 23572 4480 23624 4486
rect 23572 4422 23624 4428
rect 23584 4214 23612 4422
rect 23572 4208 23624 4214
rect 23572 4150 23624 4156
rect 23676 4078 23704 6598
rect 24412 6186 24440 6802
rect 24780 6662 24808 6870
rect 25148 6866 25176 8230
rect 25320 8016 25372 8022
rect 25320 7958 25372 7964
rect 25332 7546 25360 7958
rect 25320 7540 25372 7546
rect 25320 7482 25372 7488
rect 25136 6860 25188 6866
rect 25136 6802 25188 6808
rect 24768 6656 24820 6662
rect 24768 6598 24820 6604
rect 24780 6458 24808 6598
rect 24768 6452 24820 6458
rect 24768 6394 24820 6400
rect 25332 6390 25360 7482
rect 25412 6860 25464 6866
rect 25412 6802 25464 6808
rect 25424 6458 25452 6802
rect 25504 6656 25556 6662
rect 25504 6598 25556 6604
rect 25412 6452 25464 6458
rect 25412 6394 25464 6400
rect 25320 6384 25372 6390
rect 25320 6326 25372 6332
rect 24400 6180 24452 6186
rect 24400 6122 24452 6128
rect 24412 5914 24440 6122
rect 24400 5908 24452 5914
rect 24400 5850 24452 5856
rect 24030 5672 24086 5681
rect 24030 5607 24086 5616
rect 23940 5092 23992 5098
rect 23940 5034 23992 5040
rect 23952 4826 23980 5034
rect 23940 4820 23992 4826
rect 23940 4762 23992 4768
rect 23848 4684 23900 4690
rect 23848 4626 23900 4632
rect 23664 4072 23716 4078
rect 23664 4014 23716 4020
rect 23296 3936 23348 3942
rect 23296 3878 23348 3884
rect 23294 3768 23350 3777
rect 23676 3738 23704 4014
rect 23860 4010 23888 4626
rect 23848 4004 23900 4010
rect 23848 3946 23900 3952
rect 23294 3703 23296 3712
rect 23348 3703 23350 3712
rect 23664 3732 23716 3738
rect 23296 3674 23348 3680
rect 23664 3674 23716 3680
rect 23756 3596 23808 3602
rect 23756 3538 23808 3544
rect 23388 3392 23440 3398
rect 23388 3334 23440 3340
rect 22836 3188 22888 3194
rect 22836 3130 22888 3136
rect 23400 2854 23428 3334
rect 23768 2922 23796 3538
rect 23756 2916 23808 2922
rect 23756 2858 23808 2864
rect 23388 2848 23440 2854
rect 23388 2790 23440 2796
rect 23400 2446 23428 2790
rect 23388 2440 23440 2446
rect 23388 2382 23440 2388
rect 23860 480 23888 3946
rect 24044 2650 24072 5607
rect 24952 5568 25004 5574
rect 24952 5510 25004 5516
rect 24768 5160 24820 5166
rect 24768 5102 24820 5108
rect 24860 5160 24912 5166
rect 24860 5102 24912 5108
rect 24306 4856 24362 4865
rect 24306 4791 24308 4800
rect 24360 4791 24362 4800
rect 24308 4762 24360 4768
rect 24320 4078 24348 4762
rect 24584 4752 24636 4758
rect 24584 4694 24636 4700
rect 24308 4072 24360 4078
rect 24308 4014 24360 4020
rect 24400 3392 24452 3398
rect 24400 3334 24452 3340
rect 24412 3058 24440 3334
rect 24596 3126 24624 4694
rect 24676 4616 24728 4622
rect 24676 4558 24728 4564
rect 24688 4321 24716 4558
rect 24674 4312 24730 4321
rect 24674 4247 24730 4256
rect 24688 4146 24716 4247
rect 24676 4140 24728 4146
rect 24676 4082 24728 4088
rect 24780 4078 24808 5102
rect 24768 4072 24820 4078
rect 24768 4014 24820 4020
rect 24872 3738 24900 5102
rect 24964 4554 24992 5510
rect 25044 5024 25096 5030
rect 25042 4992 25044 5001
rect 25096 4992 25098 5001
rect 25042 4927 25098 4936
rect 25318 4992 25374 5001
rect 25318 4927 25374 4936
rect 24952 4548 25004 4554
rect 24952 4490 25004 4496
rect 24860 3732 24912 3738
rect 24860 3674 24912 3680
rect 24964 3670 24992 4490
rect 25332 3777 25360 4927
rect 25516 4826 25544 6598
rect 25608 5370 25636 8434
rect 26240 8424 26292 8430
rect 26240 8366 26292 8372
rect 26148 8356 26200 8362
rect 26148 8298 26200 8304
rect 25964 7744 26016 7750
rect 25964 7686 26016 7692
rect 25976 7546 26004 7686
rect 25964 7540 26016 7546
rect 25964 7482 26016 7488
rect 25872 6724 25924 6730
rect 25872 6666 25924 6672
rect 25596 5364 25648 5370
rect 25596 5306 25648 5312
rect 25504 4820 25556 4826
rect 25504 4762 25556 4768
rect 25608 4214 25636 5306
rect 25884 4826 25912 6666
rect 26160 6458 26188 8298
rect 26252 8090 26280 8366
rect 26240 8084 26292 8090
rect 26240 8026 26292 8032
rect 26620 7546 26648 8570
rect 26792 8356 26844 8362
rect 26792 8298 26844 8304
rect 26804 8022 26832 8298
rect 28092 8090 28120 8570
rect 27620 8084 27672 8090
rect 27620 8026 27672 8032
rect 28080 8084 28132 8090
rect 28080 8026 28132 8032
rect 26792 8016 26844 8022
rect 26792 7958 26844 7964
rect 26700 7880 26752 7886
rect 26700 7822 26752 7828
rect 26424 7540 26476 7546
rect 26424 7482 26476 7488
rect 26608 7540 26660 7546
rect 26608 7482 26660 7488
rect 26436 7342 26464 7482
rect 26424 7336 26476 7342
rect 26424 7278 26476 7284
rect 26516 7336 26568 7342
rect 26516 7278 26568 7284
rect 26148 6452 26200 6458
rect 26148 6394 26200 6400
rect 26528 6254 26556 7278
rect 26712 6730 26740 7822
rect 27632 6934 27660 8026
rect 27804 8016 27856 8022
rect 27804 7958 27856 7964
rect 27816 7546 27844 7958
rect 28736 7954 28764 8570
rect 29380 8022 29408 8774
rect 28816 8016 28868 8022
rect 28816 7958 28868 7964
rect 29368 8016 29420 8022
rect 29368 7958 29420 7964
rect 28724 7948 28776 7954
rect 28724 7890 28776 7896
rect 28736 7546 28764 7890
rect 27804 7540 27856 7546
rect 27804 7482 27856 7488
rect 28724 7540 28776 7546
rect 28724 7482 28776 7488
rect 27816 7002 27844 7482
rect 27804 6996 27856 7002
rect 27804 6938 27856 6944
rect 27620 6928 27672 6934
rect 27620 6870 27672 6876
rect 28828 6866 28856 7958
rect 29276 7404 29328 7410
rect 29276 7346 29328 7352
rect 29288 6866 29316 7346
rect 29368 7336 29420 7342
rect 29368 7278 29420 7284
rect 29380 7002 29408 7278
rect 29368 6996 29420 7002
rect 29368 6938 29420 6944
rect 27252 6860 27304 6866
rect 27252 6802 27304 6808
rect 28080 6860 28132 6866
rect 28080 6802 28132 6808
rect 28816 6860 28868 6866
rect 28816 6802 28868 6808
rect 29276 6860 29328 6866
rect 29276 6802 29328 6808
rect 26700 6724 26752 6730
rect 26700 6666 26752 6672
rect 26712 6322 26740 6666
rect 26700 6316 26752 6322
rect 26700 6258 26752 6264
rect 26516 6248 26568 6254
rect 26516 6190 26568 6196
rect 26528 5914 26556 6190
rect 27264 6118 27292 6802
rect 27344 6656 27396 6662
rect 27344 6598 27396 6604
rect 27712 6656 27764 6662
rect 27712 6598 27764 6604
rect 27252 6112 27304 6118
rect 27252 6054 27304 6060
rect 26516 5908 26568 5914
rect 26516 5850 26568 5856
rect 26792 5704 26844 5710
rect 27264 5681 27292 6054
rect 26792 5646 26844 5652
rect 27250 5672 27306 5681
rect 26804 5370 26832 5646
rect 27250 5607 27306 5616
rect 26240 5364 26292 5370
rect 26240 5306 26292 5312
rect 26792 5364 26844 5370
rect 26792 5306 26844 5312
rect 26252 4826 26280 5306
rect 27160 5160 27212 5166
rect 27160 5102 27212 5108
rect 26332 5024 26384 5030
rect 26332 4966 26384 4972
rect 25872 4820 25924 4826
rect 25872 4762 25924 4768
rect 26240 4820 26292 4826
rect 26240 4762 26292 4768
rect 25870 4584 25926 4593
rect 25870 4519 25926 4528
rect 26148 4548 26200 4554
rect 25596 4208 25648 4214
rect 25596 4150 25648 4156
rect 25504 4072 25556 4078
rect 25504 4014 25556 4020
rect 25318 3768 25374 3777
rect 25318 3703 25320 3712
rect 25372 3703 25374 3712
rect 25320 3674 25372 3680
rect 24952 3664 25004 3670
rect 25332 3643 25360 3674
rect 24952 3606 25004 3612
rect 25228 3596 25280 3602
rect 25228 3538 25280 3544
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24780 3233 24808 3334
rect 24766 3224 24822 3233
rect 25240 3194 25268 3538
rect 25516 3194 25544 4014
rect 25608 3534 25636 4150
rect 25884 4078 25912 4519
rect 26148 4490 26200 4496
rect 25872 4072 25924 4078
rect 25872 4014 25924 4020
rect 26160 3534 26188 4490
rect 26344 3738 26372 4966
rect 26516 4616 26568 4622
rect 26516 4558 26568 4564
rect 26528 4282 26556 4558
rect 26516 4276 26568 4282
rect 26516 4218 26568 4224
rect 26528 4010 26556 4218
rect 26516 4004 26568 4010
rect 26516 3946 26568 3952
rect 26332 3732 26384 3738
rect 26332 3674 26384 3680
rect 25596 3528 25648 3534
rect 25596 3470 25648 3476
rect 26148 3528 26200 3534
rect 26148 3470 26200 3476
rect 24766 3159 24822 3168
rect 25228 3188 25280 3194
rect 24584 3120 24636 3126
rect 24584 3062 24636 3068
rect 24400 3052 24452 3058
rect 24400 2994 24452 3000
rect 24780 2922 24808 3159
rect 25228 3130 25280 3136
rect 25504 3188 25556 3194
rect 25504 3130 25556 3136
rect 24768 2916 24820 2922
rect 24768 2858 24820 2864
rect 24952 2848 25004 2854
rect 24952 2790 25004 2796
rect 24490 2680 24546 2689
rect 24032 2644 24084 2650
rect 24490 2615 24492 2624
rect 24032 2586 24084 2592
rect 24544 2615 24546 2624
rect 24492 2586 24544 2592
rect 24030 2408 24086 2417
rect 24030 2343 24086 2352
rect 24044 2310 24072 2343
rect 24032 2304 24084 2310
rect 24032 2246 24084 2252
rect 24044 2145 24072 2246
rect 24030 2136 24086 2145
rect 24030 2071 24086 2080
rect 24964 480 24992 2790
rect 25962 2680 26018 2689
rect 26528 2650 26556 3946
rect 26976 3936 27028 3942
rect 26976 3878 27028 3884
rect 26988 2990 27016 3878
rect 27068 3732 27120 3738
rect 27068 3674 27120 3680
rect 27080 3602 27108 3674
rect 27068 3596 27120 3602
rect 27068 3538 27120 3544
rect 27172 3398 27200 5102
rect 27160 3392 27212 3398
rect 27160 3334 27212 3340
rect 27158 3224 27214 3233
rect 27158 3159 27160 3168
rect 27212 3159 27214 3168
rect 27160 3130 27212 3136
rect 26976 2984 27028 2990
rect 26976 2926 27028 2932
rect 25962 2615 25964 2624
rect 26016 2615 26018 2624
rect 26516 2644 26568 2650
rect 25964 2586 26016 2592
rect 26516 2586 26568 2592
rect 27172 2582 27200 3130
rect 26056 2576 26108 2582
rect 25778 2544 25834 2553
rect 26056 2518 26108 2524
rect 27160 2576 27212 2582
rect 27160 2518 27212 2524
rect 25778 2479 25780 2488
rect 25832 2479 25834 2488
rect 25780 2450 25832 2456
rect 26068 2310 26096 2518
rect 26056 2304 26108 2310
rect 26056 2246 26108 2252
rect 26068 480 26096 2246
rect 27264 480 27292 5607
rect 27356 3369 27384 6598
rect 27528 6112 27580 6118
rect 27528 6054 27580 6060
rect 27436 5024 27488 5030
rect 27436 4966 27488 4972
rect 27448 4486 27476 4966
rect 27436 4480 27488 4486
rect 27436 4422 27488 4428
rect 27540 3738 27568 6054
rect 27724 5914 27752 6598
rect 28092 6458 28120 6802
rect 28448 6792 28500 6798
rect 28448 6734 28500 6740
rect 28356 6724 28408 6730
rect 28356 6666 28408 6672
rect 28368 6458 28396 6666
rect 28080 6452 28132 6458
rect 28080 6394 28132 6400
rect 28356 6452 28408 6458
rect 28356 6394 28408 6400
rect 28460 6322 28488 6734
rect 29288 6390 29316 6802
rect 29276 6384 29328 6390
rect 29276 6326 29328 6332
rect 28448 6316 28500 6322
rect 28448 6258 28500 6264
rect 28356 6248 28408 6254
rect 28356 6190 28408 6196
rect 28368 5914 28396 6190
rect 28460 5914 28488 6258
rect 29288 6202 29316 6326
rect 29196 6174 29316 6202
rect 29644 6248 29696 6254
rect 29644 6190 29696 6196
rect 27712 5908 27764 5914
rect 27712 5850 27764 5856
rect 28356 5908 28408 5914
rect 28356 5850 28408 5856
rect 28448 5908 28500 5914
rect 28448 5850 28500 5856
rect 28368 5642 28396 5850
rect 29196 5710 29224 6174
rect 29276 6112 29328 6118
rect 29276 6054 29328 6060
rect 29288 5778 29316 6054
rect 29656 5846 29684 6190
rect 29748 5953 29776 13903
rect 30852 13870 30880 14418
rect 31300 14272 31352 14278
rect 31680 14226 31708 14894
rect 31300 14214 31352 14220
rect 31312 14074 31340 14214
rect 31588 14198 31708 14226
rect 31300 14068 31352 14074
rect 31300 14010 31352 14016
rect 31588 14006 31616 14198
rect 31772 14090 31800 15302
rect 32140 14618 32168 15506
rect 32128 14612 32180 14618
rect 32128 14554 32180 14560
rect 31680 14062 31800 14090
rect 31576 14000 31628 14006
rect 31576 13942 31628 13948
rect 31680 13938 31708 14062
rect 31668 13932 31720 13938
rect 31668 13874 31720 13880
rect 30840 13864 30892 13870
rect 30840 13806 30892 13812
rect 30852 13530 30880 13806
rect 31680 13530 31708 13874
rect 31944 13728 31996 13734
rect 31944 13670 31996 13676
rect 31956 13530 31984 13670
rect 30840 13524 30892 13530
rect 30840 13466 30892 13472
rect 31668 13524 31720 13530
rect 31668 13466 31720 13472
rect 31944 13524 31996 13530
rect 31944 13466 31996 13472
rect 32324 13410 32352 16102
rect 33060 15910 33088 16934
rect 33232 16584 33284 16590
rect 33232 16526 33284 16532
rect 33244 16250 33272 16526
rect 33232 16244 33284 16250
rect 33232 16186 33284 16192
rect 33048 15904 33100 15910
rect 33048 15846 33100 15852
rect 33060 14890 33088 15846
rect 33428 15706 33456 17138
rect 33888 16794 33916 17138
rect 33876 16788 33928 16794
rect 33876 16730 33928 16736
rect 33416 15700 33468 15706
rect 33416 15642 33468 15648
rect 33232 15564 33284 15570
rect 33232 15506 33284 15512
rect 33048 14884 33100 14890
rect 33048 14826 33100 14832
rect 33244 14822 33272 15506
rect 33692 15360 33744 15366
rect 33692 15302 33744 15308
rect 33704 14958 33732 15302
rect 33692 14952 33744 14958
rect 33690 14920 33692 14929
rect 33744 14920 33746 14929
rect 33690 14855 33746 14864
rect 32496 14816 32548 14822
rect 32496 14758 32548 14764
rect 33232 14816 33284 14822
rect 33232 14758 33284 14764
rect 33876 14816 33928 14822
rect 33876 14758 33928 14764
rect 34152 14816 34204 14822
rect 34152 14758 34204 14764
rect 32508 14618 32536 14758
rect 32496 14612 32548 14618
rect 32496 14554 32548 14560
rect 32404 13796 32456 13802
rect 32404 13738 32456 13744
rect 32416 13530 32444 13738
rect 32508 13734 32536 14554
rect 33416 14544 33468 14550
rect 33416 14486 33468 14492
rect 32588 14476 32640 14482
rect 32588 14418 32640 14424
rect 32600 14074 32628 14418
rect 33428 14278 33456 14486
rect 33784 14476 33836 14482
rect 33784 14418 33836 14424
rect 33324 14272 33376 14278
rect 33324 14214 33376 14220
rect 33416 14272 33468 14278
rect 33416 14214 33468 14220
rect 33796 14226 33824 14418
rect 33888 14414 33916 14758
rect 33876 14408 33928 14414
rect 33876 14350 33928 14356
rect 34060 14272 34112 14278
rect 32588 14068 32640 14074
rect 32588 14010 32640 14016
rect 32496 13728 32548 13734
rect 32496 13670 32548 13676
rect 33140 13728 33192 13734
rect 33140 13670 33192 13676
rect 33152 13530 33180 13670
rect 32404 13524 32456 13530
rect 32404 13466 32456 13472
rect 32864 13524 32916 13530
rect 32864 13466 32916 13472
rect 33140 13524 33192 13530
rect 33140 13466 33192 13472
rect 32220 13388 32272 13394
rect 32324 13382 32536 13410
rect 32220 13330 32272 13336
rect 30380 13252 30432 13258
rect 30380 13194 30432 13200
rect 29826 12880 29882 12889
rect 30392 12850 30420 13194
rect 30472 13184 30524 13190
rect 30472 13126 30524 13132
rect 30484 12986 30512 13126
rect 32232 12986 32260 13330
rect 30472 12980 30524 12986
rect 30472 12922 30524 12928
rect 32220 12980 32272 12986
rect 32220 12922 32272 12928
rect 29826 12815 29828 12824
rect 29880 12815 29882 12824
rect 30380 12844 30432 12850
rect 29828 12786 29880 12792
rect 30380 12786 30432 12792
rect 31944 12844 31996 12850
rect 31944 12786 31996 12792
rect 29840 12442 29868 12786
rect 30288 12708 30340 12714
rect 30288 12650 30340 12656
rect 30300 12442 30328 12650
rect 31208 12640 31260 12646
rect 31208 12582 31260 12588
rect 29828 12436 29880 12442
rect 29828 12378 29880 12384
rect 30288 12436 30340 12442
rect 30288 12378 30340 12384
rect 30472 12300 30524 12306
rect 30472 12242 30524 12248
rect 30196 12232 30248 12238
rect 30196 12174 30248 12180
rect 30208 11286 30236 12174
rect 30380 12096 30432 12102
rect 30300 12044 30380 12050
rect 30300 12038 30432 12044
rect 30300 12022 30420 12038
rect 30196 11280 30248 11286
rect 30196 11222 30248 11228
rect 30300 11098 30328 12022
rect 30380 11552 30432 11558
rect 30380 11494 30432 11500
rect 30208 11070 30328 11098
rect 30012 10464 30064 10470
rect 30012 10406 30064 10412
rect 30024 10130 30052 10406
rect 30208 10198 30236 11070
rect 30392 10690 30420 11494
rect 30484 11354 30512 12242
rect 30840 12232 30892 12238
rect 30840 12174 30892 12180
rect 30852 11898 30880 12174
rect 31220 12102 31248 12582
rect 31956 12442 31984 12786
rect 32312 12640 32364 12646
rect 32312 12582 32364 12588
rect 31944 12436 31996 12442
rect 31944 12378 31996 12384
rect 31208 12096 31260 12102
rect 31208 12038 31260 12044
rect 32324 11898 32352 12582
rect 30840 11892 30892 11898
rect 30840 11834 30892 11840
rect 32312 11892 32364 11898
rect 32312 11834 32364 11840
rect 30852 11354 30880 11834
rect 32404 11620 32456 11626
rect 32404 11562 32456 11568
rect 30472 11348 30524 11354
rect 30472 11290 30524 11296
rect 30840 11348 30892 11354
rect 30840 11290 30892 11296
rect 30300 10662 30420 10690
rect 30300 10606 30328 10662
rect 30288 10600 30340 10606
rect 30288 10542 30340 10548
rect 30300 10266 30328 10542
rect 30288 10260 30340 10266
rect 30288 10202 30340 10208
rect 30196 10192 30248 10198
rect 30196 10134 30248 10140
rect 30012 10124 30064 10130
rect 30012 10066 30064 10072
rect 30024 9722 30052 10066
rect 30196 10056 30248 10062
rect 30196 9998 30248 10004
rect 30208 9722 30236 9998
rect 30012 9716 30064 9722
rect 30012 9658 30064 9664
rect 30196 9716 30248 9722
rect 30196 9658 30248 9664
rect 30300 9654 30328 10202
rect 30852 9654 30880 11290
rect 32416 11286 32444 11562
rect 32404 11280 32456 11286
rect 32404 11222 32456 11228
rect 32128 11144 32180 11150
rect 32128 11086 32180 11092
rect 32140 10810 32168 11086
rect 32416 10810 32444 11222
rect 32508 10826 32536 13382
rect 32876 12442 32904 13466
rect 33048 13252 33100 13258
rect 33048 13194 33100 13200
rect 33060 12442 33088 13194
rect 33336 12850 33364 14214
rect 33428 13938 33456 14214
rect 33796 14198 33916 14226
rect 34060 14214 34112 14220
rect 33888 14006 33916 14198
rect 33876 14000 33928 14006
rect 33874 13968 33876 13977
rect 33928 13968 33930 13977
rect 33416 13932 33468 13938
rect 33874 13903 33930 13912
rect 33416 13874 33468 13880
rect 33416 13524 33468 13530
rect 33416 13466 33468 13472
rect 33324 12844 33376 12850
rect 33324 12786 33376 12792
rect 33428 12442 33456 13466
rect 33600 12708 33652 12714
rect 33600 12650 33652 12656
rect 33612 12442 33640 12650
rect 34072 12442 34100 14214
rect 34164 13870 34192 14758
rect 34532 14634 34560 17983
rect 34256 14606 34560 14634
rect 34152 13864 34204 13870
rect 34152 13806 34204 13812
rect 34256 12481 34284 14606
rect 34348 14482 34560 14498
rect 34348 14476 34572 14482
rect 34348 14470 34520 14476
rect 34348 13394 34376 14470
rect 34520 14418 34572 14424
rect 34520 14340 34572 14346
rect 34520 14282 34572 14288
rect 34532 13546 34560 14282
rect 34440 13518 34560 13546
rect 34440 13462 34468 13518
rect 34428 13456 34480 13462
rect 34428 13398 34480 13404
rect 34336 13388 34388 13394
rect 34336 13330 34388 13336
rect 34428 13320 34480 13326
rect 34428 13262 34480 13268
rect 34440 12850 34468 13262
rect 34428 12844 34480 12850
rect 34428 12786 34480 12792
rect 34242 12472 34298 12481
rect 32864 12436 32916 12442
rect 32864 12378 32916 12384
rect 33048 12436 33100 12442
rect 33048 12378 33100 12384
rect 33416 12436 33468 12442
rect 33416 12378 33468 12384
rect 33600 12436 33652 12442
rect 33600 12378 33652 12384
rect 34060 12436 34112 12442
rect 34242 12407 34298 12416
rect 34336 12436 34388 12442
rect 34060 12378 34112 12384
rect 34336 12378 34388 12384
rect 33876 12300 33928 12306
rect 33876 12242 33928 12248
rect 33888 11762 33916 12242
rect 34348 12238 34376 12378
rect 33968 12232 34020 12238
rect 33968 12174 34020 12180
rect 34336 12232 34388 12238
rect 34336 12174 34388 12180
rect 34440 12186 34468 12786
rect 34716 12730 34744 19110
rect 34808 12866 34836 21286
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 35268 19281 35296 24511
rect 35360 22982 35388 25214
rect 35440 25152 35492 25158
rect 35440 25094 35492 25100
rect 35452 24818 35480 25094
rect 35544 24857 35572 25638
rect 35530 24848 35586 24857
rect 35440 24812 35492 24818
rect 35530 24783 35586 24792
rect 35636 24800 35664 28999
rect 35728 27130 35756 29158
rect 35912 29073 35940 29990
rect 35992 29640 36044 29646
rect 35992 29582 36044 29588
rect 35898 29064 35954 29073
rect 35898 28999 35954 29008
rect 36004 28762 36032 29582
rect 35992 28756 36044 28762
rect 35992 28698 36044 28704
rect 35992 28620 36044 28626
rect 35992 28562 36044 28568
rect 36004 27878 36032 28562
rect 36096 28422 36124 31078
rect 36740 30326 36768 33215
rect 36832 32570 36860 34439
rect 36820 32564 36872 32570
rect 36820 32506 36872 32512
rect 37096 32224 37148 32230
rect 37096 32166 37148 32172
rect 36728 30320 36780 30326
rect 36728 30262 36780 30268
rect 36176 30116 36228 30122
rect 36176 30058 36228 30064
rect 36084 28416 36136 28422
rect 36084 28358 36136 28364
rect 36188 28234 36216 30058
rect 36268 29232 36320 29238
rect 36266 29200 36268 29209
rect 36320 29200 36322 29209
rect 36266 29135 36322 29144
rect 36728 28416 36780 28422
rect 36728 28358 36780 28364
rect 36096 28206 36216 28234
rect 36740 28218 36768 28358
rect 36728 28212 36780 28218
rect 35992 27872 36044 27878
rect 35992 27814 36044 27820
rect 35716 27124 35768 27130
rect 35716 27066 35768 27072
rect 35716 26920 35768 26926
rect 36004 26874 36032 27814
rect 35716 26862 35768 26868
rect 35728 26518 35756 26862
rect 35820 26846 36032 26874
rect 35716 26512 35768 26518
rect 35716 26454 35768 26460
rect 35636 24772 35756 24800
rect 35440 24754 35492 24760
rect 35452 24410 35480 24754
rect 35440 24404 35492 24410
rect 35440 24346 35492 24352
rect 35452 23254 35480 24346
rect 35728 24154 35756 24772
rect 35636 24126 35756 24154
rect 35440 23248 35492 23254
rect 35440 23190 35492 23196
rect 35348 22976 35400 22982
rect 35348 22918 35400 22924
rect 35440 22432 35492 22438
rect 35440 22374 35492 22380
rect 35532 22432 35584 22438
rect 35532 22374 35584 22380
rect 35452 22234 35480 22374
rect 35440 22228 35492 22234
rect 35440 22170 35492 22176
rect 35346 21584 35402 21593
rect 35346 21519 35348 21528
rect 35400 21519 35402 21528
rect 35440 21548 35492 21554
rect 35348 21490 35400 21496
rect 35440 21490 35492 21496
rect 35346 21176 35402 21185
rect 35346 21111 35402 21120
rect 35360 20924 35388 21111
rect 35452 21078 35480 21490
rect 35440 21072 35492 21078
rect 35440 21014 35492 21020
rect 35360 20896 35480 20924
rect 35348 20800 35400 20806
rect 35452 20777 35480 20896
rect 35348 20742 35400 20748
rect 35438 20768 35494 20777
rect 35360 19990 35388 20742
rect 35438 20703 35494 20712
rect 35348 19984 35400 19990
rect 35348 19926 35400 19932
rect 35360 19514 35388 19926
rect 35348 19508 35400 19514
rect 35348 19450 35400 19456
rect 35254 19272 35310 19281
rect 35254 19207 35310 19216
rect 35256 19168 35308 19174
rect 35256 19110 35308 19116
rect 35268 18970 35296 19110
rect 35256 18964 35308 18970
rect 35256 18906 35308 18912
rect 35452 18850 35480 20703
rect 35268 18822 35480 18850
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 35268 17270 35296 18822
rect 35438 18728 35494 18737
rect 35438 18663 35494 18672
rect 35452 17746 35480 18663
rect 35440 17740 35492 17746
rect 35440 17682 35492 17688
rect 35346 17504 35402 17513
rect 35346 17439 35402 17448
rect 35256 17264 35308 17270
rect 35256 17206 35308 17212
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 35360 16017 35388 17439
rect 35452 17338 35480 17682
rect 35440 17332 35492 17338
rect 35440 17274 35492 17280
rect 35346 16008 35402 16017
rect 35346 15943 35402 15952
rect 35256 15564 35308 15570
rect 35256 15506 35308 15512
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 35268 14890 35296 15506
rect 35348 15360 35400 15366
rect 35348 15302 35400 15308
rect 35360 15162 35388 15302
rect 35348 15156 35400 15162
rect 35348 15098 35400 15104
rect 35256 14884 35308 14890
rect 35256 14826 35308 14832
rect 35268 14482 35296 14826
rect 35256 14476 35308 14482
rect 35256 14418 35308 14424
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 35268 14074 35296 14418
rect 35348 14408 35400 14414
rect 35348 14350 35400 14356
rect 35256 14068 35308 14074
rect 35256 14010 35308 14016
rect 35360 13870 35388 14350
rect 35440 14272 35492 14278
rect 35440 14214 35492 14220
rect 35348 13864 35400 13870
rect 35348 13806 35400 13812
rect 35256 13728 35308 13734
rect 35256 13670 35308 13676
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 34808 12838 35112 12866
rect 34716 12702 34836 12730
rect 34520 12640 34572 12646
rect 34520 12582 34572 12588
rect 34532 12374 34560 12582
rect 34610 12472 34666 12481
rect 34610 12407 34666 12416
rect 34520 12368 34572 12374
rect 34520 12310 34572 12316
rect 34624 12238 34652 12407
rect 34612 12232 34664 12238
rect 33980 11898 34008 12174
rect 34348 11898 34376 12174
rect 34440 12158 34560 12186
rect 34612 12174 34664 12180
rect 34428 12096 34480 12102
rect 34428 12038 34480 12044
rect 33968 11892 34020 11898
rect 33968 11834 34020 11840
rect 34336 11892 34388 11898
rect 34336 11834 34388 11840
rect 33876 11756 33928 11762
rect 33876 11698 33928 11704
rect 33508 11552 33560 11558
rect 33508 11494 33560 11500
rect 33520 11354 33548 11494
rect 33508 11348 33560 11354
rect 33508 11290 33560 11296
rect 32128 10804 32180 10810
rect 32128 10746 32180 10752
rect 32404 10804 32456 10810
rect 32508 10798 32628 10826
rect 32404 10746 32456 10752
rect 32416 10690 32444 10746
rect 32416 10662 32536 10690
rect 32404 10532 32456 10538
rect 32404 10474 32456 10480
rect 31024 10464 31076 10470
rect 31024 10406 31076 10412
rect 31036 10266 31064 10406
rect 32416 10266 32444 10474
rect 32508 10266 32536 10662
rect 31024 10260 31076 10266
rect 31024 10202 31076 10208
rect 32404 10260 32456 10266
rect 32404 10202 32456 10208
rect 32496 10260 32548 10266
rect 32496 10202 32548 10208
rect 30288 9648 30340 9654
rect 30288 9590 30340 9596
rect 30840 9648 30892 9654
rect 30840 9590 30892 9596
rect 30104 7744 30156 7750
rect 30104 7686 30156 7692
rect 30116 7342 30144 7686
rect 30104 7336 30156 7342
rect 30104 7278 30156 7284
rect 30380 7200 30432 7206
rect 30380 7142 30432 7148
rect 30392 6866 30420 7142
rect 30380 6860 30432 6866
rect 30380 6802 30432 6808
rect 30392 6458 30420 6802
rect 30656 6656 30708 6662
rect 30656 6598 30708 6604
rect 30668 6458 30696 6598
rect 30380 6452 30432 6458
rect 30380 6394 30432 6400
rect 30656 6452 30708 6458
rect 30656 6394 30708 6400
rect 29920 6316 29972 6322
rect 29920 6258 29972 6264
rect 29734 5944 29790 5953
rect 29932 5914 29960 6258
rect 30668 6254 30696 6394
rect 30656 6248 30708 6254
rect 30656 6190 30708 6196
rect 29734 5879 29790 5888
rect 29920 5908 29972 5914
rect 29920 5850 29972 5856
rect 29644 5840 29696 5846
rect 29644 5782 29696 5788
rect 29276 5772 29328 5778
rect 29276 5714 29328 5720
rect 29184 5704 29236 5710
rect 29184 5646 29236 5652
rect 28356 5636 28408 5642
rect 28356 5578 28408 5584
rect 29196 5370 29224 5646
rect 30564 5568 30616 5574
rect 30564 5510 30616 5516
rect 29184 5364 29236 5370
rect 29184 5306 29236 5312
rect 28264 5228 28316 5234
rect 28264 5170 28316 5176
rect 27988 5160 28040 5166
rect 27988 5102 28040 5108
rect 28000 5030 28028 5102
rect 27620 5024 27672 5030
rect 27620 4966 27672 4972
rect 27988 5024 28040 5030
rect 27988 4966 28040 4972
rect 27632 4690 27660 4966
rect 27710 4856 27766 4865
rect 27710 4791 27766 4800
rect 27724 4758 27752 4791
rect 27712 4752 27764 4758
rect 28000 4729 28028 4966
rect 28276 4826 28304 5170
rect 28264 4820 28316 4826
rect 28264 4762 28316 4768
rect 27712 4694 27764 4700
rect 27986 4720 28042 4729
rect 27620 4684 27672 4690
rect 27620 4626 27672 4632
rect 27724 4146 27752 4694
rect 27986 4655 28042 4664
rect 27894 4584 27950 4593
rect 27894 4519 27896 4528
rect 27948 4519 27950 4528
rect 27896 4490 27948 4496
rect 28276 4282 28304 4762
rect 28632 4684 28684 4690
rect 28632 4626 28684 4632
rect 28644 4282 28672 4626
rect 29000 4480 29052 4486
rect 29000 4422 29052 4428
rect 28264 4276 28316 4282
rect 28264 4218 28316 4224
rect 28632 4276 28684 4282
rect 28632 4218 28684 4224
rect 29012 4146 29040 4422
rect 27712 4140 27764 4146
rect 27712 4082 27764 4088
rect 29000 4140 29052 4146
rect 29000 4082 29052 4088
rect 28264 4072 28316 4078
rect 28264 4014 28316 4020
rect 27528 3732 27580 3738
rect 27528 3674 27580 3680
rect 28172 3596 28224 3602
rect 28172 3538 28224 3544
rect 27342 3360 27398 3369
rect 27342 3295 27398 3304
rect 28184 2854 28212 3538
rect 28276 3398 28304 4014
rect 29196 3913 29224 5306
rect 29920 5228 29972 5234
rect 29920 5170 29972 5176
rect 29460 5092 29512 5098
rect 29460 5034 29512 5040
rect 29276 5024 29328 5030
rect 29276 4966 29328 4972
rect 29288 4758 29316 4966
rect 29276 4752 29328 4758
rect 29276 4694 29328 4700
rect 29472 4282 29500 5034
rect 29736 5024 29788 5030
rect 29736 4966 29788 4972
rect 29748 4826 29776 4966
rect 29932 4826 29960 5170
rect 30576 5114 30604 5510
rect 30668 5370 30696 6190
rect 31392 6112 31444 6118
rect 31392 6054 31444 6060
rect 31208 5568 31260 5574
rect 31208 5510 31260 5516
rect 30656 5364 30708 5370
rect 30656 5306 30708 5312
rect 30576 5086 30696 5114
rect 30668 5030 30696 5086
rect 31220 5030 31248 5510
rect 31404 5234 31432 6054
rect 31942 5944 31998 5953
rect 31942 5879 31998 5888
rect 31956 5642 31984 5879
rect 31944 5636 31996 5642
rect 31944 5578 31996 5584
rect 32496 5636 32548 5642
rect 32496 5578 32548 5584
rect 32312 5568 32364 5574
rect 32312 5510 32364 5516
rect 31392 5228 31444 5234
rect 31392 5170 31444 5176
rect 30656 5024 30708 5030
rect 30840 5024 30892 5030
rect 30656 4966 30708 4972
rect 30838 4992 30840 5001
rect 31208 5024 31260 5030
rect 30892 4992 30894 5001
rect 30668 4865 30696 4966
rect 31208 4966 31260 4972
rect 30838 4927 30894 4936
rect 30654 4856 30710 4865
rect 29736 4820 29788 4826
rect 29736 4762 29788 4768
rect 29920 4820 29972 4826
rect 30654 4791 30710 4800
rect 29920 4762 29972 4768
rect 29460 4276 29512 4282
rect 29460 4218 29512 4224
rect 29182 3904 29238 3913
rect 29182 3839 29238 3848
rect 28448 3528 28500 3534
rect 28448 3470 28500 3476
rect 28264 3392 28316 3398
rect 28264 3334 28316 3340
rect 28354 3360 28410 3369
rect 28172 2848 28224 2854
rect 28172 2790 28224 2796
rect 28184 2650 28212 2790
rect 28276 2689 28304 3334
rect 28354 3295 28410 3304
rect 28262 2680 28318 2689
rect 28172 2644 28224 2650
rect 28262 2615 28318 2624
rect 28172 2586 28224 2592
rect 28184 2553 28212 2586
rect 28170 2544 28226 2553
rect 28170 2479 28226 2488
rect 28368 480 28396 3295
rect 28460 3194 28488 3470
rect 29196 3194 29224 3839
rect 29458 3768 29514 3777
rect 29932 3738 29960 4762
rect 30380 4684 30432 4690
rect 30380 4626 30432 4632
rect 30288 4480 30340 4486
rect 30288 4422 30340 4428
rect 30012 4140 30064 4146
rect 30012 4082 30064 4088
rect 29458 3703 29514 3712
rect 29920 3732 29972 3738
rect 28448 3188 28500 3194
rect 28448 3130 28500 3136
rect 29184 3188 29236 3194
rect 29184 3130 29236 3136
rect 29196 2650 29224 3130
rect 29184 2644 29236 2650
rect 29184 2586 29236 2592
rect 29472 480 29500 3703
rect 29920 3674 29972 3680
rect 29932 2582 29960 3674
rect 30024 2990 30052 4082
rect 30300 4060 30328 4422
rect 30392 4282 30420 4626
rect 30840 4616 30892 4622
rect 31220 4593 31248 4966
rect 31404 4826 31432 5170
rect 31760 5092 31812 5098
rect 31760 5034 31812 5040
rect 31772 4978 31800 5034
rect 31680 4950 31800 4978
rect 31392 4820 31444 4826
rect 31392 4762 31444 4768
rect 31484 4752 31536 4758
rect 31298 4720 31354 4729
rect 31484 4694 31536 4700
rect 31298 4655 31354 4664
rect 30840 4558 30892 4564
rect 31206 4584 31262 4593
rect 30380 4276 30432 4282
rect 30380 4218 30432 4224
rect 30852 4214 30880 4558
rect 31206 4519 31262 4528
rect 30840 4208 30892 4214
rect 30840 4150 30892 4156
rect 30748 4140 30800 4146
rect 30748 4082 30800 4088
rect 30380 4072 30432 4078
rect 30300 4032 30380 4060
rect 30380 4014 30432 4020
rect 30760 3194 30788 4082
rect 31208 3936 31260 3942
rect 31208 3878 31260 3884
rect 31220 3466 31248 3878
rect 31312 3602 31340 4655
rect 31496 3738 31524 4694
rect 31680 4010 31708 4950
rect 32324 4826 32352 5510
rect 31760 4820 31812 4826
rect 31760 4762 31812 4768
rect 32312 4820 32364 4826
rect 32312 4762 32364 4768
rect 31772 4146 31800 4762
rect 31760 4140 31812 4146
rect 31760 4082 31812 4088
rect 31668 4004 31720 4010
rect 31668 3946 31720 3952
rect 31852 3936 31904 3942
rect 32128 3936 32180 3942
rect 31852 3878 31904 3884
rect 32126 3904 32128 3913
rect 32180 3904 32182 3913
rect 31864 3777 31892 3878
rect 32126 3839 32182 3848
rect 31850 3768 31906 3777
rect 31484 3732 31536 3738
rect 31850 3703 31906 3712
rect 31484 3674 31536 3680
rect 31300 3596 31352 3602
rect 31300 3538 31352 3544
rect 31208 3460 31260 3466
rect 31208 3402 31260 3408
rect 31312 3194 31340 3538
rect 31852 3392 31904 3398
rect 31904 3340 31984 3346
rect 31852 3334 31984 3340
rect 31864 3318 31984 3334
rect 30748 3188 30800 3194
rect 30748 3130 30800 3136
rect 31300 3188 31352 3194
rect 31300 3130 31352 3136
rect 31956 2990 31984 3318
rect 30012 2984 30064 2990
rect 31944 2984 31996 2990
rect 30012 2926 30064 2932
rect 31666 2952 31722 2961
rect 29920 2576 29972 2582
rect 29920 2518 29972 2524
rect 30024 2310 30052 2926
rect 31944 2926 31996 2932
rect 31666 2887 31722 2896
rect 30012 2304 30064 2310
rect 30012 2246 30064 2252
rect 30562 2000 30618 2009
rect 30562 1935 30618 1944
rect 30576 480 30604 1935
rect 31680 480 31708 2887
rect 31956 2650 31984 2926
rect 32140 2650 32168 3839
rect 32508 3641 32536 5578
rect 32600 3754 32628 10798
rect 32956 10464 33008 10470
rect 32956 10406 33008 10412
rect 32968 10062 32996 10406
rect 33520 10198 33548 11290
rect 33980 11286 34008 11834
rect 33968 11280 34020 11286
rect 33968 11222 34020 11228
rect 34348 11082 34376 11834
rect 34336 11076 34388 11082
rect 34336 11018 34388 11024
rect 34348 10418 34376 11018
rect 34440 10554 34468 12038
rect 34532 10742 34560 12158
rect 34612 12096 34664 12102
rect 34612 12038 34664 12044
rect 34624 11558 34652 12038
rect 34612 11552 34664 11558
rect 34612 11494 34664 11500
rect 34624 11150 34652 11494
rect 34808 11370 34836 12702
rect 34888 12640 34940 12646
rect 34888 12582 34940 12588
rect 34900 12238 34928 12582
rect 34888 12232 34940 12238
rect 34888 12174 34940 12180
rect 35084 12186 35112 12838
rect 35268 12782 35296 13670
rect 35452 13326 35480 14214
rect 35348 13320 35400 13326
rect 35348 13262 35400 13268
rect 35440 13320 35492 13326
rect 35440 13262 35492 13268
rect 35256 12776 35308 12782
rect 35256 12718 35308 12724
rect 35256 12640 35308 12646
rect 35256 12582 35308 12588
rect 35268 12322 35296 12582
rect 35360 12442 35388 13262
rect 35348 12436 35400 12442
rect 35348 12378 35400 12384
rect 35268 12294 35388 12322
rect 35084 12158 35296 12186
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 34716 11342 34836 11370
rect 34612 11144 34664 11150
rect 34612 11086 34664 11092
rect 34624 10810 34652 11086
rect 34612 10804 34664 10810
rect 34612 10746 34664 10752
rect 34520 10736 34572 10742
rect 34520 10678 34572 10684
rect 34440 10526 34652 10554
rect 34348 10390 34560 10418
rect 33508 10192 33560 10198
rect 33508 10134 33560 10140
rect 32956 10056 33008 10062
rect 32956 9998 33008 10004
rect 32968 9722 32996 9998
rect 33520 9722 33548 10134
rect 34532 9994 34560 10390
rect 34520 9988 34572 9994
rect 34520 9930 34572 9936
rect 32956 9716 33008 9722
rect 32956 9658 33008 9664
rect 33508 9716 33560 9722
rect 33508 9658 33560 9664
rect 33324 6112 33376 6118
rect 33324 6054 33376 6060
rect 32680 5704 32732 5710
rect 32680 5646 32732 5652
rect 32692 5370 32720 5646
rect 33140 5568 33192 5574
rect 33140 5510 33192 5516
rect 32680 5364 32732 5370
rect 32680 5306 32732 5312
rect 32692 5166 32720 5306
rect 33048 5228 33100 5234
rect 32968 5188 33048 5216
rect 32680 5160 32732 5166
rect 32680 5102 32732 5108
rect 32680 5024 32732 5030
rect 32680 4966 32732 4972
rect 32692 4185 32720 4966
rect 32678 4176 32734 4185
rect 32678 4111 32734 4120
rect 32968 3942 32996 5188
rect 33048 5170 33100 5176
rect 33152 5098 33180 5510
rect 33232 5296 33284 5302
rect 33232 5238 33284 5244
rect 33140 5092 33192 5098
rect 33140 5034 33192 5040
rect 33048 4548 33100 4554
rect 33048 4490 33100 4496
rect 32956 3936 33008 3942
rect 32956 3878 33008 3884
rect 32600 3726 32720 3754
rect 32494 3632 32550 3641
rect 32312 3596 32364 3602
rect 32494 3567 32550 3576
rect 32312 3538 32364 3544
rect 32324 3398 32352 3538
rect 32508 3534 32536 3567
rect 32692 3534 32720 3726
rect 33060 3534 33088 4490
rect 33244 3720 33272 5238
rect 33336 4826 33364 6054
rect 34336 5772 34388 5778
rect 33980 5710 34008 5741
rect 34336 5714 34388 5720
rect 33968 5704 34020 5710
rect 33966 5672 33968 5681
rect 34020 5672 34022 5681
rect 33966 5607 34022 5616
rect 34244 5636 34296 5642
rect 33980 5370 34008 5607
rect 34244 5578 34296 5584
rect 33968 5364 34020 5370
rect 33968 5306 34020 5312
rect 33324 4820 33376 4826
rect 33324 4762 33376 4768
rect 33784 4616 33836 4622
rect 33784 4558 33836 4564
rect 33796 3942 33824 4558
rect 33692 3936 33744 3942
rect 33692 3878 33744 3884
rect 33784 3936 33836 3942
rect 33784 3878 33836 3884
rect 33152 3692 33272 3720
rect 32496 3528 32548 3534
rect 32496 3470 32548 3476
rect 32680 3528 32732 3534
rect 33048 3528 33100 3534
rect 32680 3470 32732 3476
rect 32770 3496 32826 3505
rect 32404 3460 32456 3466
rect 32404 3402 32456 3408
rect 32312 3392 32364 3398
rect 32312 3334 32364 3340
rect 32324 2825 32352 3334
rect 32416 3058 32444 3402
rect 32508 3194 32536 3470
rect 32496 3188 32548 3194
rect 32496 3130 32548 3136
rect 32404 3052 32456 3058
rect 32404 2994 32456 3000
rect 32692 2854 32720 3470
rect 33048 3470 33100 3476
rect 32770 3431 32826 3440
rect 32680 2848 32732 2854
rect 32310 2816 32366 2825
rect 32680 2790 32732 2796
rect 32310 2751 32366 2760
rect 31944 2644 31996 2650
rect 31944 2586 31996 2592
rect 32128 2644 32180 2650
rect 32128 2586 32180 2592
rect 32784 480 32812 3431
rect 33152 3074 33180 3692
rect 33232 3596 33284 3602
rect 33232 3538 33284 3544
rect 33244 3194 33272 3538
rect 33232 3188 33284 3194
rect 33232 3130 33284 3136
rect 33060 3046 33180 3074
rect 33060 2990 33088 3046
rect 33048 2984 33100 2990
rect 33048 2926 33100 2932
rect 33704 2582 33732 3878
rect 33980 3126 34008 5306
rect 34256 5098 34284 5578
rect 34348 5370 34376 5714
rect 34520 5568 34572 5574
rect 34520 5510 34572 5516
rect 34336 5364 34388 5370
rect 34336 5306 34388 5312
rect 34244 5092 34296 5098
rect 34244 5034 34296 5040
rect 33968 3120 34020 3126
rect 33968 3062 34020 3068
rect 34256 2650 34284 5034
rect 34532 4826 34560 5510
rect 34520 4820 34572 4826
rect 34520 4762 34572 4768
rect 34428 4480 34480 4486
rect 34480 4428 34560 4434
rect 34428 4422 34560 4428
rect 34440 4406 34560 4422
rect 34532 3738 34560 4406
rect 34624 4162 34652 10526
rect 34716 7426 34744 11342
rect 34796 11280 34848 11286
rect 34796 11222 34848 11228
rect 34808 10810 34836 11222
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 34796 10804 34848 10810
rect 34796 10746 34848 10752
rect 34808 10266 34836 10746
rect 34796 10260 34848 10266
rect 34796 10202 34848 10208
rect 34794 10160 34850 10169
rect 34794 10095 34850 10104
rect 34808 9081 34836 10095
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 34794 9072 34850 9081
rect 34794 9007 34850 9016
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 35268 7546 35296 12158
rect 35256 7540 35308 7546
rect 35256 7482 35308 7488
rect 34716 7398 35296 7426
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 34794 5128 34850 5137
rect 34794 5063 34850 5072
rect 34704 5024 34756 5030
rect 34704 4966 34756 4972
rect 34716 4690 34744 4966
rect 34704 4684 34756 4690
rect 34704 4626 34756 4632
rect 34716 4282 34744 4626
rect 34808 4554 34836 5063
rect 34796 4548 34848 4554
rect 34796 4490 34848 4496
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 34704 4276 34756 4282
rect 34704 4218 34756 4224
rect 34624 4134 34744 4162
rect 34610 3768 34666 3777
rect 34520 3732 34572 3738
rect 34610 3703 34666 3712
rect 34520 3674 34572 3680
rect 34624 3670 34652 3703
rect 34612 3664 34664 3670
rect 34612 3606 34664 3612
rect 34336 3392 34388 3398
rect 34336 3334 34388 3340
rect 34348 3058 34376 3334
rect 34336 3052 34388 3058
rect 34336 2994 34388 3000
rect 34716 2961 34744 4134
rect 35164 4072 35216 4078
rect 35164 4014 35216 4020
rect 34796 3596 34848 3602
rect 34796 3538 34848 3544
rect 34808 3194 34836 3538
rect 35176 3482 35204 4014
rect 35268 4010 35296 7398
rect 35360 4185 35388 12294
rect 35438 11520 35494 11529
rect 35438 11455 35494 11464
rect 35452 10130 35480 11455
rect 35440 10124 35492 10130
rect 35440 10066 35492 10072
rect 35452 9722 35480 10066
rect 35440 9716 35492 9722
rect 35440 9658 35492 9664
rect 35544 7857 35572 22374
rect 35636 18306 35664 24126
rect 35716 24064 35768 24070
rect 35716 24006 35768 24012
rect 35728 23662 35756 24006
rect 35716 23656 35768 23662
rect 35820 23633 35848 26846
rect 35992 26512 36044 26518
rect 35992 26454 36044 26460
rect 35900 26308 35952 26314
rect 35900 26250 35952 26256
rect 35912 25838 35940 26250
rect 36004 26042 36032 26454
rect 35992 26036 36044 26042
rect 35992 25978 36044 25984
rect 35900 25832 35952 25838
rect 35900 25774 35952 25780
rect 35716 23598 35768 23604
rect 35806 23624 35862 23633
rect 35728 23322 35756 23598
rect 35806 23559 35862 23568
rect 35716 23316 35768 23322
rect 35716 23258 35768 23264
rect 35728 22642 35756 23258
rect 35716 22636 35768 22642
rect 35716 22578 35768 22584
rect 35990 22536 36046 22545
rect 35900 22500 35952 22506
rect 36096 22522 36124 28206
rect 36728 28154 36780 28160
rect 36544 27328 36596 27334
rect 36544 27270 36596 27276
rect 36452 27124 36504 27130
rect 36452 27066 36504 27072
rect 36174 26888 36230 26897
rect 36174 26823 36230 26832
rect 36188 26042 36216 26823
rect 36176 26036 36228 26042
rect 36176 25978 36228 25984
rect 36464 24290 36492 27066
rect 36556 26926 36584 27270
rect 36820 27056 36872 27062
rect 36818 27024 36820 27033
rect 36872 27024 36874 27033
rect 36818 26959 36874 26968
rect 36544 26920 36596 26926
rect 36544 26862 36596 26868
rect 36464 24262 36584 24290
rect 36452 24200 36504 24206
rect 36452 24142 36504 24148
rect 36464 22778 36492 24142
rect 36556 22778 36584 24262
rect 36818 24168 36874 24177
rect 36818 24103 36874 24112
rect 36832 23866 36860 24103
rect 36820 23860 36872 23866
rect 36820 23802 36872 23808
rect 36832 22778 36860 23802
rect 36912 22976 36964 22982
rect 36912 22918 36964 22924
rect 36452 22772 36504 22778
rect 36452 22714 36504 22720
rect 36544 22772 36596 22778
rect 36544 22714 36596 22720
rect 36820 22772 36872 22778
rect 36820 22714 36872 22720
rect 36464 22574 36492 22714
rect 36046 22494 36124 22522
rect 36452 22568 36504 22574
rect 36452 22510 36504 22516
rect 35990 22471 36046 22480
rect 35900 22442 35952 22448
rect 35912 21690 35940 22442
rect 35900 21684 35952 21690
rect 35900 21626 35952 21632
rect 36004 21570 36032 22471
rect 36556 22438 36584 22714
rect 36544 22432 36596 22438
rect 36544 22374 36596 22380
rect 36832 22234 36860 22714
rect 36924 22710 36952 22918
rect 36912 22704 36964 22710
rect 36912 22646 36964 22652
rect 36820 22228 36872 22234
rect 36820 22170 36872 22176
rect 35820 21542 36032 21570
rect 35716 19236 35768 19242
rect 35716 19178 35768 19184
rect 35728 18970 35756 19178
rect 35716 18964 35768 18970
rect 35716 18906 35768 18912
rect 35714 18320 35770 18329
rect 35636 18278 35714 18306
rect 35714 18255 35770 18264
rect 35622 17640 35678 17649
rect 35622 17575 35624 17584
rect 35676 17575 35678 17584
rect 35624 17546 35676 17552
rect 35624 17264 35676 17270
rect 35624 17206 35676 17212
rect 35636 12594 35664 17206
rect 35728 12714 35756 18255
rect 35716 12708 35768 12714
rect 35716 12650 35768 12656
rect 35636 12566 35756 12594
rect 35622 12472 35678 12481
rect 35622 12407 35678 12416
rect 35636 10606 35664 12407
rect 35624 10600 35676 10606
rect 35624 10542 35676 10548
rect 35622 10296 35678 10305
rect 35622 10231 35678 10240
rect 35530 7848 35586 7857
rect 35530 7783 35586 7792
rect 35532 7540 35584 7546
rect 35532 7482 35584 7488
rect 35440 4616 35492 4622
rect 35440 4558 35492 4564
rect 35346 4176 35402 4185
rect 35346 4111 35402 4120
rect 35256 4004 35308 4010
rect 35256 3946 35308 3952
rect 35176 3454 35296 3482
rect 35452 3466 35480 4558
rect 35544 4434 35572 7482
rect 35636 4570 35664 10231
rect 35728 6633 35756 12566
rect 35714 6624 35770 6633
rect 35714 6559 35770 6568
rect 35820 5409 35848 21542
rect 36176 20800 36228 20806
rect 37108 20777 37136 32166
rect 37188 30592 37240 30598
rect 37188 30534 37240 30540
rect 37200 29306 37228 30534
rect 37188 29300 37240 29306
rect 37188 29242 37240 29248
rect 37188 27872 37240 27878
rect 37188 27814 37240 27820
rect 37200 21185 37228 27814
rect 37844 24585 37872 34478
rect 38016 29028 38068 29034
rect 38016 28970 38068 28976
rect 37830 24576 37886 24585
rect 37830 24511 37886 24520
rect 38028 22409 38056 28970
rect 38014 22400 38070 22409
rect 38014 22335 38070 22344
rect 37186 21176 37242 21185
rect 37186 21111 37242 21120
rect 36176 20742 36228 20748
rect 37094 20768 37150 20777
rect 36188 20330 36216 20742
rect 37094 20703 37150 20712
rect 36636 20528 36688 20534
rect 36634 20496 36636 20505
rect 36688 20496 36690 20505
rect 36634 20431 36690 20440
rect 36176 20324 36228 20330
rect 36176 20266 36228 20272
rect 36188 19718 36216 20266
rect 36176 19712 36228 19718
rect 36176 19654 36228 19660
rect 36188 19378 36216 19654
rect 36176 19372 36228 19378
rect 36176 19314 36228 19320
rect 36544 15700 36596 15706
rect 36544 15642 36596 15648
rect 36556 15609 36584 15642
rect 36542 15600 36598 15609
rect 35900 15564 35952 15570
rect 36542 15535 36598 15544
rect 35900 15506 35952 15512
rect 35912 14822 35940 15506
rect 37094 15056 37150 15065
rect 37094 14991 37150 15000
rect 36818 14920 36874 14929
rect 36818 14855 36874 14864
rect 35900 14816 35952 14822
rect 35900 14758 35952 14764
rect 35912 14618 35940 14758
rect 36832 14618 36860 14855
rect 35900 14612 35952 14618
rect 35900 14554 35952 14560
rect 36820 14612 36872 14618
rect 36820 14554 36872 14560
rect 37108 14550 37136 14991
rect 37096 14544 37148 14550
rect 37096 14486 37148 14492
rect 36544 14476 36596 14482
rect 36544 14418 36596 14424
rect 35900 13796 35952 13802
rect 35900 13738 35952 13744
rect 35912 12986 35940 13738
rect 36556 13530 36584 14418
rect 37108 14074 37136 14486
rect 37096 14068 37148 14074
rect 37096 14010 37148 14016
rect 36544 13524 36596 13530
rect 36544 13466 36596 13472
rect 35992 13388 36044 13394
rect 35992 13330 36044 13336
rect 36004 13190 36032 13330
rect 35992 13184 36044 13190
rect 35992 13126 36044 13132
rect 35900 12980 35952 12986
rect 35900 12922 35952 12928
rect 36004 12782 36032 13126
rect 35992 12776 36044 12782
rect 35992 12718 36044 12724
rect 36004 12442 36032 12718
rect 36634 12608 36690 12617
rect 36634 12543 36690 12552
rect 35992 12436 36044 12442
rect 35992 12378 36044 12384
rect 36268 12300 36320 12306
rect 36268 12242 36320 12248
rect 36280 11898 36308 12242
rect 36268 11892 36320 11898
rect 36268 11834 36320 11840
rect 35992 11620 36044 11626
rect 35992 11562 36044 11568
rect 36004 11354 36032 11562
rect 35992 11348 36044 11354
rect 35992 11290 36044 11296
rect 35806 5400 35862 5409
rect 35806 5335 35862 5344
rect 35636 4542 35848 4570
rect 35716 4480 35768 4486
rect 35544 4406 35664 4434
rect 35716 4422 35768 4428
rect 35532 4004 35584 4010
rect 35532 3946 35584 3952
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 35268 3194 35296 3454
rect 35440 3460 35492 3466
rect 35440 3402 35492 3408
rect 35544 3346 35572 3946
rect 35452 3318 35572 3346
rect 34796 3188 34848 3194
rect 34796 3130 34848 3136
rect 35256 3188 35308 3194
rect 35256 3130 35308 3136
rect 34794 3088 34850 3097
rect 34794 3023 34850 3032
rect 34702 2952 34758 2961
rect 34702 2887 34758 2896
rect 34428 2848 34480 2854
rect 34426 2816 34428 2825
rect 34480 2816 34482 2825
rect 34426 2751 34482 2760
rect 34244 2644 34296 2650
rect 34244 2586 34296 2592
rect 33692 2576 33744 2582
rect 33692 2518 33744 2524
rect 33874 2408 33930 2417
rect 33874 2343 33930 2352
rect 33888 480 33916 2343
rect 34808 1850 34836 3023
rect 35268 2514 35296 3130
rect 35256 2508 35308 2514
rect 35256 2450 35308 2456
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 34808 1822 35020 1850
rect 34992 480 35020 1822
rect 35452 649 35480 3318
rect 35636 1737 35664 4406
rect 35728 4078 35756 4422
rect 35820 4162 35848 4542
rect 36084 4548 36136 4554
rect 36084 4490 36136 4496
rect 35820 4134 35940 4162
rect 35716 4072 35768 4078
rect 35716 4014 35768 4020
rect 35728 3466 35756 4014
rect 35912 3942 35940 4134
rect 35900 3936 35952 3942
rect 35900 3878 35952 3884
rect 35716 3460 35768 3466
rect 35716 3402 35768 3408
rect 35622 1728 35678 1737
rect 35622 1663 35678 1672
rect 35438 640 35494 649
rect 35438 575 35494 584
rect 36096 480 36124 4490
rect 36648 4049 36676 12543
rect 37186 4584 37242 4593
rect 37186 4519 37242 4528
rect 36634 4040 36690 4049
rect 36634 3975 36690 3984
rect 36820 3528 36872 3534
rect 36820 3470 36872 3476
rect 36544 3392 36596 3398
rect 36544 3334 36596 3340
rect 36556 2990 36584 3334
rect 36832 3194 36860 3470
rect 36820 3188 36872 3194
rect 36820 3130 36872 3136
rect 36544 2984 36596 2990
rect 36544 2926 36596 2932
rect 36556 2650 36584 2926
rect 36544 2644 36596 2650
rect 36544 2586 36596 2592
rect 37200 480 37228 4519
rect 39394 4040 39450 4049
rect 39394 3975 39450 3984
rect 37370 3632 37426 3641
rect 37370 3567 37426 3576
rect 37384 3194 37412 3567
rect 37372 3188 37424 3194
rect 37372 3130 37424 3136
rect 38290 2816 38346 2825
rect 38290 2751 38346 2760
rect 38304 480 38332 2751
rect 39408 480 39436 3975
rect 570 0 626 480
rect 1674 0 1730 480
rect 2778 0 2834 480
rect 3882 0 3938 480
rect 4986 0 5042 480
rect 6090 0 6146 480
rect 7194 0 7250 480
rect 8298 0 8354 480
rect 9402 0 9458 480
rect 10506 0 10562 480
rect 11610 0 11666 480
rect 12714 0 12770 480
rect 13910 0 13966 480
rect 15014 0 15070 480
rect 16118 0 16174 480
rect 17222 0 17278 480
rect 18326 0 18382 480
rect 19430 0 19486 480
rect 20534 0 20590 480
rect 21638 0 21694 480
rect 22742 0 22798 480
rect 23846 0 23902 480
rect 24950 0 25006 480
rect 26054 0 26110 480
rect 27250 0 27306 480
rect 28354 0 28410 480
rect 29458 0 29514 480
rect 30562 0 30618 480
rect 31666 0 31722 480
rect 32770 0 32826 480
rect 33874 0 33930 480
rect 34978 0 35034 480
rect 36082 0 36138 480
rect 37186 0 37242 480
rect 38290 0 38346 480
rect 39394 0 39450 480
<< via2 >>
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 9954 35128 10010 35184
rect 22742 35128 22798 35184
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 22374 27240 22430 27296
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 22650 26732 22652 26752
rect 22652 26732 22704 26752
rect 22704 26732 22706 26752
rect 22650 26696 22706 26732
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 9954 20576 10010 20632
rect 7378 20032 7434 20088
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 7562 16768 7618 16824
rect 5446 16632 5502 16688
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 7010 16632 7066 16688
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 9218 16632 9274 16688
rect 16486 18128 16542 18184
rect 9770 16768 9826 16824
rect 15290 16904 15346 16960
rect 11058 16632 11114 16688
rect 8942 15000 8998 15056
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 13266 13132 13268 13152
rect 13268 13132 13320 13152
rect 13320 13132 13322 13152
rect 13266 13096 13322 13132
rect 7838 9324 7840 9344
rect 7840 9324 7892 9344
rect 7892 9324 7894 9344
rect 7838 9288 7894 9324
rect 9402 9288 9458 9344
rect 8942 9152 8998 9208
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 5170 6976 5226 7032
rect 4894 6740 4896 6760
rect 4896 6740 4948 6760
rect 4948 6740 4950 6760
rect 4894 6704 4950 6740
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 7746 6996 7802 7032
rect 7746 6976 7748 6996
rect 7748 6976 7800 6996
rect 7800 6976 7802 6996
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 3054 4140 3110 4176
rect 3054 4120 3056 4140
rect 3056 4120 3108 4140
rect 3108 4120 3110 4140
rect 3330 3984 3386 4040
rect 2042 3712 2098 3768
rect 3790 3712 3846 3768
rect 3146 2644 3202 2680
rect 3146 2624 3148 2644
rect 3148 2624 3200 2644
rect 3200 2624 3202 2644
rect 2042 2508 2098 2544
rect 2042 2488 2044 2508
rect 2044 2488 2096 2508
rect 2096 2488 2098 2508
rect 5262 3848 5318 3904
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 4158 3068 4160 3088
rect 4160 3068 4212 3088
rect 4212 3068 4214 3088
rect 4158 3032 4214 3068
rect 4710 3032 4766 3088
rect 7194 5652 7196 5672
rect 7196 5652 7248 5672
rect 7248 5652 7250 5672
rect 7194 5616 7250 5652
rect 7470 5092 7526 5128
rect 7470 5072 7472 5092
rect 7472 5072 7524 5092
rect 7524 5072 7526 5092
rect 6090 4120 6146 4176
rect 5814 3440 5870 3496
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 4802 2080 4858 2136
rect 7930 4140 7986 4176
rect 7930 4120 7932 4140
rect 7932 4120 7984 4140
rect 7984 4120 7986 4140
rect 7286 3884 7288 3904
rect 7288 3884 7340 3904
rect 7340 3884 7342 3904
rect 7286 3848 7342 3884
rect 8482 4004 8538 4040
rect 8482 3984 8484 4004
rect 8484 3984 8536 4004
rect 8536 3984 8538 4004
rect 8390 3476 8392 3496
rect 8392 3476 8444 3496
rect 8444 3476 8446 3496
rect 8390 3440 8446 3476
rect 10414 9152 10470 9208
rect 9862 5228 9918 5264
rect 9862 5208 9864 5228
rect 9864 5208 9916 5228
rect 9916 5208 9918 5228
rect 9954 3984 10010 4040
rect 9770 3440 9826 3496
rect 10874 8492 10930 8528
rect 10874 8472 10876 8492
rect 10876 8472 10928 8492
rect 10928 8472 10930 8492
rect 10506 6180 10562 6216
rect 10506 6160 10508 6180
rect 10508 6160 10560 6180
rect 10560 6160 10562 6180
rect 10598 5364 10654 5400
rect 10598 5344 10600 5364
rect 10600 5344 10652 5364
rect 10652 5344 10654 5364
rect 10782 4936 10838 4992
rect 10506 4800 10562 4856
rect 10874 4664 10930 4720
rect 10506 3848 10562 3904
rect 10966 3596 11022 3632
rect 10966 3576 10968 3596
rect 10968 3576 11020 3596
rect 11020 3576 11022 3596
rect 12438 6160 12494 6216
rect 12162 5616 12218 5672
rect 12622 5208 12678 5264
rect 12530 4936 12586 4992
rect 13174 11056 13230 11112
rect 14002 13640 14058 13696
rect 13542 9696 13598 9752
rect 12898 4528 12954 4584
rect 12898 3884 12900 3904
rect 12900 3884 12952 3904
rect 12952 3884 12954 3904
rect 12898 3848 12954 3884
rect 13082 4972 13084 4992
rect 13084 4972 13136 4992
rect 13136 4972 13138 4992
rect 13082 4936 13138 4972
rect 12622 3304 12678 3360
rect 11702 2760 11758 2816
rect 12622 2488 12678 2544
rect 13818 8508 13820 8528
rect 13820 8508 13872 8528
rect 13872 8508 13874 8528
rect 13818 8472 13874 8508
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 20534 20304 20590 20360
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 20902 19896 20958 19952
rect 22466 20340 22468 20360
rect 22468 20340 22520 20360
rect 22520 20340 22522 20360
rect 22466 20304 22522 20340
rect 21362 20168 21418 20224
rect 21270 20052 21326 20088
rect 21270 20032 21272 20052
rect 21272 20032 21324 20052
rect 21324 20032 21326 20052
rect 20994 19236 21050 19272
rect 20994 19216 20996 19236
rect 20996 19216 21048 19236
rect 21048 19216 21050 19236
rect 17038 16632 17094 16688
rect 19890 18128 19946 18184
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 19982 17620 19984 17640
rect 19984 17620 20036 17640
rect 20036 17620 20038 17640
rect 19982 17584 20038 17620
rect 18418 16940 18420 16960
rect 18420 16940 18472 16960
rect 18472 16940 18474 16960
rect 18418 16904 18474 16940
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 17498 15680 17554 15736
rect 16118 15136 16174 15192
rect 14554 13640 14610 13696
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 19430 15680 19486 15736
rect 20810 16652 20866 16688
rect 20810 16632 20812 16652
rect 20812 16632 20864 16652
rect 20864 16632 20866 16652
rect 22374 18944 22430 19000
rect 35714 39344 35770 39400
rect 35622 38120 35678 38176
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 37554 36896 37610 36952
rect 33966 35672 34022 35728
rect 28354 34584 28410 34640
rect 29918 34584 29974 34640
rect 23846 27104 23902 27160
rect 26514 27276 26516 27296
rect 26516 27276 26568 27296
rect 26568 27276 26570 27296
rect 26514 27240 26570 27276
rect 26422 27124 26478 27160
rect 26422 27104 26424 27124
rect 26424 27104 26476 27124
rect 26476 27104 26478 27124
rect 26606 26732 26608 26752
rect 26608 26732 26660 26752
rect 26660 26732 26662 26752
rect 26606 26696 26662 26732
rect 27158 26324 27160 26344
rect 27160 26324 27212 26344
rect 27212 26324 27214 26344
rect 27158 26288 27214 26324
rect 24582 24792 24638 24848
rect 27618 24792 27674 24848
rect 24674 23568 24730 23624
rect 24214 21392 24270 21448
rect 24122 20168 24178 20224
rect 23846 20032 23902 20088
rect 24306 21120 24362 21176
rect 25594 21428 25596 21448
rect 25596 21428 25648 21448
rect 25648 21428 25650 21448
rect 25594 21392 25650 21428
rect 23662 19216 23718 19272
rect 25042 18964 25098 19000
rect 25042 18944 25044 18964
rect 25044 18944 25096 18964
rect 25096 18944 25098 18964
rect 22742 18400 22798 18456
rect 18786 14864 18842 14920
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 21546 16768 21602 16824
rect 22006 17584 22062 17640
rect 21914 16652 21970 16688
rect 21914 16632 21916 16652
rect 21916 16632 21968 16652
rect 21968 16632 21970 16652
rect 21638 14864 21694 14920
rect 16670 13640 16726 13696
rect 16210 13096 16266 13152
rect 17498 11056 17554 11112
rect 19154 11736 19210 11792
rect 18694 11056 18750 11112
rect 15566 9696 15622 9752
rect 17038 9580 17094 9616
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 23478 16788 23534 16824
rect 23478 16768 23480 16788
rect 23480 16768 23532 16788
rect 23532 16768 23534 16788
rect 22374 16632 22430 16688
rect 24030 16224 24086 16280
rect 23754 15988 23756 16008
rect 23756 15988 23808 16008
rect 23808 15988 23810 16008
rect 23754 15952 23810 15988
rect 26422 22480 26478 22536
rect 26698 21684 26754 21720
rect 26698 21664 26700 21684
rect 26700 21664 26752 21684
rect 26752 21664 26754 21684
rect 28078 23568 28134 23624
rect 34334 32172 34336 32192
rect 34336 32172 34388 32192
rect 34388 32172 34390 32192
rect 34334 32136 34390 32172
rect 32310 30368 32366 30424
rect 32310 29552 32366 29608
rect 32586 28464 32642 28520
rect 28722 26696 28778 26752
rect 30470 27240 30526 27296
rect 30286 26424 30342 26480
rect 29550 24112 29606 24168
rect 26514 18420 26570 18456
rect 26514 18400 26516 18420
rect 26516 18400 26568 18420
rect 26568 18400 26570 18420
rect 26514 16632 26570 16688
rect 26238 16244 26294 16280
rect 26238 16224 26240 16244
rect 26240 16224 26292 16244
rect 26292 16224 26294 16244
rect 25686 16088 25742 16144
rect 26054 15680 26110 15736
rect 27250 17856 27306 17912
rect 27158 16768 27214 16824
rect 28446 21392 28502 21448
rect 27986 20204 27988 20224
rect 27988 20204 28040 20224
rect 28040 20204 28042 20224
rect 27986 20168 28042 20204
rect 28078 19488 28134 19544
rect 27802 19216 27858 19272
rect 25594 13948 25596 13968
rect 25596 13948 25648 13968
rect 25648 13948 25650 13968
rect 25594 13912 25650 13948
rect 21914 12960 21970 13016
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 21730 12280 21786 12336
rect 20626 11736 20682 11792
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 20810 11076 20866 11112
rect 17038 9560 17040 9580
rect 17040 9560 17092 9580
rect 17092 9560 17094 9580
rect 20810 11056 20812 11076
rect 20812 11056 20864 11076
rect 20864 11056 20866 11076
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 20626 9560 20682 9616
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 17038 7248 17094 7304
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 13450 3848 13506 3904
rect 13358 3712 13414 3768
rect 13358 3304 13414 3360
rect 12990 2896 13046 2952
rect 12990 2624 13046 2680
rect 13910 2760 13966 2816
rect 14462 4528 14518 4584
rect 19154 7384 19210 7440
rect 17130 6432 17186 6488
rect 14922 4936 14978 4992
rect 15290 3848 15346 3904
rect 15658 4528 15714 4584
rect 16118 5344 16174 5400
rect 16946 5616 17002 5672
rect 15842 4392 15898 4448
rect 15750 4256 15806 4312
rect 17590 5344 17646 5400
rect 16394 4800 16450 4856
rect 16762 4800 16818 4856
rect 16302 4548 16358 4584
rect 16302 4528 16304 4548
rect 16304 4528 16356 4548
rect 16356 4528 16358 4548
rect 16578 4664 16634 4720
rect 16762 4020 16764 4040
rect 16764 4020 16816 4040
rect 16816 4020 16818 4040
rect 16762 3984 16818 4020
rect 16854 3848 16910 3904
rect 16946 3576 17002 3632
rect 17406 4256 17462 4312
rect 17222 3440 17278 3496
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 20074 7248 20130 7304
rect 19430 6452 19486 6488
rect 19430 6432 19432 6452
rect 19432 6432 19484 6452
rect 19484 6432 19486 6452
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 19430 5616 19486 5672
rect 17498 3188 17554 3224
rect 17498 3168 17500 3188
rect 17500 3168 17552 3188
rect 17552 3168 17554 3188
rect 18234 4800 18290 4856
rect 18694 4564 18696 4584
rect 18696 4564 18748 4584
rect 18748 4564 18750 4584
rect 18694 4528 18750 4564
rect 19338 4800 19394 4856
rect 20626 5364 20682 5400
rect 21546 9560 21602 9616
rect 26698 15000 26754 15056
rect 26882 13504 26938 13560
rect 25686 12980 25742 13016
rect 25686 12960 25688 12980
rect 25688 12960 25740 12980
rect 25740 12960 25742 12980
rect 24398 12552 24454 12608
rect 27434 12824 27490 12880
rect 29734 23588 29790 23624
rect 29734 23568 29736 23588
rect 29736 23568 29788 23588
rect 29788 23568 29790 23588
rect 30470 26288 30526 26344
rect 32126 26696 32182 26752
rect 32310 26424 32366 26480
rect 33598 29144 33654 29200
rect 34518 30368 34574 30424
rect 34702 29688 34758 29744
rect 30930 25880 30986 25936
rect 30654 24656 30710 24712
rect 29274 21664 29330 21720
rect 33874 26832 33930 26888
rect 34426 26968 34482 27024
rect 34702 27512 34758 27568
rect 33046 23568 33102 23624
rect 31758 21800 31814 21856
rect 30194 20712 30250 20768
rect 30746 20596 30802 20632
rect 30746 20576 30748 20596
rect 30748 20576 30800 20596
rect 30800 20576 30802 20596
rect 30562 18300 30564 18320
rect 30564 18300 30616 18320
rect 30616 18300 30618 18320
rect 30562 18264 30618 18300
rect 27894 16108 27950 16144
rect 27894 16088 27896 16108
rect 27896 16088 27948 16108
rect 27948 16088 27950 16108
rect 27802 15136 27858 15192
rect 27710 12280 27766 12336
rect 21086 7384 21142 7440
rect 20902 5652 20904 5672
rect 20904 5652 20956 5672
rect 20956 5652 20958 5672
rect 20902 5616 20958 5652
rect 20626 5344 20628 5364
rect 20628 5344 20680 5364
rect 20680 5344 20682 5364
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 19706 4392 19762 4448
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 20350 4428 20352 4448
rect 20352 4428 20404 4448
rect 20404 4428 20406 4448
rect 20350 4392 20406 4428
rect 19246 3032 19302 3088
rect 20074 3168 20130 3224
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 21730 8336 21786 8392
rect 21546 5344 21602 5400
rect 21086 2624 21142 2680
rect 29366 16788 29422 16824
rect 29366 16768 29368 16788
rect 29368 16768 29420 16788
rect 29420 16768 29422 16788
rect 29550 16652 29606 16688
rect 29550 16632 29552 16652
rect 29552 16632 29604 16652
rect 29604 16632 29606 16652
rect 31482 17856 31538 17912
rect 32126 21528 32182 21584
rect 31850 20712 31906 20768
rect 34334 21800 34390 21856
rect 32770 20440 32826 20496
rect 32126 19488 32182 19544
rect 33138 19252 33140 19272
rect 33140 19252 33192 19272
rect 33192 19252 33194 19272
rect 33138 19216 33194 19252
rect 32218 18028 32220 18048
rect 32220 18028 32272 18048
rect 32272 18028 32274 18048
rect 32218 17992 32274 18028
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 35346 32136 35402 32192
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 36818 34448 36874 34504
rect 36726 33224 36782 33280
rect 35990 32000 36046 32056
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 35530 30776 35586 30832
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 35346 27240 35402 27296
rect 35714 29552 35770 29608
rect 35622 29008 35678 29064
rect 35254 24656 35310 24712
rect 34886 24556 34888 24576
rect 34888 24556 34940 24576
rect 34940 24556 34942 24576
rect 34886 24520 34942 24556
rect 35254 24520 35310 24576
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 34518 17992 34574 18048
rect 31666 15564 31722 15600
rect 31666 15544 31668 15564
rect 31668 15544 31720 15564
rect 31720 15544 31722 15564
rect 29734 13912 29790 13968
rect 29458 13524 29514 13560
rect 29458 13504 29460 13524
rect 29460 13504 29512 13524
rect 29512 13504 29514 13524
rect 23662 9596 23664 9616
rect 23664 9596 23716 9616
rect 23716 9596 23718 9616
rect 23662 9560 23718 9596
rect 24030 8336 24086 8392
rect 22006 4800 22062 4856
rect 22190 4392 22246 4448
rect 22650 4256 22706 4312
rect 22374 2796 22376 2816
rect 22376 2796 22428 2816
rect 22428 2796 22430 2816
rect 22374 2760 22430 2796
rect 23110 4936 23166 4992
rect 24030 5616 24086 5672
rect 23294 3732 23350 3768
rect 23294 3712 23296 3732
rect 23296 3712 23348 3732
rect 23348 3712 23350 3732
rect 24306 4820 24362 4856
rect 24306 4800 24308 4820
rect 24308 4800 24360 4820
rect 24360 4800 24362 4820
rect 24674 4256 24730 4312
rect 25042 4972 25044 4992
rect 25044 4972 25096 4992
rect 25096 4972 25098 4992
rect 25042 4936 25098 4972
rect 25318 4936 25374 4992
rect 27250 5616 27306 5672
rect 25870 4528 25926 4584
rect 25318 3732 25374 3768
rect 25318 3712 25320 3732
rect 25320 3712 25372 3732
rect 25372 3712 25374 3732
rect 24766 3168 24822 3224
rect 24490 2644 24546 2680
rect 24490 2624 24492 2644
rect 24492 2624 24544 2644
rect 24544 2624 24546 2644
rect 24030 2352 24086 2408
rect 24030 2080 24086 2136
rect 25962 2644 26018 2680
rect 27158 3188 27214 3224
rect 27158 3168 27160 3188
rect 27160 3168 27212 3188
rect 27212 3168 27214 3188
rect 25962 2624 25964 2644
rect 25964 2624 26016 2644
rect 26016 2624 26018 2644
rect 25778 2508 25834 2544
rect 25778 2488 25780 2508
rect 25780 2488 25832 2508
rect 25832 2488 25834 2508
rect 33690 14900 33692 14920
rect 33692 14900 33744 14920
rect 33744 14900 33746 14920
rect 33690 14864 33746 14900
rect 29826 12844 29882 12880
rect 29826 12824 29828 12844
rect 29828 12824 29880 12844
rect 29880 12824 29882 12844
rect 33874 13948 33876 13968
rect 33876 13948 33928 13968
rect 33928 13948 33930 13968
rect 33874 13912 33930 13948
rect 34242 12416 34298 12472
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 35530 24792 35586 24848
rect 35898 29008 35954 29064
rect 36266 29180 36268 29200
rect 36268 29180 36320 29200
rect 36320 29180 36322 29200
rect 36266 29144 36322 29180
rect 35346 21548 35402 21584
rect 35346 21528 35348 21548
rect 35348 21528 35400 21548
rect 35400 21528 35402 21548
rect 35346 21120 35402 21176
rect 35438 20712 35494 20768
rect 35254 19216 35310 19272
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 35438 18672 35494 18728
rect 35346 17448 35402 17504
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 35346 15952 35402 16008
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 34610 12416 34666 12472
rect 29734 5888 29790 5944
rect 27710 4800 27766 4856
rect 27986 4664 28042 4720
rect 27894 4548 27950 4584
rect 27894 4528 27896 4548
rect 27896 4528 27948 4548
rect 27948 4528 27950 4548
rect 27342 3304 27398 3360
rect 31942 5888 31998 5944
rect 30838 4972 30840 4992
rect 30840 4972 30892 4992
rect 30892 4972 30894 4992
rect 30838 4936 30894 4972
rect 30654 4800 30710 4856
rect 29182 3848 29238 3904
rect 28354 3304 28410 3360
rect 28262 2624 28318 2680
rect 28170 2488 28226 2544
rect 29458 3712 29514 3768
rect 31298 4664 31354 4720
rect 31206 4528 31262 4584
rect 32126 3884 32128 3904
rect 32128 3884 32180 3904
rect 32180 3884 32182 3904
rect 32126 3848 32182 3884
rect 31850 3712 31906 3768
rect 31666 2896 31722 2952
rect 30562 1944 30618 2000
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 32678 4120 32734 4176
rect 32494 3576 32550 3632
rect 33966 5652 33968 5672
rect 33968 5652 34020 5672
rect 34020 5652 34022 5672
rect 33966 5616 34022 5652
rect 32770 3440 32826 3496
rect 32310 2760 32366 2816
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 34794 10104 34850 10160
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 34794 9016 34850 9072
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 34794 5072 34850 5128
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 34610 3712 34666 3768
rect 35438 11464 35494 11520
rect 35806 23568 35862 23624
rect 35990 22480 36046 22536
rect 36174 26832 36230 26888
rect 36818 27004 36820 27024
rect 36820 27004 36872 27024
rect 36872 27004 36874 27024
rect 36818 26968 36874 27004
rect 36818 24112 36874 24168
rect 35714 18264 35770 18320
rect 35622 17604 35678 17640
rect 35622 17584 35624 17604
rect 35624 17584 35676 17604
rect 35676 17584 35678 17604
rect 35622 12416 35678 12472
rect 35622 10240 35678 10296
rect 35530 7792 35586 7848
rect 35346 4120 35402 4176
rect 35714 6568 35770 6624
rect 37830 24520 37886 24576
rect 38014 22344 38070 22400
rect 37186 21120 37242 21176
rect 37094 20712 37150 20768
rect 36634 20476 36636 20496
rect 36636 20476 36688 20496
rect 36688 20476 36690 20496
rect 36634 20440 36690 20476
rect 36542 15544 36598 15600
rect 37094 15000 37150 15056
rect 36818 14864 36874 14920
rect 36634 12552 36690 12608
rect 35806 5344 35862 5400
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 34794 3032 34850 3088
rect 34702 2896 34758 2952
rect 34426 2796 34428 2816
rect 34428 2796 34480 2816
rect 34480 2796 34482 2816
rect 34426 2760 34482 2796
rect 33874 2352 33930 2408
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
rect 35622 1672 35678 1728
rect 35438 584 35494 640
rect 37186 4528 37242 4584
rect 36634 3984 36690 4040
rect 39394 3984 39450 4040
rect 37370 3576 37426 3632
rect 38290 2760 38346 2816
<< metal3 >>
rect 35709 39402 35775 39405
rect 39520 39402 40000 39432
rect 35709 39400 40000 39402
rect 35709 39344 35714 39400
rect 35770 39344 40000 39400
rect 35709 39342 40000 39344
rect 35709 39339 35775 39342
rect 39520 39312 40000 39342
rect 35617 38178 35683 38181
rect 39520 38178 40000 38208
rect 35617 38176 40000 38178
rect 35617 38120 35622 38176
rect 35678 38120 40000 38176
rect 35617 38118 40000 38120
rect 35617 38115 35683 38118
rect 39520 38088 40000 38118
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 37549 36954 37615 36957
rect 39520 36954 40000 36984
rect 37549 36952 40000 36954
rect 37549 36896 37554 36952
rect 37610 36896 40000 36952
rect 37549 36894 40000 36896
rect 37549 36891 37615 36894
rect 39520 36864 40000 36894
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 35871 35248 35872
rect 33961 35730 34027 35733
rect 39520 35730 40000 35760
rect 33961 35728 40000 35730
rect 33961 35672 33966 35728
rect 34022 35672 40000 35728
rect 33961 35670 40000 35672
rect 33961 35667 34027 35670
rect 39520 35640 40000 35670
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 9949 35186 10015 35189
rect 22737 35186 22803 35189
rect 9949 35184 22803 35186
rect 9949 35128 9954 35184
rect 10010 35128 22742 35184
rect 22798 35128 22803 35184
rect 9949 35126 22803 35128
rect 9949 35123 10015 35126
rect 22737 35123 22803 35126
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 28349 34642 28415 34645
rect 29913 34642 29979 34645
rect 28349 34640 29979 34642
rect 28349 34584 28354 34640
rect 28410 34584 29918 34640
rect 29974 34584 29979 34640
rect 28349 34582 29979 34584
rect 28349 34579 28415 34582
rect 29913 34579 29979 34582
rect 36813 34506 36879 34509
rect 39520 34506 40000 34536
rect 36813 34504 40000 34506
rect 36813 34448 36818 34504
rect 36874 34448 40000 34504
rect 36813 34446 40000 34448
rect 36813 34443 36879 34446
rect 39520 34416 40000 34446
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 0 33328 480 33448
rect 36721 33282 36787 33285
rect 39520 33282 40000 33312
rect 36721 33280 40000 33282
rect 36721 33224 36726 33280
rect 36782 33224 40000 33280
rect 36721 33222 40000 33224
rect 36721 33219 36787 33222
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 39520 33192 40000 33222
rect 19568 33151 19888 33152
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 34329 32194 34395 32197
rect 35341 32194 35407 32197
rect 34329 32192 35407 32194
rect 34329 32136 34334 32192
rect 34390 32136 35346 32192
rect 35402 32136 35407 32192
rect 34329 32134 35407 32136
rect 34329 32131 34395 32134
rect 35341 32131 35407 32134
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 35985 32058 36051 32061
rect 39520 32058 40000 32088
rect 35985 32056 40000 32058
rect 35985 32000 35990 32056
rect 36046 32000 40000 32056
rect 35985 31998 40000 32000
rect 35985 31995 36051 31998
rect 39520 31968 40000 31998
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 31519 35248 31520
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 35525 30834 35591 30837
rect 39520 30834 40000 30864
rect 35525 30832 40000 30834
rect 35525 30776 35530 30832
rect 35586 30776 40000 30832
rect 35525 30774 40000 30776
rect 35525 30771 35591 30774
rect 39520 30744 40000 30774
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 32305 30426 32371 30429
rect 34513 30426 34579 30429
rect 32305 30424 34579 30426
rect 32305 30368 32310 30424
rect 32366 30368 34518 30424
rect 34574 30368 34579 30424
rect 32305 30366 34579 30368
rect 32305 30363 32371 30366
rect 34513 30363 34579 30366
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 34697 29746 34763 29749
rect 34697 29744 36002 29746
rect 34697 29688 34702 29744
rect 34758 29688 36002 29744
rect 34697 29686 36002 29688
rect 34697 29683 34763 29686
rect 32305 29610 32371 29613
rect 35709 29610 35775 29613
rect 32305 29608 35775 29610
rect 32305 29552 32310 29608
rect 32366 29552 35714 29608
rect 35770 29552 35775 29608
rect 32305 29550 35775 29552
rect 35942 29610 36002 29686
rect 39520 29610 40000 29640
rect 35942 29550 40000 29610
rect 32305 29547 32371 29550
rect 35709 29547 35775 29550
rect 39520 29520 40000 29550
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 33593 29202 33659 29205
rect 36261 29202 36327 29205
rect 33593 29200 36327 29202
rect 33593 29144 33598 29200
rect 33654 29144 36266 29200
rect 36322 29144 36327 29200
rect 33593 29142 36327 29144
rect 33593 29139 33659 29142
rect 36261 29139 36327 29142
rect 35617 29066 35683 29069
rect 35893 29066 35959 29069
rect 35617 29064 35959 29066
rect 35617 29008 35622 29064
rect 35678 29008 35898 29064
rect 35954 29008 35959 29064
rect 35617 29006 35959 29008
rect 35617 29003 35683 29006
rect 35893 29003 35959 29006
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 32581 28522 32647 28525
rect 32581 28520 35404 28522
rect 32581 28464 32586 28520
rect 32642 28464 35404 28520
rect 32581 28462 35404 28464
rect 32581 28459 32647 28462
rect 35344 28386 35404 28462
rect 39520 28386 40000 28416
rect 35344 28326 40000 28386
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 39520 28296 40000 28326
rect 34928 28255 35248 28256
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 34697 27570 34763 27573
rect 34654 27568 34763 27570
rect 34654 27512 34702 27568
rect 34758 27512 34763 27568
rect 34654 27507 34763 27512
rect 22369 27298 22435 27301
rect 26509 27298 26575 27301
rect 22369 27296 26575 27298
rect 22369 27240 22374 27296
rect 22430 27240 26514 27296
rect 26570 27240 26575 27296
rect 22369 27238 26575 27240
rect 22369 27235 22435 27238
rect 26509 27235 26575 27238
rect 30465 27298 30531 27301
rect 34654 27298 34714 27507
rect 30465 27296 34714 27298
rect 30465 27240 30470 27296
rect 30526 27240 34714 27296
rect 30465 27238 34714 27240
rect 35341 27298 35407 27301
rect 39520 27298 40000 27328
rect 35341 27296 40000 27298
rect 35341 27240 35346 27296
rect 35402 27240 40000 27296
rect 35341 27238 40000 27240
rect 30465 27235 30531 27238
rect 35341 27235 35407 27238
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 39520 27208 40000 27238
rect 34928 27167 35248 27168
rect 23841 27162 23907 27165
rect 26417 27162 26483 27165
rect 23841 27160 26483 27162
rect 23841 27104 23846 27160
rect 23902 27104 26422 27160
rect 26478 27104 26483 27160
rect 23841 27102 26483 27104
rect 23841 27099 23907 27102
rect 26417 27099 26483 27102
rect 34421 27026 34487 27029
rect 36813 27026 36879 27029
rect 34421 27024 36879 27026
rect 34421 26968 34426 27024
rect 34482 26968 36818 27024
rect 36874 26968 36879 27024
rect 34421 26966 36879 26968
rect 34421 26963 34487 26966
rect 36813 26963 36879 26966
rect 33869 26890 33935 26893
rect 36169 26890 36235 26893
rect 33869 26888 36235 26890
rect 33869 26832 33874 26888
rect 33930 26832 36174 26888
rect 36230 26832 36235 26888
rect 33869 26830 36235 26832
rect 33869 26827 33935 26830
rect 36169 26827 36235 26830
rect 22645 26754 22711 26757
rect 26601 26754 26667 26757
rect 22645 26752 26667 26754
rect 22645 26696 22650 26752
rect 22706 26696 26606 26752
rect 26662 26696 26667 26752
rect 22645 26694 26667 26696
rect 22645 26691 22711 26694
rect 26601 26691 26667 26694
rect 28717 26754 28783 26757
rect 32121 26754 32187 26757
rect 28717 26752 32187 26754
rect 28717 26696 28722 26752
rect 28778 26696 32126 26752
rect 32182 26696 32187 26752
rect 28717 26694 32187 26696
rect 28717 26691 28783 26694
rect 32121 26691 32187 26694
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 30281 26482 30347 26485
rect 32305 26482 32371 26485
rect 30281 26480 32371 26482
rect 30281 26424 30286 26480
rect 30342 26424 32310 26480
rect 32366 26424 32371 26480
rect 30281 26422 32371 26424
rect 30281 26419 30347 26422
rect 32305 26419 32371 26422
rect 27153 26346 27219 26349
rect 30465 26346 30531 26349
rect 27153 26344 30531 26346
rect 27153 26288 27158 26344
rect 27214 26288 30470 26344
rect 30526 26288 30531 26344
rect 27153 26286 30531 26288
rect 27153 26283 27219 26286
rect 30465 26283 30531 26286
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 26079 35248 26080
rect 39520 26074 40000 26104
rect 35574 26014 40000 26074
rect 30925 25938 30991 25941
rect 35574 25938 35634 26014
rect 39520 25984 40000 26014
rect 30925 25936 35634 25938
rect 30925 25880 30930 25936
rect 30986 25880 35634 25936
rect 30925 25878 35634 25880
rect 30925 25875 30991 25878
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 24577 24850 24643 24853
rect 27613 24850 27679 24853
rect 24577 24848 27679 24850
rect 24577 24792 24582 24848
rect 24638 24792 27618 24848
rect 27674 24792 27679 24848
rect 24577 24790 27679 24792
rect 24577 24787 24643 24790
rect 27613 24787 27679 24790
rect 35525 24850 35591 24853
rect 39520 24850 40000 24880
rect 35525 24848 40000 24850
rect 35525 24792 35530 24848
rect 35586 24792 40000 24848
rect 35525 24790 40000 24792
rect 35525 24787 35591 24790
rect 39520 24760 40000 24790
rect 30649 24714 30715 24717
rect 35249 24714 35315 24717
rect 30649 24712 35315 24714
rect 30649 24656 30654 24712
rect 30710 24656 35254 24712
rect 35310 24656 35315 24712
rect 30649 24654 35315 24656
rect 30649 24651 30715 24654
rect 35249 24651 35315 24654
rect 34881 24578 34947 24581
rect 35249 24578 35315 24581
rect 37825 24578 37891 24581
rect 34881 24576 37891 24578
rect 34881 24520 34886 24576
rect 34942 24520 35254 24576
rect 35310 24520 37830 24576
rect 37886 24520 37891 24576
rect 34881 24518 37891 24520
rect 34881 24515 34947 24518
rect 35249 24515 35315 24518
rect 37825 24515 37891 24518
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 29545 24170 29611 24173
rect 36813 24170 36879 24173
rect 29545 24168 36879 24170
rect 29545 24112 29550 24168
rect 29606 24112 36818 24168
rect 36874 24112 36879 24168
rect 29545 24110 36879 24112
rect 29545 24107 29611 24110
rect 36813 24107 36879 24110
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 24669 23626 24735 23629
rect 28073 23626 28139 23629
rect 24669 23624 28139 23626
rect 24669 23568 24674 23624
rect 24730 23568 28078 23624
rect 28134 23568 28139 23624
rect 24669 23566 28139 23568
rect 24669 23563 24735 23566
rect 28073 23563 28139 23566
rect 29729 23626 29795 23629
rect 33041 23626 33107 23629
rect 29729 23624 33107 23626
rect 29729 23568 29734 23624
rect 29790 23568 33046 23624
rect 33102 23568 33107 23624
rect 29729 23566 33107 23568
rect 29729 23563 29795 23566
rect 33041 23563 33107 23566
rect 35801 23626 35867 23629
rect 39520 23626 40000 23656
rect 35801 23624 40000 23626
rect 35801 23568 35806 23624
rect 35862 23568 40000 23624
rect 35801 23566 40000 23568
rect 35801 23563 35867 23566
rect 39520 23536 40000 23566
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 22815 35248 22816
rect 26417 22538 26483 22541
rect 35985 22538 36051 22541
rect 26417 22536 36051 22538
rect 26417 22480 26422 22536
rect 26478 22480 35990 22536
rect 36046 22480 36051 22536
rect 26417 22478 36051 22480
rect 26417 22475 26483 22478
rect 35985 22475 36051 22478
rect 38009 22402 38075 22405
rect 39520 22402 40000 22432
rect 38009 22400 40000 22402
rect 38009 22344 38014 22400
rect 38070 22344 40000 22400
rect 38009 22342 40000 22344
rect 38009 22339 38075 22342
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 39520 22312 40000 22342
rect 19568 22271 19888 22272
rect 31753 21858 31819 21861
rect 34329 21858 34395 21861
rect 31753 21856 34395 21858
rect 31753 21800 31758 21856
rect 31814 21800 34334 21856
rect 34390 21800 34395 21856
rect 31753 21798 34395 21800
rect 31753 21795 31819 21798
rect 34329 21795 34395 21798
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 21727 35248 21728
rect 26693 21722 26759 21725
rect 29269 21722 29335 21725
rect 26693 21720 29335 21722
rect 26693 21664 26698 21720
rect 26754 21664 29274 21720
rect 29330 21664 29335 21720
rect 26693 21662 29335 21664
rect 26693 21659 26759 21662
rect 29269 21659 29335 21662
rect 32121 21586 32187 21589
rect 35341 21586 35407 21589
rect 32121 21584 35407 21586
rect 32121 21528 32126 21584
rect 32182 21528 35346 21584
rect 35402 21528 35407 21584
rect 32121 21526 35407 21528
rect 32121 21523 32187 21526
rect 35341 21523 35407 21526
rect 24209 21450 24275 21453
rect 25589 21450 25655 21453
rect 28441 21450 28507 21453
rect 24209 21448 28507 21450
rect 24209 21392 24214 21448
rect 24270 21392 25594 21448
rect 25650 21392 28446 21448
rect 28502 21392 28507 21448
rect 24209 21390 28507 21392
rect 24209 21387 24275 21390
rect 25589 21387 25655 21390
rect 28441 21387 28507 21390
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 24301 21178 24367 21181
rect 35341 21178 35407 21181
rect 24301 21176 35407 21178
rect 24301 21120 24306 21176
rect 24362 21120 35346 21176
rect 35402 21120 35407 21176
rect 24301 21118 35407 21120
rect 24301 21115 24367 21118
rect 35341 21115 35407 21118
rect 37181 21178 37247 21181
rect 39520 21178 40000 21208
rect 37181 21176 40000 21178
rect 37181 21120 37186 21176
rect 37242 21120 40000 21176
rect 37181 21118 40000 21120
rect 37181 21115 37247 21118
rect 39520 21088 40000 21118
rect 30189 20770 30255 20773
rect 31845 20770 31911 20773
rect 30189 20768 31911 20770
rect 30189 20712 30194 20768
rect 30250 20712 31850 20768
rect 31906 20712 31911 20768
rect 30189 20710 31911 20712
rect 30189 20707 30255 20710
rect 31845 20707 31911 20710
rect 35433 20770 35499 20773
rect 37089 20770 37155 20773
rect 35433 20768 37155 20770
rect 35433 20712 35438 20768
rect 35494 20712 37094 20768
rect 37150 20712 37155 20768
rect 35433 20710 37155 20712
rect 35433 20707 35499 20710
rect 37089 20707 37155 20710
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 9949 20634 10015 20637
rect 30741 20634 30807 20637
rect 9949 20632 30807 20634
rect 9949 20576 9954 20632
rect 10010 20576 30746 20632
rect 30802 20576 30807 20632
rect 9949 20574 30807 20576
rect 9949 20571 10015 20574
rect 30741 20571 30807 20574
rect 32765 20498 32831 20501
rect 36629 20498 36695 20501
rect 32765 20496 36695 20498
rect 32765 20440 32770 20496
rect 32826 20440 36634 20496
rect 36690 20440 36695 20496
rect 32765 20438 36695 20440
rect 32765 20435 32831 20438
rect 36629 20435 36695 20438
rect 20529 20362 20595 20365
rect 22461 20362 22527 20365
rect 20529 20360 22527 20362
rect 20529 20304 20534 20360
rect 20590 20304 22466 20360
rect 22522 20304 22527 20360
rect 20529 20302 22527 20304
rect 20529 20299 20595 20302
rect 22461 20299 22527 20302
rect 21357 20226 21423 20229
rect 24117 20226 24183 20229
rect 27981 20226 28047 20229
rect 21357 20224 28047 20226
rect 21357 20168 21362 20224
rect 21418 20168 24122 20224
rect 24178 20168 27986 20224
rect 28042 20168 28047 20224
rect 21357 20166 28047 20168
rect 21357 20163 21423 20166
rect 24117 20163 24183 20166
rect 27981 20163 28047 20166
rect 19568 20160 19888 20161
rect 0 20090 480 20120
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 7373 20090 7439 20093
rect 0 20088 7439 20090
rect 0 20032 7378 20088
rect 7434 20032 7439 20088
rect 0 20030 7439 20032
rect 0 20000 480 20030
rect 7373 20027 7439 20030
rect 21265 20090 21331 20093
rect 23841 20090 23907 20093
rect 21265 20088 23907 20090
rect 21265 20032 21270 20088
rect 21326 20032 23846 20088
rect 23902 20032 23907 20088
rect 21265 20030 23907 20032
rect 21265 20027 21331 20030
rect 23841 20027 23907 20030
rect 20897 19954 20963 19957
rect 39520 19954 40000 19984
rect 20897 19952 22386 19954
rect 20897 19896 20902 19952
rect 20958 19896 22386 19952
rect 20897 19894 22386 19896
rect 20897 19891 20963 19894
rect 22326 19818 22386 19894
rect 34286 19894 40000 19954
rect 31526 19818 31770 19852
rect 34286 19818 34346 19894
rect 39520 19864 40000 19894
rect 22326 19792 34346 19818
rect 22326 19758 31586 19792
rect 31710 19758 34346 19792
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 28073 19546 28139 19549
rect 32121 19546 32187 19549
rect 28073 19544 32187 19546
rect 28073 19488 28078 19544
rect 28134 19488 32126 19544
rect 32182 19488 32187 19544
rect 28073 19486 32187 19488
rect 28073 19483 28139 19486
rect 32121 19483 32187 19486
rect 20989 19274 21055 19277
rect 23657 19274 23723 19277
rect 20989 19272 23723 19274
rect 20989 19216 20994 19272
rect 21050 19216 23662 19272
rect 23718 19216 23723 19272
rect 20989 19214 23723 19216
rect 20989 19211 21055 19214
rect 23657 19211 23723 19214
rect 27797 19274 27863 19277
rect 33133 19274 33199 19277
rect 27797 19272 33199 19274
rect 27797 19216 27802 19272
rect 27858 19216 33138 19272
rect 33194 19216 33199 19272
rect 27797 19214 33199 19216
rect 27797 19211 27863 19214
rect 33133 19211 33199 19214
rect 34646 19212 34652 19276
rect 34716 19274 34722 19276
rect 35249 19274 35315 19277
rect 34716 19272 35315 19274
rect 34716 19216 35254 19272
rect 35310 19216 35315 19272
rect 34716 19214 35315 19216
rect 34716 19212 34722 19214
rect 35249 19211 35315 19214
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 22369 19002 22435 19005
rect 25037 19002 25103 19005
rect 22369 19000 25103 19002
rect 22369 18944 22374 19000
rect 22430 18944 25042 19000
rect 25098 18944 25103 19000
rect 22369 18942 25103 18944
rect 22369 18939 22435 18942
rect 25037 18939 25103 18942
rect 35433 18730 35499 18733
rect 39520 18730 40000 18760
rect 35433 18728 40000 18730
rect 35433 18672 35438 18728
rect 35494 18672 40000 18728
rect 35433 18670 40000 18672
rect 35433 18667 35499 18670
rect 39520 18640 40000 18670
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 22737 18458 22803 18461
rect 26509 18458 26575 18461
rect 22737 18456 26575 18458
rect 22737 18400 22742 18456
rect 22798 18400 26514 18456
rect 26570 18400 26575 18456
rect 22737 18398 26575 18400
rect 22737 18395 22803 18398
rect 26509 18395 26575 18398
rect 30557 18322 30623 18325
rect 35709 18322 35775 18325
rect 30557 18320 35775 18322
rect 30557 18264 30562 18320
rect 30618 18264 35714 18320
rect 35770 18264 35775 18320
rect 30557 18262 35775 18264
rect 30557 18259 30623 18262
rect 35709 18259 35775 18262
rect 16481 18186 16547 18189
rect 19885 18186 19951 18189
rect 16481 18184 19951 18186
rect 16481 18128 16486 18184
rect 16542 18128 19890 18184
rect 19946 18128 19951 18184
rect 16481 18126 19951 18128
rect 16481 18123 16547 18126
rect 19885 18123 19951 18126
rect 32213 18050 32279 18053
rect 34513 18050 34579 18053
rect 32213 18048 34579 18050
rect 32213 17992 32218 18048
rect 32274 17992 34518 18048
rect 34574 17992 34579 18048
rect 32213 17990 34579 17992
rect 32213 17987 32279 17990
rect 34513 17987 34579 17990
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 27245 17914 27311 17917
rect 31477 17914 31543 17917
rect 27245 17912 31543 17914
rect 27245 17856 27250 17912
rect 27306 17856 31482 17912
rect 31538 17856 31543 17912
rect 27245 17854 31543 17856
rect 27245 17851 27311 17854
rect 31477 17851 31543 17854
rect 19977 17642 20043 17645
rect 22001 17642 22067 17645
rect 35617 17642 35683 17645
rect 19977 17640 35683 17642
rect 19977 17584 19982 17640
rect 20038 17584 22006 17640
rect 22062 17584 35622 17640
rect 35678 17584 35683 17640
rect 19977 17582 35683 17584
rect 19977 17579 20043 17582
rect 22001 17579 22067 17582
rect 35617 17579 35683 17582
rect 35341 17506 35407 17509
rect 39520 17506 40000 17536
rect 35341 17504 40000 17506
rect 35341 17448 35346 17504
rect 35402 17448 40000 17504
rect 35341 17446 40000 17448
rect 35341 17443 35407 17446
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 39520 17416 40000 17446
rect 34928 17375 35248 17376
rect 15285 16962 15351 16965
rect 18413 16962 18479 16965
rect 15285 16960 18479 16962
rect 15285 16904 15290 16960
rect 15346 16904 18418 16960
rect 18474 16904 18479 16960
rect 15285 16902 18479 16904
rect 15285 16899 15351 16902
rect 18413 16899 18479 16902
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 7557 16826 7623 16829
rect 9765 16826 9831 16829
rect 7557 16824 9831 16826
rect 7557 16768 7562 16824
rect 7618 16768 9770 16824
rect 9826 16768 9831 16824
rect 7557 16766 9831 16768
rect 7557 16763 7623 16766
rect 9765 16763 9831 16766
rect 21541 16826 21607 16829
rect 23473 16826 23539 16829
rect 21541 16824 23539 16826
rect 21541 16768 21546 16824
rect 21602 16768 23478 16824
rect 23534 16768 23539 16824
rect 21541 16766 23539 16768
rect 21541 16763 21607 16766
rect 23473 16763 23539 16766
rect 27153 16826 27219 16829
rect 29361 16826 29427 16829
rect 27153 16824 29427 16826
rect 27153 16768 27158 16824
rect 27214 16768 29366 16824
rect 29422 16768 29427 16824
rect 27153 16766 29427 16768
rect 27153 16763 27219 16766
rect 29361 16763 29427 16766
rect 5441 16690 5507 16693
rect 7005 16690 7071 16693
rect 5441 16688 7071 16690
rect 5441 16632 5446 16688
rect 5502 16632 7010 16688
rect 7066 16632 7071 16688
rect 5441 16630 7071 16632
rect 5441 16627 5507 16630
rect 7005 16627 7071 16630
rect 9213 16690 9279 16693
rect 11053 16690 11119 16693
rect 9213 16688 11119 16690
rect 9213 16632 9218 16688
rect 9274 16632 11058 16688
rect 11114 16632 11119 16688
rect 9213 16630 11119 16632
rect 9213 16627 9279 16630
rect 11053 16627 11119 16630
rect 17033 16690 17099 16693
rect 20805 16690 20871 16693
rect 17033 16688 20871 16690
rect 17033 16632 17038 16688
rect 17094 16632 20810 16688
rect 20866 16632 20871 16688
rect 17033 16630 20871 16632
rect 17033 16627 17099 16630
rect 20805 16627 20871 16630
rect 21909 16690 21975 16693
rect 22369 16690 22435 16693
rect 21909 16688 22435 16690
rect 21909 16632 21914 16688
rect 21970 16632 22374 16688
rect 22430 16632 22435 16688
rect 21909 16630 22435 16632
rect 21909 16627 21975 16630
rect 22369 16627 22435 16630
rect 26509 16690 26575 16693
rect 29545 16690 29611 16693
rect 26509 16688 29611 16690
rect 26509 16632 26514 16688
rect 26570 16632 29550 16688
rect 29606 16632 29611 16688
rect 26509 16630 29611 16632
rect 26509 16627 26575 16630
rect 29545 16627 29611 16630
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 16287 35248 16288
rect 24025 16282 24091 16285
rect 26233 16282 26299 16285
rect 39520 16282 40000 16312
rect 24025 16280 26299 16282
rect 24025 16224 24030 16280
rect 24086 16224 26238 16280
rect 26294 16224 26299 16280
rect 24025 16222 26299 16224
rect 24025 16219 24091 16222
rect 26233 16219 26299 16222
rect 35574 16222 40000 16282
rect 25681 16146 25747 16149
rect 27889 16146 27955 16149
rect 25681 16144 27955 16146
rect 25681 16088 25686 16144
rect 25742 16088 27894 16144
rect 27950 16088 27955 16144
rect 25681 16086 27955 16088
rect 25681 16083 25747 16086
rect 27889 16083 27955 16086
rect 23749 16010 23815 16013
rect 35341 16010 35407 16013
rect 23749 16008 35407 16010
rect 23749 15952 23754 16008
rect 23810 15952 35346 16008
rect 35402 15952 35407 16008
rect 23749 15950 35407 15952
rect 23749 15947 23815 15950
rect 35341 15947 35407 15950
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 17493 15738 17559 15741
rect 19425 15738 19491 15741
rect 17493 15736 19491 15738
rect 17493 15680 17498 15736
rect 17554 15680 19430 15736
rect 19486 15680 19491 15736
rect 17493 15678 19491 15680
rect 17493 15675 17559 15678
rect 19425 15675 19491 15678
rect 26049 15738 26115 15741
rect 35574 15738 35634 16222
rect 39520 16192 40000 16222
rect 26049 15736 35634 15738
rect 26049 15680 26054 15736
rect 26110 15680 35634 15736
rect 26049 15678 35634 15680
rect 26049 15675 26115 15678
rect 31661 15602 31727 15605
rect 36537 15602 36603 15605
rect 31661 15600 36603 15602
rect 31661 15544 31666 15600
rect 31722 15544 36542 15600
rect 36598 15544 36603 15600
rect 31661 15542 36603 15544
rect 31661 15539 31727 15542
rect 36537 15539 36603 15542
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 15199 35248 15200
rect 16113 15194 16179 15197
rect 27797 15194 27863 15197
rect 16113 15192 27863 15194
rect 16113 15136 16118 15192
rect 16174 15136 27802 15192
rect 27858 15136 27863 15192
rect 16113 15134 27863 15136
rect 16113 15131 16179 15134
rect 27797 15131 27863 15134
rect 8937 15058 9003 15061
rect 26693 15058 26759 15061
rect 8937 15056 26759 15058
rect 8937 15000 8942 15056
rect 8998 15000 26698 15056
rect 26754 15000 26759 15056
rect 8937 14998 26759 15000
rect 8937 14995 9003 14998
rect 26693 14995 26759 14998
rect 37089 15058 37155 15061
rect 39520 15058 40000 15088
rect 37089 15056 40000 15058
rect 37089 15000 37094 15056
rect 37150 15000 40000 15056
rect 37089 14998 40000 15000
rect 37089 14995 37155 14998
rect 39520 14968 40000 14998
rect 18781 14922 18847 14925
rect 21633 14922 21699 14925
rect 18781 14920 21699 14922
rect 18781 14864 18786 14920
rect 18842 14864 21638 14920
rect 21694 14864 21699 14920
rect 18781 14862 21699 14864
rect 18781 14859 18847 14862
rect 21633 14859 21699 14862
rect 33685 14922 33751 14925
rect 36813 14922 36879 14925
rect 33685 14920 36879 14922
rect 33685 14864 33690 14920
rect 33746 14864 36818 14920
rect 36874 14864 36879 14920
rect 33685 14862 36879 14864
rect 33685 14859 33751 14862
rect 36813 14859 36879 14862
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 14111 35248 14112
rect 25589 13970 25655 13973
rect 29729 13970 29795 13973
rect 25589 13968 29795 13970
rect 25589 13912 25594 13968
rect 25650 13912 29734 13968
rect 29790 13912 29795 13968
rect 25589 13910 29795 13912
rect 25589 13907 25655 13910
rect 29729 13907 29795 13910
rect 33869 13970 33935 13973
rect 39520 13970 40000 14000
rect 33869 13968 40000 13970
rect 33869 13912 33874 13968
rect 33930 13912 40000 13968
rect 33869 13910 40000 13912
rect 33869 13907 33935 13910
rect 39520 13880 40000 13910
rect 13997 13698 14063 13701
rect 14549 13698 14615 13701
rect 16665 13698 16731 13701
rect 13997 13696 16731 13698
rect 13997 13640 14002 13696
rect 14058 13640 14554 13696
rect 14610 13640 16670 13696
rect 16726 13640 16731 13696
rect 13997 13638 16731 13640
rect 13997 13635 14063 13638
rect 14549 13635 14615 13638
rect 16665 13635 16731 13638
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 26877 13562 26943 13565
rect 29453 13562 29519 13565
rect 26877 13560 29519 13562
rect 26877 13504 26882 13560
rect 26938 13504 29458 13560
rect 29514 13504 29519 13560
rect 26877 13502 29519 13504
rect 26877 13499 26943 13502
rect 29453 13499 29519 13502
rect 13261 13154 13327 13157
rect 16205 13154 16271 13157
rect 13261 13152 16271 13154
rect 13261 13096 13266 13152
rect 13322 13096 16210 13152
rect 16266 13096 16271 13152
rect 13261 13094 16271 13096
rect 13261 13091 13327 13094
rect 16205 13091 16271 13094
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 13023 35248 13024
rect 21909 13018 21975 13021
rect 25681 13018 25747 13021
rect 21909 13016 25747 13018
rect 21909 12960 21914 13016
rect 21970 12960 25686 13016
rect 25742 12960 25747 13016
rect 21909 12958 25747 12960
rect 21909 12955 21975 12958
rect 25681 12955 25747 12958
rect 27429 12882 27495 12885
rect 29821 12882 29887 12885
rect 27429 12880 29887 12882
rect 27429 12824 27434 12880
rect 27490 12824 29826 12880
rect 29882 12824 29887 12880
rect 27429 12822 29887 12824
rect 27429 12819 27495 12822
rect 29821 12819 29887 12822
rect 39520 12746 40000 12776
rect 37414 12686 40000 12746
rect 24393 12610 24459 12613
rect 36629 12610 36695 12613
rect 24393 12608 36695 12610
rect 24393 12552 24398 12608
rect 24454 12552 36634 12608
rect 36690 12552 36695 12608
rect 24393 12550 36695 12552
rect 24393 12547 24459 12550
rect 36629 12547 36695 12550
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 34237 12474 34303 12477
rect 34605 12474 34671 12477
rect 34237 12472 34671 12474
rect 34237 12416 34242 12472
rect 34298 12416 34610 12472
rect 34666 12416 34671 12472
rect 34237 12414 34671 12416
rect 34237 12411 34303 12414
rect 34605 12411 34671 12414
rect 35617 12474 35683 12477
rect 37414 12474 37474 12686
rect 39520 12656 40000 12686
rect 35617 12472 37474 12474
rect 35617 12416 35622 12472
rect 35678 12416 37474 12472
rect 35617 12414 37474 12416
rect 35617 12411 35683 12414
rect 21725 12338 21791 12341
rect 27705 12338 27771 12341
rect 21725 12336 27771 12338
rect 21725 12280 21730 12336
rect 21786 12280 27710 12336
rect 27766 12280 27771 12336
rect 21725 12278 27771 12280
rect 21725 12275 21791 12278
rect 27705 12275 27771 12278
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 11935 35248 11936
rect 19149 11794 19215 11797
rect 20621 11794 20687 11797
rect 19149 11792 20687 11794
rect 19149 11736 19154 11792
rect 19210 11736 20626 11792
rect 20682 11736 20687 11792
rect 19149 11734 20687 11736
rect 19149 11731 19215 11734
rect 20621 11731 20687 11734
rect 35433 11522 35499 11525
rect 39520 11522 40000 11552
rect 35433 11520 40000 11522
rect 35433 11464 35438 11520
rect 35494 11464 40000 11520
rect 35433 11462 40000 11464
rect 35433 11459 35499 11462
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 39520 11432 40000 11462
rect 19568 11391 19888 11392
rect 13169 11114 13235 11117
rect 13302 11114 13308 11116
rect 13169 11112 13308 11114
rect 13169 11056 13174 11112
rect 13230 11056 13308 11112
rect 13169 11054 13308 11056
rect 13169 11051 13235 11054
rect 13302 11052 13308 11054
rect 13372 11052 13378 11116
rect 17493 11114 17559 11117
rect 18689 11114 18755 11117
rect 20805 11114 20871 11117
rect 17493 11112 20871 11114
rect 17493 11056 17498 11112
rect 17554 11056 18694 11112
rect 18750 11056 20810 11112
rect 20866 11056 20871 11112
rect 17493 11054 20871 11056
rect 17493 11051 17559 11054
rect 18689 11051 18755 11054
rect 20805 11051 20871 11054
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 10847 35248 10848
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 35617 10298 35683 10301
rect 39520 10298 40000 10328
rect 35617 10296 40000 10298
rect 35617 10240 35622 10296
rect 35678 10240 40000 10296
rect 35617 10238 40000 10240
rect 35617 10235 35683 10238
rect 39520 10208 40000 10238
rect 34646 10100 34652 10164
rect 34716 10162 34722 10164
rect 34789 10162 34855 10165
rect 34716 10160 34855 10162
rect 34716 10104 34794 10160
rect 34850 10104 34855 10160
rect 34716 10102 34855 10104
rect 34716 10100 34722 10102
rect 34789 10099 34855 10102
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 13537 9754 13603 9757
rect 15561 9754 15627 9757
rect 13537 9752 15627 9754
rect 13537 9696 13542 9752
rect 13598 9696 15566 9752
rect 15622 9696 15627 9752
rect 13537 9694 15627 9696
rect 13537 9691 13603 9694
rect 15561 9691 15627 9694
rect 17033 9618 17099 9621
rect 20621 9618 20687 9621
rect 17033 9616 20687 9618
rect 17033 9560 17038 9616
rect 17094 9560 20626 9616
rect 20682 9560 20687 9616
rect 17033 9558 20687 9560
rect 17033 9555 17099 9558
rect 20621 9555 20687 9558
rect 21541 9618 21607 9621
rect 23657 9618 23723 9621
rect 21541 9616 23723 9618
rect 21541 9560 21546 9616
rect 21602 9560 23662 9616
rect 23718 9560 23723 9616
rect 21541 9558 23723 9560
rect 21541 9555 21607 9558
rect 23657 9555 23723 9558
rect 7833 9346 7899 9349
rect 9397 9346 9463 9349
rect 7833 9344 9463 9346
rect 7833 9288 7838 9344
rect 7894 9288 9402 9344
rect 9458 9288 9463 9344
rect 7833 9286 9463 9288
rect 7833 9283 7899 9286
rect 9397 9283 9463 9286
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 8937 9210 9003 9213
rect 10409 9210 10475 9213
rect 8937 9208 10475 9210
rect 8937 9152 8942 9208
rect 8998 9152 10414 9208
rect 10470 9152 10475 9208
rect 8937 9150 10475 9152
rect 8937 9147 9003 9150
rect 10409 9147 10475 9150
rect 34789 9074 34855 9077
rect 39520 9074 40000 9104
rect 34789 9072 40000 9074
rect 34789 9016 34794 9072
rect 34850 9016 40000 9072
rect 34789 9014 40000 9016
rect 34789 9011 34855 9014
rect 39520 8984 40000 9014
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 10869 8530 10935 8533
rect 13813 8530 13879 8533
rect 10869 8528 13879 8530
rect 10869 8472 10874 8528
rect 10930 8472 13818 8528
rect 13874 8472 13879 8528
rect 10869 8470 13879 8472
rect 10869 8467 10935 8470
rect 13813 8467 13879 8470
rect 21725 8394 21791 8397
rect 24025 8394 24091 8397
rect 21725 8392 24091 8394
rect 21725 8336 21730 8392
rect 21786 8336 24030 8392
rect 24086 8336 24091 8392
rect 21725 8334 24091 8336
rect 21725 8331 21791 8334
rect 24025 8331 24091 8334
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 35525 7850 35591 7853
rect 39520 7850 40000 7880
rect 35525 7848 40000 7850
rect 35525 7792 35530 7848
rect 35586 7792 40000 7848
rect 35525 7790 40000 7792
rect 35525 7787 35591 7790
rect 39520 7760 40000 7790
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 19149 7442 19215 7445
rect 21081 7442 21147 7445
rect 19149 7440 21147 7442
rect 19149 7384 19154 7440
rect 19210 7384 21086 7440
rect 21142 7384 21147 7440
rect 19149 7382 21147 7384
rect 19149 7379 19215 7382
rect 21081 7379 21147 7382
rect 17033 7306 17099 7309
rect 20069 7306 20135 7309
rect 17033 7304 20135 7306
rect 17033 7248 17038 7304
rect 17094 7248 20074 7304
rect 20130 7248 20135 7304
rect 17033 7246 20135 7248
rect 17033 7243 17099 7246
rect 20069 7243 20135 7246
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 5165 7034 5231 7037
rect 7741 7034 7807 7037
rect 5165 7032 7807 7034
rect 5165 6976 5170 7032
rect 5226 6976 7746 7032
rect 7802 6976 7807 7032
rect 5165 6974 7807 6976
rect 5165 6971 5231 6974
rect 7741 6971 7807 6974
rect 0 6762 480 6792
rect 4889 6762 4955 6765
rect 0 6760 4955 6762
rect 0 6704 4894 6760
rect 4950 6704 4955 6760
rect 0 6702 4955 6704
rect 0 6672 480 6702
rect 4889 6699 4955 6702
rect 35709 6626 35775 6629
rect 39520 6626 40000 6656
rect 35709 6624 40000 6626
rect 35709 6568 35714 6624
rect 35770 6568 40000 6624
rect 35709 6566 40000 6568
rect 35709 6563 35775 6566
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 39520 6536 40000 6566
rect 34928 6495 35248 6496
rect 17125 6490 17191 6493
rect 19425 6490 19491 6493
rect 17125 6488 19491 6490
rect 17125 6432 17130 6488
rect 17186 6432 19430 6488
rect 19486 6432 19491 6488
rect 17125 6430 19491 6432
rect 17125 6427 17191 6430
rect 19425 6427 19491 6430
rect 10501 6218 10567 6221
rect 12433 6218 12499 6221
rect 10501 6216 12499 6218
rect 10501 6160 10506 6216
rect 10562 6160 12438 6216
rect 12494 6160 12499 6216
rect 10501 6158 12499 6160
rect 10501 6155 10567 6158
rect 12433 6155 12499 6158
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 29729 5946 29795 5949
rect 31937 5946 32003 5949
rect 29729 5944 32003 5946
rect 29729 5888 29734 5944
rect 29790 5888 31942 5944
rect 31998 5888 32003 5944
rect 29729 5886 32003 5888
rect 29729 5883 29795 5886
rect 31937 5883 32003 5886
rect 7189 5674 7255 5677
rect 12157 5674 12223 5677
rect 7189 5672 12223 5674
rect 7189 5616 7194 5672
rect 7250 5616 12162 5672
rect 12218 5616 12223 5672
rect 7189 5614 12223 5616
rect 7189 5611 7255 5614
rect 12157 5611 12223 5614
rect 16941 5674 17007 5677
rect 19425 5674 19491 5677
rect 16941 5672 19491 5674
rect 16941 5616 16946 5672
rect 17002 5616 19430 5672
rect 19486 5616 19491 5672
rect 16941 5614 19491 5616
rect 16941 5611 17007 5614
rect 19425 5611 19491 5614
rect 20897 5674 20963 5677
rect 24025 5674 24091 5677
rect 20897 5672 24091 5674
rect 20897 5616 20902 5672
rect 20958 5616 24030 5672
rect 24086 5616 24091 5672
rect 20897 5614 24091 5616
rect 20897 5611 20963 5614
rect 24025 5611 24091 5614
rect 27245 5674 27311 5677
rect 33961 5674 34027 5677
rect 27245 5672 34027 5674
rect 27245 5616 27250 5672
rect 27306 5616 33966 5672
rect 34022 5616 34027 5672
rect 27245 5614 34027 5616
rect 27245 5611 27311 5614
rect 33961 5611 34027 5614
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 10593 5402 10659 5405
rect 16113 5402 16179 5405
rect 10593 5400 16179 5402
rect 10593 5344 10598 5400
rect 10654 5344 16118 5400
rect 16174 5344 16179 5400
rect 10593 5342 16179 5344
rect 10593 5339 10659 5342
rect 16113 5339 16179 5342
rect 17585 5402 17651 5405
rect 20621 5402 20687 5405
rect 21541 5402 21607 5405
rect 17585 5400 21607 5402
rect 17585 5344 17590 5400
rect 17646 5344 20626 5400
rect 20682 5344 21546 5400
rect 21602 5344 21607 5400
rect 17585 5342 21607 5344
rect 17585 5339 17651 5342
rect 20621 5339 20687 5342
rect 21541 5339 21607 5342
rect 35801 5402 35867 5405
rect 39520 5402 40000 5432
rect 35801 5400 40000 5402
rect 35801 5344 35806 5400
rect 35862 5344 40000 5400
rect 35801 5342 40000 5344
rect 35801 5339 35867 5342
rect 39520 5312 40000 5342
rect 9857 5266 9923 5269
rect 12617 5266 12683 5269
rect 9857 5264 12683 5266
rect 9857 5208 9862 5264
rect 9918 5208 12622 5264
rect 12678 5208 12683 5264
rect 9857 5206 12683 5208
rect 9857 5203 9923 5206
rect 12617 5203 12683 5206
rect 7465 5130 7531 5133
rect 34789 5130 34855 5133
rect 7465 5128 34855 5130
rect 7465 5072 7470 5128
rect 7526 5072 34794 5128
rect 34850 5072 34855 5128
rect 7465 5070 34855 5072
rect 7465 5067 7531 5070
rect 34789 5067 34855 5070
rect 10777 4994 10843 4997
rect 12525 4994 12591 4997
rect 10777 4992 12591 4994
rect 10777 4936 10782 4992
rect 10838 4936 12530 4992
rect 12586 4936 12591 4992
rect 10777 4934 12591 4936
rect 10777 4931 10843 4934
rect 12525 4931 12591 4934
rect 13077 4994 13143 4997
rect 14917 4994 14983 4997
rect 13077 4992 14983 4994
rect 13077 4936 13082 4992
rect 13138 4936 14922 4992
rect 14978 4936 14983 4992
rect 13077 4934 14983 4936
rect 13077 4931 13143 4934
rect 14917 4931 14983 4934
rect 23105 4994 23171 4997
rect 25037 4994 25103 4997
rect 23105 4992 25103 4994
rect 23105 4936 23110 4992
rect 23166 4936 25042 4992
rect 25098 4936 25103 4992
rect 23105 4934 25103 4936
rect 23105 4931 23171 4934
rect 25037 4931 25103 4934
rect 25313 4994 25379 4997
rect 30833 4994 30899 4997
rect 25313 4992 30899 4994
rect 25313 4936 25318 4992
rect 25374 4936 30838 4992
rect 30894 4936 30899 4992
rect 25313 4934 30899 4936
rect 25313 4931 25379 4934
rect 30833 4931 30899 4934
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 10501 4858 10567 4861
rect 16389 4858 16455 4861
rect 10501 4856 16455 4858
rect 10501 4800 10506 4856
rect 10562 4800 16394 4856
rect 16450 4800 16455 4856
rect 10501 4798 16455 4800
rect 10501 4795 10567 4798
rect 16389 4795 16455 4798
rect 16757 4858 16823 4861
rect 18229 4858 18295 4861
rect 19333 4858 19399 4861
rect 16757 4856 19399 4858
rect 16757 4800 16762 4856
rect 16818 4800 18234 4856
rect 18290 4800 19338 4856
rect 19394 4800 19399 4856
rect 16757 4798 19399 4800
rect 16757 4795 16823 4798
rect 18229 4795 18295 4798
rect 19333 4795 19399 4798
rect 22001 4858 22067 4861
rect 24301 4858 24367 4861
rect 22001 4856 24367 4858
rect 22001 4800 22006 4856
rect 22062 4800 24306 4856
rect 24362 4800 24367 4856
rect 22001 4798 24367 4800
rect 22001 4795 22067 4798
rect 24301 4795 24367 4798
rect 27705 4858 27771 4861
rect 30649 4858 30715 4861
rect 27705 4856 30715 4858
rect 27705 4800 27710 4856
rect 27766 4800 30654 4856
rect 30710 4800 30715 4856
rect 27705 4798 30715 4800
rect 27705 4795 27771 4798
rect 30649 4795 30715 4798
rect 10869 4722 10935 4725
rect 16573 4722 16639 4725
rect 10869 4720 16639 4722
rect 10869 4664 10874 4720
rect 10930 4664 16578 4720
rect 16634 4664 16639 4720
rect 10869 4662 16639 4664
rect 10869 4659 10935 4662
rect 16573 4659 16639 4662
rect 27981 4722 28047 4725
rect 31293 4722 31359 4725
rect 27981 4720 31359 4722
rect 27981 4664 27986 4720
rect 28042 4664 31298 4720
rect 31354 4664 31359 4720
rect 27981 4662 31359 4664
rect 27981 4659 28047 4662
rect 31293 4659 31359 4662
rect 12893 4586 12959 4589
rect 14457 4586 14523 4589
rect 15653 4586 15719 4589
rect 12893 4584 15719 4586
rect 12893 4528 12898 4584
rect 12954 4528 14462 4584
rect 14518 4528 15658 4584
rect 15714 4528 15719 4584
rect 12893 4526 15719 4528
rect 12893 4523 12959 4526
rect 14457 4523 14523 4526
rect 15653 4523 15719 4526
rect 16297 4586 16363 4589
rect 18689 4586 18755 4589
rect 16297 4584 18755 4586
rect 16297 4528 16302 4584
rect 16358 4528 18694 4584
rect 18750 4528 18755 4584
rect 16297 4526 18755 4528
rect 16297 4523 16363 4526
rect 18689 4523 18755 4526
rect 25865 4586 25931 4589
rect 27889 4586 27955 4589
rect 31201 4586 31267 4589
rect 37181 4586 37247 4589
rect 25865 4584 31267 4586
rect 25865 4528 25870 4584
rect 25926 4528 27894 4584
rect 27950 4528 31206 4584
rect 31262 4528 31267 4584
rect 25865 4526 31267 4528
rect 25865 4523 25931 4526
rect 27889 4523 27955 4526
rect 31201 4523 31267 4526
rect 33872 4584 37247 4586
rect 33872 4528 37186 4584
rect 37242 4528 37247 4584
rect 33872 4526 37247 4528
rect 15837 4450 15903 4453
rect 19701 4450 19767 4453
rect 15837 4448 19767 4450
rect 15837 4392 15842 4448
rect 15898 4392 19706 4448
rect 19762 4392 19767 4448
rect 15837 4390 19767 4392
rect 15837 4387 15903 4390
rect 19701 4387 19767 4390
rect 20345 4450 20411 4453
rect 22185 4450 22251 4453
rect 20345 4448 22251 4450
rect 20345 4392 20350 4448
rect 20406 4392 22190 4448
rect 22246 4392 22251 4448
rect 20345 4390 22251 4392
rect 20345 4387 20411 4390
rect 22185 4387 22251 4390
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 15745 4314 15811 4317
rect 17401 4314 17467 4317
rect 15745 4312 17467 4314
rect 15745 4256 15750 4312
rect 15806 4256 17406 4312
rect 17462 4256 17467 4312
rect 15745 4254 17467 4256
rect 15745 4251 15811 4254
rect 17401 4251 17467 4254
rect 22645 4314 22711 4317
rect 24669 4314 24735 4317
rect 22645 4312 24735 4314
rect 22645 4256 22650 4312
rect 22706 4256 24674 4312
rect 24730 4256 24735 4312
rect 22645 4254 24735 4256
rect 22645 4251 22711 4254
rect 24669 4251 24735 4254
rect 3049 4178 3115 4181
rect 6085 4178 6151 4181
rect 3049 4176 6151 4178
rect 3049 4120 3054 4176
rect 3110 4120 6090 4176
rect 6146 4120 6151 4176
rect 3049 4118 6151 4120
rect 3049 4115 3115 4118
rect 6085 4115 6151 4118
rect 7925 4178 7991 4181
rect 32673 4178 32739 4181
rect 33872 4178 33932 4526
rect 37181 4523 37247 4526
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 4319 35248 4320
rect 7925 4176 33932 4178
rect 7925 4120 7930 4176
rect 7986 4120 32678 4176
rect 32734 4120 33932 4176
rect 7925 4118 33932 4120
rect 35341 4178 35407 4181
rect 39520 4178 40000 4208
rect 35341 4176 40000 4178
rect 35341 4120 35346 4176
rect 35402 4120 40000 4176
rect 35341 4118 40000 4120
rect 7925 4115 7991 4118
rect 32673 4115 32739 4118
rect 35341 4115 35407 4118
rect 39520 4088 40000 4118
rect 3325 4042 3391 4045
rect 8477 4042 8543 4045
rect 3325 4040 8543 4042
rect 3325 3984 3330 4040
rect 3386 3984 8482 4040
rect 8538 3984 8543 4040
rect 3325 3982 8543 3984
rect 3325 3979 3391 3982
rect 8477 3979 8543 3982
rect 9949 4042 10015 4045
rect 16757 4042 16823 4045
rect 9949 4040 16823 4042
rect 9949 3984 9954 4040
rect 10010 3984 16762 4040
rect 16818 3984 16823 4040
rect 9949 3982 16823 3984
rect 9949 3979 10015 3982
rect 16757 3979 16823 3982
rect 36629 4042 36695 4045
rect 39389 4042 39455 4045
rect 36629 4040 39455 4042
rect 36629 3984 36634 4040
rect 36690 3984 39394 4040
rect 39450 3984 39455 4040
rect 36629 3982 39455 3984
rect 36629 3979 36695 3982
rect 39389 3979 39455 3982
rect 5257 3906 5323 3909
rect 7281 3906 7347 3909
rect 5257 3904 7347 3906
rect 5257 3848 5262 3904
rect 5318 3848 7286 3904
rect 7342 3848 7347 3904
rect 5257 3846 7347 3848
rect 5257 3843 5323 3846
rect 7281 3843 7347 3846
rect 10501 3906 10567 3909
rect 12893 3906 12959 3909
rect 10501 3904 12959 3906
rect 10501 3848 10506 3904
rect 10562 3848 12898 3904
rect 12954 3848 12959 3904
rect 10501 3846 12959 3848
rect 10501 3843 10567 3846
rect 12893 3843 12959 3846
rect 13445 3906 13511 3909
rect 15285 3906 15351 3909
rect 16849 3906 16915 3909
rect 13445 3904 16915 3906
rect 13445 3848 13450 3904
rect 13506 3848 15290 3904
rect 15346 3848 16854 3904
rect 16910 3848 16915 3904
rect 13445 3846 16915 3848
rect 13445 3843 13511 3846
rect 15285 3843 15351 3846
rect 16849 3843 16915 3846
rect 29177 3906 29243 3909
rect 32121 3906 32187 3909
rect 29177 3904 32187 3906
rect 29177 3848 29182 3904
rect 29238 3848 32126 3904
rect 32182 3848 32187 3904
rect 29177 3846 32187 3848
rect 29177 3843 29243 3846
rect 32121 3843 32187 3846
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 2037 3772 2103 3773
rect 2037 3770 2084 3772
rect 1992 3768 2084 3770
rect 1992 3712 2042 3768
rect 1992 3710 2084 3712
rect 2037 3708 2084 3710
rect 2148 3708 2154 3772
rect 3785 3770 3851 3773
rect 13353 3770 13419 3773
rect 3785 3768 13419 3770
rect 3785 3712 3790 3768
rect 3846 3712 13358 3768
rect 13414 3712 13419 3768
rect 3785 3710 13419 3712
rect 2037 3707 2103 3708
rect 3785 3707 3851 3710
rect 13353 3707 13419 3710
rect 23289 3770 23355 3773
rect 25313 3770 25379 3773
rect 23289 3768 25379 3770
rect 23289 3712 23294 3768
rect 23350 3712 25318 3768
rect 25374 3712 25379 3768
rect 23289 3710 25379 3712
rect 23289 3707 23355 3710
rect 25313 3707 25379 3710
rect 28942 3708 28948 3772
rect 29012 3770 29018 3772
rect 29453 3770 29519 3773
rect 29012 3768 29519 3770
rect 29012 3712 29458 3768
rect 29514 3712 29519 3768
rect 29012 3710 29519 3712
rect 29012 3708 29018 3710
rect 29453 3707 29519 3710
rect 31845 3770 31911 3773
rect 34605 3770 34671 3773
rect 31845 3768 34671 3770
rect 31845 3712 31850 3768
rect 31906 3712 34610 3768
rect 34666 3712 34671 3768
rect 31845 3710 34671 3712
rect 31845 3707 31911 3710
rect 34605 3707 34671 3710
rect 10961 3634 11027 3637
rect 16941 3634 17007 3637
rect 10961 3632 17007 3634
rect 10961 3576 10966 3632
rect 11022 3576 16946 3632
rect 17002 3576 17007 3632
rect 10961 3574 17007 3576
rect 10961 3571 11027 3574
rect 16941 3571 17007 3574
rect 32489 3634 32555 3637
rect 37365 3634 37431 3637
rect 32489 3632 37431 3634
rect 32489 3576 32494 3632
rect 32550 3576 37370 3632
rect 37426 3576 37431 3632
rect 32489 3574 37431 3576
rect 32489 3571 32555 3574
rect 37365 3571 37431 3574
rect 5809 3498 5875 3501
rect 8385 3498 8451 3501
rect 5809 3496 8451 3498
rect 5809 3440 5814 3496
rect 5870 3440 8390 3496
rect 8446 3440 8451 3496
rect 5809 3438 8451 3440
rect 5809 3435 5875 3438
rect 8385 3435 8451 3438
rect 9765 3498 9831 3501
rect 17217 3498 17283 3501
rect 32765 3498 32831 3501
rect 9765 3496 17283 3498
rect 9765 3440 9770 3496
rect 9826 3440 17222 3496
rect 17278 3440 17283 3496
rect 9765 3438 17283 3440
rect 9765 3435 9831 3438
rect 17217 3435 17283 3438
rect 27110 3496 32831 3498
rect 27110 3440 32770 3496
rect 32826 3440 32831 3496
rect 27110 3438 32831 3440
rect 12617 3362 12683 3365
rect 12750 3362 12756 3364
rect 12617 3360 12756 3362
rect 12617 3304 12622 3360
rect 12678 3304 12756 3360
rect 12617 3302 12756 3304
rect 12617 3299 12683 3302
rect 12750 3300 12756 3302
rect 12820 3300 12826 3364
rect 13353 3362 13419 3365
rect 27110 3362 27170 3438
rect 32765 3435 32831 3438
rect 13353 3360 27170 3362
rect 13353 3304 13358 3360
rect 13414 3304 27170 3360
rect 13353 3302 27170 3304
rect 27337 3362 27403 3365
rect 28349 3362 28415 3365
rect 27337 3360 28415 3362
rect 27337 3304 27342 3360
rect 27398 3304 28354 3360
rect 28410 3304 28415 3360
rect 27337 3302 28415 3304
rect 13353 3299 13419 3302
rect 27337 3299 27403 3302
rect 28349 3299 28415 3302
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 3231 35248 3232
rect 17493 3226 17559 3229
rect 20069 3226 20135 3229
rect 17493 3224 20135 3226
rect 17493 3168 17498 3224
rect 17554 3168 20074 3224
rect 20130 3168 20135 3224
rect 17493 3166 20135 3168
rect 17493 3163 17559 3166
rect 20069 3163 20135 3166
rect 24761 3226 24827 3229
rect 27153 3226 27219 3229
rect 24761 3224 27219 3226
rect 24761 3168 24766 3224
rect 24822 3168 27158 3224
rect 27214 3168 27219 3224
rect 24761 3166 27219 3168
rect 24761 3163 24827 3166
rect 27153 3163 27219 3166
rect 4153 3090 4219 3093
rect 4705 3090 4771 3093
rect 19241 3092 19307 3093
rect 4838 3090 4844 3092
rect 4153 3088 4844 3090
rect 4153 3032 4158 3088
rect 4214 3032 4710 3088
rect 4766 3032 4844 3088
rect 4153 3030 4844 3032
rect 4153 3027 4219 3030
rect 4705 3027 4771 3030
rect 4838 3028 4844 3030
rect 4908 3028 4914 3092
rect 19190 3028 19196 3092
rect 19260 3090 19307 3092
rect 34789 3090 34855 3093
rect 19260 3088 34855 3090
rect 19302 3032 34794 3088
rect 34850 3032 34855 3088
rect 19260 3030 34855 3032
rect 19260 3028 19307 3030
rect 19241 3027 19307 3028
rect 34789 3027 34855 3030
rect 12985 2954 13051 2957
rect 31661 2954 31727 2957
rect 12985 2952 31727 2954
rect 12985 2896 12990 2952
rect 13046 2896 31666 2952
rect 31722 2896 31727 2952
rect 12985 2894 31727 2896
rect 12985 2891 13051 2894
rect 31661 2891 31727 2894
rect 34697 2954 34763 2957
rect 39520 2954 40000 2984
rect 34697 2952 40000 2954
rect 34697 2896 34702 2952
rect 34758 2896 40000 2952
rect 34697 2894 40000 2896
rect 34697 2891 34763 2894
rect 39520 2864 40000 2894
rect 11697 2818 11763 2821
rect 13905 2818 13971 2821
rect 11697 2816 13971 2818
rect 11697 2760 11702 2816
rect 11758 2760 13910 2816
rect 13966 2760 13971 2816
rect 11697 2758 13971 2760
rect 11697 2755 11763 2758
rect 13905 2755 13971 2758
rect 22369 2818 22435 2821
rect 32305 2818 32371 2821
rect 22369 2816 32371 2818
rect 22369 2760 22374 2816
rect 22430 2760 32310 2816
rect 32366 2760 32371 2816
rect 22369 2758 32371 2760
rect 22369 2755 22435 2758
rect 32305 2755 32371 2758
rect 34421 2818 34487 2821
rect 38285 2818 38351 2821
rect 34421 2816 38351 2818
rect 34421 2760 34426 2816
rect 34482 2760 38290 2816
rect 38346 2760 38351 2816
rect 34421 2758 38351 2760
rect 34421 2755 34487 2758
rect 38285 2755 38351 2758
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 3141 2682 3207 2685
rect 12985 2682 13051 2685
rect 3141 2680 13051 2682
rect 3141 2624 3146 2680
rect 3202 2624 12990 2680
rect 13046 2624 13051 2680
rect 3141 2622 13051 2624
rect 3141 2619 3207 2622
rect 12985 2619 13051 2622
rect 21081 2682 21147 2685
rect 24485 2682 24551 2685
rect 21081 2680 24551 2682
rect 21081 2624 21086 2680
rect 21142 2624 24490 2680
rect 24546 2624 24551 2680
rect 21081 2622 24551 2624
rect 21081 2619 21147 2622
rect 24485 2619 24551 2622
rect 25957 2682 26023 2685
rect 28257 2682 28323 2685
rect 25957 2680 28323 2682
rect 25957 2624 25962 2680
rect 26018 2624 28262 2680
rect 28318 2624 28323 2680
rect 25957 2622 28323 2624
rect 25957 2619 26023 2622
rect 28257 2619 28323 2622
rect 2037 2546 2103 2549
rect 12617 2546 12683 2549
rect 2037 2544 12683 2546
rect 2037 2488 2042 2544
rect 2098 2488 12622 2544
rect 12678 2488 12683 2544
rect 2037 2486 12683 2488
rect 2037 2483 2103 2486
rect 12617 2483 12683 2486
rect 25773 2546 25839 2549
rect 28165 2546 28231 2549
rect 25773 2544 28231 2546
rect 25773 2488 25778 2544
rect 25834 2488 28170 2544
rect 28226 2488 28231 2544
rect 25773 2486 28231 2488
rect 25773 2483 25839 2486
rect 28165 2483 28231 2486
rect 24025 2410 24091 2413
rect 33869 2410 33935 2413
rect 24025 2408 33935 2410
rect 24025 2352 24030 2408
rect 24086 2352 33874 2408
rect 33930 2352 33935 2408
rect 24025 2350 33935 2352
rect 24025 2347 24091 2350
rect 33869 2347 33935 2350
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2143 35248 2144
rect 4797 2138 4863 2141
rect 24025 2138 24091 2141
rect 4797 2136 24091 2138
rect 4797 2080 4802 2136
rect 4858 2080 24030 2136
rect 24086 2080 24091 2136
rect 4797 2078 24091 2080
rect 4797 2075 4863 2078
rect 24025 2075 24091 2078
rect 12382 1940 12388 2004
rect 12452 2002 12458 2004
rect 13302 2002 13308 2004
rect 12452 1942 13308 2002
rect 12452 1940 12458 1942
rect 13302 1940 13308 1942
rect 13372 2002 13378 2004
rect 30557 2002 30623 2005
rect 13372 2000 30623 2002
rect 13372 1944 30562 2000
rect 30618 1944 30623 2000
rect 13372 1942 30623 1944
rect 13372 1940 13378 1942
rect 30557 1939 30623 1942
rect 35617 1730 35683 1733
rect 39520 1730 40000 1760
rect 35617 1728 40000 1730
rect 35617 1672 35622 1728
rect 35678 1672 40000 1728
rect 35617 1670 40000 1672
rect 35617 1667 35683 1670
rect 39520 1640 40000 1670
rect 35433 642 35499 645
rect 39520 642 40000 672
rect 35433 640 40000 642
rect 35433 584 35438 640
rect 35494 584 40000 640
rect 35433 582 40000 584
rect 35433 579 35499 582
rect 39520 552 40000 582
<< via3 >>
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 34652 19212 34716 19276
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 13308 11052 13372 11116
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 34652 10100 34716 10164
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 2084 3768 2148 3772
rect 2084 3712 2098 3768
rect 2098 3712 2148 3768
rect 2084 3708 2148 3712
rect 28948 3708 29012 3772
rect 12756 3300 12820 3364
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 4844 3028 4908 3092
rect 19196 3088 19260 3092
rect 19196 3032 19246 3088
rect 19246 3032 19260 3088
rect 19196 3028 19260 3032
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
rect 12388 1940 12452 2004
rect 13308 1940 13372 2004
<< metal4 >>
rect 4208 37024 4528 37584
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 19568 37568 19888 37584
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 34928 37024 35248 37584
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 22880 35248 23904
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34651 19276 34717 19277
rect 34651 19212 34652 19276
rect 34716 19212 34717 19276
rect 34651 19211 34717 19212
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 13307 11116 13373 11117
rect 13307 11052 13308 11116
rect 13372 11052 13373 11116
rect 13307 11051 13373 11052
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 12170 3710 12450 3770
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 12390 2005 12450 3710
rect 12758 3365 12818 3622
rect 12755 3364 12821 3365
rect 12755 3300 12756 3364
rect 12820 3300 12821 3364
rect 12755 3299 12821 3300
rect 13310 2005 13370 11051
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 34654 10165 34714 19211
rect 34928 18528 35248 19552
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34651 10164 34717 10165
rect 34651 10100 34652 10164
rect 34716 10100 34717 10164
rect 34651 10099 34717 10100
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5472 35248 6496
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 4384 35248 5408
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2128 19888 2688
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2128 35248 2144
rect 12387 2004 12453 2005
rect 12387 1940 12388 2004
rect 12452 1940 12453 2004
rect 12387 1939 12453 1940
rect 13307 2004 13373 2005
rect 13307 1940 13308 2004
rect 13372 1940 13373 2004
rect 13307 1939 13373 1940
<< via4 >>
rect 1998 3772 2234 3858
rect 1998 3708 2084 3772
rect 2084 3708 2148 3772
rect 2148 3708 2234 3772
rect 1998 3622 2234 3708
rect 11934 3622 12170 3858
rect 4758 3092 4994 3178
rect 4758 3028 4844 3092
rect 4844 3028 4908 3092
rect 4908 3028 4994 3092
rect 4758 2942 4994 3028
rect 12670 3622 12906 3858
rect 19110 3092 19346 3178
rect 19110 3028 19196 3092
rect 19196 3028 19260 3092
rect 19260 3028 19346 3092
rect 19110 2942 19346 3028
rect 28862 3772 29098 3858
rect 28862 3708 28948 3772
rect 28948 3708 29012 3772
rect 29012 3708 29098 3772
rect 28862 3622 29098 3708
<< metal5 >>
rect 1956 3858 12212 3900
rect 1956 3622 1998 3858
rect 2234 3622 11934 3858
rect 12170 3622 12212 3858
rect 1956 3580 12212 3622
rect 12628 3858 29140 3900
rect 12628 3622 12670 3858
rect 12906 3622 28862 3858
rect 29098 3622 29140 3858
rect 12628 3580 29140 3622
rect 4716 3178 19388 3220
rect 4716 2942 4758 3178
rect 4994 2942 19110 3178
rect 19346 2942 19388 3178
rect 4716 2900 19388 2942
use sky130_fd_sc_hd__fill_2  FILLER_1_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7
timestamp 1604666999
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604666999
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _65_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604666999
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_11 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 2116 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11
timestamp 1604666999
transform 1 0 2116 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 2300 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604666999
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604666999
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604666999
transform 1 0 2484 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_19
timestamp 1604666999
transform 1 0 2852 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1604666999
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19
timestamp 1604666999
transform 1 0 2852 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604666999
transform 1 0 3036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604666999
transform 1 0 3128 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604666999
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604666999
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604666999
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1604666999
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_26
timestamp 1604666999
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604666999
transform 1 0 4140 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604666999
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 4048 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_30
timestamp 1604666999
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37
timestamp 1604666999
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41
timestamp 1604666999
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
timestamp 1604666999
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604666999
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 4232 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
timestamp 1604666999
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1604666999
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1604666999
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
timestamp 1604666999
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 1604666999
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1604666999
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604666999
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
timestamp 1604666999
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
timestamp 1604666999
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604666999
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63
timestamp 1604666999
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
timestamp 1604666999
transform 1 0 7176 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
timestamp 1604666999
transform 1 0 6808 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_85 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 8924 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_81
timestamp 1604666999
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604666999
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604666999
transform 1 0 8740 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_91
timestamp 1604666999
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1604666999
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
timestamp 1604666999
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 9292 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
timestamp 1604666999
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604666999
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 9844 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
timestamp 1604666999
transform 1 0 9752 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1604666999
transform 1 0 11500 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604666999
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604666999
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1604666999
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
timestamp 1604666999
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_123
timestamp 1604666999
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121
timestamp 1604666999
transform 1 0 12236 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604666999
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604666999
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_127
timestamp 1604666999
transform 1 0 12788 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_125
timestamp 1604666999
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 12604 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604666999
transform 1 0 12972 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_142
timestamp 1604666999
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_138
timestamp 1604666999
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1604666999
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCD
timestamp 1604666999
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCE
timestamp 1604666999
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 12880 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 14536 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 15456 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604666999
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCD
timestamp 1604666999
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1604666999
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_170
timestamp 1604666999
transform 1 0 16744 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCE
timestamp 1604666999
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_175
timestamp 1604666999
transform 1 0 17204 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_175
timestamp 1604666999
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604666999
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_179
timestamp 1604666999
transform 1 0 17572 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_183
timestamp 1604666999
transform 1 0 17940 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_179
timestamp 1604666999
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604666999
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp 1604666999
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 18584 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 18032 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_207
timestamp 1604666999
transform 1 0 20148 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_203
timestamp 1604666999
transform 1 0 19780 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1604666999
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCD
timestamp 1604666999
transform 1 0 19964 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__D
timestamp 1604666999
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCE
timestamp 1604666999
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_218
timestamp 1604666999
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_213
timestamp 1604666999
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604666999
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 21252 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_
timestamp 1604666999
transform 1 0 20516 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_2  FILLER_1_235
timestamp 1604666999
transform 1 0 22724 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_238
timestamp 1604666999
transform 1 0 23000 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 22908 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_239
timestamp 1604666999
transform 1 0 23092 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 23276 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_245
timestamp 1604666999
transform 1 0 23644 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_243
timestamp 1604666999
transform 1 0 23460 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_244
timestamp 1604666999
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604666999
transform 1 0 23828 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604666999
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604666999
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_260
timestamp 1604666999
transform 1 0 25024 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_249
timestamp 1604666999
transform 1 0 24012 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_258
timestamp 1604666999
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604666999
transform 1 0 24196 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604666999
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_264
timestamp 1604666999
transform 1 0 25392 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_271
timestamp 1604666999
transform 1 0 26036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_262
timestamp 1604666999
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
timestamp 1604666999
transform 1 0 25208 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604666999
transform 1 0 25392 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
timestamp 1604666999
transform 1 0 25576 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604666999
transform 1 0 26220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 25576 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
timestamp 1604666999
transform 1 0 25760 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_0_275
timestamp 1604666999
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
timestamp 1604666999
transform 1 0 26588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604666999
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_295
timestamp 1604666999
transform 1 0 28244 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_291
timestamp 1604666999
transform 1 0 27876 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_287
timestamp 1604666999
transform 1 0 27508 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
timestamp 1604666999
transform 1 0 27692 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 28060 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 28428 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
timestamp 1604666999
transform 1 0 26864 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_0_299
timestamp 1604666999
transform 1 0 28612 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_299
timestamp 1604666999
transform 1 0 28612 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604666999
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 28980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 29072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_303
timestamp 1604666999
transform 1 0 28980 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1604666999
transform 1 0 29256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_306
timestamp 1604666999
transform 1 0 29256 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604666999
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 29440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_311
timestamp 1604666999
transform 1 0 29716 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 29348 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 29808 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_330
timestamp 1604666999
transform 1 0 31464 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_326
timestamp 1604666999
transform 1 0 31096 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_331
timestamp 1604666999
transform 1 0 31556 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604666999
transform 1 0 31280 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__D
timestamp 1604666999
transform 1 0 31832 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCE
timestamp 1604666999
transform 1 0 31648 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_342
timestamp 1604666999
transform 1 0 32568 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_336
timestamp 1604666999
transform 1 0 32016 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 32292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604666999
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 32844 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_
timestamp 1604666999
transform 1 0 31832 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_2  FILLER_1_362
timestamp 1604666999
transform 1 0 34408 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_358
timestamp 1604666999
transform 1 0 34040 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCE
timestamp 1604666999
transform 1 0 34224 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_367
timestamp 1604666999
transform 1 0 34868 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_364
timestamp 1604666999
transform 1 0 34592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 34776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 34592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604666999
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_368
timestamp 1604666999
transform 1 0 34960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 35144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 35236 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604666999
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 35420 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 35420 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 37352 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 37352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_392
timestamp 1604666999
transform 1 0 37168 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_396 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 37536 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_392
timestamp 1604666999
transform 1 0 37168 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_396
timestamp 1604666999
transform 1 0 37536 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604666999
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604666999
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604666999
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_402
timestamp 1604666999
transform 1 0 38088 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_404
timestamp 1604666999
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_404
timestamp 1604666999
transform 1 0 38272 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604666999
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604666999
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_32
timestamp 1604666999
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1604666999
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604666999
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604666999
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604666999
transform 1 0 4232 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_42
timestamp 1604666999
transform 1 0 4968 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_38
timestamp 1604666999
transform 1 0 4600 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604666999
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
timestamp 1604666999
transform 1 0 4784 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
timestamp 1604666999
transform 1 0 5336 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604666999
transform 1 0 7820 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
timestamp 1604666999
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604666999
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_65
timestamp 1604666999
transform 1 0 7084 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_69
timestamp 1604666999
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604666999
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 9844 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604666999
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1604666999
transform 1 0 8648 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_86
timestamp 1604666999
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1604666999
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1604666999
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_97
timestamp 1604666999
transform 1 0 10028 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10488 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 12328 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 10304 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 11500 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 11868 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_111
timestamp 1604666999
transform 1 0 11316 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_115
timestamp 1604666999
transform 1 0 11684 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_119
timestamp 1604666999
transform 1 0 12052 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__D
timestamp 1604666999
transform 1 0 14536 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1604666999
transform 1 0 14076 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_145
timestamp 1604666999
transform 1 0 14444 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_148
timestamp 1604666999
transform 1 0 14720 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_158
timestamp 1604666999
transform 1 0 15640 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_154
timestamp 1604666999
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1604666999
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 14904 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 15456 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604666999
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 15824 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_173
timestamp 1604666999
transform 1 0 17020 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_169
timestamp 1604666999
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 16836 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_
timestamp 1604666999
transform 1 0 17388 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 17204 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 20976 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604666999
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 20148 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_201
timestamp 1604666999
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_205
timestamp 1604666999
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_209
timestamp 1604666999
transform 1 0 20332 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_215
timestamp 1604666999
transform 1 0 20884 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604666999
transform 1 0 23736 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 23552 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 23184 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_235
timestamp 1604666999
transform 1 0 22724 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_239
timestamp 1604666999
transform 1 0 23092 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_242
timestamp 1604666999
transform 1 0 23368 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604666999
transform 1 0 24840 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604666999
transform 1 0 24288 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604666999
transform 1 0 24656 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 26220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 25852 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1604666999
transform 1 0 24104 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_254
timestamp 1604666999
transform 1 0 24472 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_267
timestamp 1604666999
transform 1 0 25668 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_271
timestamp 1604666999
transform 1 0 26036 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604666999
transform 1 0 26496 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 28428 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604666999
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 27508 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 27876 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604666999
transform 1 0 28244 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_285
timestamp 1604666999
transform 1 0 27324 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_289
timestamp 1604666999
transform 1 0 27692 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_293
timestamp 1604666999
transform 1 0 28060 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 30728 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 30360 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_316
timestamp 1604666999
transform 1 0 30176 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_320
timestamp 1604666999
transform 1 0 30544 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604666999
transform 1 0 30912 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_
timestamp 1604666999
transform 1 0 32476 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604666999
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCD
timestamp 1604666999
transform 1 0 32292 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCD
timestamp 1604666999
transform 1 0 31832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 31464 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_328
timestamp 1604666999
transform 1 0 31280 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_332
timestamp 1604666999
transform 1 0 31648 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_337
timestamp 1604666999
transform 1 0 32108 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 35236 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 34868 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1604666999
transform 1 0 34684 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_369
timestamp 1604666999
transform 1 0 35052 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 35420 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604666999
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 36432 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 36800 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_382
timestamp 1604666999
transform 1 0 36248 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_386
timestamp 1604666999
transform 1 0 36616 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_390
timestamp 1604666999
transform 1 0 36984 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_396
timestamp 1604666999
transform 1 0 37536 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604666999
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_398
timestamp 1604666999
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_406
timestamp 1604666999
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604666999
transform 1 0 3128 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604666999
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604666999
transform 1 0 2944 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604666999
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1604666999
transform 1 0 2484 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_19
timestamp 1604666999
transform 1 0 2852 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
timestamp 1604666999
transform 1 0 4232 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
timestamp 1604666999
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604666999
transform 1 0 3680 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_26
timestamp 1604666999
transform 1 0 3496 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_30
timestamp 1604666999
transform 1 0 3864 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604666999
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604666999
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604666999
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_53
timestamp 1604666999
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1604666999
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_71
timestamp 1604666999
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604666999
transform 1 0 8372 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604666999
transform 1 0 9936 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604666999
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604666999
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_75
timestamp 1604666999
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_88
timestamp 1604666999
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_92
timestamp 1604666999
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_109
timestamp 1604666999
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_105
timestamp 1604666999
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604666999
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_113
timestamp 1604666999
transform 1 0 11500 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 11316 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604666999
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 14260 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 14076 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_132
timestamp 1604666999
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_136
timestamp 1604666999
transform 1 0 13616 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_140
timestamp 1604666999
transform 1 0 13984 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604666999
transform 1 0 16744 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 16560 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_162
timestamp 1604666999
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1604666999
transform 1 0 16376 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 18584 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604666999
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 17664 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604666999
transform 1 0 17296 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_174
timestamp 1604666999
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_178
timestamp 1604666999
transform 1 0 17480 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_182
timestamp 1604666999
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_184
timestamp 1604666999
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604666999
transform 1 0 21068 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_209
timestamp 1604666999
transform 1 0 20332 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_213
timestamp 1604666999
transform 1 0 20700 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_230
timestamp 1604666999
transform 1 0 22264 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_226
timestamp 1604666999
transform 1 0 21896 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 22448 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 22080 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_238
timestamp 1604666999
transform 1 0 23000 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_234
timestamp 1604666999
transform 1 0 22632 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604666999
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604666999
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604666999
transform 1 0 23644 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
timestamp 1604666999
transform 1 0 25576 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
timestamp 1604666999
transform 1 0 25392 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
timestamp 1604666999
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_254
timestamp 1604666999
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_258
timestamp 1604666999
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_262
timestamp 1604666999
transform 1 0 25208 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604666999
transform 1 0 28060 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
timestamp 1604666999
transform 1 0 27508 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
timestamp 1604666999
transform 1 0 27876 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_285
timestamp 1604666999
transform 1 0 27324 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_289
timestamp 1604666999
transform 1 0 27692 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_297
timestamp 1604666999
transform 1 0 28428 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_301
timestamp 1604666999
transform 1 0 28796 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604666999
transform 1 0 28612 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604666999
transform 1 0 28980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604666999
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604666999
transform 1 0 29256 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_315
timestamp 1604666999
transform 1 0 30084 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_310
timestamp 1604666999
transform 1 0 29624 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 29900 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 30268 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_319
timestamp 1604666999
transform 1 0 30452 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 30728 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 32292 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 32108 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 31740 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_331
timestamp 1604666999
transform 1 0 31556 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_335
timestamp 1604666999
transform 1 0 31924 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604666999
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 34224 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 35236 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 34592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_358
timestamp 1604666999
transform 1 0 34040 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_362
timestamp 1604666999
transform 1 0 34408 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_367
timestamp 1604666999
transform 1 0 34868 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 35420 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_3_392
timestamp 1604666999
transform 1 0 37168 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604666999
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_404
timestamp 1604666999
transform 1 0 38272 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604666999
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604666999
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604666999
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604666999
transform 1 0 4508 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604666999
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
timestamp 1604666999
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604666999
transform 1 0 5612 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604666999
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_32
timestamp 1604666999
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_36
timestamp 1604666999
transform 1 0 4416 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_46
timestamp 1604666999
transform 1 0 5336 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604666999
transform 1 0 7728 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604666999
transform 1 0 6072 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_51
timestamp 1604666999
transform 1 0 5796 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_63
timestamp 1604666999
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_67
timestamp 1604666999
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_71
timestamp 1604666999
transform 1 0 7636 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_76
timestamp 1604666999
transform 1 0 8096 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp 1604666999
transform 1 0 8924 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_81
timestamp 1604666999
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_89
timestamp 1604666999
transform 1 0 9292 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604666999
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_93
timestamp 1604666999
transform 1 0 9660 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604666999
transform 1 0 9752 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_4_99
timestamp 1604666999
transform 1 0 10212 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 10948 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 10396 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_103
timestamp 1604666999
transform 1 0 10580 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 13432 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_126
timestamp 1604666999
transform 1 0 12696 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_130
timestamp 1604666999
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_143
timestamp 1604666999
transform 1 0 14260 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_147
timestamp 1604666999
transform 1 0 14628 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604666999
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604666999
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 16652 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_163
timestamp 1604666999
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_167
timestamp 1604666999
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_171
timestamp 1604666999
transform 1 0 16836 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 19228 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 17664 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 17480 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 18676 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__D
timestamp 1604666999
transform 1 0 17112 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 19044 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_176
timestamp 1604666999
transform 1 0 17296 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_189
timestamp 1604666999
transform 1 0 18492 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_193
timestamp 1604666999
transform 1 0 18860 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 20884 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604666999
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_206
timestamp 1604666999
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_210
timestamp 1604666999
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604666999
transform 1 0 23368 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 23920 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 23000 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_234
timestamp 1604666999
transform 1 0 22632 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_240
timestamp 1604666999
transform 1 0 23184 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_246
timestamp 1604666999
transform 1 0 23736 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604666999
transform 1 0 24840 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 24656 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 24288 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604666999
transform 1 0 25852 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 26220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1604666999
transform 1 0 24104 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_254
timestamp 1604666999
transform 1 0 24472 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_267
timestamp 1604666999
transform 1 0 25668 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_271
timestamp 1604666999
transform 1 0 26036 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
timestamp 1604666999
transform 1 0 26496 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604666999
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 28428 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_295
timestamp 1604666999
transform 1 0 28244 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604666999
transform 1 0 28980 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 30268 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 29532 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 29900 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_299
timestamp 1604666999
transform 1 0 28612 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_307
timestamp 1604666999
transform 1 0 29348 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_311
timestamp 1604666999
transform 1 0 29716 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_315
timestamp 1604666999
transform 1 0 30084 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_326
timestamp 1604666999
transform 1 0 31096 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_330
timestamp 1604666999
transform 1 0 31464 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604666999
transform 1 0 31280 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_334
timestamp 1604666999
transform 1 0 31832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 31648 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604666999
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _47_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 32108 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_340
timestamp 1604666999
transform 1 0 32384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__D
timestamp 1604666999
transform 1 0 32568 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_344
timestamp 1604666999
transform 1 0 32752 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 32936 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604666999
transform 1 0 34684 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 33120 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 34500 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 34132 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_357
timestamp 1604666999
transform 1 0 33948 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_361
timestamp 1604666999
transform 1 0 34316 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604666999
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 35696 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_374
timestamp 1604666999
transform 1 0 35512 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_378
timestamp 1604666999
transform 1 0 35880 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_390
timestamp 1604666999
transform 1 0 36984 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_396
timestamp 1604666999
transform 1 0 37536 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604666999
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_398
timestamp 1604666999
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_406
timestamp 1604666999
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604666999
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604666999
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604666999
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
timestamp 1604666999
transform 1 0 4232 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
timestamp 1604666999
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1604666999
transform 1 0 3588 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_31
timestamp 1604666999
transform 1 0 3956 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_53
timestamp 1604666999
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1604666999
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604666999
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604666999
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604666999
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604666999
transform 1 0 6808 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_66
timestamp 1604666999
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604666999
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_70
timestamp 1604666999
transform 1 0 7544 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 7728 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604666999
transform 1 0 7912 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604666999
transform 1 0 9384 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604666999
transform 1 0 8464 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604666999
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_78
timestamp 1604666999
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_82
timestamp 1604666999
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_86
timestamp 1604666999
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_99
timestamp 1604666999
transform 1 0 10212 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604666999
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604666999
transform 1 0 10948 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604666999
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604666999
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604666999
transform 1 0 10488 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_104
timestamp 1604666999
transform 1 0 10672 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_111
timestamp 1604666999
transform 1 0 11316 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_116
timestamp 1604666999
transform 1 0 11776 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 13892 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604666999
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_127
timestamp 1604666999
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_131
timestamp 1604666999
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_135
timestamp 1604666999
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604666999
transform 1 0 16376 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604666999
transform 1 0 16928 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_158
timestamp 1604666999
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_162
timestamp 1604666999
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_170
timestamp 1604666999
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604666999
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_174
timestamp 1604666999
transform 1 0 17112 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_179
timestamp 1604666999
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_193
timestamp 1604666999
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_197
timestamp 1604666999
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604666999
transform 1 0 19596 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_205
timestamp 1604666999
transform 1 0 19964 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604666999
transform 1 0 20148 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_209
timestamp 1604666999
transform 1 0 20332 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 20516 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604666999
transform 1 0 20700 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_217
timestamp 1604666999
transform 1 0 21068 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_221
timestamp 1604666999
transform 1 0 21436 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604666999
transform 1 0 21252 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604666999
transform 1 0 21988 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 23644 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604666999
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604666999
transform 1 0 21804 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_236
timestamp 1604666999
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_240
timestamp 1604666999
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604666999
transform 1 0 26128 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 25576 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 25944 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_264
timestamp 1604666999
transform 1 0 25392 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_268
timestamp 1604666999
transform 1 0 25760 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604666999
transform 1 0 27600 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604666999
transform 1 0 26680 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 27416 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 27048 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_276
timestamp 1604666999
transform 1 0 26496 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_280
timestamp 1604666999
transform 1 0 26864 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_284
timestamp 1604666999
transform 1 0 27232 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_297
timestamp 1604666999
transform 1 0 28428 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 29256 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604666999
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
timestamp 1604666999
transform 1 0 28980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 28612 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
timestamp 1604666999
transform 1 0 30268 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604666999
transform 1 0 30636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_301
timestamp 1604666999
transform 1 0 28796 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_315
timestamp 1604666999
transform 1 0 30084 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_319
timestamp 1604666999
transform 1 0 30452 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604666999
transform 1 0 30820 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 32568 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 32384 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 32016 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_332
timestamp 1604666999
transform 1 0 31648 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_338
timestamp 1604666999
transform 1 0 32200 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_359
timestamp 1604666999
transform 1 0 34132 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_355
timestamp 1604666999
transform 1 0 33764 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_351
timestamp 1604666999
transform 1 0 33396 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 33580 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 33948 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_363
timestamp 1604666999
transform 1 0 34500 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 34316 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604666999
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _49_
timestamp 1604666999
transform 1 0 34868 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_370
timestamp 1604666999
transform 1 0 35144 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_382
timestamp 1604666999
transform 1 0 36248 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_394
timestamp 1604666999
transform 1 0 37352 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604666999
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_406
timestamp 1604666999
transform 1 0 38456 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604666999
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604666999
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604666999
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604666999
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604666999
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604666999
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1604666999
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604666999
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
timestamp 1604666999
transform 1 0 4232 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604666999
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_43
timestamp 1604666999
transform 1 0 5060 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_39
timestamp 1604666999
transform 1 0 4692 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_48
timestamp 1604666999
transform 1 0 5520 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
timestamp 1604666999
transform 1 0 5244 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
timestamp 1604666999
transform 1 0 4876 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604666999
transform 1 0 5612 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_7_47
timestamp 1604666999
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604666999
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_36
timestamp 1604666999
transform 1 0 4416 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_58
timestamp 1604666999
transform 1 0 6440 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
timestamp 1604666999
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
timestamp 1604666999
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604666999
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_73
timestamp 1604666999
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_69
timestamp 1604666999
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_64
timestamp 1604666999
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 7636 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1604666999
transform 1 0 7176 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
timestamp 1604666999
transform 1 0 6808 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_81
timestamp 1604666999
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_81
timestamp 1604666999
transform 1 0 8556 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 8740 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 8004 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604666999
transform 1 0 8188 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_91
timestamp 1604666999
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_85
timestamp 1604666999
transform 1 0 8924 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1604666999
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_89
timestamp 1604666999
transform 1 0 9292 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604666999
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_97
timestamp 1604666999
transform 1 0 10028 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604666999
transform 1 0 9844 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_104
timestamp 1604666999
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_110
timestamp 1604666999
transform 1 0 11224 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_106
timestamp 1604666999
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604666999
transform 1 0 11040 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 10304 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604666999
transform 1 0 10488 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_118
timestamp 1604666999
transform 1 0 11960 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604666999
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604666999
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604666999
transform 1 0 11592 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604666999
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_108
timestamp 1604666999
transform 1 0 11040 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCD
timestamp 1604666999
transform 1 0 12972 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 13064 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 12696 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_128
timestamp 1604666999
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_127
timestamp 1604666999
transform 1 0 12788 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 13340 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_132
timestamp 1604666999
transform 1 0 13248 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_131
timestamp 1604666999
transform 1 0 13156 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_135
timestamp 1604666999
transform 1 0 13524 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_149
timestamp 1604666999
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_145
timestamp 1604666999
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__D
timestamp 1604666999
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCE
timestamp 1604666999
transform 1 0 13708 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_
timestamp 1604666999
transform 1 0 13892 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604666999
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_7_163
timestamp 1604666999
transform 1 0 16100 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_6_167
timestamp 1604666999
transform 1 0 16468 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_163
timestamp 1604666999
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_169
timestamp 1604666999
transform 1 0 16652 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 16744 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604666999
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1604666999
transform 1 0 16928 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1604666999
transform 1 0 16928 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 17388 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_175
timestamp 1604666999
transform 1 0 17204 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_179
timestamp 1604666999
transform 1 0 17572 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_175
timestamp 1604666999
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_179
timestamp 1604666999
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604666999
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 17756 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_197
timestamp 1604666999
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1604666999
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 17940 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_6_206
timestamp 1604666999
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_202
timestamp 1604666999
transform 1 0 19688 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 19872 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 19596 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_217
timestamp 1604666999
transform 1 0 21068 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_214
timestamp 1604666999
transform 1 0 20792 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_210
timestamp 1604666999
transform 1 0 20424 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_218
timestamp 1604666999
transform 1 0 21160 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_210
timestamp 1604666999
transform 1 0 20424 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604666999
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604666999
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604666999
transform 1 0 21160 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1604666999
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1604666999
transform 1 0 21528 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_222
timestamp 1604666999
transform 1 0 21528 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604666999
transform 1 0 21344 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_226
timestamp 1604666999
transform 1 0 21896 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_234
timestamp 1604666999
transform 1 0 22632 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_230
timestamp 1604666999
transform 1 0 22264 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 21712 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604666999
transform 1 0 22264 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 22448 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604666999
transform 1 0 21712 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604666999
transform 1 0 21896 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604666999
transform 1 0 22448 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_240
timestamp 1604666999
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_236
timestamp 1604666999
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 22816 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604666999
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 23644 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 23000 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_6_257
timestamp 1604666999
transform 1 0 24748 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_268
timestamp 1604666999
transform 1 0 25760 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1604666999
transform 1 0 25392 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_261
timestamp 1604666999
transform 1 0 25116 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 24932 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604666999
transform 1 0 25576 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_269
timestamp 1604666999
transform 1 0 25852 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 26128 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 25944 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604666999
transform 1 0 26128 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1604666999
transform 1 0 26956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_281
timestamp 1604666999
transform 1 0 26956 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_276
timestamp 1604666999
transform 1 0 26496 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_274
timestamp 1604666999
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 26772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 27140 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604666999
transform 1 0 27140 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604666999
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_285
timestamp 1604666999
transform 1 0 27324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604666999
transform 1 0 27508 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604666999
transform 1 0 27692 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604666999
transform 1 0 27324 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_297
timestamp 1604666999
transform 1 0 28428 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_293
timestamp 1604666999
transform 1 0 28060 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_298
timestamp 1604666999
transform 1 0 28520 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_294
timestamp 1604666999
transform 1 0 28152 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604666999
transform 1 0 28336 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604666999
transform 1 0 28244 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_301
timestamp 1604666999
transform 1 0 28796 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_302
timestamp 1604666999
transform 1 0 28888 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604666999
transform 1 0 28704 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
timestamp 1604666999
transform 1 0 28612 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
timestamp 1604666999
transform 1 0 28980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604666999
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604666999
transform 1 0 29256 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_319
timestamp 1604666999
transform 1 0 30452 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_315
timestamp 1604666999
transform 1 0 30084 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604666999
transform 1 0 30636 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604666999
transform 1 0 30268 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
timestamp 1604666999
transform 1 0 29164 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_323
timestamp 1604666999
transform 1 0 30820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_328
timestamp 1604666999
transform 1 0 31280 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_324
timestamp 1604666999
transform 1 0 30912 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 31832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604666999
transform 1 0 31004 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604666999
transform 1 0 31096 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_347
timestamp 1604666999
transform 1 0 33028 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_339
timestamp 1604666999
transform 1 0 32292 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_346
timestamp 1604666999
transform 1 0 32936 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_341
timestamp 1604666999
transform 1 0 32476 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_337
timestamp 1604666999
transform 1 0 32108 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 32292 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604666999
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _48_
timestamp 1604666999
transform 1 0 32660 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_327
timestamp 1604666999
transform 1 0 31188 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_356
timestamp 1604666999
transform 1 0 33856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_350
timestamp 1604666999
transform 1 0 33304 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 33120 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604666999
transform 1 0 33948 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _50_
timestamp 1604666999
transform 1 0 33304 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_365
timestamp 1604666999
transform 1 0 34684 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604666999
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_367
timestamp 1604666999
transform 1 0 34868 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_353
timestamp 1604666999
transform 1 0 33580 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_366
timestamp 1604666999
transform 1 0 34776 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604666999
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_378
timestamp 1604666999
transform 1 0 35880 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_390
timestamp 1604666999
transform 1 0 36984 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_396
timestamp 1604666999
transform 1 0 37536 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_379
timestamp 1604666999
transform 1 0 35972 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_391
timestamp 1604666999
transform 1 0 37076 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604666999
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604666999
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_398
timestamp 1604666999
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_406
timestamp 1604666999
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_403
timestamp 1604666999
transform 1 0 38180 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604666999
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604666999
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604666999
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
timestamp 1604666999
transform 1 0 4876 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604666999
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604666999
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_32
timestamp 1604666999
transform 1 0 4048 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_40
timestamp 1604666999
transform 1 0 4784 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604666999
transform 1 0 7360 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_60
timestamp 1604666999
transform 1 0 6624 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_81
timestamp 1604666999
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_77
timestamp 1604666999
transform 1 0 8188 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_85
timestamp 1604666999
transform 1 0 8924 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_93
timestamp 1604666999
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1604666999
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604666999
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_97
timestamp 1604666999
transform 1 0 10028 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 10120 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 10304 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_8_119
timestamp 1604666999
transform 1 0 12052 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 13432 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_131
timestamp 1604666999
transform 1 0 13156 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_145
timestamp 1604666999
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1604666999
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1604666999
transform 1 0 15916 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604666999
transform 1 0 16928 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604666999
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 15456 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_154
timestamp 1604666999
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_158
timestamp 1604666999
transform 1 0 15640 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_164
timestamp 1604666999
transform 1 0 16192 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 18032 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 17848 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_176
timestamp 1604666999
transform 1 0 17296 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_180
timestamp 1604666999
transform 1 0 17664 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604666999
transform 1 0 20884 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604666999
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 19964 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_203
timestamp 1604666999
transform 1 0 19780 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_207
timestamp 1604666999
transform 1 0 20148 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1604666999
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_220
timestamp 1604666999
transform 1 0 21344 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604666999
transform 1 0 23644 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 23460 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 23092 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 22724 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_232
timestamp 1604666999
transform 1 0 22448 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_237
timestamp 1604666999
transform 1 0 22908 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_241
timestamp 1604666999
transform 1 0 23276 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604666999
transform 1 0 25300 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604666999
transform 1 0 24656 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 26220 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 25852 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_254
timestamp 1604666999
transform 1 0 24472 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_258
timestamp 1604666999
transform 1 0 24840 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_262
timestamp 1604666999
transform 1 0 25208 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_267
timestamp 1604666999
transform 1 0 25668 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_271
timestamp 1604666999
transform 1 0 26036 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604666999
transform 1 0 26588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604666999
transform 1 0 27692 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604666999
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 27140 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 27508 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604666999
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_281
timestamp 1604666999
transform 1 0 26956 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_285
timestamp 1604666999
transform 1 0 27324 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_298
timestamp 1604666999
transform 1 0 28520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
timestamp 1604666999
transform 1 0 29256 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
timestamp 1604666999
transform 1 0 28704 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
timestamp 1604666999
transform 1 0 29072 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_302
timestamp 1604666999
transform 1 0 28888 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604666999
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_325
timestamp 1604666999
transform 1 0 31004 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_333
timestamp 1604666999
transform 1 0 31740 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_337
timestamp 1604666999
transform 1 0 32108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_349
timestamp 1604666999
transform 1 0 33212 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_361
timestamp 1604666999
transform 1 0 34316 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604666999
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_373
timestamp 1604666999
transform 1 0 35420 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_385
timestamp 1604666999
transform 1 0 36524 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604666999
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_398
timestamp 1604666999
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_406
timestamp 1604666999
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604666999
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604666999
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604666999
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604666999
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
timestamp 1604666999
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_27
timestamp 1604666999
transform 1 0 3588 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_33
timestamp 1604666999
transform 1 0 4140 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_36
timestamp 1604666999
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_40
timestamp 1604666999
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_53
timestamp 1604666999
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1604666999
transform 1 0 6348 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
timestamp 1604666999
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1604666999
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604666999
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_69
timestamp 1604666999
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_66
timestamp 1604666999
transform 1 0 7176 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_73
timestamp 1604666999
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604666999
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604666999
transform 1 0 8188 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604666999
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_96
timestamp 1604666999
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_100
timestamp 1604666999
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604666999
transform 1 0 10672 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_117
timestamp 1604666999
transform 1 0 11868 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1604666999
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 12052 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1604666999
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604666999
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604666999
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 13892 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 13708 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604666999
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 13340 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_127
timestamp 1604666999
transform 1 0 12788 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_131
timestamp 1604666999
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_135
timestamp 1604666999
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604666999
transform 1 0 16836 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_158
timestamp 1604666999
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_162
timestamp 1604666999
transform 1 0 16008 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_170
timestamp 1604666999
transform 1 0 16744 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_184
timestamp 1604666999
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_179
timestamp 1604666999
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_175
timestamp 1604666999
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604666999
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604666999
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604666999
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_189
timestamp 1604666999
transform 1 0 18492 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 18308 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 18676 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 18860 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
timestamp 1604666999
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 20792 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_212
timestamp 1604666999
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_216
timestamp 1604666999
transform 1 0 20976 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_220
timestamp 1604666999
transform 1 0 21344 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_223
timestamp 1604666999
transform 1 0 21620 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604666999
transform 1 0 23920 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604666999
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
timestamp 1604666999
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604666999
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
timestamp 1604666999
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_227
timestamp 1604666999
transform 1 0 21988 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_235
timestamp 1604666999
transform 1 0 22724 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_240
timestamp 1604666999
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_245
timestamp 1604666999
transform 1 0 23644 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
timestamp 1604666999
transform 1 0 26220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
timestamp 1604666999
transform 1 0 25852 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_267
timestamp 1604666999
transform 1 0 25668 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_271
timestamp 1604666999
transform 1 0 26036 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
timestamp 1604666999
transform 1 0 26404 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
timestamp 1604666999
transform 1 0 28336 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_294
timestamp 1604666999
transform 1 0 28152 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_298
timestamp 1604666999
transform 1 0 28520 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
timestamp 1604666999
transform 1 0 29256 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604666999
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
timestamp 1604666999
transform 1 0 28704 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_302
timestamp 1604666999
transform 1 0 28888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_325
timestamp 1604666999
transform 1 0 31004 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1604666999
transform 1 0 32108 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604666999
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1604666999
transform 1 0 33212 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_361
timestamp 1604666999
transform 1 0 34316 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_365
timestamp 1604666999
transform 1 0 34684 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_367
timestamp 1604666999
transform 1 0 34868 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_379
timestamp 1604666999
transform 1 0 35972 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_391
timestamp 1604666999
transform 1 0 37076 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604666999
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_403
timestamp 1604666999
transform 1 0 38180 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604666999
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604666999
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604666999
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
timestamp 1604666999
transform 1 0 5428 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604666999
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604666999
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1604666999
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_46
timestamp 1604666999
transform 1 0 5336 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604666999
transform 1 0 7912 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
timestamp 1604666999
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_66
timestamp 1604666999
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_70
timestamp 1604666999
transform 1 0 7544 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 9936 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604666999
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_83
timestamp 1604666999
transform 1 0 8740 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1604666999
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_93
timestamp 1604666999
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_115
timestamp 1604666999
transform 1 0 11684 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1604666999
transform 1 0 12696 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1604666999
transform 1 0 13708 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 13156 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 13524 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_125
timestamp 1604666999
transform 1 0 12604 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_129
timestamp 1604666999
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_133
timestamp 1604666999
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_140
timestamp 1604666999
transform 1 0 13984 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 15272 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604666999
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1604666999
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_173
timestamp 1604666999
transform 1 0 17020 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604666999
transform 1 0 19228 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604666999
transform 1 0 17756 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 18860 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 17204 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_177
timestamp 1604666999
transform 1 0 17388 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_185
timestamp 1604666999
transform 1 0 18124 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_195
timestamp 1604666999
transform 1 0 19044 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
timestamp 1604666999
transform 1 0 21436 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604666999
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 21068 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_206
timestamp 1604666999
transform 1 0 20056 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_215
timestamp 1604666999
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_219
timestamp 1604666999
transform 1 0 21252 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
timestamp 1604666999
transform 1 0 23920 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
timestamp 1604666999
transform 1 0 23736 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_240
timestamp 1604666999
transform 1 0 23184 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_267
timestamp 1604666999
transform 1 0 25668 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604666999
transform 1 0 26864 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604666999
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
timestamp 1604666999
transform 1 0 26680 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
timestamp 1604666999
transform 1 0 27968 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_276
timestamp 1604666999
transform 1 0 26496 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_289
timestamp 1604666999
transform 1 0 27692 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_294
timestamp 1604666999
transform 1 0 28152 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
timestamp 1604666999
transform 1 0 28704 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_10_319
timestamp 1604666999
transform 1 0 30452 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604666999
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_331
timestamp 1604666999
transform 1 0 31556 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_335
timestamp 1604666999
transform 1 0 31924 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_337
timestamp 1604666999
transform 1 0 32108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_349
timestamp 1604666999
transform 1 0 33212 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_361
timestamp 1604666999
transform 1 0 34316 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604666999
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_373
timestamp 1604666999
transform 1 0 35420 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_385
timestamp 1604666999
transform 1 0 36524 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604666999
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_398
timestamp 1604666999
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_406
timestamp 1604666999
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604666999
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604666999
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604666999
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1604666999
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1604666999
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
timestamp 1604666999
transform 1 0 6808 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604666999
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
timestamp 1604666999
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
timestamp 1604666999
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1604666999
transform 1 0 5796 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1604666999
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_81
timestamp 1604666999
transform 1 0 8556 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_89
timestamp 1604666999
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_93
timestamp 1604666999
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_97
timestamp 1604666999
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10396 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 12420 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604666999
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1604666999
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_114
timestamp 1604666999
transform 1 0 11592 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_142
timestamp 1604666999
transform 1 0 14168 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_146
timestamp 1604666999
transform 1 0 14536 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1604666999
transform 1 0 14904 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604666999
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_153
timestamp 1604666999
transform 1 0 15180 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_158
timestamp 1604666999
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_162
timestamp 1604666999
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_175
timestamp 1604666999
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_179
timestamp 1604666999
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604666999
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604666999
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_188
timestamp 1604666999
transform 1 0 18400 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604666999
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_192
timestamp 1604666999
transform 1 0 18768 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_195
timestamp 1604666999
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_203
timestamp 1604666999
transform 1 0 19780 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604666999
transform 1 0 19412 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_207
timestamp 1604666999
transform 1 0 20148 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 19964 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604666999
transform 1 0 20516 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604666999
transform 1 0 20700 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_217
timestamp 1604666999
transform 1 0 21068 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1604666999
transform 1 0 21436 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 21252 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 21620 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604666999
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
timestamp 1604666999
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
timestamp 1604666999
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_225
timestamp 1604666999
transform 1 0 21804 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_233
timestamp 1604666999
transform 1 0 22540 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_236
timestamp 1604666999
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_240
timestamp 1604666999
transform 1 0 23184 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_245
timestamp 1604666999
transform 1 0 23644 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604666999
transform 1 0 25116 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 24932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 24564 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_253
timestamp 1604666999
transform 1 0 24380 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_257
timestamp 1604666999
transform 1 0 24748 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_270
timestamp 1604666999
transform 1 0 25944 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
timestamp 1604666999
transform 1 0 26680 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
timestamp 1604666999
transform 1 0 26496 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_297
timestamp 1604666999
transform 1 0 28428 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604666999
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
timestamp 1604666999
transform 1 0 28612 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_301
timestamp 1604666999
transform 1 0 28796 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_306
timestamp 1604666999
transform 1 0 29256 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_318
timestamp 1604666999
transform 1 0 30360 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_330
timestamp 1604666999
transform 1 0 31464 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_342
timestamp 1604666999
transform 1 0 32568 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604666999
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_354
timestamp 1604666999
transform 1 0 33672 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_367
timestamp 1604666999
transform 1 0 34868 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_379
timestamp 1604666999
transform 1 0 35972 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_391
timestamp 1604666999
transform 1 0 37076 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604666999
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_403
timestamp 1604666999
transform 1 0 38180 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604666999
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604666999
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604666999
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604666999
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604666999
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1604666999
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1604666999
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
timestamp 1604666999
transform 1 0 6992 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
timestamp 1604666999
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_56
timestamp 1604666999
transform 1 0 6256 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604666999
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_83
timestamp 1604666999
transform 1 0 8740 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1604666999
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_93
timestamp 1604666999
transform 1 0 9660 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 10580 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10396 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_122
timestamp 1604666999
transform 1 0 12328 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604666999
transform 1 0 13064 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 12880 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_139
timestamp 1604666999
transform 1 0 13892 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 16192 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604666999
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1604666999
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_154
timestamp 1604666999
transform 1 0 15272 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_162
timestamp 1604666999
transform 1 0 16008 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604666999
transform 1 0 18860 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 18124 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 18492 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_183
timestamp 1604666999
transform 1 0 17940 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_187
timestamp 1604666999
transform 1 0 18308 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_191
timestamp 1604666999
transform 1 0 18676 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604666999
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604666999
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604666999
transform 1 0 19872 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_202
timestamp 1604666999
transform 1 0 19688 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_206
timestamp 1604666999
transform 1 0 20056 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
timestamp 1604666999
transform 1 0 22632 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_12_224
timestamp 1604666999
transform 1 0 21712 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_232
timestamp 1604666999
transform 1 0 22448 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 25116 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_253
timestamp 1604666999
transform 1 0 24380 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_263
timestamp 1604666999
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
timestamp 1604666999
transform 1 0 27968 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604666999
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_276
timestamp 1604666999
transform 1 0 26496 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_288
timestamp 1604666999
transform 1 0 27600 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_311
timestamp 1604666999
transform 1 0 29716 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604666999
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_323
timestamp 1604666999
transform 1 0 30820 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_335
timestamp 1604666999
transform 1 0 31924 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_337
timestamp 1604666999
transform 1 0 32108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_349
timestamp 1604666999
transform 1 0 33212 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_361
timestamp 1604666999
transform 1 0 34316 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604666999
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_373
timestamp 1604666999
transform 1 0 35420 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_385
timestamp 1604666999
transform 1 0 36524 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604666999
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_398
timestamp 1604666999
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_406
timestamp 1604666999
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604666999
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604666999
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604666999
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604666999
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604666999
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604666999
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_36
timestamp 1604666999
transform 1 0 4416 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 1604666999
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604666999
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
timestamp 1604666999
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604666999
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_41
timestamp 1604666999
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_45
timestamp 1604666999
transform 1 0 5244 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_39
timestamp 1604666999
transform 1 0 4692 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
timestamp 1604666999
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604666999
transform 1 0 4692 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
timestamp 1604666999
transform 1 0 5060 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_49
timestamp 1604666999
transform 1 0 5612 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1604666999
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
timestamp 1604666999
transform 1 0 5060 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_14_66
timestamp 1604666999
transform 1 0 7176 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_62
timestamp 1604666999
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1604666999
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604666999
transform 1 0 6992 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
timestamp 1604666999
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604666999
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604666999
transform 1 0 7176 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_74
timestamp 1604666999
transform 1 0 7912 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_70
timestamp 1604666999
transform 1 0 7544 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604666999
transform 1 0 7728 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604666999
transform 1 0 7912 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_14_83
timestamp 1604666999
transform 1 0 8740 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_82
timestamp 1604666999
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604666999
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604666999
transform 1 0 8280 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1604666999
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_90
timestamp 1604666999
transform 1 0 9384 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_86
timestamp 1604666999
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604666999
transform 1 0 9200 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604666999
transform 1 0 8832 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604666999
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_97
timestamp 1604666999
transform 1 0 10028 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_95
timestamp 1604666999
transform 1 0 9844 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604666999
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604666999
transform 1 0 9660 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_107
timestamp 1604666999
transform 1 0 10948 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_103
timestamp 1604666999
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604666999
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604666999
transform 1 0 10764 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_121
timestamp 1604666999
transform 1 0 12236 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_123
timestamp 1604666999
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_118
timestamp 1604666999
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_115
timestamp 1604666999
transform 1 0 11684 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604666999
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1604666999
transform 1 0 11132 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_125
timestamp 1604666999
transform 1 0 12604 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604666999
transform 1 0 12880 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1604666999
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_145
timestamp 1604666999
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_148
timestamp 1604666999
transform 1 0 14720 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_141
timestamp 1604666999
transform 1 0 14076 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_137
timestamp 1604666999
transform 1 0 13708 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCD
timestamp 1604666999
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1604666999
transform 1 0 14444 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 12696 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_13_158
timestamp 1604666999
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604666999
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_168
timestamp 1604666999
transform 1 0 16560 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_162
timestamp 1604666999
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 16376 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604666999
transform 1 0 16376 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1604666999
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 16836 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_13_179
timestamp 1604666999
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_175
timestamp 1604666999
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604666999
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_190
timestamp 1604666999
transform 1 0 18584 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_193
timestamp 1604666999
transform 1 0 18860 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 18768 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604666999
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_194
timestamp 1604666999
transform 1 0 18952 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_197
timestamp 1604666999
transform 1 0 19228 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604666999
transform 1 0 19320 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604666999
transform 1 0 19320 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_208
timestamp 1604666999
transform 1 0 20240 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_200
timestamp 1604666999
transform 1 0 19504 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 20516 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604666999
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604666999
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604666999
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_213
timestamp 1604666999
transform 1 0 20700 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_217
timestamp 1604666999
transform 1 0 21068 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 21252 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 21436 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_219
timestamp 1604666999
transform 1 0 21252 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_223
timestamp 1604666999
transform 1 0 21620 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604666999
transform 1 0 21436 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_14_202
timestamp 1604666999
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_233
timestamp 1604666999
transform 1 0 22540 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_229
timestamp 1604666999
transform 1 0 22172 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_230
timestamp 1604666999
transform 1 0 22264 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604666999
transform 1 0 22356 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604666999
transform 1 0 21988 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_243
timestamp 1604666999
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_239
timestamp 1604666999
transform 1 0 23092 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_236
timestamp 1604666999
transform 1 0 22816 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
timestamp 1604666999
transform 1 0 22908 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
timestamp 1604666999
transform 1 0 23092 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
timestamp 1604666999
transform 1 0 23276 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604666999
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604666999
transform 1 0 23644 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
timestamp 1604666999
transform 1 0 23276 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604666999
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604666999
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604666999
transform 1 0 25392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_254
timestamp 1604666999
transform 1 0 24472 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_258
timestamp 1604666999
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_262
timestamp 1604666999
transform 1 0 25208 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_266
timestamp 1604666999
transform 1 0 25576 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_260
timestamp 1604666999
transform 1 0 25024 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_272
timestamp 1604666999
transform 1 0 26128 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604666999
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_278
timestamp 1604666999
transform 1 0 26680 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_290
timestamp 1604666999
transform 1 0 27784 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_276
timestamp 1604666999
transform 1 0 26496 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_288
timestamp 1604666999
transform 1 0 27600 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_308
timestamp 1604666999
transform 1 0 29440 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_300
timestamp 1604666999
transform 1 0 28704 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_306
timestamp 1604666999
transform 1 0 29256 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_302
timestamp 1604666999
transform 1 0 28888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 29624 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604666999
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604666999
transform 1 0 29624 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_316
timestamp 1604666999
transform 1 0 30176 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_312
timestamp 1604666999
transform 1 0 29808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 30360 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 29992 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_319
timestamp 1604666999
transform 1 0 30452 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_320
timestamp 1604666999
transform 1 0 30544 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_335
timestamp 1604666999
transform 1 0 31924 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_331
timestamp 1604666999
transform 1 0 31556 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_345
timestamp 1604666999
transform 1 0 32844 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_341
timestamp 1604666999
transform 1 0 32476 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_337
timestamp 1604666999
transform 1 0 32108 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_344
timestamp 1604666999
transform 1 0 32752 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
timestamp 1604666999
transform 1 0 32660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
timestamp 1604666999
transform 1 0 32292 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
timestamp 1604666999
transform 1 0 32936 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604666999
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_332
timestamp 1604666999
transform 1 0 31648 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
timestamp 1604666999
transform 1 0 32936 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604666999
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
timestamp 1604666999
transform 1 0 33304 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_348
timestamp 1604666999
transform 1 0 33120 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_352
timestamp 1604666999
transform 1 0 33488 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_364
timestamp 1604666999
transform 1 0 34592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_367
timestamp 1604666999
transform 1 0 34868 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_365
timestamp 1604666999
transform 1 0 34684 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604666999
transform 1 0 35420 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604666999
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604666999
transform 1 0 35420 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_375
timestamp 1604666999
transform 1 0 35604 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_387
timestamp 1604666999
transform 1 0 36708 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1604666999
transform 1 0 35788 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_389
timestamp 1604666999
transform 1 0 36892 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604666999
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604666999
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_399
timestamp 1604666999
transform 1 0 37812 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_398
timestamp 1604666999
transform 1 0 37720 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_406
timestamp 1604666999
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604666999
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1604666999
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1604666999
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
timestamp 1604666999
transform 1 0 4232 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
timestamp 1604666999
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604666999
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_27
timestamp 1604666999
transform 1 0 3588 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_30
timestamp 1604666999
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604666999
transform 1 0 7084 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604666999
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
timestamp 1604666999
transform 1 0 6256 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604666999
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1604666999
transform 1 0 5980 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_58
timestamp 1604666999
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_62
timestamp 1604666999
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_69
timestamp 1604666999
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_73
timestamp 1604666999
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
timestamp 1604666999
transform 1 0 8188 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
timestamp 1604666999
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
timestamp 1604666999
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_96
timestamp 1604666999
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_104
timestamp 1604666999
transform 1 0 10672 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_100
timestamp 1604666999
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
timestamp 1604666999
transform 1 0 10488 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_108
timestamp 1604666999
transform 1 0 11040 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604666999
transform 1 0 11132 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1604666999
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_117
timestamp 1604666999
transform 1 0 11868 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604666999
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_123
timestamp 1604666999
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604666999
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_
timestamp 1604666999
transform 1 0 13708 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCE
timestamp 1604666999
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 12696 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__D
timestamp 1604666999
transform 1 0 13156 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_128
timestamp 1604666999
transform 1 0 12880 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_133
timestamp 1604666999
transform 1 0 13340 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604666999
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_161
timestamp 1604666999
transform 1 0 15916 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 18032 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604666999
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604666999
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1604666999
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 1604666999
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 21252 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 20516 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_203
timestamp 1604666999
transform 1 0 19780 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_213
timestamp 1604666999
transform 1 0 20700 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_217
timestamp 1604666999
transform 1 0 21068 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_221
timestamp 1604666999
transform 1 0 21436 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604666999
transform 1 0 21988 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
timestamp 1604666999
transform 1 0 23644 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604666999
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
timestamp 1604666999
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
timestamp 1604666999
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604666999
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_236
timestamp 1604666999
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_240
timestamp 1604666999
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_264
timestamp 1604666999
transform 1 0 25392 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
timestamp 1604666999
transform 1 0 28152 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
timestamp 1604666999
transform 1 0 28520 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_276
timestamp 1604666999
transform 1 0 26496 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_288
timestamp 1604666999
transform 1 0 27600 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_296
timestamp 1604666999
transform 1 0 28336 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
timestamp 1604666999
transform 1 0 29624 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604666999
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
timestamp 1604666999
transform 1 0 29440 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
timestamp 1604666999
transform 1 0 28980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_300
timestamp 1604666999
transform 1 0 28704 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_306
timestamp 1604666999
transform 1 0 29256 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
timestamp 1604666999
transform 1 0 32108 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
timestamp 1604666999
transform 1 0 31924 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
timestamp 1604666999
transform 1 0 31556 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_329
timestamp 1604666999
transform 1 0 31372 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_333
timestamp 1604666999
transform 1 0 31740 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604666999
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
timestamp 1604666999
transform 1 0 34592 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
timestamp 1604666999
transform 1 0 35052 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_356
timestamp 1604666999
transform 1 0 33856 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_367
timestamp 1604666999
transform 1 0 34868 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_371
timestamp 1604666999
transform 1 0 35236 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604666999
transform 1 0 35420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604666999
transform 1 0 35972 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_377
timestamp 1604666999
transform 1 0 35788 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_381
timestamp 1604666999
transform 1 0 36156 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1604666999
transform 1 0 37260 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604666999
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1604666999
transform 1 0 38364 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604666999
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1604666999
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1604666999
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604666999
transform 1 0 4692 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604666999
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604666999
transform 1 0 4508 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1604666999
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_32
timestamp 1604666999
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_36
timestamp 1604666999
transform 1 0 4416 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_48
timestamp 1604666999
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
timestamp 1604666999
transform 1 0 6256 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 5704 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 6072 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_52
timestamp 1604666999
transform 1 0 5888 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_83
timestamp 1604666999
transform 1 0 8740 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_79
timestamp 1604666999
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_75
timestamp 1604666999
transform 1 0 8004 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 8556 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
timestamp 1604666999
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
timestamp 1604666999
transform 1 0 8188 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_88
timestamp 1604666999
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604666999
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
timestamp 1604666999
transform 1 0 9660 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_16_112
timestamp 1604666999
transform 1 0 11408 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_124
timestamp 1604666999
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 12696 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_16_145
timestamp 1604666999
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604666999
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1604666999
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1604666999
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604666999
transform 1 0 17848 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_16_178
timestamp 1604666999
transform 1 0 17480 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604666999
transform 1 0 21252 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604666999
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
timestamp 1604666999
transform 1 0 19780 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604666999
transform 1 0 21068 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604666999
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_201
timestamp 1604666999
transform 1 0 19596 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_205
timestamp 1604666999
transform 1 0 19964 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_211
timestamp 1604666999
transform 1 0 20516 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_215
timestamp 1604666999
transform 1 0 20884 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
timestamp 1604666999
transform 1 0 23460 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
timestamp 1604666999
transform 1 0 23276 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
timestamp 1604666999
transform 1 0 22908 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
timestamp 1604666999
transform 1 0 22540 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_228
timestamp 1604666999
transform 1 0 22080 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_232
timestamp 1604666999
transform 1 0 22448 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_235
timestamp 1604666999
transform 1 0 22724 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_239
timestamp 1604666999
transform 1 0 23092 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_262
timestamp 1604666999
transform 1 0 25208 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
timestamp 1604666999
transform 1 0 28152 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604666999
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604666999
transform 1 0 27600 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 26680 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604666999
transform 1 0 27968 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_274
timestamp 1604666999
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_276
timestamp 1604666999
transform 1 0 26496 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_280
timestamp 1604666999
transform 1 0 26864 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_290
timestamp 1604666999
transform 1 0 27784 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 30084 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 30452 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_313
timestamp 1604666999
transform 1 0 29900 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_317
timestamp 1604666999
transform 1 0 30268 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_321
timestamp 1604666999
transform 1 0 30636 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
timestamp 1604666999
transform 1 0 32108 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604666999
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 30820 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_325
timestamp 1604666999
transform 1 0 31004 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_333
timestamp 1604666999
transform 1 0 31740 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
timestamp 1604666999
transform 1 0 34592 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604666999
transform 1 0 34040 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_356
timestamp 1604666999
transform 1 0 33856 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_360
timestamp 1604666999
transform 1 0 34224 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604666999
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_383
timestamp 1604666999
transform 1 0 36340 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_395
timestamp 1604666999
transform 1 0 37444 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604666999
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_398
timestamp 1604666999
transform 1 0 37720 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_406
timestamp 1604666999
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604666999
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1604666999
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_15
timestamp 1604666999
transform 1 0 2484 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_23
timestamp 1604666999
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
timestamp 1604666999
transform 1 0 3956 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
timestamp 1604666999
transform 1 0 3772 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
timestamp 1604666999
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_27
timestamp 1604666999
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604666999
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604666999
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604666999
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604666999
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_50
timestamp 1604666999
transform 1 0 5704 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_54
timestamp 1604666999
transform 1 0 6072 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1604666999
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_71
timestamp 1604666999
transform 1 0 7636 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
timestamp 1604666999
transform 1 0 9016 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
timestamp 1604666999
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_77
timestamp 1604666999
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_81
timestamp 1604666999
transform 1 0 8556 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604666999
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604666999
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604666999
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_105
timestamp 1604666999
transform 1 0 10764 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_109
timestamp 1604666999
transform 1 0 11132 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_112
timestamp 1604666999
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_116
timestamp 1604666999
transform 1 0 11776 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_123
timestamp 1604666999
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 13156 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 12972 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 12604 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_127
timestamp 1604666999
transform 1 0 12788 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 16652 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_150
timestamp 1604666999
transform 1 0 14904 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_162
timestamp 1604666999
transform 1 0 16008 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_168
timestamp 1604666999
transform 1 0 16560 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_171
timestamp 1604666999
transform 1 0 16836 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_184
timestamp 1604666999
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_179
timestamp 1604666999
transform 1 0 17572 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1604666999
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
timestamp 1604666999
transform 1 0 18216 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604666999
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_192
timestamp 1604666999
transform 1 0 18768 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_188
timestamp 1604666999
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
timestamp 1604666999
transform 1 0 18584 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
timestamp 1604666999
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
timestamp 1604666999
transform 1 0 19228 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604666999
transform 1 0 21528 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604666999
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_216
timestamp 1604666999
transform 1 0 20976 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_220
timestamp 1604666999
transform 1 0 21344 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604666999
transform 1 0 21988 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
timestamp 1604666999
transform 1 0 23644 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604666999
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 21712 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
timestamp 1604666999
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
timestamp 1604666999
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_236
timestamp 1604666999
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_240
timestamp 1604666999
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_264
timestamp 1604666999
transform 1 0 25392 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 26680 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 26496 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_297
timestamp 1604666999
transform 1 0 28428 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
timestamp 1604666999
transform 1 0 29256 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604666999
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
timestamp 1604666999
transform 1 0 28980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
timestamp 1604666999
transform 1 0 28612 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_301
timestamp 1604666999
transform 1 0 28796 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604666999
transform 1 0 32292 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604666999
transform 1 0 32108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604666999
transform 1 0 31740 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604666999
transform 1 0 31372 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_325
timestamp 1604666999
transform 1 0 31004 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_331
timestamp 1604666999
transform 1 0 31556 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_335
timestamp 1604666999
transform 1 0 31924 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_358
timestamp 1604666999
transform 1 0 34040 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_354
timestamp 1604666999
transform 1 0 33672 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_348
timestamp 1604666999
transform 1 0 33120 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604666999
transform 1 0 33856 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
timestamp 1604666999
transform 1 0 34224 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604666999
transform 1 0 33488 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_362
timestamp 1604666999
transform 1 0 34408 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
timestamp 1604666999
transform 1 0 34592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604666999
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
timestamp 1604666999
transform 1 0 34868 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
timestamp 1604666999
transform 1 0 36800 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_386
timestamp 1604666999
transform 1 0 36616 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_390
timestamp 1604666999
transform 1 0 36984 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604666999
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_402
timestamp 1604666999
transform 1 0 38088 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_406
timestamp 1604666999
transform 1 0 38456 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604666999
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1604666999
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1604666999
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604666999
transform 1 0 5152 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604666999
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604666999
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604666999
transform 1 0 4968 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 4232 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1604666999
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_32
timestamp 1604666999
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_36
timestamp 1604666999
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_40
timestamp 1604666999
transform 1 0 4784 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604666999
transform 1 0 6716 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604666999
transform 1 0 7268 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604666999
transform 1 0 7636 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_53
timestamp 1604666999
transform 1 0 5980 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_65
timestamp 1604666999
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_69
timestamp 1604666999
transform 1 0 7452 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_73
timestamp 1604666999
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604666999
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604666999
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_84
timestamp 1604666999
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_88
timestamp 1604666999
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604666999
transform 1 0 11224 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1604666999
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_106
timestamp 1604666999
transform 1 0 10856 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_115
timestamp 1604666999
transform 1 0 11684 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_123
timestamp 1604666999
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 13156 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_127
timestamp 1604666999
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_140
timestamp 1604666999
transform 1 0 13984 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_148
timestamp 1604666999
transform 1 0 14720 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1604666999
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604666999
transform 1 0 16652 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604666999
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 15732 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_157
timestamp 1604666999
transform 1 0 15548 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_161
timestamp 1604666999
transform 1 0 15916 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_165
timestamp 1604666999
transform 1 0 16284 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
timestamp 1604666999
transform 1 0 18216 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
timestamp 1604666999
transform 1 0 18032 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_178
timestamp 1604666999
transform 1 0 17480 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604666999
transform 1 0 21068 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604666999
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
timestamp 1604666999
transform 1 0 20516 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_205
timestamp 1604666999
transform 1 0 19964 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1604666999
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_215
timestamp 1604666999
transform 1 0 20884 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
timestamp 1604666999
transform 1 0 22632 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604666999
transform 1 0 22080 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604666999
transform 1 0 22448 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_226
timestamp 1604666999
transform 1 0 21896 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_230
timestamp 1604666999
transform 1 0 22264 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1604666999
transform 1 0 24380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_265
timestamp 1604666999
transform 1 0 25484 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_273
timestamp 1604666999
transform 1 0 26220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604666999
transform 1 0 27600 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604666999
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 26680 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 27048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 27416 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_276
timestamp 1604666999
transform 1 0 26496 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_280
timestamp 1604666999
transform 1 0 26864 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_284
timestamp 1604666999
transform 1 0 27232 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604666999
transform 1 0 30084 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 29532 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 29900 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_307
timestamp 1604666999
transform 1 0 29348 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_311
timestamp 1604666999
transform 1 0 29716 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_324
timestamp 1604666999
transform 1 0 30912 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 31096 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_332
timestamp 1604666999
transform 1 0 31648 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_328
timestamp 1604666999
transform 1 0 31280 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 31464 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_337
timestamp 1604666999
transform 1 0 32108 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 31832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604666999
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604666999
transform 1 0 32384 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_344
timestamp 1604666999
transform 1 0 32752 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604666999
transform 1 0 32936 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604666999
transform 1 0 33488 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
timestamp 1604666999
transform 1 0 35144 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
timestamp 1604666999
transform 1 0 34868 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 33304 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604666999
transform 1 0 34500 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_348
timestamp 1604666999
transform 1 0 33120 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_361
timestamp 1604666999
transform 1 0 34316 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1604666999
transform 1 0 34684 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_369
timestamp 1604666999
transform 1 0 35052 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604666999
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_389
timestamp 1604666999
transform 1 0 36892 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604666999
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_398
timestamp 1604666999
transform 1 0 37720 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_406
timestamp 1604666999
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604666999
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604666999
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
timestamp 1604666999
transform 1 0 3312 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1604666999
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_15
timestamp 1604666999
transform 1 0 2484 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_23
timestamp 1604666999
transform 1 0 3220 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1604666999
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1604666999
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_36
timestamp 1604666999
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_32
timestamp 1604666999
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1604666999
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_26
timestamp 1604666999
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
timestamp 1604666999
transform 1 0 4232 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
timestamp 1604666999
transform 1 0 3680 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604666999
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_49
timestamp 1604666999
transform 1 0 5612 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604666999
transform 1 0 4600 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_20_47
timestamp 1604666999
transform 1 0 5428 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
timestamp 1604666999
transform 1 0 3864 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_20_59
timestamp 1604666999
transform 1 0 6532 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_53
timestamp 1604666999
transform 1 0 5980 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604666999
transform 1 0 5796 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_69
timestamp 1604666999
transform 1 0 7452 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_64
timestamp 1604666999
transform 1 0 6992 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_62
timestamp 1604666999
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604666999
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 7084 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604666999
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604666999
transform 1 0 7268 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_20_84
timestamp 1604666999
transform 1 0 8832 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_77
timestamp 1604666999
transform 1 0 8188 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_82
timestamp 1604666999
transform 1 0 8648 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_76
timestamp 1604666999
transform 1 0 8096 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604666999
transform 1 0 8280 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604666999
transform 1 0 8464 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604666999
transform 1 0 8464 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_91
timestamp 1604666999
transform 1 0 9476 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_87
timestamp 1604666999
transform 1 0 9108 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 9292 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604666999
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 9844 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_20_107
timestamp 1604666999
transform 1 0 10948 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_102
timestamp 1604666999
transform 1 0 10488 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_123
timestamp 1604666999
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_118
timestamp 1604666999
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_114
timestamp 1604666999
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604666999
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 11224 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_20_133
timestamp 1604666999
transform 1 0 13340 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_129
timestamp 1604666999
transform 1 0 12972 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_128
timestamp 1604666999
transform 1 0 12880 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12696 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 13524 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 13156 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 13064 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_148
timestamp 1604666999
transform 1 0 14720 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_144
timestamp 1604666999
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_137
timestamp 1604666999
transform 1 0 13708 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 14536 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1604666999
transform 1 0 14076 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 13248 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1604666999
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_156
timestamp 1604666999
transform 1 0 15456 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_151
timestamp 1604666999
transform 1 0 14996 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604666999
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 15732 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_173
timestamp 1604666999
transform 1 0 17020 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_172
timestamp 1604666999
transform 1 0 16928 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_168
timestamp 1604666999
transform 1 0 16560 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 15272 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604666999
transform 1 0 18584 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
timestamp 1604666999
transform 1 0 18032 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604666999
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
timestamp 1604666999
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 18400 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_180
timestamp 1604666999
transform 1 0 17664 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_181
timestamp 1604666999
transform 1 0 17756 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_186
timestamp 1604666999
transform 1 0 18216 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_211
timestamp 1604666999
transform 1 0 20516 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_207
timestamp 1604666999
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_203
timestamp 1604666999
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 19964 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
timestamp 1604666999
transform 1 0 20332 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_223
timestamp 1604666999
transform 1 0 21620 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_215
timestamp 1604666999
transform 1 0 20884 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604666999
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_199
timestamp 1604666999
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
timestamp 1604666999
transform 1 0 20516 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_19_234
timestamp 1604666999
transform 1 0 22632 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_230
timestamp 1604666999
transform 1 0 22264 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_clk_A
timestamp 1604666999
transform 1 0 21712 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
timestamp 1604666999
transform 1 0 22448 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_245
timestamp 1604666999
transform 1 0 23644 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_238
timestamp 1604666999
transform 1 0 23000 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
timestamp 1604666999
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604666999
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_245
timestamp 1604666999
transform 1 0 23644 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
timestamp 1604666999
transform 1 0 21896 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 24380 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1604666999
transform 1 0 24196 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_273
timestamp 1604666999
transform 1 0 26220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_257
timestamp 1604666999
transform 1 0 24748 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_269
timestamp 1604666999
transform 1 0 25852 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 26496 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 26588 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604666999
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 26404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_296
timestamp 1604666999
transform 1 0 28336 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_295
timestamp 1604666999
transform 1 0 28244 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_301
timestamp 1604666999
transform 1 0 28796 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 28796 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 28612 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 28980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604666999
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604666999
transform 1 0 28980 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604666999
transform 1 0 29256 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_20_312
timestamp 1604666999
transform 1 0 29808 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_315
timestamp 1604666999
transform 1 0 30084 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 30268 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_319
timestamp 1604666999
transform 1 0 30452 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604666999
transform 1 0 30360 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 30636 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604666999
transform 1 0 30544 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_329
timestamp 1604666999
transform 1 0 31372 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_324
timestamp 1604666999
transform 1 0 30912 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_332
timestamp 1604666999
transform 1 0 31648 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 31188 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604666999
transform 1 0 30820 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604666999
transform 1 0 32016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 31832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 31832 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_336
timestamp 1604666999
transform 1 0 32016 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_333
timestamp 1604666999
transform 1 0 31740 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_337
timestamp 1604666999
transform 1 0 32108 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604666999
transform 1 0 32200 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604666999
transform 1 0 32200 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_340
timestamp 1604666999
transform 1 0 32384 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_342
timestamp 1604666999
transform 1 0 32568 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604666999
transform 1 0 32568 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_346
timestamp 1604666999
transform 1 0 32936 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 32752 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_359
timestamp 1604666999
transform 1 0 34132 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_359
timestamp 1604666999
transform 1 0 34132 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_355
timestamp 1604666999
transform 1 0 33764 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_351
timestamp 1604666999
transform 1 0 33396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 33120 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 33580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604666999
transform 1 0 34224 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604666999
transform 1 0 33304 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_363
timestamp 1604666999
transform 1 0 34500 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_367
timestamp 1604666999
transform 1 0 34868 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_362
timestamp 1604666999
transform 1 0 34408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604666999
transform 1 0 34316 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604666999
transform 1 0 34684 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
timestamp 1604666999
transform 1 0 34592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604666999
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604666999
transform 1 0 34868 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
timestamp 1604666999
transform 1 0 35144 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604666999
transform 1 0 37628 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604666999
transform 1 0 36432 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
timestamp 1604666999
transform 1 0 35880 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_389
timestamp 1604666999
transform 1 0 36892 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_376
timestamp 1604666999
transform 1 0 35696 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_380
timestamp 1604666999
transform 1 0 36064 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_386
timestamp 1604666999
transform 1 0 36616 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_394
timestamp 1604666999
transform 1 0 37352 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604666999
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604666999
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_401
timestamp 1604666999
transform 1 0 37996 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_398
timestamp 1604666999
transform 1 0 37720 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_406
timestamp 1604666999
transform 1 0 38456 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604666999
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
timestamp 1604666999
transform 1 0 3036 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604666999
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_15
timestamp 1604666999
transform 1 0 2484 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_23
timestamp 1604666999
transform 1 0 3220 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
timestamp 1604666999
transform 1 0 3956 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
timestamp 1604666999
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
timestamp 1604666999
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_27
timestamp 1604666999
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_54
timestamp 1604666999
transform 1 0 6072 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_50
timestamp 1604666999
transform 1 0 5704 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1604666999
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604666999
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604666999
transform 1 0 6808 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_66
timestamp 1604666999
transform 1 0 7176 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 7360 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_70
timestamp 1604666999
transform 1 0 7544 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604666999
transform 1 0 8372 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604666999
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_75
timestamp 1604666999
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_88
timestamp 1604666999
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_92
timestamp 1604666999
transform 1 0 9568 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_97
timestamp 1604666999
transform 1 0 10028 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604666999
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1604666999
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604666999
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1604666999
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_
timestamp 1604666999
transform 1 0 14352 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 12788 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCE
timestamp 1604666999
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 12604 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCD
timestamp 1604666999
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_136
timestamp 1604666999
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_140
timestamp 1604666999
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_168
timestamp 1604666999
transform 1 0 16560 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604666999
transform 1 0 19136 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604666999
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 18952 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 18584 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_180
timestamp 1604666999
transform 1 0 17664 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_184
timestamp 1604666999
transform 1 0 18032 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_192
timestamp 1604666999
transform 1 0 18768 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 21252 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 21620 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1604666999
transform 1 0 19964 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_217
timestamp 1604666999
transform 1 0 21068 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1604666999
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604666999
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 21988 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1604666999
transform 1 0 21804 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_229
timestamp 1604666999
transform 1 0 22172 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_241
timestamp 1604666999
transform 1 0 23276 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_245
timestamp 1604666999
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk
timestamp 1604666999
transform 1 0 25576 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_clk_A
timestamp 1604666999
transform 1 0 25392 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_257
timestamp 1604666999
transform 1 0 24748 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_263
timestamp 1604666999
transform 1 0 25300 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_269
timestamp 1604666999
transform 1 0 25852 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_273
timestamp 1604666999
transform 1 0 26220 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604666999
transform 1 0 26864 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 26680 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 26312 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_276
timestamp 1604666999
transform 1 0 26496 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_289
timestamp 1604666999
transform 1 0 27692 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_297
timestamp 1604666999
transform 1 0 28428 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_301
timestamp 1604666999
transform 1 0 28796 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604666999
transform 1 0 28612 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604666999
transform 1 0 28980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604666999
transform 1 0 29164 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604666999
transform 1 0 29256 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_310
timestamp 1604666999
transform 1 0 29624 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_317
timestamp 1604666999
transform 1 0 30268 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_314
timestamp 1604666999
transform 1 0 29992 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 30084 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_321
timestamp 1604666999
transform 1 0 30636 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 30452 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604666999
transform 1 0 32752 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 31188 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 31004 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 32568 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 32200 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_336
timestamp 1604666999
transform 1 0 32016 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_340
timestamp 1604666999
transform 1 0 32384 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
timestamp 1604666999
transform 1 0 35052 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604666999
transform 1 0 34776 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
timestamp 1604666999
transform 1 0 34592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604666999
transform 1 0 33764 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
timestamp 1604666999
transform 1 0 34224 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_353
timestamp 1604666999
transform 1 0 33580 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_357
timestamp 1604666999
transform 1 0 33948 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_362
timestamp 1604666999
transform 1 0 34408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_367
timestamp 1604666999
transform 1 0 34868 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604666999
transform 1 0 36984 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_388
timestamp 1604666999
transform 1 0 36800 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_392
timestamp 1604666999
transform 1 0 37168 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604666999
transform -1 0 38824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_404
timestamp 1604666999
transform 1 0 38272 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604666999
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604666999
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604666999
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
timestamp 1604666999
transform 1 0 4232 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604666999
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1604666999
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_32
timestamp 1604666999
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604666999
transform 1 0 6716 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604666999
transform 1 0 7728 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_53
timestamp 1604666999
transform 1 0 5980 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_70
timestamp 1604666999
transform 1 0 7544 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_74
timestamp 1604666999
transform 1 0 7912 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604666999
transform 1 0 9844 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604666999
transform 1 0 8280 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604666999
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 8096 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1604666999
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_86
timestamp 1604666999
transform 1 0 9016 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1604666999
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_99
timestamp 1604666999
transform 1 0 10212 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1604666999
transform 1 0 11500 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 12512 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 10764 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_107
timestamp 1604666999
transform 1 0 10948 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_116
timestamp 1604666999
transform 1 0 11776 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__D
timestamp 1604666999
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_143
timestamp 1604666999
transform 1 0 14260 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_147
timestamp 1604666999
transform 1 0 14628 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604666999
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1604666999
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1604666999
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 19136 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1604666999
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_190
timestamp 1604666999
transform 1 0 18584 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_198
timestamp 1604666999
transform 1 0 19320 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604666999
transform 1 0 21252 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604666999
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
timestamp 1604666999
transform 1 0 21068 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_210
timestamp 1604666999
transform 1 0 20424 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1604666999
transform 1 0 20884 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 23920 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_228
timestamp 1604666999
transform 1 0 22080 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_240
timestamp 1604666999
transform 1 0 23184 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 24288 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1604666999
transform 1 0 24104 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_254
timestamp 1604666999
transform 1 0 24472 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_266
timestamp 1604666999
transform 1 0 25576 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604666999
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 26864 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_274
timestamp 1604666999
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_276
timestamp 1604666999
transform 1 0 26496 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_282
timestamp 1604666999
transform 1 0 27048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_294
timestamp 1604666999
transform 1 0 28152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604666999
transform 1 0 30452 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604666999
transform 1 0 29348 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 30268 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_306
timestamp 1604666999
transform 1 0 29256 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_311
timestamp 1604666999
transform 1 0 29716 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604666999
transform 1 0 32108 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604666999
transform 1 0 32016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 31832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 31464 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_328
timestamp 1604666999
transform 1 0 31280 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_332
timestamp 1604666999
transform 1 0 31648 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_346
timestamp 1604666999
transform 1 0 32936 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604666999
transform 1 0 34868 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604666999
transform 1 0 33672 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604666999
transform 1 0 34684 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604666999
transform 1 0 34316 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 33304 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_352
timestamp 1604666999
transform 1 0 33488 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_358
timestamp 1604666999
transform 1 0 34040 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_363
timestamp 1604666999
transform 1 0 34500 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604666999
transform 1 0 36432 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604666999
transform 1 0 37628 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 35880 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_376
timestamp 1604666999
transform 1 0 35696 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_380
timestamp 1604666999
transform 1 0 36064 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_389
timestamp 1604666999
transform 1 0 36892 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604666999
transform -1 0 38824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_398
timestamp 1604666999
transform 1 0 37720 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_406
timestamp 1604666999
transform 1 0 38456 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604666999
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604666999
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604666999
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
timestamp 1604666999
transform 1 0 4232 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
timestamp 1604666999
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_27
timestamp 1604666999
transform 1 0 3588 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_31
timestamp 1604666999
transform 1 0 3956 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_62
timestamp 1604666999
transform 1 0 6808 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604666999
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1604666999
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
timestamp 1604666999
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
timestamp 1604666999
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1604666999
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_68
timestamp 1604666999
transform 1 0 7360 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 7176 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604666999
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604666999
transform 1 0 7728 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_23_91
timestamp 1604666999
transform 1 0 9476 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1604666999
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_103
timestamp 1604666999
transform 1 0 10580 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_115
timestamp 1604666999
transform 1 0 11684 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1604666999
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_123
timestamp 1604666999
transform 1 0 12420 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 13892 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 13708 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_131
timestamp 1604666999
transform 1 0 13156 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_135
timestamp 1604666999
transform 1 0 13524 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_148
timestamp 1604666999
transform 1 0 14720 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_160
timestamp 1604666999
transform 1 0 15824 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_172
timestamp 1604666999
transform 1 0 16928 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1604666999
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
timestamp 1604666999
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
timestamp 1604666999
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_177
timestamp 1604666999
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1604666999
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1604666999
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_196
timestamp 1604666999
transform 1 0 19136 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
timestamp 1604666999
transform 1 0 21068 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
timestamp 1604666999
transform 1 0 20884 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
timestamp 1604666999
transform 1 0 20516 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
timestamp 1604666999
transform 1 0 20148 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_204
timestamp 1604666999
transform 1 0 19872 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_209
timestamp 1604666999
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_213
timestamp 1604666999
transform 1 0 20700 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604666999
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1604666999
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_236
timestamp 1604666999
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_240
timestamp 1604666999
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604666999
transform 1 0 25392 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604666999
transform 1 0 25944 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_254
timestamp 1604666999
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_258
timestamp 1604666999
transform 1 0 24840 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_268
timestamp 1604666999
transform 1 0 25760 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_272
timestamp 1604666999
transform 1 0 26128 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 26496 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 26864 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 27324 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1604666999
transform 1 0 26680 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_282
timestamp 1604666999
transform 1 0 27048 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_287
timestamp 1604666999
transform 1 0 27508 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_299
timestamp 1604666999
transform 1 0 28612 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_310
timestamp 1604666999
transform 1 0 29624 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_306
timestamp 1604666999
transform 1 0 29256 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 29440 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1604666999
transform 1 0 29164 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_317
timestamp 1604666999
transform 1 0 30268 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 29808 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _51_
timestamp 1604666999
transform 1 0 29992 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_321
timestamp 1604666999
transform 1 0 30636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 30452 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 31004 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 30820 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_344
timestamp 1604666999
transform 1 0 32752 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_358
timestamp 1604666999
transform 1 0 34040 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_351
timestamp 1604666999
transform 1 0 33396 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_348
timestamp 1604666999
transform 1 0 33120 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604666999
transform 1 0 33212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
timestamp 1604666999
transform 1 0 34224 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604666999
transform 1 0 33672 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_367
timestamp 1604666999
transform 1 0 34868 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_362
timestamp 1604666999
transform 1 0 34408 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 34592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1604666999
transform 1 0 34776 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
timestamp 1604666999
transform 1 0 35144 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_23_389
timestamp 1604666999
transform 1 0 36892 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604666999
transform -1 0 38824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_401
timestamp 1604666999
transform 1 0 37996 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604666999
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604666999
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604666999
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
timestamp 1604666999
transform 1 0 4968 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1604666999
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
timestamp 1604666999
transform 1 0 4232 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604666999
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_32
timestamp 1604666999
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_36
timestamp 1604666999
transform 1 0 4416 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_61
timestamp 1604666999
transform 1 0 6716 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_67
timestamp 1604666999
transform 1 0 7268 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_71
timestamp 1604666999
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604666999
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1604666999
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_84
timestamp 1604666999
transform 1 0 8832 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_93
timestamp 1604666999
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1604666999
transform 1 0 10028 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1604666999
transform 1 0 11132 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1604666999
transform 1 0 12236 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 13892 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1604666999
transform 1 0 13340 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1604666999
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1604666999
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
timestamp 1604666999
transform 1 0 16836 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604666999
transform 1 0 16376 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604666999
transform 1 0 16008 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_154
timestamp 1604666999
transform 1 0 15272 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_164
timestamp 1604666999
transform 1 0 16192 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_168
timestamp 1604666999
transform 1 0 16560 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_173
timestamp 1604666999
transform 1 0 17020 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
timestamp 1604666999
transform 1 0 17204 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_24_194
timestamp 1604666999
transform 1 0 18952 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
timestamp 1604666999
transform 1 0 21068 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1604666999
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
timestamp 1604666999
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_206
timestamp 1604666999
transform 1 0 20056 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1604666999
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 23920 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 23552 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_236
timestamp 1604666999
transform 1 0 22816 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_246
timestamp 1604666999
transform 1 0 23736 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 26220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_267
timestamp 1604666999
transform 1 0 25668 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 26496 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1604666999
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_295
timestamp 1604666999
transform 1 0 28244 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 30176 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 29532 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 29900 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_307
timestamp 1604666999
transform 1 0 29348 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_311
timestamp 1604666999
transform 1 0 29716 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_315
timestamp 1604666999
transform 1 0 30084 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_325
timestamp 1604666999
transform 1 0 31004 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 31188 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_329
timestamp 1604666999
transform 1 0 31372 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 31556 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_333
timestamp 1604666999
transform 1 0 31740 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1604666999
transform 1 0 32016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604666999
transform 1 0 32108 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_341
timestamp 1604666999
transform 1 0 32476 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_345
timestamp 1604666999
transform 1 0 32844 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604666999
transform 1 0 32660 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604666999
transform 1 0 33212 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 35144 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
timestamp 1604666999
transform 1 0 34960 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604666999
transform 1 0 33764 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_353
timestamp 1604666999
transform 1 0 33580 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_357
timestamp 1604666999
transform 1 0 33948 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_365
timestamp 1604666999
transform 1 0 34684 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1604666999
transform 1 0 37628 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_389
timestamp 1604666999
transform 1 0 36892 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604666999
transform -1 0 38824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_398
timestamp 1604666999
transform 1 0 37720 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_406
timestamp 1604666999
transform 1 0 38456 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604666999
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604666999
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604666999
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604666999
transform 1 0 4876 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 4692 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 4324 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_27
timestamp 1604666999
transform 1 0 3588 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_37
timestamp 1604666999
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604666999
transform 1 0 7084 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1604666999
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 5888 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 6256 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_50
timestamp 1604666999
transform 1 0 5704 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1604666999
transform 1 0 6072 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_58
timestamp 1604666999
transform 1 0 6440 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_62
timestamp 1604666999
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_74
timestamp 1604666999
transform 1 0 7912 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 8648 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 8464 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 8096 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_78
timestamp 1604666999
transform 1 0 8280 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1604666999
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_101
timestamp 1604666999
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_105
timestamp 1604666999
transform 1 0 10764 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_117
timestamp 1604666999
transform 1 0 11868 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1604666999
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1604666999
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1604666999
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_147
timestamp 1604666999
transform 1 0 14628 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604666999
transform 1 0 16376 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604666999
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604666999
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604666999
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604666999
transform 1 0 14904 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_152
timestamp 1604666999
transform 1 0 15088 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_156
timestamp 1604666999
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_160
timestamp 1604666999
transform 1 0 15824 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
timestamp 1604666999
transform 1 0 18032 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1604666999
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
timestamp 1604666999
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
timestamp 1604666999
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1604666999
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_179
timestamp 1604666999
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604666999
transform 1 0 21068 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
timestamp 1604666999
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604666999
transform 1 0 20516 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604666999
transform 1 0 20148 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_203
timestamp 1604666999
transform 1 0 19780 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_209
timestamp 1604666999
transform 1 0 20332 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_213
timestamp 1604666999
transform 1 0 20700 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604666999
transform 1 0 23736 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1604666999
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604666999
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_236
timestamp 1604666999
transform 1 0 22816 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_245
timestamp 1604666999
transform 1 0 23644 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 24840 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 24288 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 24656 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_250
timestamp 1604666999
transform 1 0 24104 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_254
timestamp 1604666999
transform 1 0 24472 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 27324 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 26772 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 27140 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 28336 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_277
timestamp 1604666999
transform 1 0 26588 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1604666999
transform 1 0 26956 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_294
timestamp 1604666999
transform 1 0 28152 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_298
timestamp 1604666999
transform 1 0 28520 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 29348 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1604666999
transform 1 0 29164 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 30728 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 30360 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 28980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_302
timestamp 1604666999
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_306
timestamp 1604666999
transform 1 0 29256 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_316
timestamp 1604666999
transform 1 0 30176 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_320
timestamp 1604666999
transform 1 0 30544 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 30912 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 32844 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_343
timestamp 1604666999
transform 1 0 32660 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_347
timestamp 1604666999
transform 1 0 33028 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1604666999
transform 1 0 34776 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 33212 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_351
timestamp 1604666999
transform 1 0 33396 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_363
timestamp 1604666999
transform 1 0 34500 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_367
timestamp 1604666999
transform 1 0 34868 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_379
timestamp 1604666999
transform 1 0 35972 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_391
timestamp 1604666999
transform 1 0 37076 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604666999
transform -1 0 38824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_403
timestamp 1604666999
transform 1 0 38180 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604666999
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604666999
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604666999
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604666999
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604666999
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604666999
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_32
timestamp 1604666999
transform 1 0 4048 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1604666999
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1604666999
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_43
timestamp 1604666999
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_40
timestamp 1604666999
transform 1 0 4784 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 5244 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604666999
transform 1 0 5428 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1604666999
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1604666999
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604666999
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1604666999
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_56
timestamp 1604666999
transform 1 0 6256 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1604666999
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_74
timestamp 1604666999
transform 1 0 7912 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_71
timestamp 1604666999
transform 1 0 7636 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_67
timestamp 1604666999
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_64
timestamp 1604666999
transform 1 0 6992 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 7084 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604666999
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604666999
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 9660 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 8372 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1604666999
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_84
timestamp 1604666999
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1604666999
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1604666999
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_112
timestamp 1604666999
transform 1 0 11408 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_124
timestamp 1604666999
transform 1 0 12512 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1604666999
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1604666999
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_136
timestamp 1604666999
transform 1 0 13616 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_148
timestamp 1604666999
transform 1 0 14720 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1604666999
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_147
timestamp 1604666999
transform 1 0 14628 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_153
timestamp 1604666999
transform 1 0 15180 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1604666999
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
timestamp 1604666999
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1604666999
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604666999
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_169
timestamp 1604666999
transform 1 0 16652 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1604666999
transform 1 0 16100 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
timestamp 1604666999
transform 1 0 16468 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
timestamp 1604666999
transform 1 0 15456 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
timestamp 1604666999
transform 1 0 16836 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_179
timestamp 1604666999
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1604666999
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
timestamp 1604666999
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1604666999
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604666999
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_197
timestamp 1604666999
transform 1 0 19228 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_193
timestamp 1604666999
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_190
timestamp 1604666999
transform 1 0 18584 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604666999
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
timestamp 1604666999
transform 1 0 18768 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_194
timestamp 1604666999
transform 1 0 18952 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_209
timestamp 1604666999
transform 1 0 20332 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_205
timestamp 1604666999
transform 1 0 19964 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_206
timestamp 1604666999
transform 1 0 20056 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604666999
transform 1 0 20148 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604666999
transform 1 0 19596 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_213
timestamp 1604666999
transform 1 0 20700 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_215
timestamp 1604666999
transform 1 0 20884 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 20792 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1604666999
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604666999
transform 1 0 20976 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
timestamp 1604666999
transform 1 0 21068 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_27_233
timestamp 1604666999
transform 1 0 22540 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_229
timestamp 1604666999
transform 1 0 22172 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1604666999
transform 1 0 21804 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 22356 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 21988 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604666999
transform 1 0 23000 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 23368 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_236
timestamp 1604666999
transform 1 0 22816 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_240
timestamp 1604666999
transform 1 0 23184 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_237
timestamp 1604666999
transform 1 0 22908 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_240
timestamp 1604666999
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1604666999
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604666999
transform 1 0 23644 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 23552 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 25576 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 25392 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 25576 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 24840 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_263
timestamp 1604666999
transform 1 0 25300 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_268
timestamp 1604666999
transform 1 0 25760 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_254
timestamp 1604666999
transform 1 0 24472 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_260
timestamp 1604666999
transform 1 0 25024 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_285
timestamp 1604666999
transform 1 0 27324 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_274
timestamp 1604666999
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1604666999
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_298
timestamp 1604666999
transform 1 0 28520 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_294
timestamp 1604666999
transform 1 0 28152 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_290
timestamp 1604666999
transform 1 0 27784 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 27600 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCD
timestamp 1604666999
transform 1 0 28336 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCE
timestamp 1604666999
transform 1 0 27968 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_295
timestamp 1604666999
transform 1 0 28244 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 26496 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_27_310
timestamp 1604666999
transform 1 0 29624 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_306
timestamp 1604666999
transform 1 0 29256 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_302
timestamp 1604666999
transform 1 0 28888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__D
timestamp 1604666999
transform 1 0 28704 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 29348 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1604666999
transform 1 0 29164 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_313
timestamp 1604666999
transform 1 0 29900 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__D
timestamp 1604666999
transform 1 0 29716 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCE
timestamp 1604666999
transform 1 0 30084 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 29532 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_
timestamp 1604666999
transform 1 0 30268 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_2  FILLER_26_332
timestamp 1604666999
transform 1 0 31648 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_328
timestamp 1604666999
transform 1 0 31280 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 31832 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 31464 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_345
timestamp 1604666999
transform 1 0 32844 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_341
timestamp 1604666999
transform 1 0 32476 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 33028 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 32660 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1604666999
transform 1 0 32016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 32108 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_358
timestamp 1604666999
transform 1 0 34040 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_356
timestamp 1604666999
transform 1 0 33856 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 34040 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 34224 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604666999
transform 1 0 33212 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_27_367
timestamp 1604666999
transform 1 0 34868 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_362
timestamp 1604666999
transform 1 0 34408 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1604666999
transform 1 0 34776 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_372
timestamp 1604666999
transform 1 0 35328 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_360
timestamp 1604666999
transform 1 0 34224 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1604666999
transform 1 0 37628 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604666999
transform 1 0 35420 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_384
timestamp 1604666999
transform 1 0 36432 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_396
timestamp 1604666999
transform 1 0 37536 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_375
timestamp 1604666999
transform 1 0 35604 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_387
timestamp 1604666999
transform 1 0 36708 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604666999
transform -1 0 38824 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604666999
transform -1 0 38824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_398
timestamp 1604666999
transform 1 0 37720 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_406
timestamp 1604666999
transform 1 0 38456 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_399
timestamp 1604666999
transform 1 0 37812 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604666999
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604666999
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604666999
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1604666999
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1604666999
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1604666999
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1604666999
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 7544 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1604666999
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_68
timestamp 1604666999
transform 1 0 7360 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_72
timestamp 1604666999
transform 1 0 7728 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1604666999
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 8372 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_78
timestamp 1604666999
transform 1 0 8280 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_81
timestamp 1604666999
transform 1 0 8556 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_89
timestamp 1604666999
transform 1 0 9292 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1604666999
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1604666999
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1604666999
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604666999
transform 1 0 14812 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1604666999
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_141
timestamp 1604666999
transform 1 0 14076 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
timestamp 1604666999
transform 1 0 16468 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1604666999
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
timestamp 1604666999
transform 1 0 15456 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
timestamp 1604666999
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1604666999
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_154
timestamp 1604666999
transform 1 0 15272 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_158
timestamp 1604666999
transform 1 0 15640 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_162
timestamp 1604666999
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_165
timestamp 1604666999
transform 1 0 16284 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604666999
transform 1 0 18952 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 18400 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 18768 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_186
timestamp 1604666999
transform 1 0 18216 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_190
timestamp 1604666999
transform 1 0 18584 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_198
timestamp 1604666999
transform 1 0 19320 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604666999
transform 1 0 21252 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1604666999
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 19504 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 21068 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 19872 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_202
timestamp 1604666999
transform 1 0 19688 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_206
timestamp 1604666999
transform 1 0 20056 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_215
timestamp 1604666999
transform 1 0 20884 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604666999
transform 1 0 22816 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 23644 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_228
timestamp 1604666999
transform 1 0 22080 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_240
timestamp 1604666999
transform 1 0 23184 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_244
timestamp 1604666999
transform 1 0 23552 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_247
timestamp 1604666999
transform 1 0 23828 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604666999
transform 1 0 24288 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 24104 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_261
timestamp 1604666999
transform 1 0 25116 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_273
timestamp 1604666999
transform 1 0 26220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _54_
timestamp 1604666999
transform 1 0 26588 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_
timestamp 1604666999
transform 1 0 27968 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1604666999
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604666999
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_280
timestamp 1604666999
transform 1 0 26864 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCD
timestamp 1604666999
transform 1 0 30360 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 30728 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_316
timestamp 1604666999
transform 1 0 30176 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_320
timestamp 1604666999
transform 1 0 30544 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _52_
timestamp 1604666999
transform 1 0 30912 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 32108 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1604666999
transform 1 0 32016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_327
timestamp 1604666999
transform 1 0 31188 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_335
timestamp 1604666999
transform 1 0 31924 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_356
timestamp 1604666999
transform 1 0 33856 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_368
timestamp 1604666999
transform 1 0 34960 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_372
timestamp 1604666999
transform 1 0 35328 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604666999
transform 1 0 35420 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1604666999
transform 1 0 37628 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1604666999
transform 1 0 35788 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_389
timestamp 1604666999
transform 1 0 36892 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604666999
transform -1 0 38824 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_398
timestamp 1604666999
transform 1 0 37720 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_406
timestamp 1604666999
transform 1 0 38456 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604666999
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604666999
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604666999
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1604666999
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1604666999
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 7544 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1604666999
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 7360 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1604666999
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1604666999
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_62
timestamp 1604666999
transform 1 0 6808 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9660 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_89
timestamp 1604666999
transform 1 0 9292 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_95
timestamp 1604666999
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_99
timestamp 1604666999
transform 1 0 10212 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1604666999
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_111
timestamp 1604666999
transform 1 0 11316 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_119
timestamp 1604666999
transform 1 0 12052 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1604666999
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604666999
transform 1 0 14812 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604666999
transform 1 0 14628 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1604666999
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604666999
transform 1 0 16376 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
timestamp 1604666999
transform 1 0 16100 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_158
timestamp 1604666999
transform 1 0 15640 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_162
timestamp 1604666999
transform 1 0 16008 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_165
timestamp 1604666999
transform 1 0 16284 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
timestamp 1604666999
transform 1 0 18032 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1604666999
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
timestamp 1604666999
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
timestamp 1604666999
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_175
timestamp 1604666999
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_179
timestamp 1604666999
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604666999
transform 1 0 21344 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604666999
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604666999
transform 1 0 20516 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 19964 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_203
timestamp 1604666999
transform 1 0 19780 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_207
timestamp 1604666999
transform 1 0 20148 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_213
timestamp 1604666999
transform 1 0 20700 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_217
timestamp 1604666999
transform 1 0 21068 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1604666999
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 22356 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604666999
transform 1 0 22724 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_229
timestamp 1604666999
transform 1 0 22172 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_233
timestamp 1604666999
transform 1 0 22540 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_237
timestamp 1604666999
transform 1 0 22908 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_243
timestamp 1604666999
transform 1 0 23460 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_245
timestamp 1604666999
transform 1 0 23644 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 26128 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 24288 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_251
timestamp 1604666999
transform 1 0 24196 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_254
timestamp 1604666999
transform 1 0 24472 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_266
timestamp 1604666999
transform 1 0 25576 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 26680 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 26496 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_274
timestamp 1604666999
transform 1 0 26312 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_287
timestamp 1604666999
transform 1 0 27508 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 30544 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1604666999
transform 1 0 29164 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 30360 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 29992 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_299
timestamp 1604666999
transform 1 0 28612 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_306
timestamp 1604666999
transform 1 0 29256 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_316
timestamp 1604666999
transform 1 0 30176 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604666999
transform 1 0 32108 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 31924 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 31556 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_329
timestamp 1604666999
transform 1 0 31372 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_333
timestamp 1604666999
transform 1 0 31740 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_346
timestamp 1604666999
transform 1 0 32936 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1604666999
transform 1 0 34776 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_358
timestamp 1604666999
transform 1 0 34040 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_367
timestamp 1604666999
transform 1 0 34868 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_379
timestamp 1604666999
transform 1 0 35972 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_391
timestamp 1604666999
transform 1 0 37076 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604666999
transform -1 0 38824 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_403
timestamp 1604666999
transform 1 0 38180 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604666999
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604666999
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604666999
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1604666999
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1604666999
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1604666999
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1604666999
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1604666999
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1604666999
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 9660 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1604666999
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1604666999
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_112
timestamp 1604666999
transform 1 0 11408 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_124
timestamp 1604666999
transform 1 0 12512 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604666999
transform 1 0 14812 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_136
timestamp 1604666999
transform 1 0 13616 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_148
timestamp 1604666999
transform 1 0 14720 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
timestamp 1604666999
transform 1 0 16100 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1604666999
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 15916 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 15548 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_151
timestamp 1604666999
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_154
timestamp 1604666999
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_159
timestamp 1604666999
transform 1 0 15732 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604666999
transform 1 0 19228 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
timestamp 1604666999
transform 1 0 18308 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
timestamp 1604666999
transform 1 0 18676 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_182
timestamp 1604666999
transform 1 0 17848 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_186
timestamp 1604666999
transform 1 0 18216 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_189
timestamp 1604666999
transform 1 0 18492 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_193
timestamp 1604666999
transform 1 0 18860 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604666999
transform 1 0 20884 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1604666999
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 21528 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 20516 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_206
timestamp 1604666999
transform 1 0 20056 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_210
timestamp 1604666999
transform 1 0 20424 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_213
timestamp 1604666999
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_220
timestamp 1604666999
transform 1 0 21344 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604666999
transform 1 0 22080 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 21896 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 23736 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_224
timestamp 1604666999
transform 1 0 21712 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_232
timestamp 1604666999
transform 1 0 22448 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_244
timestamp 1604666999
transform 1 0 23552 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_248
timestamp 1604666999
transform 1 0 23920 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 25024 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_262
timestamp 1604666999
transform 1 0 25208 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1604666999
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 26680 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 27048 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 27416 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_274
timestamp 1604666999
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_276
timestamp 1604666999
transform 1 0 26496 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_280
timestamp 1604666999
transform 1 0 26864 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_284
timestamp 1604666999
transform 1 0 27232 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_288
timestamp 1604666999
transform 1 0 27600 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 30544 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_300
timestamp 1604666999
transform 1 0 28704 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_312
timestamp 1604666999
transform 1 0 29808 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_322
timestamp 1604666999
transform 1 0 30728 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _53_
timestamp 1604666999
transform 1 0 32108 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1604666999
transform 1 0 32016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 32568 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_334
timestamp 1604666999
transform 1 0 31832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_340
timestamp 1604666999
transform 1 0 32384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_344
timestamp 1604666999
transform 1 0 32752 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1604666999
transform 1 0 35236 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 35052 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 33212 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 33580 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_348
timestamp 1604666999
transform 1 0 33120 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_351
timestamp 1604666999
transform 1 0 33396 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_355
timestamp 1604666999
transform 1 0 33764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_367
timestamp 1604666999
transform 1 0 34868 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1604666999
transform 1 0 37628 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 35696 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_374
timestamp 1604666999
transform 1 0 35512 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_378
timestamp 1604666999
transform 1 0 35880 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_390
timestamp 1604666999
transform 1 0 36984 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_396
timestamp 1604666999
transform 1 0 37536 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604666999
transform -1 0 38824 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_398
timestamp 1604666999
transform 1 0 37720 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_406
timestamp 1604666999
transform 1 0 38456 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604666999
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604666999
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604666999
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1604666999
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1604666999
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1604666999
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1604666999
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604666999
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1604666999
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1604666999
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1604666999
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1604666999
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1604666999
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1604666999
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1604666999
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1604666999
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1604666999
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604666999
transform 1 0 16376 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604666999
transform 1 0 16192 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604666999
transform 1 0 15824 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_159
timestamp 1604666999
transform 1 0 15732 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_162
timestamp 1604666999
transform 1 0 16008 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
timestamp 1604666999
transform 1 0 18032 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1604666999
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
timestamp 1604666999
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_175
timestamp 1604666999
transform 1 0 17204 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604666999
transform 1 0 20516 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 21528 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 20332 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 19964 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_203
timestamp 1604666999
transform 1 0 19780 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_207
timestamp 1604666999
transform 1 0 20148 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_220
timestamp 1604666999
transform 1 0 21344 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_228
timestamp 1604666999
transform 1 0 22080 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_224
timestamp 1604666999
transform 1 0 21712 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 21896 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_233
timestamp 1604666999
transform 1 0 22540 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604666999
transform 1 0 22172 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_237
timestamp 1604666999
transform 1 0 22908 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604666999
transform 1 0 22724 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_241
timestamp 1604666999
transform 1 0 23276 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604666999
transform 1 0 23092 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_245
timestamp 1604666999
transform 1 0 23644 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 23828 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1604666999
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604666999
transform 1 0 25024 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 24840 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 26128 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 24196 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_249
timestamp 1604666999
transform 1 0 24012 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_253
timestamp 1604666999
transform 1 0 24380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_257
timestamp 1604666999
transform 1 0 24748 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_269
timestamp 1604666999
transform 1 0 25852 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 26680 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 27692 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 26496 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 28060 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_274
timestamp 1604666999
transform 1 0 26312 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_287
timestamp 1604666999
transform 1 0 27508 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_291
timestamp 1604666999
transform 1 0 27876 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_295
timestamp 1604666999
transform 1 0 28244 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1604666999
transform 1 0 29164 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_303
timestamp 1604666999
transform 1 0 28980 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_306
timestamp 1604666999
transform 1 0 29256 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_318
timestamp 1604666999
transform 1 0 30360 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 32292 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 33028 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 32660 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 31832 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_330
timestamp 1604666999
transform 1 0 31464 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_336
timestamp 1604666999
transform 1 0 32016 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_341
timestamp 1604666999
transform 1 0 32476 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_345
timestamp 1604666999
transform 1 0 32844 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604666999
transform 1 0 33212 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604666999
transform 1 0 35052 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1604666999
transform 1 0 34776 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 34592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 34224 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_358
timestamp 1604666999
transform 1 0 34040 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_362
timestamp 1604666999
transform 1 0 34408 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_367
timestamp 1604666999
transform 1 0 34868 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 36064 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_378
timestamp 1604666999
transform 1 0 35880 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_382
timestamp 1604666999
transform 1 0 36248 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_394
timestamp 1604666999
transform 1 0 37352 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604666999
transform -1 0 38824 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_406
timestamp 1604666999
transform 1 0 38456 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604666999
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604666999
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604666999
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1604666999
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1604666999
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604666999
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1604666999
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1604666999
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1604666999
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1604666999
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1604666999
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1604666999
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1604666999
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1604666999
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1604666999
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1604666999
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1604666999
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604666999
transform 1 0 16376 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 16744 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1604666999
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_168
timestamp 1604666999
transform 1 0 16560 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_172
timestamp 1604666999
transform 1 0 16928 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
timestamp 1604666999
transform 1 0 18308 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
timestamp 1604666999
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_186
timestamp 1604666999
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 20884 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1604666999
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 20516 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_206
timestamp 1604666999
transform 1 0 20056 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_210
timestamp 1604666999
transform 1 0 20424 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1604666999
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604666999
transform 1 0 22448 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 23736 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 23368 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_224
timestamp 1604666999
transform 1 0 21712 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_236
timestamp 1604666999
transform 1 0 22816 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_244
timestamp 1604666999
transform 1 0 23552 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _57_
timestamp 1604666999
transform 1 0 25392 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__D
timestamp 1604666999
transform 1 0 26220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 25024 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_255
timestamp 1604666999
transform 1 0 24564 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_259
timestamp 1604666999
transform 1 0 24932 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_262
timestamp 1604666999
transform 1 0 25208 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_267
timestamp 1604666999
transform 1 0 25668 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 27048 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1604666999
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCD
timestamp 1604666999
transform 1 0 26680 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_276
timestamp 1604666999
transform 1 0 26496 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_280
timestamp 1604666999
transform 1 0 26864 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1604666999
transform 1 0 29900 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 30360 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 30728 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 29348 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 29716 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1604666999
transform 1 0 28796 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1604666999
transform 1 0 29532 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_316
timestamp 1604666999
transform 1 0 30176 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_320
timestamp 1604666999
transform 1 0 30544 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 32292 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1604666999
transform 1 0 32016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__D
timestamp 1604666999
transform 1 0 31832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 31464 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_324
timestamp 1604666999
transform 1 0 30912 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_332
timestamp 1604666999
transform 1 0 31648 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_337
timestamp 1604666999
transform 1 0 32108 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 34776 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_32_358
timestamp 1604666999
transform 1 0 34040 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1604666999
transform 1 0 37628 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_385
timestamp 1604666999
transform 1 0 36524 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604666999
transform -1 0 38824 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_398
timestamp 1604666999
transform 1 0 37720 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_406
timestamp 1604666999
transform 1 0 38456 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604666999
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604666999
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604666999
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604666999
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604666999
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604666999
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1604666999
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1604666999
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1604666999
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604666999
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604666999
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604666999
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1604666999
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1604666999
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1604666999
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1604666999
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1604666999
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604666999
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1604666999
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1604666999
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_86
timestamp 1604666999
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_98
timestamp 1604666999
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1604666999
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604666999
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1604666999
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_110
timestamp 1604666999
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1604666999
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604666999
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1604666999
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_135
timestamp 1604666999
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_147
timestamp 1604666999
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1604666999
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1604666999
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1604666999
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_159
timestamp 1604666999
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_171
timestamp 1604666999
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604666999
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1604666999
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1604666999
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604666999
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_196
timestamp 1604666999
transform 1 0 19136 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1604666999
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1604666999
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 19964 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 20884 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1604666999
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 19780 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 19964 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_202
timestamp 1604666999
transform 1 0 19688 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_202
timestamp 1604666999
transform 1 0 19688 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_207
timestamp 1604666999
transform 1 0 20148 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_213
timestamp 1604666999
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_234
timestamp 1604666999
transform 1 0 22632 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_228
timestamp 1604666999
transform 1 0 22080 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_224
timestamp 1604666999
transform 1 0 21712 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 22264 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 21896 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604666999
transform 1 0 22448 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_240
timestamp 1604666999
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_236
timestamp 1604666999
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604666999
transform 1 0 23000 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1604666999
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604666999
transform 1 0 23644 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 23368 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_33_257
timestamp 1604666999
transform 1 0 24748 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_253
timestamp 1604666999
transform 1 0 24380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_249
timestamp 1604666999
transform 1 0 24012 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604666999
transform 1 0 24196 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 24840 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_269
timestamp 1604666999
transform 1 0 25852 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_265
timestamp 1604666999
transform 1 0 25484 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_261
timestamp 1604666999
transform 1 0 25116 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 26220 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 25668 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__D
timestamp 1604666999
transform 1 0 25300 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 25024 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604666999
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_283
timestamp 1604666999
transform 1 0 27140 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_279
timestamp 1604666999
transform 1 0 26772 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 27324 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCE
timestamp 1604666999
transform 1 0 26956 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1604666999
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_296
timestamp 1604666999
transform 1 0 28336 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 28520 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 27508 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_
timestamp 1604666999
transform 1 0 26588 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 29348 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 29900 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1604666999
transform 1 0 29164 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 28980 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_300
timestamp 1604666999
transform 1 0 28704 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_306
timestamp 1604666999
transform 1 0 29256 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_301
timestamp 1604666999
transform 1 0 28796 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_322
timestamp 1604666999
transform 1 0 30728 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_332
timestamp 1604666999
transform 1 0 31648 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_326
timestamp 1604666999
transform 1 0 31096 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_330
timestamp 1604666999
transform 1 0 31464 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_326
timestamp 1604666999
transform 1 0 31096 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 31464 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__D
timestamp 1604666999
transform 1 0 30912 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCD
timestamp 1604666999
transform 1 0 31832 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 31280 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCE
timestamp 1604666999
transform 1 0 31648 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_346
timestamp 1604666999
transform 1 0 32936 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1604666999
transform 1 0 32016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 32108 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_
timestamp 1604666999
transform 1 0 31832 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_1  FILLER_34_354
timestamp 1604666999
transform 1 0 33672 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_358
timestamp 1604666999
transform 1 0 34040 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 33764 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 34224 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_367
timestamp 1604666999
transform 1 0 34868 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_362
timestamp 1604666999
transform 1 0 34408 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 34592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 35052 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1604666999
transform 1 0 34776 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 35236 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 33948 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1604666999
transform 1 0 37628 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 35880 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_390
timestamp 1604666999
transform 1 0 36984 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_376
timestamp 1604666999
transform 1 0 35696 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_380
timestamp 1604666999
transform 1 0 36064 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_392
timestamp 1604666999
transform 1 0 37168 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_396
timestamp 1604666999
transform 1 0 37536 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604666999
transform -1 0 38824 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604666999
transform -1 0 38824 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_402
timestamp 1604666999
transform 1 0 38088 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_406
timestamp 1604666999
transform 1 0 38456 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_398
timestamp 1604666999
transform 1 0 37720 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_406
timestamp 1604666999
transform 1 0 38456 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604666999
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604666999
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604666999
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1604666999
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1604666999
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1604666999
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1604666999
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1604666999
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1604666999
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_74
timestamp 1604666999
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_86
timestamp 1604666999
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_98
timestamp 1604666999
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1604666999
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_110
timestamp 1604666999
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_123
timestamp 1604666999
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_135
timestamp 1604666999
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_147
timestamp 1604666999
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_159
timestamp 1604666999
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_171
timestamp 1604666999
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1604666999
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1604666999
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1604666999
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _55_
timestamp 1604666999
transform 1 0 20332 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 21344 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 21160 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 20792 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_208
timestamp 1604666999
transform 1 0 20240 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_212
timestamp 1604666999
transform 1 0 20608 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_216
timestamp 1604666999
transform 1 0 20976 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_233
timestamp 1604666999
transform 1 0 22540 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_229
timestamp 1604666999
transform 1 0 22172 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 22356 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_237
timestamp 1604666999
transform 1 0 22908 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 22724 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_241
timestamp 1604666999
transform 1 0 23276 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1604666999
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _56_
timestamp 1604666999
transform 1 0 23644 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_248
timestamp 1604666999
transform 1 0 23920 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_
timestamp 1604666999
transform 1 0 24840 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCE
timestamp 1604666999
transform 1 0 24656 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 24288 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_254
timestamp 1604666999
transform 1 0 24472 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _58_
timestamp 1604666999
transform 1 0 27784 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 27232 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 27600 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_282
timestamp 1604666999
transform 1 0 27048 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_286
timestamp 1604666999
transform 1 0 27416 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1604666999
transform 1 0 28060 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_
timestamp 1604666999
transform 1 0 30544 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1604666999
transform 1 0 29164 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCE
timestamp 1604666999
transform 1 0 30360 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604666999
transform 1 0 29992 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_306
timestamp 1604666999
transform 1 0 29256 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_316
timestamp 1604666999
transform 1 0 30176 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 32936 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_344
timestamp 1604666999
transform 1 0 32752 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_355
timestamp 1604666999
transform 1 0 33764 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_348
timestamp 1604666999
transform 1 0 33120 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 33304 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 33948 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604666999
transform 1 0 33488 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_363
timestamp 1604666999
transform 1 0 34500 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_359
timestamp 1604666999
transform 1 0 34132 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCE
timestamp 1604666999
transform 1 0 34316 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1604666999
transform 1 0 34776 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 34868 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__D
timestamp 1604666999
transform 1 0 35880 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 36248 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 36616 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_376
timestamp 1604666999
transform 1 0 35696 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_380
timestamp 1604666999
transform 1 0 36064 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_384
timestamp 1604666999
transform 1 0 36432 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_388
timestamp 1604666999
transform 1 0 36800 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604666999
transform -1 0 38824 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_400
timestamp 1604666999
transform 1 0 37904 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_406
timestamp 1604666999
transform 1 0 38456 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604666999
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1604666999
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1604666999
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1604666999
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1604666999
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1604666999
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1604666999
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1604666999
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1604666999
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1604666999
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_80
timestamp 1604666999
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_93
timestamp 1604666999
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_105
timestamp 1604666999
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_117
timestamp 1604666999
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_129
timestamp 1604666999
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1604666999
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1604666999
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_154
timestamp 1604666999
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_166
timestamp 1604666999
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_178
timestamp 1604666999
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_190
timestamp 1604666999
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1604666999
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 21344 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_202
timestamp 1604666999
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_215
timestamp 1604666999
transform 1 0 20884 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_219
timestamp 1604666999
transform 1 0 21252 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_222
timestamp 1604666999
transform 1 0 21528 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 21804 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 23920 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_244
timestamp 1604666999
transform 1 0 23552 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 24288 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCD
timestamp 1604666999
transform 1 0 25300 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 25668 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 26036 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1604666999
transform 1 0 24104 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_261
timestamp 1604666999
transform 1 0 25116 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_265
timestamp 1604666999
transform 1 0 25484 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_269
timestamp 1604666999
transform 1 0 25852 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_273
timestamp 1604666999
transform 1 0 26220 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 26496 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1604666999
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 28520 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_295
timestamp 1604666999
transform 1 0 28244 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_300
timestamp 1604666999
transform 1 0 28704 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 28888 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_304
timestamp 1604666999
transform 1 0 29072 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCD
timestamp 1604666999
transform 1 0 29256 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_312
timestamp 1604666999
transform 1 0 29808 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_308
timestamp 1604666999
transform 1 0 29440 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__D
timestamp 1604666999
transform 1 0 29624 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604666999
transform 1 0 29992 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_322
timestamp 1604666999
transform 1 0 30728 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_318
timestamp 1604666999
transform 1 0 30360 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCD
timestamp 1604666999
transform 1 0 30544 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 32108 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1604666999
transform 1 0 32016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 31832 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 30912 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_326
timestamp 1604666999
transform 1 0 31096 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_346
timestamp 1604666999
transform 1 0 32936 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_
timestamp 1604666999
transform 1 0 34316 0 -1 22304
box -38 -48 2246 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCD
timestamp 1604666999
transform 1 0 34132 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_358
timestamp 1604666999
transform 1 0 34040 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1604666999
transform 1 0 37628 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 36708 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_385
timestamp 1604666999
transform 1 0 36524 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_389
timestamp 1604666999
transform 1 0 36892 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604666999
transform -1 0 38824 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_398
timestamp 1604666999
transform 1 0 37720 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_406
timestamp 1604666999
transform 1 0 38456 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604666999
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1604666999
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1604666999
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1604666999
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1604666999
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1604666999
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_51
timestamp 1604666999
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1604666999
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1604666999
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_74
timestamp 1604666999
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_86
timestamp 1604666999
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_98
timestamp 1604666999
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1604666999
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_110
timestamp 1604666999
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_123
timestamp 1604666999
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_135
timestamp 1604666999
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_147
timestamp 1604666999
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_159
timestamp 1604666999
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_171
timestamp 1604666999
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1604666999
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1604666999
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_196
timestamp 1604666999
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_208
timestamp 1604666999
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_220
timestamp 1604666999
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 23920 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1604666999
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_232
timestamp 1604666999
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_245
timestamp 1604666999
transform 1 0 23644 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 26220 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 25852 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_267
timestamp 1604666999
transform 1 0 25668 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_271
timestamp 1604666999
transform 1 0 26036 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604666999
transform 1 0 26404 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 28520 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 28152 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_284
timestamp 1604666999
transform 1 0 27232 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_292
timestamp 1604666999
transform 1 0 27968 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_296
timestamp 1604666999
transform 1 0 28336 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_
timestamp 1604666999
transform 1 0 29256 0 1 22304
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1604666999
transform 1 0 29164 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCE
timestamp 1604666999
transform 1 0 28980 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_300
timestamp 1604666999
transform 1 0 28704 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 32936 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_330
timestamp 1604666999
transform 1 0 31464 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_342
timestamp 1604666999
transform 1 0 32568 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_356
timestamp 1604666999
transform 1 0 33856 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_352
timestamp 1604666999
transform 1 0 33488 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_348
timestamp 1604666999
transform 1 0 33120 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 33672 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 33304 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_367
timestamp 1604666999
transform 1 0 34868 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_362
timestamp 1604666999
transform 1 0 34408 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 34224 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 34592 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1604666999
transform 1 0 34776 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604666999
transform 1 0 34960 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604666999
transform 1 0 36524 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 36340 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 35972 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_377
timestamp 1604666999
transform 1 0 35788 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_381
timestamp 1604666999
transform 1 0 36156 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_394
timestamp 1604666999
transform 1 0 37352 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604666999
transform -1 0 38824 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_406
timestamp 1604666999
transform 1 0 38456 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604666999
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1604666999
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1604666999
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1604666999
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1604666999
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1604666999
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1604666999
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1604666999
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1604666999
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1604666999
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_80
timestamp 1604666999
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_93
timestamp 1604666999
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_105
timestamp 1604666999
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_117
timestamp 1604666999
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_129
timestamp 1604666999
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1604666999
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1604666999
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_154
timestamp 1604666999
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_166
timestamp 1604666999
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_178
timestamp 1604666999
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_190
timestamp 1604666999
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1604666999
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_202
timestamp 1604666999
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_215
timestamp 1604666999
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 23920 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_227
timestamp 1604666999
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_239
timestamp 1604666999
transform 1 0 23092 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_247
timestamp 1604666999
transform 1 0 23828 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_250
timestamp 1604666999
transform 1 0 24104 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_262
timestamp 1604666999
transform 1 0 25208 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 28520 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1604666999
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 26680 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_274
timestamp 1604666999
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_276
timestamp 1604666999
transform 1 0 26496 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_280
timestamp 1604666999
transform 1 0 26864 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_292
timestamp 1604666999
transform 1 0 27968 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _63_
timestamp 1604666999
transform 1 0 30176 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 29532 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 29900 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_307
timestamp 1604666999
transform 1 0 29348 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_311
timestamp 1604666999
transform 1 0 29716 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_315
timestamp 1604666999
transform 1 0 30084 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_319
timestamp 1604666999
transform 1 0 30452 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1604666999
transform 1 0 32016 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 31004 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_327
timestamp 1604666999
transform 1 0 31188 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_335
timestamp 1604666999
transform 1 0 31924 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_337
timestamp 1604666999
transform 1 0 32108 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 34960 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 33304 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 34776 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 34408 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_349
timestamp 1604666999
transform 1 0 33212 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_359
timestamp 1604666999
transform 1 0 34132 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_364
timestamp 1604666999
transform 1 0 34592 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1604666999
transform 1 0 37628 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 36892 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_387
timestamp 1604666999
transform 1 0 36708 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_391
timestamp 1604666999
transform 1 0 37076 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604666999
transform -1 0 38824 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_398
timestamp 1604666999
transform 1 0 37720 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_406
timestamp 1604666999
transform 1 0 38456 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604666999
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604666999
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1604666999
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1604666999
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604666999
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1604666999
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1604666999
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1604666999
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1604666999
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1604666999
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1604666999
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1604666999
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1604666999
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_51
timestamp 1604666999
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1604666999
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1604666999
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_74
timestamp 1604666999
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1604666999
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1604666999
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1604666999
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_86
timestamp 1604666999
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_98
timestamp 1604666999
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1604666999
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_93
timestamp 1604666999
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1604666999
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_110
timestamp 1604666999
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1604666999
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_105
timestamp 1604666999
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_117
timestamp 1604666999
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_135
timestamp 1604666999
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_147
timestamp 1604666999
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_129
timestamp 1604666999
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1604666999
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1604666999
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_159
timestamp 1604666999
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_171
timestamp 1604666999
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_154
timestamp 1604666999
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_166
timestamp 1604666999
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1604666999
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_184
timestamp 1604666999
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_196
timestamp 1604666999
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_178
timestamp 1604666999
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_190
timestamp 1604666999
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1604666999
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_208
timestamp 1604666999
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_220
timestamp 1604666999
transform 1 0 21344 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_202
timestamp 1604666999
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1604666999
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1604666999
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 23920 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_232
timestamp 1604666999
transform 1 0 22448 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_245
timestamp 1604666999
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_227
timestamp 1604666999
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_239
timestamp 1604666999
transform 1 0 23092 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_247
timestamp 1604666999
transform 1 0 23828 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_250
timestamp 1604666999
transform 1 0 24104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_257
timestamp 1604666999
transform 1 0 24748 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_253
timestamp 1604666999
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 24564 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 24380 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604666999
transform 1 0 24564 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_40_272
timestamp 1604666999
transform 1 0 26128 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_264
timestamp 1604666999
transform 1 0 25392 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_261
timestamp 1604666999
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 25300 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_265
timestamp 1604666999
transform 1 0 25484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _62_
timestamp 1604666999
transform 1 0 28152 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 28152 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1604666999
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 27968 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_277
timestamp 1604666999
transform 1 0 26588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_289
timestamp 1604666999
transform 1 0 27692 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_297
timestamp 1604666999
transform 1 0 28428 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_276
timestamp 1604666999
transform 1 0 26496 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_288
timestamp 1604666999
transform 1 0 27600 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_301
timestamp 1604666999
transform 1 0 28796 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 28980 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 28612 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1604666999
transform 1 0 29164 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 29256 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_317
timestamp 1604666999
transform 1 0 30268 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_313
timestamp 1604666999
transform 1 0 29900 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_315
timestamp 1604666999
transform 1 0 30084 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 30084 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_321
timestamp 1604666999
transform 1 0 30636 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 30452 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604666999
transform 1 0 30452 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604666999
transform 1 0 30636 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 31004 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1604666999
transform 1 0 32016 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 30820 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 31740 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_344
timestamp 1604666999
transform 1 0 32752 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_325
timestamp 1604666999
transform 1 0 31004 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_335
timestamp 1604666999
transform 1 0 31924 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_337
timestamp 1604666999
transform 1 0 32108 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_349
timestamp 1604666999
transform 1 0 33212 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_358
timestamp 1604666999
transform 1 0 34040 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_352
timestamp 1604666999
transform 1 0 33488 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 34224 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _60_
timestamp 1604666999
transform 1 0 33764 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_367
timestamp 1604666999
transform 1 0 34868 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_362
timestamp 1604666999
transform 1 0 34408 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 34592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 35236 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1604666999
transform 1 0 34776 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 33948 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__conb_1  _61_
timestamp 1604666999
transform 1 0 36432 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 35420 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1604666999
transform 1 0 37628 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 35880 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_392
timestamp 1604666999
transform 1 0 37168 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_376
timestamp 1604666999
transform 1 0 35696 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_380
timestamp 1604666999
transform 1 0 36064 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_387
timestamp 1604666999
transform 1 0 36708 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_395
timestamp 1604666999
transform 1 0 37444 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604666999
transform -1 0 38824 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604666999
transform -1 0 38824 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_404
timestamp 1604666999
transform 1 0 38272 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_398
timestamp 1604666999
transform 1 0 37720 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_406
timestamp 1604666999
transform 1 0 38456 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604666999
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1604666999
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1604666999
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1604666999
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1604666999
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1604666999
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_51
timestamp 1604666999
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_59
timestamp 1604666999
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1604666999
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_74
timestamp 1604666999
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_86
timestamp 1604666999
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_98
timestamp 1604666999
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1604666999
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_110
timestamp 1604666999
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1604666999
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_135
timestamp 1604666999
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_147
timestamp 1604666999
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_159
timestamp 1604666999
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_171
timestamp 1604666999
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1604666999
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1604666999
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1604666999
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1604666999
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_220
timestamp 1604666999
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1604666999
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 23920 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_232
timestamp 1604666999
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_245
timestamp 1604666999
transform 1 0 23644 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 24472 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 24288 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_250
timestamp 1604666999
transform 1 0 24104 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_273
timestamp 1604666999
transform 1 0 26220 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604666999
transform 1 0 28060 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 26496 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 26864 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604666999
transform 1 0 27876 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1604666999
transform 1 0 26680 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_282
timestamp 1604666999
transform 1 0 27048 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_290
timestamp 1604666999
transform 1 0 27784 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_297
timestamp 1604666999
transform 1 0 28428 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 29256 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1604666999
transform 1 0 29164 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 28980 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 28612 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_301
timestamp 1604666999
transform 1 0 28796 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 31740 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604666999
transform 1 0 31188 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 31556 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_325
timestamp 1604666999
transform 1 0 31004 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_329
timestamp 1604666999
transform 1 0 31372 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_342
timestamp 1604666999
transform 1 0 32568 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_350
timestamp 1604666999
transform 1 0 33304 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 33488 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 33120 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604666999
transform 1 0 33672 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_362
timestamp 1604666999
transform 1 0 34408 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_358
timestamp 1604666999
transform 1 0 34040 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604666999
transform 1 0 34224 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 34592 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1604666999
transform 1 0 34776 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 34868 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 35880 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_376
timestamp 1604666999
transform 1 0 35696 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_380
timestamp 1604666999
transform 1 0 36064 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_392
timestamp 1604666999
transform 1 0 37168 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604666999
transform -1 0 38824 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_404
timestamp 1604666999
transform 1 0 38272 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604666999
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604666999
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1604666999
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1604666999
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604666999
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1604666999
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1604666999
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_56
timestamp 1604666999
transform 1 0 6256 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_68
timestamp 1604666999
transform 1 0 7360 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1604666999
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_80
timestamp 1604666999
transform 1 0 8464 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_93
timestamp 1604666999
transform 1 0 9660 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_105
timestamp 1604666999
transform 1 0 10764 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_117
timestamp 1604666999
transform 1 0 11868 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_129
timestamp 1604666999
transform 1 0 12972 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1604666999
transform 1 0 14076 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1604666999
transform 1 0 15180 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_154
timestamp 1604666999
transform 1 0 15272 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_166
timestamp 1604666999
transform 1 0 16376 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_178
timestamp 1604666999
transform 1 0 17480 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_190
timestamp 1604666999
transform 1 0 18584 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1604666999
transform 1 0 20792 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_202
timestamp 1604666999
transform 1 0 19688 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_215
timestamp 1604666999
transform 1 0 20884 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 23920 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 23736 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_227
timestamp 1604666999
transform 1 0 21988 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_239
timestamp 1604666999
transform 1 0 23092 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_245
timestamp 1604666999
transform 1 0 23644 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 26220 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 25852 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_267
timestamp 1604666999
transform 1 0 25668 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_271
timestamp 1604666999
transform 1 0 26036 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 26496 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1604666999
transform 1 0 26404 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604666999
transform 1 0 28428 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_295
timestamp 1604666999
transform 1 0 28244 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 29348 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 29164 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 30360 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 28796 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 30728 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_299
timestamp 1604666999
transform 1 0 28612 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_303
timestamp 1604666999
transform 1 0 28980 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_316
timestamp 1604666999
transform 1 0 30176 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_320
timestamp 1604666999
transform 1 0 30544 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604666999
transform 1 0 30912 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_332
timestamp 1604666999
transform 1 0 31648 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_328
timestamp 1604666999
transform 1 0 31280 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_335
timestamp 1604666999
transform 1 0 31924 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 31740 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1604666999
transform 1 0 32016 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _59_
timestamp 1604666999
transform 1 0 32108 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_340
timestamp 1604666999
transform 1 0 32384 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_347
timestamp 1604666999
transform 1 0 33028 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_344
timestamp 1604666999
transform 1 0 32752 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 32844 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 33120 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 35052 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_367
timestamp 1604666999
transform 1 0 34868 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_371
timestamp 1604666999
transform 1 0 35236 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1604666999
transform 1 0 37628 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_383
timestamp 1604666999
transform 1 0 36340 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_395
timestamp 1604666999
transform 1 0 37444 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604666999
transform -1 0 38824 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_398
timestamp 1604666999
transform 1 0 37720 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_406
timestamp 1604666999
transform 1 0 38456 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1604666999
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1604666999
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1604666999
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1604666999
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1604666999
transform 1 0 4692 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1604666999
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_51
timestamp 1604666999
transform 1 0 5796 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_59
timestamp 1604666999
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_62
timestamp 1604666999
transform 1 0 6808 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_74
timestamp 1604666999
transform 1 0 7912 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_86
timestamp 1604666999
transform 1 0 9016 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_98
timestamp 1604666999
transform 1 0 10120 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1604666999
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_110
timestamp 1604666999
transform 1 0 11224 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_123
timestamp 1604666999
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_135
timestamp 1604666999
transform 1 0 13524 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_147
timestamp 1604666999
transform 1 0 14628 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_159
timestamp 1604666999
transform 1 0 15732 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_171
timestamp 1604666999
transform 1 0 16836 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1604666999
transform 1 0 17940 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_184
timestamp 1604666999
transform 1 0 18032 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_196
timestamp 1604666999
transform 1 0 19136 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_208
timestamp 1604666999
transform 1 0 20240 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_220
timestamp 1604666999
transform 1 0 21344 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1604666999
transform 1 0 23552 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604666999
transform 1 0 23828 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 23368 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604666999
transform 1 0 23000 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_232
timestamp 1604666999
transform 1 0 22448 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_240
timestamp 1604666999
transform 1 0 23184 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_245
timestamp 1604666999
transform 1 0 23644 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 24012 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 25944 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_268
timestamp 1604666999
transform 1 0 25760 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_272
timestamp 1604666999
transform 1 0 26128 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604666999
transform 1 0 26496 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604666999
transform 1 0 28060 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 26312 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 27876 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 27508 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_285
timestamp 1604666999
transform 1 0 27324 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_289
timestamp 1604666999
transform 1 0 27692 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_297
timestamp 1604666999
transform 1 0 28428 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 29900 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1604666999
transform 1 0 29164 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 29716 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 28612 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 28980 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_301
timestamp 1604666999
transform 1 0 28796 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_306
timestamp 1604666999
transform 1 0 29256 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_310
timestamp 1604666999
transform 1 0 29624 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 32844 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 32660 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 32292 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 31924 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_332
timestamp 1604666999
transform 1 0 31648 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_337
timestamp 1604666999
transform 1 0 32108 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_341
timestamp 1604666999
transform 1 0 32476 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604666999
transform 1 0 34868 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1604666999
transform 1 0 34776 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604666999
transform 1 0 34592 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 33856 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_354
timestamp 1604666999
transform 1 0 33672 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_358
timestamp 1604666999
transform 1 0 34040 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_371
timestamp 1604666999
transform 1 0 35236 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604666999
transform 1 0 35972 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604666999
transform 1 0 35420 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604666999
transform 1 0 35788 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604666999
transform 1 0 36524 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_375
timestamp 1604666999
transform 1 0 35604 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_383
timestamp 1604666999
transform 1 0 36340 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_387
timestamp 1604666999
transform 1 0 36708 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1604666999
transform -1 0 38824 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_399
timestamp 1604666999
transform 1 0 37812 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1604666999
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1604666999
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1604666999
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1604666999
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_27
timestamp 1604666999
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_32
timestamp 1604666999
transform 1 0 4048 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_44
timestamp 1604666999
transform 1 0 5152 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_56
timestamp 1604666999
transform 1 0 6256 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_68
timestamp 1604666999
transform 1 0 7360 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1604666999
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_80
timestamp 1604666999
transform 1 0 8464 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_93
timestamp 1604666999
transform 1 0 9660 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_105
timestamp 1604666999
transform 1 0 10764 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_117
timestamp 1604666999
transform 1 0 11868 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_129
timestamp 1604666999
transform 1 0 12972 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1604666999
transform 1 0 14076 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1604666999
transform 1 0 15180 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_154
timestamp 1604666999
transform 1 0 15272 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_166
timestamp 1604666999
transform 1 0 16376 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_178
timestamp 1604666999
transform 1 0 17480 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_190
timestamp 1604666999
transform 1 0 18584 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1604666999
transform 1 0 20792 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_202
timestamp 1604666999
transform 1 0 19688 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_215
timestamp 1604666999
transform 1 0 20884 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604666999
transform 1 0 23552 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 23368 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_227
timestamp 1604666999
transform 1 0 21988 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_239
timestamp 1604666999
transform 1 0 23092 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 26220 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 25852 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_263
timestamp 1604666999
transform 1 0 25300 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_271
timestamp 1604666999
transform 1 0 26036 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604666999
transform 1 0 26496 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604666999
transform 1 0 28060 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1604666999
transform 1 0 26404 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 27508 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_285
timestamp 1604666999
transform 1 0 27324 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_289
timestamp 1604666999
transform 1 0 27692 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604666999
transform 1 0 29624 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604666999
transform 1 0 30636 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604666999
transform 1 0 29072 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 29440 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_302
timestamp 1604666999
transform 1 0 28888 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1604666999
transform 1 0 29256 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_319
timestamp 1604666999
transform 1 0 30452 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 32936 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1604666999
transform 1 0 32016 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 32752 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 32384 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604666999
transform 1 0 31832 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_323
timestamp 1604666999
transform 1 0 30820 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_331
timestamp 1604666999
transform 1 0 31556 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_337
timestamp 1604666999
transform 1 0 32108 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_342
timestamp 1604666999
transform 1 0 32568 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
timestamp 1604666999
transform 1 0 35144 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_365
timestamp 1604666999
transform 1 0 34684 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_369
timestamp 1604666999
transform 1 0 35052 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_372
timestamp 1604666999
transform 1 0 35328 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604666999
transform 1 0 35420 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1604666999
transform 1 0 37628 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_378
timestamp 1604666999
transform 1 0 35880 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_390
timestamp 1604666999
transform 1 0 36984 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_396
timestamp 1604666999
transform 1 0 37536 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1604666999
transform -1 0 38824 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_398
timestamp 1604666999
transform 1 0 37720 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_406
timestamp 1604666999
transform 1 0 38456 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1604666999
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1604666999
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1604666999
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1604666999
transform 1 0 3588 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1604666999
transform 1 0 4692 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1604666999
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_51
timestamp 1604666999
transform 1 0 5796 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_59
timestamp 1604666999
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_62
timestamp 1604666999
transform 1 0 6808 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_74
timestamp 1604666999
transform 1 0 7912 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_86
timestamp 1604666999
transform 1 0 9016 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_98
timestamp 1604666999
transform 1 0 10120 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1604666999
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_110
timestamp 1604666999
transform 1 0 11224 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_123
timestamp 1604666999
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_135
timestamp 1604666999
transform 1 0 13524 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_147
timestamp 1604666999
transform 1 0 14628 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_159
timestamp 1604666999
transform 1 0 15732 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_171
timestamp 1604666999
transform 1 0 16836 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1604666999
transform 1 0 17940 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_184
timestamp 1604666999
transform 1 0 18032 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_196
timestamp 1604666999
transform 1 0 19136 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_208
timestamp 1604666999
transform 1 0 20240 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_220
timestamp 1604666999
transform 1 0 21344 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604666999
transform 1 0 22448 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
timestamp 1604666999
transform 1 0 23644 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1604666999
transform 1 0 23552 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
timestamp 1604666999
transform 1 0 23368 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
timestamp 1604666999
transform 1 0 23000 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604666999
transform 1 0 22264 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_228
timestamp 1604666999
transform 1 0 22080 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_236
timestamp 1604666999
transform 1 0 22816 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_240
timestamp 1604666999
transform 1 0 23184 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 25576 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 26220 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_264
timestamp 1604666999
transform 1 0 25392 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_268
timestamp 1604666999
transform 1 0 25760 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_272
timestamp 1604666999
transform 1 0 26128 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604666999
transform 1 0 27140 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604666999
transform 1 0 28244 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 26956 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 26588 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_275
timestamp 1604666999
transform 1 0 26404 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_279
timestamp 1604666999
transform 1 0 26772 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_292
timestamp 1604666999
transform 1 0 27968 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_297
timestamp 1604666999
transform 1 0 28428 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 29532 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1604666999
transform 1 0 29164 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 28980 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604666999
transform 1 0 28612 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_301
timestamp 1604666999
transform 1 0 28796 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_306
timestamp 1604666999
transform 1 0 29256 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604666999
transform 1 0 32108 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 33028 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 32660 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604666999
transform 1 0 31924 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604666999
transform 1 0 31464 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_328
timestamp 1604666999
transform 1 0 31280 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_332
timestamp 1604666999
transform 1 0 31648 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_341
timestamp 1604666999
transform 1 0 32476 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_345
timestamp 1604666999
transform 1 0 32844 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604666999
transform 1 0 33212 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1604666999
transform 1 0 34776 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 35236 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 34592 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
timestamp 1604666999
transform 1 0 34224 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_358
timestamp 1604666999
transform 1 0 34040 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_362
timestamp 1604666999
transform 1 0 34408 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_367
timestamp 1604666999
transform 1 0 34868 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 35420 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_45_392
timestamp 1604666999
transform 1 0 37168 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1604666999
transform -1 0 38824 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_404
timestamp 1604666999
transform 1 0 38272 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1604666999
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1604666999
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1604666999
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1604666999
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1604666999
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1604666999
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1604666999
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_27
timestamp 1604666999
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_32
timestamp 1604666999
transform 1 0 4048 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_44
timestamp 1604666999
transform 1 0 5152 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1604666999
transform 1 0 3588 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1604666999
transform 1 0 4692 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1604666999
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_56
timestamp 1604666999
transform 1 0 6256 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_68
timestamp 1604666999
transform 1 0 7360 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_51
timestamp 1604666999
transform 1 0 5796 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_59
timestamp 1604666999
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_62
timestamp 1604666999
transform 1 0 6808 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_74
timestamp 1604666999
transform 1 0 7912 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1604666999
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_80
timestamp 1604666999
transform 1 0 8464 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_93
timestamp 1604666999
transform 1 0 9660 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_86
timestamp 1604666999
transform 1 0 9016 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_98
timestamp 1604666999
transform 1 0 10120 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1604666999
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_105
timestamp 1604666999
transform 1 0 10764 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_117
timestamp 1604666999
transform 1 0 11868 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_110
timestamp 1604666999
transform 1 0 11224 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_123
timestamp 1604666999
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_129
timestamp 1604666999
transform 1 0 12972 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1604666999
transform 1 0 14076 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_135
timestamp 1604666999
transform 1 0 13524 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_147
timestamp 1604666999
transform 1 0 14628 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1604666999
transform 1 0 15180 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_154
timestamp 1604666999
transform 1 0 15272 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_166
timestamp 1604666999
transform 1 0 16376 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_159
timestamp 1604666999
transform 1 0 15732 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_171
timestamp 1604666999
transform 1 0 16836 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1604666999
transform 1 0 17940 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_178
timestamp 1604666999
transform 1 0 17480 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_190
timestamp 1604666999
transform 1 0 18584 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_184
timestamp 1604666999
transform 1 0 18032 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_196
timestamp 1604666999
transform 1 0 19136 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1604666999
transform 1 0 20792 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_202
timestamp 1604666999
transform 1 0 19688 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_215
timestamp 1604666999
transform 1 0 20884 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_208
timestamp 1604666999
transform 1 0 20240 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_220
timestamp 1604666999
transform 1 0 21344 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_232
timestamp 1604666999
transform 1 0 22448 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
timestamp 1604666999
transform 1 0 22632 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
timestamp 1604666999
transform 1 0 23368 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
timestamp 1604666999
transform 1 0 23000 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 23276 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_239
timestamp 1604666999
transform 1 0 23092 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_236
timestamp 1604666999
transform 1 0 22816 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_240
timestamp 1604666999
transform 1 0 23184 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1604666999
transform 1 0 23552 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
timestamp 1604666999
transform 1 0 23644 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_243
timestamp 1604666999
transform 1 0 23460 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604666999
transform 1 0 23828 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_46_227
timestamp 1604666999
transform 1 0 21988 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
timestamp 1604666999
transform 1 0 23644 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604666999
transform 1 0 26128 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604666999
transform 1 0 25944 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 25576 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 26220 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_256
timestamp 1604666999
transform 1 0 24656 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_268
timestamp 1604666999
transform 1 0 25760 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_272
timestamp 1604666999
transform 1 0 26128 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_264
timestamp 1604666999
transform 1 0 25392 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_268
timestamp 1604666999
transform 1 0 25760 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_280
timestamp 1604666999
transform 1 0 26864 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_276
timestamp 1604666999
transform 1 0 26496 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 27048 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 26680 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1604666999
transform 1 0 26404 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604666999
transform 1 0 26496 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_284
timestamp 1604666999
transform 1 0 27232 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_290
timestamp 1604666999
transform 1 0 27784 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_285
timestamp 1604666999
transform 1 0 27324 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 27600 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 27416 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604666999
transform 1 0 27600 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_297
timestamp 1604666999
transform 1 0 28428 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_295
timestamp 1604666999
transform 1 0 28244 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604666999
transform 1 0 28060 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_306
timestamp 1604666999
transform 1 0 29256 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_301
timestamp 1604666999
transform 1 0 28796 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_299
timestamp 1604666999
transform 1 0 28612 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
timestamp 1604666999
transform 1 0 28704 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
timestamp 1604666999
transform 1 0 28612 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
timestamp 1604666999
transform 1 0 28980 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1604666999
transform 1 0 29164 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604666999
transform 1 0 28888 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_46_315
timestamp 1604666999
transform 1 0 30084 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_311
timestamp 1604666999
transform 1 0 29716 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
timestamp 1604666999
transform 1 0 30268 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 29900 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604666999
transform 1 0 30452 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
timestamp 1604666999
transform 1 0 29440 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_47_327
timestamp 1604666999
transform 1 0 31188 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 31740 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604666999
transform 1 0 31924 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_343
timestamp 1604666999
transform 1 0 32660 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_339
timestamp 1604666999
transform 1 0 32292 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_346
timestamp 1604666999
transform 1 0 32936 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_341
timestamp 1604666999
transform 1 0 32476 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 32752 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604666999
transform 1 0 32476 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
timestamp 1604666999
transform 1 0 33028 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1604666999
transform 1 0 32016 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604666999
transform 1 0 32108 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_324
timestamp 1604666999
transform 1 0 30912 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_358
timestamp 1604666999
transform 1 0 34040 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_359
timestamp 1604666999
transform 1 0 34132 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 33120 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
timestamp 1604666999
transform 1 0 34224 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 33304 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604666999
transform 1 0 33212 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_47_367
timestamp 1604666999
transform 1 0 34868 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_362
timestamp 1604666999
transform 1 0 34408 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_369
timestamp 1604666999
transform 1 0 35052 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_363
timestamp 1604666999
transform 1 0 34500 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 34316 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 34592 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604666999
transform 1 0 35236 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1604666999
transform 1 0 34776 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
timestamp 1604666999
transform 1 0 35144 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_47_381
timestamp 1604666999
transform 1 0 36156 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_377
timestamp 1604666999
transform 1 0 35788 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604666999
transform 1 0 35972 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604666999
transform 1 0 35420 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_389
timestamp 1604666999
transform 1 0 36892 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_389
timestamp 1604666999
transform 1 0 36892 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604666999
transform 1 0 37076 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1604666999
transform 1 0 37628 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604666999
transform 1 0 36524 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1604666999
transform 1 0 37260 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1604666999
transform -1 0 38824 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1604666999
transform -1 0 38824 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_398
timestamp 1604666999
transform 1 0 37720 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_406
timestamp 1604666999
transform 1 0 38456 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1604666999
transform 1 0 38364 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1604666999
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1604666999
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1604666999
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1604666999
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_27
timestamp 1604666999
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_32
timestamp 1604666999
transform 1 0 4048 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_44
timestamp 1604666999
transform 1 0 5152 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_56
timestamp 1604666999
transform 1 0 6256 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_68
timestamp 1604666999
transform 1 0 7360 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1604666999
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_80
timestamp 1604666999
transform 1 0 8464 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_93
timestamp 1604666999
transform 1 0 9660 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_105
timestamp 1604666999
transform 1 0 10764 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_117
timestamp 1604666999
transform 1 0 11868 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_129
timestamp 1604666999
transform 1 0 12972 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1604666999
transform 1 0 14076 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1604666999
transform 1 0 15180 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_154
timestamp 1604666999
transform 1 0 15272 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_166
timestamp 1604666999
transform 1 0 16376 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_178
timestamp 1604666999
transform 1 0 17480 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_190
timestamp 1604666999
transform 1 0 18584 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1604666999
transform 1 0 20792 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_202
timestamp 1604666999
transform 1 0 19688 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_215
timestamp 1604666999
transform 1 0 20884 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
timestamp 1604666999
transform 1 0 23368 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_48_227
timestamp 1604666999
transform 1 0 21988 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_239
timestamp 1604666999
transform 1 0 23092 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 26220 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_261
timestamp 1604666999
transform 1 0 25116 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604666999
transform 1 0 26496 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604666999
transform 1 0 28060 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1604666999
transform 1 0 26404 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 27600 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_285
timestamp 1604666999
transform 1 0 27324 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_290
timestamp 1604666999
transform 1 0 27784 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_297
timestamp 1604666999
transform 1 0 28428 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
timestamp 1604666999
transform 1 0 29164 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
timestamp 1604666999
transform 1 0 28980 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1604666999
transform 1 0 32016 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
timestamp 1604666999
transform 1 0 32844 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604666999
transform 1 0 32476 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_324
timestamp 1604666999
transform 1 0 30912 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_337
timestamp 1604666999
transform 1 0 32108 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_343
timestamp 1604666999
transform 1 0 32660 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_347
timestamp 1604666999
transform 1 0 33028 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
timestamp 1604666999
transform 1 0 33212 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 35328 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_368
timestamp 1604666999
transform 1 0 34960 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604666999
transform 1 0 35696 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1604666999
transform 1 0 37628 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 36248 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_374
timestamp 1604666999
transform 1 0 35512 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_380
timestamp 1604666999
transform 1 0 36064 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_384
timestamp 1604666999
transform 1 0 36432 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_396
timestamp 1604666999
transform 1 0 37536 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1604666999
transform -1 0 38824 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_398
timestamp 1604666999
transform 1 0 37720 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_406
timestamp 1604666999
transform 1 0 38456 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1604666999
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1604666999
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1604666999
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1604666999
transform 1 0 3588 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1604666999
transform 1 0 4692 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1604666999
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_51
timestamp 1604666999
transform 1 0 5796 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_59
timestamp 1604666999
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_62
timestamp 1604666999
transform 1 0 6808 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_74
timestamp 1604666999
transform 1 0 7912 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_86
timestamp 1604666999
transform 1 0 9016 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_98
timestamp 1604666999
transform 1 0 10120 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1604666999
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_110
timestamp 1604666999
transform 1 0 11224 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_123
timestamp 1604666999
transform 1 0 12420 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_135
timestamp 1604666999
transform 1 0 13524 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_147
timestamp 1604666999
transform 1 0 14628 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_159
timestamp 1604666999
transform 1 0 15732 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_171
timestamp 1604666999
transform 1 0 16836 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1604666999
transform 1 0 17940 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_184
timestamp 1604666999
transform 1 0 18032 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_196
timestamp 1604666999
transform 1 0 19136 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_208
timestamp 1604666999
transform 1 0 20240 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_220
timestamp 1604666999
transform 1 0 21344 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
timestamp 1604666999
transform 1 0 23920 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1604666999
transform 1 0 23552 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
timestamp 1604666999
transform 1 0 23368 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
timestamp 1604666999
transform 1 0 23000 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_232
timestamp 1604666999
transform 1 0 22448 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_240
timestamp 1604666999
transform 1 0 23184 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_245
timestamp 1604666999
transform 1 0 23644 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
timestamp 1604666999
transform 1 0 26220 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
timestamp 1604666999
transform 1 0 25852 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_267
timestamp 1604666999
transform 1 0 25668 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_271
timestamp 1604666999
transform 1 0 26036 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604666999
transform 1 0 26404 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604666999
transform 1 0 27968 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604666999
transform 1 0 27784 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 27416 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_284
timestamp 1604666999
transform 1 0 27232 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_288
timestamp 1604666999
transform 1 0 27600 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_296
timestamp 1604666999
transform 1 0 28336 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
timestamp 1604666999
transform 1 0 29256 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1604666999
transform 1 0 29164 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
timestamp 1604666999
transform 1 0 28980 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
timestamp 1604666999
transform 1 0 28612 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_301
timestamp 1604666999
transform 1 0 28796 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604666999
transform 1 0 32108 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
timestamp 1604666999
transform 1 0 32844 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604666999
transform 1 0 31924 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_325
timestamp 1604666999
transform 1 0 31004 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_333
timestamp 1604666999
transform 1 0 31740 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_341
timestamp 1604666999
transform 1 0 32476 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_347
timestamp 1604666999
transform 1 0 33028 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604666999
transform 1 0 33212 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
timestamp 1604666999
transform 1 0 34868 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1604666999
transform 1 0 34776 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
timestamp 1604666999
transform 1 0 34592 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604666999
transform 1 0 34224 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_358
timestamp 1604666999
transform 1 0 34040 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_362
timestamp 1604666999
transform 1 0 34408 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604666999
transform 1 0 37352 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 36800 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_386
timestamp 1604666999
transform 1 0 36616 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_390
timestamp 1604666999
transform 1 0 36984 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1604666999
transform -1 0 38824 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604666999
transform 1 0 37904 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_398
timestamp 1604666999
transform 1 0 37720 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_402
timestamp 1604666999
transform 1 0 38088 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_406
timestamp 1604666999
transform 1 0 38456 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1604666999
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1604666999
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1604666999
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1604666999
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_27
timestamp 1604666999
transform 1 0 3588 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_32
timestamp 1604666999
transform 1 0 4048 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_44
timestamp 1604666999
transform 1 0 5152 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_56
timestamp 1604666999
transform 1 0 6256 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_68
timestamp 1604666999
transform 1 0 7360 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1604666999
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_80
timestamp 1604666999
transform 1 0 8464 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_93
timestamp 1604666999
transform 1 0 9660 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_105
timestamp 1604666999
transform 1 0 10764 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_117
timestamp 1604666999
transform 1 0 11868 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_129
timestamp 1604666999
transform 1 0 12972 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1604666999
transform 1 0 14076 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1604666999
transform 1 0 15180 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_154
timestamp 1604666999
transform 1 0 15272 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_166
timestamp 1604666999
transform 1 0 16376 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_178
timestamp 1604666999
transform 1 0 17480 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_190
timestamp 1604666999
transform 1 0 18584 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1604666999
transform 1 0 20792 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_202
timestamp 1604666999
transform 1 0 19688 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_215
timestamp 1604666999
transform 1 0 20884 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
timestamp 1604666999
transform 1 0 23920 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
timestamp 1604666999
transform 1 0 23736 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_227
timestamp 1604666999
transform 1 0 21988 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_239
timestamp 1604666999
transform 1 0 23092 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_245
timestamp 1604666999
transform 1 0 23644 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 26220 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_267
timestamp 1604666999
transform 1 0 25668 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
timestamp 1604666999
transform 1 0 26496 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1604666999
transform 1 0 26404 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_295
timestamp 1604666999
transform 1 0 28244 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
timestamp 1604666999
transform 1 0 28980 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
timestamp 1604666999
transform 1 0 28796 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_322
timestamp 1604666999
transform 1 0 30728 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
timestamp 1604666999
transform 1 0 32844 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1604666999
transform 1 0 32016 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604666999
transform 1 0 32660 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_334
timestamp 1604666999
transform 1 0 31832 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_337
timestamp 1604666999
transform 1 0 32108 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604666999
transform 1 0 35328 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
timestamp 1604666999
transform 1 0 34868 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_364
timestamp 1604666999
transform 1 0 34592 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_369
timestamp 1604666999
transform 1 0 35052 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1604666999
transform 1 0 37628 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_381
timestamp 1604666999
transform 1 0 36156 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_393
timestamp 1604666999
transform 1 0 37260 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1604666999
transform -1 0 38824 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_398
timestamp 1604666999
transform 1 0 37720 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_406
timestamp 1604666999
transform 1 0 38456 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1604666999
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1604666999
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1604666999
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1604666999
transform 1 0 3588 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1604666999
transform 1 0 4692 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1604666999
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_51
timestamp 1604666999
transform 1 0 5796 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_59
timestamp 1604666999
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_62
timestamp 1604666999
transform 1 0 6808 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_74
timestamp 1604666999
transform 1 0 7912 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_86
timestamp 1604666999
transform 1 0 9016 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_98
timestamp 1604666999
transform 1 0 10120 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1604666999
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_110
timestamp 1604666999
transform 1 0 11224 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_123
timestamp 1604666999
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_135
timestamp 1604666999
transform 1 0 13524 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_147
timestamp 1604666999
transform 1 0 14628 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_159
timestamp 1604666999
transform 1 0 15732 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_171
timestamp 1604666999
transform 1 0 16836 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1604666999
transform 1 0 17940 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_184
timestamp 1604666999
transform 1 0 18032 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_196
timestamp 1604666999
transform 1 0 19136 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_208
timestamp 1604666999
transform 1 0 20240 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_220
timestamp 1604666999
transform 1 0 21344 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1604666999
transform 1 0 23552 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
timestamp 1604666999
transform 1 0 23920 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_232
timestamp 1604666999
transform 1 0 22448 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_245
timestamp 1604666999
transform 1 0 23644 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
timestamp 1604666999
transform 1 0 24932 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
timestamp 1604666999
transform 1 0 24748 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604666999
transform 1 0 24380 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_250
timestamp 1604666999
transform 1 0 24104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_255
timestamp 1604666999
transform 1 0 24564 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604666999
transform 1 0 27416 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
timestamp 1604666999
transform 1 0 26864 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604666999
transform 1 0 27232 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
timestamp 1604666999
transform 1 0 28428 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_278
timestamp 1604666999
transform 1 0 26680 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_282
timestamp 1604666999
transform 1 0 27048 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_295
timestamp 1604666999
transform 1 0 28244 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604666999
transform 1 0 29256 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1604666999
transform 1 0 29164 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604666999
transform 1 0 28796 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604666999
transform 1 0 30268 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_299
timestamp 1604666999
transform 1 0 28612 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_303
timestamp 1604666999
transform 1 0 28980 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_315
timestamp 1604666999
transform 1 0 30084 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_319
timestamp 1604666999
transform 1 0 30452 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
timestamp 1604666999
transform 1 0 32936 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
timestamp 1604666999
transform 1 0 32568 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604666999
transform 1 0 32200 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604666999
transform 1 0 31832 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_331
timestamp 1604666999
transform 1 0 31556 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_336
timestamp 1604666999
transform 1 0 32016 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_340
timestamp 1604666999
transform 1 0 32384 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_344
timestamp 1604666999
transform 1 0 32752 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604666999
transform 1 0 33120 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604666999
transform 1 0 34868 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1604666999
transform 1 0 34776 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604666999
transform 1 0 34132 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 34592 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_357
timestamp 1604666999
transform 1 0 33948 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_361
timestamp 1604666999
transform 1 0 34316 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604666999
transform 1 0 36432 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1604666999
transform 1 0 35880 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1604666999
transform 1 0 36984 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 36248 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_376
timestamp 1604666999
transform 1 0 35696 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_380
timestamp 1604666999
transform 1 0 36064 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_388
timestamp 1604666999
transform 1 0 36800 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_392
timestamp 1604666999
transform 1 0 37168 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1604666999
transform -1 0 38824 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_404
timestamp 1604666999
transform 1 0 38272 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1604666999
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1604666999
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1604666999
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1604666999
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1604666999
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1604666999
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1604666999
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_27
timestamp 1604666999
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_32
timestamp 1604666999
transform 1 0 4048 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_44
timestamp 1604666999
transform 1 0 5152 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1604666999
transform 1 0 3588 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1604666999
transform 1 0 4692 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1604666999
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_56
timestamp 1604666999
transform 1 0 6256 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_68
timestamp 1604666999
transform 1 0 7360 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_51
timestamp 1604666999
transform 1 0 5796 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_59
timestamp 1604666999
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_62
timestamp 1604666999
transform 1 0 6808 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_74
timestamp 1604666999
transform 1 0 7912 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1604666999
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_80
timestamp 1604666999
transform 1 0 8464 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_93
timestamp 1604666999
transform 1 0 9660 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_86
timestamp 1604666999
transform 1 0 9016 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_98
timestamp 1604666999
transform 1 0 10120 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1604666999
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_105
timestamp 1604666999
transform 1 0 10764 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_117
timestamp 1604666999
transform 1 0 11868 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_110
timestamp 1604666999
transform 1 0 11224 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_123
timestamp 1604666999
transform 1 0 12420 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_129
timestamp 1604666999
transform 1 0 12972 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1604666999
transform 1 0 14076 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_135
timestamp 1604666999
transform 1 0 13524 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_147
timestamp 1604666999
transform 1 0 14628 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1604666999
transform 1 0 15180 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_154
timestamp 1604666999
transform 1 0 15272 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_166
timestamp 1604666999
transform 1 0 16376 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_159
timestamp 1604666999
transform 1 0 15732 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_171
timestamp 1604666999
transform 1 0 16836 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1604666999
transform 1 0 17940 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_178
timestamp 1604666999
transform 1 0 17480 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_190
timestamp 1604666999
transform 1 0 18584 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_184
timestamp 1604666999
transform 1 0 18032 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_196
timestamp 1604666999
transform 1 0 19136 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1604666999
transform 1 0 20792 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_202
timestamp 1604666999
transform 1 0 19688 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_215
timestamp 1604666999
transform 1 0 20884 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_208
timestamp 1604666999
transform 1 0 20240 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_220
timestamp 1604666999
transform 1 0 21344 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1604666999
transform 1 0 23552 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_227
timestamp 1604666999
transform 1 0 21988 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_239
timestamp 1604666999
transform 1 0 23092 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_232
timestamp 1604666999
transform 1 0 22448 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_245
timestamp 1604666999
transform 1 0 23644 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_257
timestamp 1604666999
transform 1 0 24748 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_254
timestamp 1604666999
transform 1 0 24472 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1604666999
transform 1 0 24196 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604666999
transform 1 0 24288 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604666999
transform 1 0 24840 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
timestamp 1604666999
transform 1 0 24656 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604666999
transform 1 0 24840 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_52_267
timestamp 1604666999
transform 1 0 25668 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_272
timestamp 1604666999
transform 1 0 26128 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_260
timestamp 1604666999
transform 1 0 25024 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
timestamp 1604666999
transform 1 0 26864 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1604666999
transform 1 0 26404 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 28244 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604666999
transform 1 0 27416 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_276
timestamp 1604666999
transform 1 0 26496 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_284
timestamp 1604666999
transform 1 0 27232 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_288
timestamp 1604666999
transform 1 0 27600 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_294
timestamp 1604666999
transform 1 0 28152 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_297
timestamp 1604666999
transform 1 0 28428 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_301
timestamp 1604666999
transform 1 0 28796 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_308
timestamp 1604666999
transform 1 0 29440 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_305
timestamp 1604666999
transform 1 0 29164 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_299
timestamp 1604666999
transform 1 0 28612 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604666999
transform 1 0 29624 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604666999
transform 1 0 29256 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 28612 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1604666999
transform 1 0 29164 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_318
timestamp 1604666999
transform 1 0 30360 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_306
timestamp 1604666999
transform 1 0 29256 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_312
timestamp 1604666999
transform 1 0 29808 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_332
timestamp 1604666999
transform 1 0 31648 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_326
timestamp 1604666999
transform 1 0 31096 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604666999
transform 1 0 30912 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604666999
transform 1 0 31464 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 31832 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604666999
transform 1 0 32016 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604666999
transform 1 0 32108 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1604666999
transform 1 0 32016 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_340
timestamp 1604666999
transform 1 0 32384 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 32568 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 32660 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_341
timestamp 1604666999
transform 1 0 32476 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_344
timestamp 1604666999
transform 1 0 32752 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 32936 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604666999
transform 1 0 33028 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_345
timestamp 1604666999
transform 1 0 32844 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_324
timestamp 1604666999
transform 1 0 30912 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_357
timestamp 1604666999
transform 1 0 33948 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604666999
transform 1 0 34224 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604666999
transform 1 0 33120 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_367
timestamp 1604666999
transform 1 0 34868 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_362
timestamp 1604666999
transform 1 0 34408 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_372
timestamp 1604666999
transform 1 0 35328 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_368
timestamp 1604666999
transform 1 0 34960 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
timestamp 1604666999
transform 1 0 34592 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
timestamp 1604666999
transform 1 0 35144 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1604666999
transform 1 0 34776 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604666999
transform 1 0 35052 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
timestamp 1604666999
transform 1 0 33212 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_53_378
timestamp 1604666999
transform 1 0 35880 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_380
timestamp 1604666999
transform 1 0 36064 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 36248 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604666999
transform 1 0 36064 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604666999
transform 1 0 35512 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604666999
transform 1 0 35696 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_396
timestamp 1604666999
transform 1 0 37536 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1604666999
transform 1 0 37628 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_394
timestamp 1604666999
transform 1 0 37352 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_382
timestamp 1604666999
transform 1 0 36248 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_384
timestamp 1604666999
transform 1 0 36432 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1604666999
transform -1 0 38824 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1604666999
transform -1 0 38824 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_398
timestamp 1604666999
transform 1 0 37720 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_406
timestamp 1604666999
transform 1 0 38456 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_406
timestamp 1604666999
transform 1 0 38456 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1604666999
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1604666999
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1604666999
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1604666999
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_27
timestamp 1604666999
transform 1 0 3588 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_32
timestamp 1604666999
transform 1 0 4048 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_44
timestamp 1604666999
transform 1 0 5152 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_56
timestamp 1604666999
transform 1 0 6256 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_68
timestamp 1604666999
transform 1 0 7360 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1604666999
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_80
timestamp 1604666999
transform 1 0 8464 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_93
timestamp 1604666999
transform 1 0 9660 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_105
timestamp 1604666999
transform 1 0 10764 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_117
timestamp 1604666999
transform 1 0 11868 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_129
timestamp 1604666999
transform 1 0 12972 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1604666999
transform 1 0 14076 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1604666999
transform 1 0 15180 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_154
timestamp 1604666999
transform 1 0 15272 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_166
timestamp 1604666999
transform 1 0 16376 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_178
timestamp 1604666999
transform 1 0 17480 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_190
timestamp 1604666999
transform 1 0 18584 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1604666999
transform 1 0 20792 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_202
timestamp 1604666999
transform 1 0 19688 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_215
timestamp 1604666999
transform 1 0 20884 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_227
timestamp 1604666999
transform 1 0 21988 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_239
timestamp 1604666999
transform 1 0 23092 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_251
timestamp 1604666999
transform 1 0 24196 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_263
timestamp 1604666999
transform 1 0 25300 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 28244 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1604666999
transform 1 0 26404 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_276
timestamp 1604666999
transform 1 0 26496 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_288
timestamp 1604666999
transform 1 0 27600 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_294
timestamp 1604666999
transform 1 0 28152 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 30360 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 30728 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_314
timestamp 1604666999
transform 1 0 29992 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_320
timestamp 1604666999
transform 1 0 30544 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604666999
transform 1 0 32660 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604666999
transform 1 0 30912 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1604666999
transform 1 0 32016 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 32476 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 31832 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_328
timestamp 1604666999
transform 1 0 31280 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_337
timestamp 1604666999
transform 1 0 32108 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
timestamp 1604666999
transform 1 0 35144 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604666999
transform 1 0 34960 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604666999
transform 1 0 34592 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 33672 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 34040 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_352
timestamp 1604666999
transform 1 0 33488 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_356
timestamp 1604666999
transform 1 0 33856 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_360
timestamp 1604666999
transform 1 0 34224 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_366
timestamp 1604666999
transform 1 0 34776 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1604666999
transform 1 0 37628 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_389
timestamp 1604666999
transform 1 0 36892 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1604666999
transform -1 0 38824 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_398
timestamp 1604666999
transform 1 0 37720 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_406
timestamp 1604666999
transform 1 0 38456 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1604666999
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1604666999
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1604666999
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1604666999
transform 1 0 3588 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1604666999
transform 1 0 4692 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1604666999
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_51
timestamp 1604666999
transform 1 0 5796 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_59
timestamp 1604666999
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_62
timestamp 1604666999
transform 1 0 6808 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_74
timestamp 1604666999
transform 1 0 7912 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_86
timestamp 1604666999
transform 1 0 9016 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_98
timestamp 1604666999
transform 1 0 10120 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1604666999
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_110
timestamp 1604666999
transform 1 0 11224 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_123
timestamp 1604666999
transform 1 0 12420 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_135
timestamp 1604666999
transform 1 0 13524 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_147
timestamp 1604666999
transform 1 0 14628 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_159
timestamp 1604666999
transform 1 0 15732 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_171
timestamp 1604666999
transform 1 0 16836 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1604666999
transform 1 0 17940 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_184
timestamp 1604666999
transform 1 0 18032 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_196
timestamp 1604666999
transform 1 0 19136 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_208
timestamp 1604666999
transform 1 0 20240 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_220
timestamp 1604666999
transform 1 0 21344 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1604666999
transform 1 0 23552 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_232
timestamp 1604666999
transform 1 0 22448 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_245
timestamp 1604666999
transform 1 0 23644 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_257
timestamp 1604666999
transform 1 0 24748 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_269
timestamp 1604666999
transform 1 0 25852 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1604666999
transform 1 0 26956 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1604666999
transform 1 0 28060 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604666999
transform 1 0 30360 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1604666999
transform 1 0 29164 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 29440 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 29808 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 30176 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_306
timestamp 1604666999
transform 1 0 29256 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_310
timestamp 1604666999
transform 1 0 29624 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_314
timestamp 1604666999
transform 1 0 29992 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604666999
transform 1 0 31924 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 31740 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 31372 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_327
timestamp 1604666999
transform 1 0 31188 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_331
timestamp 1604666999
transform 1 0 31556 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_344
timestamp 1604666999
transform 1 0 32752 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_350
timestamp 1604666999
transform 1 0 33304 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 33120 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 33488 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604666999
transform 1 0 33672 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_367
timestamp 1604666999
transform 1 0 34868 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_362
timestamp 1604666999
transform 1 0 34408 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_358
timestamp 1604666999
transform 1 0 34040 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1604666999
transform 1 0 34224 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
timestamp 1604666999
transform 1 0 34592 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1604666999
transform 1 0 34776 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604666999
transform 1 0 35052 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604666999
transform 1 0 36616 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1604666999
transform 1 0 37168 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604666999
transform 1 0 36064 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
timestamp 1604666999
transform 1 0 36432 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_378
timestamp 1604666999
transform 1 0 35880 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_382
timestamp 1604666999
transform 1 0 36248 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_390
timestamp 1604666999
transform 1 0 36984 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_394
timestamp 1604666999
transform 1 0 37352 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1604666999
transform -1 0 38824 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_55_406
timestamp 1604666999
transform 1 0 38456 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1604666999
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1604666999
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1604666999
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1604666999
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_27
timestamp 1604666999
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_32
timestamp 1604666999
transform 1 0 4048 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_44
timestamp 1604666999
transform 1 0 5152 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_56
timestamp 1604666999
transform 1 0 6256 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_68
timestamp 1604666999
transform 1 0 7360 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1604666999
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_80
timestamp 1604666999
transform 1 0 8464 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_93
timestamp 1604666999
transform 1 0 9660 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_105
timestamp 1604666999
transform 1 0 10764 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_117
timestamp 1604666999
transform 1 0 11868 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_129
timestamp 1604666999
transform 1 0 12972 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1604666999
transform 1 0 14076 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1604666999
transform 1 0 15180 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_154
timestamp 1604666999
transform 1 0 15272 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_166
timestamp 1604666999
transform 1 0 16376 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_178
timestamp 1604666999
transform 1 0 17480 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_190
timestamp 1604666999
transform 1 0 18584 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1604666999
transform 1 0 20792 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_202
timestamp 1604666999
transform 1 0 19688 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_215
timestamp 1604666999
transform 1 0 20884 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_227
timestamp 1604666999
transform 1 0 21988 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_239
timestamp 1604666999
transform 1 0 23092 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_251
timestamp 1604666999
transform 1 0 24196 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_263
timestamp 1604666999
transform 1 0 25300 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1604666999
transform 1 0 26404 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_276
timestamp 1604666999
transform 1 0 26496 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_288
timestamp 1604666999
transform 1 0 27600 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 29440 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_56_300
timestamp 1604666999
transform 1 0 28704 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1604666999
transform 1 0 32016 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 32476 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604666999
transform 1 0 32844 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_327
timestamp 1604666999
transform 1 0 31188 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_335
timestamp 1604666999
transform 1 0 31924 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_337
timestamp 1604666999
transform 1 0 32108 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_343
timestamp 1604666999
transform 1 0 32660 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_347
timestamp 1604666999
transform 1 0 33028 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604666999
transform 1 0 33488 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
timestamp 1604666999
transform 1 0 35144 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
timestamp 1604666999
transform 1 0 34960 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 33212 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_351
timestamp 1604666999
transform 1 0 33396 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_361
timestamp 1604666999
transform 1 0 34316 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_367
timestamp 1604666999
transform 1 0 34868 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1604666999
transform 1 0 37628 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_389
timestamp 1604666999
transform 1 0 36892 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1604666999
transform -1 0 38824 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_398
timestamp 1604666999
transform 1 0 37720 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_406
timestamp 1604666999
transform 1 0 38456 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1604666999
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1604666999
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1604666999
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1604666999
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1604666999
transform 1 0 4692 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1604666999
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_51
timestamp 1604666999
transform 1 0 5796 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_59
timestamp 1604666999
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_62
timestamp 1604666999
transform 1 0 6808 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_74
timestamp 1604666999
transform 1 0 7912 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_86
timestamp 1604666999
transform 1 0 9016 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_98
timestamp 1604666999
transform 1 0 10120 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1604666999
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_110
timestamp 1604666999
transform 1 0 11224 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_123
timestamp 1604666999
transform 1 0 12420 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_135
timestamp 1604666999
transform 1 0 13524 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_147
timestamp 1604666999
transform 1 0 14628 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_159
timestamp 1604666999
transform 1 0 15732 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_171
timestamp 1604666999
transform 1 0 16836 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1604666999
transform 1 0 17940 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_184
timestamp 1604666999
transform 1 0 18032 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_196
timestamp 1604666999
transform 1 0 19136 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_208
timestamp 1604666999
transform 1 0 20240 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_220
timestamp 1604666999
transform 1 0 21344 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1604666999
transform 1 0 23552 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_232
timestamp 1604666999
transform 1 0 22448 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_245
timestamp 1604666999
transform 1 0 23644 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_257
timestamp 1604666999
transform 1 0 24748 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_269
timestamp 1604666999
transform 1 0 25852 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1604666999
transform 1 0 26956 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1604666999
transform 1 0 28060 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 29992 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1604666999
transform 1 0 29164 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 29808 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_306
timestamp 1604666999
transform 1 0 29256 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604666999
transform 1 0 32476 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604666999
transform 1 0 32108 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_333
timestamp 1604666999
transform 1 0 31740 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_339
timestamp 1604666999
transform 1 0 32292 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_354
timestamp 1604666999
transform 1 0 33672 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_350
timestamp 1604666999
transform 1 0 33304 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
timestamp 1604666999
transform 1 0 34224 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 33488 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_367
timestamp 1604666999
transform 1 0 34868 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_362
timestamp 1604666999
transform 1 0 34408 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
timestamp 1604666999
transform 1 0 34592 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
timestamp 1604666999
transform 1 0 35052 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1604666999
transform 1 0 34776 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
timestamp 1604666999
transform 1 0 35236 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_57_390
timestamp 1604666999
transform 1 0 36984 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1604666999
transform -1 0 38824 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_402
timestamp 1604666999
transform 1 0 38088 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_406
timestamp 1604666999
transform 1 0 38456 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1604666999
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1604666999
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1604666999
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1604666999
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_27
timestamp 1604666999
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_32
timestamp 1604666999
transform 1 0 4048 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_44
timestamp 1604666999
transform 1 0 5152 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_56
timestamp 1604666999
transform 1 0 6256 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_68
timestamp 1604666999
transform 1 0 7360 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1604666999
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_80
timestamp 1604666999
transform 1 0 8464 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_93
timestamp 1604666999
transform 1 0 9660 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_105
timestamp 1604666999
transform 1 0 10764 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_117
timestamp 1604666999
transform 1 0 11868 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_129
timestamp 1604666999
transform 1 0 12972 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1604666999
transform 1 0 14076 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1604666999
transform 1 0 15180 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_154
timestamp 1604666999
transform 1 0 15272 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_166
timestamp 1604666999
transform 1 0 16376 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_178
timestamp 1604666999
transform 1 0 17480 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_190
timestamp 1604666999
transform 1 0 18584 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1604666999
transform 1 0 20792 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_202
timestamp 1604666999
transform 1 0 19688 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_215
timestamp 1604666999
transform 1 0 20884 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_227
timestamp 1604666999
transform 1 0 21988 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_239
timestamp 1604666999
transform 1 0 23092 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_251
timestamp 1604666999
transform 1 0 24196 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_263
timestamp 1604666999
transform 1 0 25300 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1604666999
transform 1 0 26404 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_276
timestamp 1604666999
transform 1 0 26496 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_288
timestamp 1604666999
transform 1 0 27600 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 29992 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 30452 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_300
timestamp 1604666999
transform 1 0 28704 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_312
timestamp 1604666999
transform 1 0 29808 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_316
timestamp 1604666999
transform 1 0 30176 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_321
timestamp 1604666999
transform 1 0 30636 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604666999
transform 1 0 32108 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1604666999
transform 1 0 32016 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_333
timestamp 1604666999
transform 1 0 31740 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
timestamp 1604666999
transform 1 0 34592 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
timestamp 1604666999
transform 1 0 34408 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 34040 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_356
timestamp 1604666999
transform 1 0 33856 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_360
timestamp 1604666999
transform 1 0 34224 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1604666999
transform 1 0 37628 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_383
timestamp 1604666999
transform 1 0 36340 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_395
timestamp 1604666999
transform 1 0 37444 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1604666999
transform -1 0 38824 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_398
timestamp 1604666999
transform 1 0 37720 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_406
timestamp 1604666999
transform 1 0 38456 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1604666999
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1604666999
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1604666999
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1604666999
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1604666999
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1604666999
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1604666999
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1604666999
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1604666999
transform 1 0 4692 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_27
timestamp 1604666999
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_32
timestamp 1604666999
transform 1 0 4048 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_44
timestamp 1604666999
transform 1 0 5152 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1604666999
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_51
timestamp 1604666999
transform 1 0 5796 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_59
timestamp 1604666999
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_62
timestamp 1604666999
transform 1 0 6808 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_74
timestamp 1604666999
transform 1 0 7912 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_56
timestamp 1604666999
transform 1 0 6256 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_68
timestamp 1604666999
transform 1 0 7360 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1604666999
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_86
timestamp 1604666999
transform 1 0 9016 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_98
timestamp 1604666999
transform 1 0 10120 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_80
timestamp 1604666999
transform 1 0 8464 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_93
timestamp 1604666999
transform 1 0 9660 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1604666999
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_110
timestamp 1604666999
transform 1 0 11224 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_123
timestamp 1604666999
transform 1 0 12420 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_105
timestamp 1604666999
transform 1 0 10764 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_117
timestamp 1604666999
transform 1 0 11868 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_135
timestamp 1604666999
transform 1 0 13524 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_147
timestamp 1604666999
transform 1 0 14628 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_129
timestamp 1604666999
transform 1 0 12972 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1604666999
transform 1 0 14076 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1604666999
transform 1 0 15180 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_159
timestamp 1604666999
transform 1 0 15732 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_171
timestamp 1604666999
transform 1 0 16836 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_154
timestamp 1604666999
transform 1 0 15272 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_166
timestamp 1604666999
transform 1 0 16376 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1604666999
transform 1 0 17940 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_184
timestamp 1604666999
transform 1 0 18032 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_196
timestamp 1604666999
transform 1 0 19136 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_178
timestamp 1604666999
transform 1 0 17480 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_190
timestamp 1604666999
transform 1 0 18584 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1604666999
transform 1 0 20792 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_208
timestamp 1604666999
transform 1 0 20240 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_220
timestamp 1604666999
transform 1 0 21344 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_202
timestamp 1604666999
transform 1 0 19688 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_215
timestamp 1604666999
transform 1 0 20884 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1604666999
transform 1 0 23552 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_232
timestamp 1604666999
transform 1 0 22448 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_245
timestamp 1604666999
transform 1 0 23644 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_227
timestamp 1604666999
transform 1 0 21988 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_239
timestamp 1604666999
transform 1 0 23092 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_257
timestamp 1604666999
transform 1 0 24748 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_269
timestamp 1604666999
transform 1 0 25852 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_251
timestamp 1604666999
transform 1 0 24196 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_263
timestamp 1604666999
transform 1 0 25300 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1604666999
transform 1 0 26404 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1604666999
transform 1 0 26956 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1604666999
transform 1 0 28060 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_276
timestamp 1604666999
transform 1 0 26496 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_288
timestamp 1604666999
transform 1 0 27600 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 30452 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1604666999
transform 1 0 29164 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 30268 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_306
timestamp 1604666999
transform 1 0 29256 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_314
timestamp 1604666999
transform 1 0 29992 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_300
timestamp 1604666999
transform 1 0 28704 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_312
timestamp 1604666999
transform 1 0 29808 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604666999
transform 1 0 32936 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
timestamp 1604666999
transform 1 0 32108 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1604666999
transform 1 0 32016 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
timestamp 1604666999
transform 1 0 32384 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
timestamp 1604666999
transform 1 0 32752 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_338
timestamp 1604666999
transform 1 0 32200 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_342
timestamp 1604666999
transform 1 0 32568 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_324
timestamp 1604666999
transform 1 0 30912 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_356
timestamp 1604666999
transform 1 0 33856 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_359
timestamp 1604666999
transform 1 0 34132 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_355
timestamp 1604666999
transform 1 0 33764 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
timestamp 1604666999
transform 1 0 34224 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_362
timestamp 1604666999
transform 1 0 34408 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
timestamp 1604666999
transform 1 0 34408 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
timestamp 1604666999
transform 1 0 34592 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1604666999
transform 1 0 34776 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
timestamp 1604666999
transform 1 0 34592 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
timestamp 1604666999
transform 1 0 34868 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604666999
transform 1 0 37352 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1604666999
transform 1 0 37628 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_386
timestamp 1604666999
transform 1 0 36616 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_383
timestamp 1604666999
transform 1 0 36340 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_395
timestamp 1604666999
transform 1 0 37444 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1604666999
transform -1 0 38824 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1604666999
transform -1 0 38824 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1604666999
transform 1 0 37904 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_398
timestamp 1604666999
transform 1 0 37720 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_402
timestamp 1604666999
transform 1 0 38088 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_406
timestamp 1604666999
transform 1 0 38456 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_398
timestamp 1604666999
transform 1 0 37720 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_406
timestamp 1604666999
transform 1 0 38456 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1604666999
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1604666999
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1604666999
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1604666999
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1604666999
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1604666999
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_51
timestamp 1604666999
transform 1 0 5796 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_59
timestamp 1604666999
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_62
timestamp 1604666999
transform 1 0 6808 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_74
timestamp 1604666999
transform 1 0 7912 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_86
timestamp 1604666999
transform 1 0 9016 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_98
timestamp 1604666999
transform 1 0 10120 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1604666999
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_110
timestamp 1604666999
transform 1 0 11224 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_123
timestamp 1604666999
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_135
timestamp 1604666999
transform 1 0 13524 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_147
timestamp 1604666999
transform 1 0 14628 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_159
timestamp 1604666999
transform 1 0 15732 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_171
timestamp 1604666999
transform 1 0 16836 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1604666999
transform 1 0 17940 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_184
timestamp 1604666999
transform 1 0 18032 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_196
timestamp 1604666999
transform 1 0 19136 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_208
timestamp 1604666999
transform 1 0 20240 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_220
timestamp 1604666999
transform 1 0 21344 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1604666999
transform 1 0 23552 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_232
timestamp 1604666999
transform 1 0 22448 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_245
timestamp 1604666999
transform 1 0 23644 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_257
timestamp 1604666999
transform 1 0 24748 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_269
timestamp 1604666999
transform 1 0 25852 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1604666999
transform 1 0 26956 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1604666999
transform 1 0 28060 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1604666999
transform 1 0 29164 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_306
timestamp 1604666999
transform 1 0 29256 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_318
timestamp 1604666999
transform 1 0 30360 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 32936 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_330
timestamp 1604666999
transform 1 0 31464 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_342
timestamp 1604666999
transform 1 0 32568 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1604666999
transform 1 0 34776 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A
timestamp 1604666999
transform 1 0 35236 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 33304 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_348
timestamp 1604666999
transform 1 0 33120 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_352
timestamp 1604666999
transform 1 0 33488 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_364
timestamp 1604666999
transform 1 0 34592 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_367
timestamp 1604666999
transform 1 0 34868 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1604666999
transform 1 0 35420 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1604666999
transform 1 0 35972 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_377
timestamp 1604666999
transform 1 0 35788 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_381
timestamp 1604666999
transform 1 0 36156 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1604666999
transform 1 0 37260 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1604666999
transform -1 0 38824 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1604666999
transform 1 0 38364 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1604666999
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1604666999
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1604666999
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1604666999
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_27
timestamp 1604666999
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_32
timestamp 1604666999
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_44
timestamp 1604666999
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_56
timestamp 1604666999
transform 1 0 6256 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_68
timestamp 1604666999
transform 1 0 7360 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1604666999
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_80
timestamp 1604666999
transform 1 0 8464 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_93
timestamp 1604666999
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_105
timestamp 1604666999
transform 1 0 10764 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_117
timestamp 1604666999
transform 1 0 11868 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_129
timestamp 1604666999
transform 1 0 12972 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1604666999
transform 1 0 14076 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1604666999
transform 1 0 15180 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_154
timestamp 1604666999
transform 1 0 15272 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_166
timestamp 1604666999
transform 1 0 16376 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_178
timestamp 1604666999
transform 1 0 17480 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_190
timestamp 1604666999
transform 1 0 18584 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1604666999
transform 1 0 20792 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_202
timestamp 1604666999
transform 1 0 19688 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_215
timestamp 1604666999
transform 1 0 20884 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_227
timestamp 1604666999
transform 1 0 21988 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_239
timestamp 1604666999
transform 1 0 23092 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_251
timestamp 1604666999
transform 1 0 24196 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_263
timestamp 1604666999
transform 1 0 25300 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1604666999
transform 1 0 26404 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_276
timestamp 1604666999
transform 1 0 26496 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_288
timestamp 1604666999
transform 1 0 27600 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_300
timestamp 1604666999
transform 1 0 28704 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_312
timestamp 1604666999
transform 1 0 29808 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1604666999
transform 1 0 32016 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_324
timestamp 1604666999
transform 1 0 30912 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_337
timestamp 1604666999
transform 1 0 32108 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_349
timestamp 1604666999
transform 1 0 33212 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_361
timestamp 1604666999
transform 1 0 34316 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1604666999
transform 1 0 35420 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1604666999
transform 1 0 37628 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1604666999
transform 1 0 35788 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_389
timestamp 1604666999
transform 1 0 36892 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1604666999
transform -1 0 38824 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_398
timestamp 1604666999
transform 1 0 37720 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_406
timestamp 1604666999
transform 1 0 38456 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1604666999
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1604666999
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1604666999
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1604666999
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1604666999
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1604666999
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_51
timestamp 1604666999
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_59
timestamp 1604666999
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_62
timestamp 1604666999
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_74
timestamp 1604666999
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_86
timestamp 1604666999
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_98
timestamp 1604666999
transform 1 0 10120 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1604666999
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_110
timestamp 1604666999
transform 1 0 11224 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_123
timestamp 1604666999
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_135
timestamp 1604666999
transform 1 0 13524 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_147
timestamp 1604666999
transform 1 0 14628 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_159
timestamp 1604666999
transform 1 0 15732 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_171
timestamp 1604666999
transform 1 0 16836 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1604666999
transform 1 0 17940 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_184
timestamp 1604666999
transform 1 0 18032 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_196
timestamp 1604666999
transform 1 0 19136 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_208
timestamp 1604666999
transform 1 0 20240 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_220
timestamp 1604666999
transform 1 0 21344 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1604666999
transform 1 0 23552 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_232
timestamp 1604666999
transform 1 0 22448 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_245
timestamp 1604666999
transform 1 0 23644 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_257
timestamp 1604666999
transform 1 0 24748 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_269
timestamp 1604666999
transform 1 0 25852 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1604666999
transform 1 0 26956 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1604666999
transform 1 0 28060 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1604666999
transform 1 0 29164 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_306
timestamp 1604666999
transform 1 0 29256 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_318
timestamp 1604666999
transform 1 0 30360 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_330
timestamp 1604666999
transform 1 0 31464 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_342
timestamp 1604666999
transform 1 0 32568 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1604666999
transform 1 0 34776 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_354
timestamp 1604666999
transform 1 0 33672 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_367
timestamp 1604666999
transform 1 0 34868 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_379
timestamp 1604666999
transform 1 0 35972 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_391
timestamp 1604666999
transform 1 0 37076 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1604666999
transform -1 0 38824 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_403
timestamp 1604666999
transform 1 0 38180 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1604666999
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1604666999
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1604666999
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1604666999
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_27
timestamp 1604666999
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_32
timestamp 1604666999
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_44
timestamp 1604666999
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1604666999
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_56
timestamp 1604666999
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_63
timestamp 1604666999
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1604666999
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_75
timestamp 1604666999
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_87
timestamp 1604666999
transform 1 0 9108 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_94
timestamp 1604666999
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1604666999
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_106
timestamp 1604666999
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_118
timestamp 1604666999
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_125
timestamp 1604666999
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_137
timestamp 1604666999
transform 1 0 13708 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_149
timestamp 1604666999
transform 1 0 14812 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1604666999
transform 1 0 15364 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_156
timestamp 1604666999
transform 1 0 15456 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_168
timestamp 1604666999
transform 1 0 16560 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1604666999
transform 1 0 18216 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_180
timestamp 1604666999
transform 1 0 17664 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_187
timestamp 1604666999
transform 1 0 18308 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1604666999
transform 1 0 21068 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_199
timestamp 1604666999
transform 1 0 19412 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_211
timestamp 1604666999
transform 1 0 20516 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_218
timestamp 1604666999
transform 1 0 21160 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1604666999
transform 1 0 23920 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_230
timestamp 1604666999
transform 1 0 22264 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_242
timestamp 1604666999
transform 1 0 23368 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_249
timestamp 1604666999
transform 1 0 24012 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_261
timestamp 1604666999
transform 1 0 25116 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_273
timestamp 1604666999
transform 1 0 26220 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1604666999
transform 1 0 26772 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_280
timestamp 1604666999
transform 1 0 26864 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_292
timestamp 1604666999
transform 1 0 27968 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1604666999
transform 1 0 29624 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_304
timestamp 1604666999
transform 1 0 29072 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_311
timestamp 1604666999
transform 1 0 29716 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1604666999
transform 1 0 32476 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_323
timestamp 1604666999
transform 1 0 30820 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_335
timestamp 1604666999
transform 1 0 31924 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_342
timestamp 1604666999
transform 1 0 32568 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1604666999
transform 1 0 35328 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_354
timestamp 1604666999
transform 1 0 33672 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_366
timestamp 1604666999
transform 1 0 34776 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_373
timestamp 1604666999
transform 1 0 35420 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_385
timestamp 1604666999
transform 1 0 36524 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_397
timestamp 1604666999
transform 1 0 37628 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1604666999
transform -1 0 38824 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1604666999
transform 1 0 38180 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_404
timestamp 1604666999
transform 1 0 38272 0 -1 37536
box -38 -48 314 592
<< labels >>
rlabel metal2 s 38290 0 38346 480 6 Test_en
port 0 nsew default input
rlabel metal2 s 9402 0 9458 480 6 bottom_width_0_height_0__pin_16_
port 1 nsew default input
rlabel metal2 s 10506 0 10562 480 6 bottom_width_0_height_0__pin_17_
port 2 nsew default input
rlabel metal2 s 11610 0 11666 480 6 bottom_width_0_height_0__pin_18_
port 3 nsew default input
rlabel metal2 s 12714 0 12770 480 6 bottom_width_0_height_0__pin_19_
port 4 nsew default input
rlabel metal2 s 13910 0 13966 480 6 bottom_width_0_height_0__pin_20_
port 5 nsew default input
rlabel metal2 s 15014 0 15070 480 6 bottom_width_0_height_0__pin_21_
port 6 nsew default input
rlabel metal2 s 16118 0 16174 480 6 bottom_width_0_height_0__pin_22_
port 7 nsew default input
rlabel metal2 s 17222 0 17278 480 6 bottom_width_0_height_0__pin_23_
port 8 nsew default input
rlabel metal2 s 18326 0 18382 480 6 bottom_width_0_height_0__pin_24_
port 9 nsew default input
rlabel metal2 s 19430 0 19486 480 6 bottom_width_0_height_0__pin_25_
port 10 nsew default input
rlabel metal2 s 20534 0 20590 480 6 bottom_width_0_height_0__pin_26_
port 11 nsew default input
rlabel metal2 s 21638 0 21694 480 6 bottom_width_0_height_0__pin_27_
port 12 nsew default input
rlabel metal2 s 22742 0 22798 480 6 bottom_width_0_height_0__pin_28_
port 13 nsew default input
rlabel metal2 s 23846 0 23902 480 6 bottom_width_0_height_0__pin_29_
port 14 nsew default input
rlabel metal2 s 24950 0 25006 480 6 bottom_width_0_height_0__pin_30_
port 15 nsew default input
rlabel metal2 s 26054 0 26110 480 6 bottom_width_0_height_0__pin_31_
port 16 nsew default input
rlabel metal2 s 29458 0 29514 480 6 bottom_width_0_height_0__pin_42_lower
port 17 nsew default tristate
rlabel metal2 s 570 0 626 480 6 bottom_width_0_height_0__pin_42_upper
port 18 nsew default tristate
rlabel metal2 s 30562 0 30618 480 6 bottom_width_0_height_0__pin_43_lower
port 19 nsew default tristate
rlabel metal2 s 1674 0 1730 480 6 bottom_width_0_height_0__pin_43_upper
port 20 nsew default tristate
rlabel metal2 s 31666 0 31722 480 6 bottom_width_0_height_0__pin_44_lower
port 21 nsew default tristate
rlabel metal2 s 2778 0 2834 480 6 bottom_width_0_height_0__pin_44_upper
port 22 nsew default tristate
rlabel metal2 s 32770 0 32826 480 6 bottom_width_0_height_0__pin_45_lower
port 23 nsew default tristate
rlabel metal2 s 3882 0 3938 480 6 bottom_width_0_height_0__pin_45_upper
port 24 nsew default tristate
rlabel metal2 s 33874 0 33930 480 6 bottom_width_0_height_0__pin_46_lower
port 25 nsew default tristate
rlabel metal2 s 4986 0 5042 480 6 bottom_width_0_height_0__pin_46_upper
port 26 nsew default tristate
rlabel metal2 s 34978 0 35034 480 6 bottom_width_0_height_0__pin_47_lower
port 27 nsew default tristate
rlabel metal2 s 6090 0 6146 480 6 bottom_width_0_height_0__pin_47_upper
port 28 nsew default tristate
rlabel metal2 s 36082 0 36138 480 6 bottom_width_0_height_0__pin_48_lower
port 29 nsew default tristate
rlabel metal2 s 7194 0 7250 480 6 bottom_width_0_height_0__pin_48_upper
port 30 nsew default tristate
rlabel metal2 s 37186 0 37242 480 6 bottom_width_0_height_0__pin_49_lower
port 31 nsew default tristate
rlabel metal2 s 8298 0 8354 480 6 bottom_width_0_height_0__pin_49_upper
port 32 nsew default tristate
rlabel metal2 s 27250 0 27306 480 6 bottom_width_0_height_0__pin_50_
port 33 nsew default tristate
rlabel metal2 s 28354 0 28410 480 6 bottom_width_0_height_0__pin_51_
port 34 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 ccff_head
port 35 nsew default input
rlabel metal3 s 39520 10208 40000 10328 6 ccff_tail
port 36 nsew default tristate
rlabel metal2 s 39394 0 39450 480 6 clk
port 37 nsew default input
rlabel metal3 s 0 33328 480 33448 6 left_width_0_height_0__pin_52_
port 38 nsew default input
rlabel metal3 s 0 6672 480 6792 6 prog_clk
port 39 nsew default input
rlabel metal3 s 39520 11432 40000 11552 6 right_width_0_height_0__pin_0_
port 40 nsew default input
rlabel metal3 s 39520 23536 40000 23656 6 right_width_0_height_0__pin_10_
port 41 nsew default input
rlabel metal3 s 39520 24760 40000 24880 6 right_width_0_height_0__pin_11_
port 42 nsew default input
rlabel metal3 s 39520 25984 40000 26104 6 right_width_0_height_0__pin_12_
port 43 nsew default input
rlabel metal3 s 39520 27208 40000 27328 6 right_width_0_height_0__pin_13_
port 44 nsew default input
rlabel metal3 s 39520 28296 40000 28416 6 right_width_0_height_0__pin_14_
port 45 nsew default input
rlabel metal3 s 39520 29520 40000 29640 6 right_width_0_height_0__pin_15_
port 46 nsew default input
rlabel metal3 s 39520 12656 40000 12776 6 right_width_0_height_0__pin_1_
port 47 nsew default input
rlabel metal3 s 39520 13880 40000 14000 6 right_width_0_height_0__pin_2_
port 48 nsew default input
rlabel metal3 s 39520 2864 40000 2984 6 right_width_0_height_0__pin_34_lower
port 49 nsew default tristate
rlabel metal3 s 39520 30744 40000 30864 6 right_width_0_height_0__pin_34_upper
port 50 nsew default tristate
rlabel metal3 s 39520 4088 40000 4208 6 right_width_0_height_0__pin_35_lower
port 51 nsew default tristate
rlabel metal3 s 39520 31968 40000 32088 6 right_width_0_height_0__pin_35_upper
port 52 nsew default tristate
rlabel metal3 s 39520 5312 40000 5432 6 right_width_0_height_0__pin_36_lower
port 53 nsew default tristate
rlabel metal3 s 39520 33192 40000 33312 6 right_width_0_height_0__pin_36_upper
port 54 nsew default tristate
rlabel metal3 s 39520 6536 40000 6656 6 right_width_0_height_0__pin_37_lower
port 55 nsew default tristate
rlabel metal3 s 39520 34416 40000 34536 6 right_width_0_height_0__pin_37_upper
port 56 nsew default tristate
rlabel metal3 s 39520 7760 40000 7880 6 right_width_0_height_0__pin_38_lower
port 57 nsew default tristate
rlabel metal3 s 39520 35640 40000 35760 6 right_width_0_height_0__pin_38_upper
port 58 nsew default tristate
rlabel metal3 s 39520 8984 40000 9104 6 right_width_0_height_0__pin_39_lower
port 59 nsew default tristate
rlabel metal3 s 39520 36864 40000 36984 6 right_width_0_height_0__pin_39_upper
port 60 nsew default tristate
rlabel metal3 s 39520 14968 40000 15088 6 right_width_0_height_0__pin_3_
port 61 nsew default input
rlabel metal3 s 39520 552 40000 672 6 right_width_0_height_0__pin_40_lower
port 62 nsew default tristate
rlabel metal3 s 39520 38088 40000 38208 6 right_width_0_height_0__pin_40_upper
port 63 nsew default tristate
rlabel metal3 s 39520 1640 40000 1760 6 right_width_0_height_0__pin_41_lower
port 64 nsew default tristate
rlabel metal3 s 39520 39312 40000 39432 6 right_width_0_height_0__pin_41_upper
port 65 nsew default tristate
rlabel metal3 s 39520 16192 40000 16312 6 right_width_0_height_0__pin_4_
port 66 nsew default input
rlabel metal3 s 39520 17416 40000 17536 6 right_width_0_height_0__pin_5_
port 67 nsew default input
rlabel metal3 s 39520 18640 40000 18760 6 right_width_0_height_0__pin_6_
port 68 nsew default input
rlabel metal3 s 39520 19864 40000 19984 6 right_width_0_height_0__pin_7_
port 69 nsew default input
rlabel metal3 s 39520 21088 40000 21208 6 right_width_0_height_0__pin_8_
port 70 nsew default input
rlabel metal3 s 39520 22312 40000 22432 6 right_width_0_height_0__pin_9_
port 71 nsew default input
rlabel metal2 s 9954 39520 10010 40000 6 top_width_0_height_0__pin_32_
port 72 nsew default input
rlabel metal2 s 29918 39520 29974 40000 6 top_width_0_height_0__pin_33_
port 73 nsew default input
rlabel metal4 s 4208 2128 4528 37584 6 VPWR
port 74 nsew default input
rlabel metal4 s 19568 2128 19888 37584 6 VGND
port 75 nsew default input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
