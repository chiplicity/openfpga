* NGSPICE file created from cbx_1__0_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_4 abstract view
.subckt sky130_fd_sc_hd__ebufn_4 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

.subckt cbx_1__0_ IO_ISOL_N SC_IN_BOT SC_IN_TOP SC_OUT_BOT SC_OUT_TOP bottom_grid_pin_0_
+ bottom_grid_pin_10_ bottom_grid_pin_12_ bottom_grid_pin_14_ bottom_grid_pin_16_
+ bottom_grid_pin_2_ bottom_grid_pin_4_ bottom_grid_pin_6_ bottom_grid_pin_8_ ccff_head
+ ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11] chanx_left_in[12]
+ chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16] chanx_left_in[17]
+ chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3]
+ chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8]
+ chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11] chanx_left_out[12]
+ chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16] chanx_left_out[17]
+ chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3]
+ chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8]
+ chanx_left_out[9] chanx_right_in[0] chanx_right_in[10] chanx_right_in[11] chanx_right_in[12]
+ chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16] chanx_right_in[17]
+ chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11] chanx_right_out[12]
+ chanx_right_out[13] chanx_right_out[14] chanx_right_out[15] chanx_right_out[16]
+ chanx_right_out[17] chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chanx_right_out[9] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8] prog_clk_0_N_in prog_clk_0_W_out top_width_0_height_0__pin_0_
+ top_width_0_height_0__pin_10_ top_width_0_height_0__pin_11_lower top_width_0_height_0__pin_11_upper
+ top_width_0_height_0__pin_12_ top_width_0_height_0__pin_13_lower top_width_0_height_0__pin_13_upper
+ top_width_0_height_0__pin_14_ top_width_0_height_0__pin_15_lower top_width_0_height_0__pin_15_upper
+ top_width_0_height_0__pin_16_ top_width_0_height_0__pin_17_lower top_width_0_height_0__pin_17_upper
+ top_width_0_height_0__pin_1_lower top_width_0_height_0__pin_1_upper top_width_0_height_0__pin_2_
+ top_width_0_height_0__pin_3_lower top_width_0_height_0__pin_3_upper top_width_0_height_0__pin_4_
+ top_width_0_height_0__pin_5_lower top_width_0_height_0__pin_5_upper top_width_0_height_0__pin_6_
+ top_width_0_height_0__pin_7_lower top_width_0_height_0__pin_7_upper top_width_0_height_0__pin_8_
+ top_width_0_height_0__pin_9_lower top_width_0_height_0__pin_9_upper VPWR VGND
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_top_ipin_7.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_1.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_83_ chanx_right_in[1] VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_2
XFILLER_8_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_66_ _66_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4] sky130_fd_sc_hd__buf_2
XFILLER_5_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_6.mux_l2_in_0_ mux_top_ipin_6.mux_l1_in_1_/X mux_top_ipin_6.mux_l1_in_0_/X
+ mux_top_ipin_6.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_49_ chanx_left_in[16] VGND VGND VPWR VPWR chanx_right_out[16] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_6.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_6.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_1.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_82_ chanx_right_in[0] VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_2
XFILLER_10_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_65_ _65_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3] sky130_fd_sc_hd__buf_2
X_48_ chanx_left_in[15] VGND VGND VPWR VPWR chanx_right_out[15] sky130_fd_sc_hd__buf_2
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_6.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_6.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_81_ SC_IN_BOT VGND VGND VPWR VPWR SC_OUT_TOP sky130_fd_sc_hd__buf_2
XFILLER_12_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_64_ _64_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2] sky130_fd_sc_hd__buf_2
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xlogical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _58_/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
XFILLER_4_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_4.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_8_ sky130_fd_sc_hd__buf_4
XFILLER_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_47_ chanx_left_in[14] VGND VGND VPWR VPWR chanx_right_out[14] sky130_fd_sc_hd__buf_2
XFILLER_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_80_ SC_IN_TOP VGND VGND VPWR VPWR SC_OUT_BOT sky130_fd_sc_hd__buf_2
XFILLER_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_63_ _63_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1] sky130_fd_sc_hd__buf_2
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xprog_clk_0_FTB00 prog_clk_0_N_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
XFILLER_0_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_46_ chanx_left_in[13] VGND VGND VPWR VPWR chanx_right_out[13] sky130_fd_sc_hd__buf_2
XFILLER_9_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29_ chanx_right_in[16] VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_2
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xlogical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_/CLK logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xlogical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N VGND VGND VPWR VPWR _58_/A sky130_fd_sc_hd__or2b_4
Xmux_top_ipin_2.mux_l2_in_3_ _11_/HI chanx_right_in[18] mux_top_ipin_2.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_62_ _62_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0] sky130_fd_sc_hd__buf_2
XFILLER_5_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_2.mux_l4_in_0_ mux_top_ipin_2.mux_l3_in_1_/X mux_top_ipin_2.mux_l3_in_0_/X
+ mux_top_ipin_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_45_ chanx_left_in[12] VGND VGND VPWR VPWR chanx_right_out[12] sky130_fd_sc_hd__buf_2
X_28_ chanx_right_in[15] VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_7.mux_l2_in_3_ _16_/HI chanx_right_in[17] mux_top_ipin_7.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_2.mux_l3_in_1_ mux_top_ipin_2.mux_l2_in_3_/X mux_top_ipin_2.mux_l2_in_2_/X
+ mux_top_ipin_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_2.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[12] mux_top_ipin_2.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_7.mux_l4_in_0_ mux_top_ipin_7.mux_l3_in_1_/X mux_top_ipin_7.mux_l3_in_0_/X
+ mux_top_ipin_7.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_61_ _61_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8] sky130_fd_sc_hd__buf_2
XFILLER_5_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_7.mux_l3_in_1_ mux_top_ipin_7.mux_l2_in_3_/X mux_top_ipin_7.mux_l2_in_2_/X
+ mux_top_ipin_7.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_44_ chanx_left_in[11] VGND VGND VPWR VPWR chanx_right_out[11] sky130_fd_sc_hd__buf_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27_ chanx_right_in[14] VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_7.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[11] mux_top_ipin_7.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xlogical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_/CLK logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_2.mux_l3_in_0_ mux_top_ipin_2.mux_l2_in_1_/X mux_top_ipin_2.mux_l2_in_0_/X
+ mux_top_ipin_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_2.mux_l2_in_1_ chanx_left_in[12] mux_top_ipin_2.mux_l1_in_2_/X mux_top_ipin_2.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_60_ _60_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_2.mux_l1_in_2_ chanx_right_in[6] chanx_left_in[6] mux_top_ipin_2.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_7.mux_l3_in_0_ mux_top_ipin_7.mux_l2_in_1_/X mux_top_ipin_7.mux_l2_in_0_/X
+ mux_top_ipin_7.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_7.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_14_ sky130_fd_sc_hd__buf_4
X_43_ chanx_left_in[10] VGND VGND VPWR VPWR chanx_right_out[10] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_7.mux_l2_in_1_ chanx_left_in[11] mux_top_ipin_7.mux_l1_in_2_/X mux_top_ipin_7.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26_ chanx_right_in[13] VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_2
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09_ VGND VGND VPWR VPWR _09_/HI _09_/LO sky130_fd_sc_hd__conb_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_7.mux_l1_in_2_ chanx_right_in[7] chanx_left_in[7] mux_top_ipin_7.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_2.mux_l2_in_0_ mux_top_ipin_2.mux_l1_in_1_/X mux_top_ipin_2.mux_l1_in_0_/X
+ mux_top_ipin_2.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _53_/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
XFILLER_5_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_2.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_2.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_1.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_42_ chanx_left_in[9] VGND VGND VPWR VPWR chanx_right_out[9] sky130_fd_sc_hd__buf_2
XFILLER_20_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_7.mux_l2_in_0_ mux_top_ipin_7.mux_l1_in_1_/X mux_top_ipin_7.mux_l1_in_0_/X
+ mux_top_ipin_7.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_25_ chanx_right_in[12] VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_2
XFILLER_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_7.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_7.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xlogical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N VGND VGND VPWR VPWR _56_/A sky130_fd_sc_hd__or2b_4
XFILLER_7_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_top_ipin_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ sky130_fd_sc_hd__clkbuf_1
Xmux_top_ipin_2.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_2.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_1.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_41_ chanx_left_in[8] VGND VGND VPWR VPWR chanx_right_out[8] sky130_fd_sc_hd__buf_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24_ chanx_right_in[11] VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_2
XFILLER_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_top_ipin_7.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_0.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_0_ sky130_fd_sc_hd__buf_4
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_7.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_7.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xlogical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
+ logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR top_width_0_height_0__pin_13_lower sky130_fd_sc_hd__ebufn_4
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_4.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_1.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_40_ chanx_left_in[7] VGND VGND VPWR VPWR chanx_right_out[7] sky130_fd_sc_hd__buf_2
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23_ chanx_right_in[10] VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_2
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_top_ipin_7.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xlogical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
+ logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR top_width_0_height_0__pin_7_lower sky130_fd_sc_hd__ebufn_4
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_4.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xlogical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_/CLK logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ sky130_fd_sc_hd__dfxtp_1
Xlogical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _57_/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22_ chanx_right_in[9] VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_2
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_top_ipin_7.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
+ logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR top_width_0_height_0__pin_1_lower sky130_fd_sc_hd__ebufn_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_3.mux_l2_in_3_ _12_/HI chanx_right_in[19] mux_top_ipin_3.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21_ chanx_right_in[8] VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_2
XFILLER_1_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_top_ipin_6.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_3.mux_l4_in_0_ mux_top_ipin_3.mux_l3_in_1_/X mux_top_ipin_3.mux_l3_in_0_/X
+ mux_top_ipin_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_8.mux_l2_in_3_ _17_/HI chanx_right_in[18] mux_top_ipin_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xlogical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N VGND VGND VPWR VPWR _54_/A sky130_fd_sc_hd__or2b_4
Xmux_top_ipin_3.mux_l3_in_1_ mux_top_ipin_3.mux_l2_in_3_/X mux_top_ipin_3.mux_l2_in_2_/X
+ mux_top_ipin_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_3.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[13] mux_top_ipin_3.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_8.mux_l4_in_0_ mux_top_ipin_8.mux_l3_in_1_/X mux_top_ipin_8.mux_l3_in_0_/X
+ mux_top_ipin_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20_ chanx_right_in[7] VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_8.mux_l3_in_1_ mux_top_ipin_8.mux_l2_in_3_/X mux_top_ipin_8.mux_l2_in_2_/X
+ mux_top_ipin_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_8.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[12] mux_top_ipin_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_3.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_6_ sky130_fd_sc_hd__buf_4
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_3.mux_l3_in_0_ mux_top_ipin_3.mux_l2_in_1_/X mux_top_ipin_3.mux_l2_in_0_/X
+ mux_top_ipin_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_3.mux_l2_in_1_ chanx_left_in[13] mux_top_ipin_3.mux_l1_in_2_/X mux_top_ipin_3.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_3.mux_l1_in_2_ chanx_right_in[7] chanx_left_in[7] mux_top_ipin_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xlogical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _61_/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
X_79_ top_width_0_height_0__pin_9_lower VGND VGND VPWR VPWR top_width_0_height_0__pin_9_upper
+ sky130_fd_sc_hd__buf_2
Xmux_top_ipin_8.mux_l3_in_0_ mux_top_ipin_8.mux_l2_in_1_/X mux_top_ipin_8.mux_l2_in_0_/X
+ mux_top_ipin_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_8.mux_l2_in_1_ chanx_left_in[12] mux_top_ipin_8.mux_l1_in_2_/X mux_top_ipin_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_8.mux_l1_in_2_ chanx_right_in[8] chanx_left_in[8] mux_top_ipin_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_3.mux_l2_in_0_ mux_top_ipin_3.mux_l1_in_1_/X mux_top_ipin_3.mux_l1_in_0_/X
+ mux_top_ipin_3.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_78_ top_width_0_height_0__pin_7_lower VGND VGND VPWR VPWR top_width_0_height_0__pin_7_upper
+ sky130_fd_sc_hd__buf_2
Xmux_top_ipin_3.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_2_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_8.mux_l2_in_0_ mux_top_ipin_8.mux_l1_in_1_/X mux_top_ipin_8.mux_l1_in_0_/X
+ mux_top_ipin_8.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xlogical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_/CLK logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ sky130_fd_sc_hd__dfxtp_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_8.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_77_ top_width_0_height_0__pin_5_lower VGND VGND VPWR VPWR top_width_0_height_0__pin_5_upper
+ sky130_fd_sc_hd__buf_2
Xmux_top_ipin_3.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xlogical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE ccff_tail
+ IO_ISOL_N VGND VGND VPWR VPWR _61_/A sky130_fd_sc_hd__or2b_4
XFILLER_21_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_8.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_76_ top_width_0_height_0__pin_3_lower VGND VGND VPWR VPWR top_width_0_height_0__pin_3_upper
+ sky130_fd_sc_hd__buf_2
XFILLER_19_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_59_ _59_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6] sky130_fd_sc_hd__buf_2
XFILLER_16_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_6.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_12_ sky130_fd_sc_hd__buf_4
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_75_ top_width_0_height_0__pin_1_lower VGND VGND VPWR VPWR top_width_0_height_0__pin_1_upper
+ sky130_fd_sc_hd__buf_2
XFILLER_19_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_58_ _58_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5] sky130_fd_sc_hd__buf_2
XFILLER_2_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xlogical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _56_/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
X_74_ top_width_0_height_0__pin_17_lower VGND VGND VPWR VPWR top_width_0_height_0__pin_17_upper
+ sky130_fd_sc_hd__buf_2
Xmux_top_ipin_4.mux_l2_in_3_ _13_/HI chanx_right_in[14] mux_top_ipin_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_57_ _57_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4] sky130_fd_sc_hd__buf_2
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_0_
+ _53_/A VGND VGND VPWR VPWR _62_/A sky130_fd_sc_hd__ebufn_4
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_4.mux_l4_in_0_ mux_top_ipin_4.mux_l3_in_1_/X mux_top_ipin_4.mux_l3_in_0_/X
+ mux_top_ipin_4.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_4.mux_l3_in_1_ mux_top_ipin_4.mux_l2_in_3_/X mux_top_ipin_4.mux_l2_in_2_/X
+ mux_top_ipin_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xlogical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_/CLK logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_73_ top_width_0_height_0__pin_15_lower VGND VGND VPWR VPWR top_width_0_height_0__pin_15_upper
+ sky130_fd_sc_hd__buf_2
Xmux_top_ipin_4.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[8] mux_top_ipin_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xprog_clk_0_W_FTB01 prog_clk_0_N_in VGND VGND VPWR VPWR prog_clk_0_W_out sky130_fd_sc_hd__buf_4
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_/CLK sky130_fd_sc_hd__clkbuf_1
X_56_ _56_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3] sky130_fd_sc_hd__buf_2
XFILLER_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xlogical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N VGND VGND VPWR VPWR _59_/A sky130_fd_sc_hd__or2b_4
X_39_ chanx_left_in[6] VGND VGND VPWR VPWR chanx_right_out[6] sky130_fd_sc_hd__buf_2
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_0.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_4.mux_l3_in_0_ mux_top_ipin_4.mux_l2_in_1_/X mux_top_ipin_4.mux_l2_in_0_/X
+ mux_top_ipin_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xlogical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
+ logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR top_width_0_height_0__pin_17_lower sky130_fd_sc_hd__ebufn_4
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_top_ipin_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_72_ top_width_0_height_0__pin_13_lower VGND VGND VPWR VPWR top_width_0_height_0__pin_13_upper
+ sky130_fd_sc_hd__buf_2
Xmux_top_ipin_4.mux_l2_in_1_ chanx_left_in[8] mux_top_ipin_4.mux_l1_in_2_/X mux_top_ipin_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_3.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
X_55_ _55_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2] sky130_fd_sc_hd__buf_2
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_4.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_top_ipin_4.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xlogical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_2_
+ _54_/A VGND VGND VPWR VPWR _63_/A sky130_fd_sc_hd__ebufn_4
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_38_ chanx_left_in[5] VGND VGND VPWR VPWR chanx_right_out[5] sky130_fd_sc_hd__buf_2
XFILLER_22_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_0.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xlogical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
+ logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR top_width_0_height_0__pin_11_lower sky130_fd_sc_hd__ebufn_4
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_6.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_71_ top_width_0_height_0__pin_11_lower VGND VGND VPWR VPWR top_width_0_height_0__pin_11_upper
+ sky130_fd_sc_hd__buf_2
Xmux_top_ipin_4.mux_l2_in_0_ mux_top_ipin_4.mux_l1_in_1_/X mux_top_ipin_4.mux_l1_in_0_/X
+ mux_top_ipin_4.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_3.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xlogical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _60_/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
XFILLER_2_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_54_ _54_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1] sky130_fd_sc_hd__buf_2
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_4.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_4.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ prog_clk_0_FTB00/X VGND VGND VPWR VPWR clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_37_ chanx_left_in[4] VGND VGND VPWR VPWR chanx_right_out[4] sky130_fd_sc_hd__buf_2
XFILLER_11_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ ccff_head VGND VGND VPWR VPWR mux_top_ipin_0.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_17_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xlogical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
+ logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR top_width_0_height_0__pin_5_lower sky130_fd_sc_hd__ebufn_4
XFILLER_3_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_6.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_70_ _70_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8] sky130_fd_sc_hd__buf_2
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xlogical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_4_
+ _55_/A VGND VGND VPWR VPWR _64_/A sky130_fd_sc_hd__ebufn_4
X_53_ _53_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0] sky130_fd_sc_hd__buf_2
XFILLER_2_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_4.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_4.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_36_ chanx_left_in[3] VGND VGND VPWR VPWR chanx_right_out[3] sky130_fd_sc_hd__buf_2
XFILLER_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19_ chanx_right_in[6] VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_2
XFILLER_4_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_2.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_4_ sky130_fd_sc_hd__buf_4
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_52_ chanx_left_in[19] VGND VGND VPWR VPWR chanx_right_out[19] sky130_fd_sc_hd__buf_2
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xlogical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N VGND VGND VPWR VPWR _57_/A sky130_fd_sc_hd__or2b_4
X_35_ chanx_left_in[2] VGND VGND VPWR VPWR chanx_right_out[2] sky130_fd_sc_hd__buf_2
XFILLER_22_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_/CLK mux_top_ipin_8.mux_l4_in_0_/S VGND
+ VGND VPWR VPWR logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18_ chanx_right_in[5] VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_2
XFILLER_17_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xlogical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_6_
+ _56_/A VGND VGND VPWR VPWR _65_/A sky130_fd_sc_hd__ebufn_4
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_51_ chanx_left_in[18] VGND VGND VPWR VPWR chanx_right_out[18] sky130_fd_sc_hd__buf_2
XFILLER_2_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34_ chanx_left_in[1] VGND VGND VPWR VPWR chanx_right_out[1] sky130_fd_sc_hd__buf_2
Xclkbuf_2_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17_ VGND VGND VPWR VPWR _17_/HI _17_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_0.mux_l2_in_3_ _09_/HI chanx_right_in[16] mux_top_ipin_0.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_0.mux_l4_in_0_ mux_top_ipin_0.mux_l3_in_1_/X mux_top_ipin_0.mux_l3_in_0_/X
+ mux_top_ipin_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_50_ chanx_left_in[17] VGND VGND VPWR VPWR chanx_right_out[17] sky130_fd_sc_hd__buf_2
XFILLER_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33_ chanx_left_in[0] VGND VGND VPWR VPWR chanx_right_out[0] sky130_fd_sc_hd__buf_2
Xlogical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_/CLK logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_5.mux_l2_in_3_ _14_/HI chanx_right_in[15] mux_top_ipin_5.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_0.mux_l3_in_1_ mux_top_ipin_0.mux_l2_in_3_/X mux_top_ipin_0.mux_l2_in_2_/X
+ mux_top_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_16_ VGND VGND VPWR VPWR _16_/HI _16_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_5.mux_l4_in_0_ mux_top_ipin_5.mux_l3_in_1_/X mux_top_ipin_5.mux_l3_in_0_/X
+ mux_top_ipin_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_0.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[10] mux_top_ipin_0.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xlogical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_8_
+ _57_/A VGND VGND VPWR VPWR _66_/A sky130_fd_sc_hd__ebufn_4
Xmux_top_ipin_5.mux_l3_in_1_ mux_top_ipin_5.mux_l2_in_3_/X mux_top_ipin_5.mux_l2_in_2_/X
+ mux_top_ipin_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xlogical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _55_/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
XFILLER_14_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_32_ chanx_right_in[19] VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_5.mux_l2_in_2_ chanx_left_in[15] chanx_right_in[9] mux_top_ipin_5.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_0.mux_l3_in_0_ mux_top_ipin_0.mux_l2_in_1_/X mux_top_ipin_0.mux_l2_in_0_/X
+ mux_top_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15_ VGND VGND VPWR VPWR _15_/HI _15_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_0.mux_l2_in_1_ chanx_left_in[10] mux_top_ipin_0.mux_l1_in_2_/X mux_top_ipin_0.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_0.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_top_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_5.mux_l3_in_0_ mux_top_ipin_5.mux_l2_in_1_/X mux_top_ipin_5.mux_l2_in_0_/X
+ mux_top_ipin_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_5.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_10_ sky130_fd_sc_hd__buf_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xlogical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N VGND VGND VPWR VPWR _55_/A sky130_fd_sc_hd__or2b_4
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_31_ chanx_right_in[18] VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_5.mux_l2_in_1_ chanx_left_in[9] mux_top_ipin_5.mux_l1_in_2_/X mux_top_ipin_5.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14_ VGND VGND VPWR VPWR _14_/HI _14_/LO sky130_fd_sc_hd__conb_1
Xmux_top_ipin_5.mux_l1_in_2_ chanx_right_in[5] chanx_left_in[5] mux_top_ipin_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_0.mux_l2_in_0_ mux_top_ipin_0.mux_l1_in_1_/X mux_top_ipin_0.mux_l1_in_0_/X
+ mux_top_ipin_0.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xlogical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_10_
+ _58_/A VGND VGND VPWR VPWR _67_/A sky130_fd_sc_hd__ebufn_4
Xmux_top_ipin_0.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_5.mux_l2_in_0_ mux_top_ipin_5.mux_l1_in_1_/X mux_top_ipin_5.mux_l1_in_0_/X
+ mux_top_ipin_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_30_ chanx_right_in[17] VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_2
XFILLER_3_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13_ VGND VGND VPWR VPWR _13_/HI _13_/LO sky130_fd_sc_hd__conb_1
XFILLER_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_5.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_0.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xlogical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _59_/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
XFILLER_9_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12_ VGND VGND VPWR VPWR _12_/HI _12_/LO sky130_fd_sc_hd__conb_1
Xclkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_6_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_5.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xlogical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_12_
+ _59_/A VGND VGND VPWR VPWR _68_/A sky130_fd_sc_hd__ebufn_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xlogical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_/CLK logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ sky130_fd_sc_hd__dfxtp_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11_ VGND VGND VPWR VPWR _11_/HI _11_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_8.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_16_ sky130_fd_sc_hd__buf_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N VGND VGND VPWR VPWR _53_/A sky130_fd_sc_hd__or2b_4
XFILLER_12_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10_ VGND VGND VPWR VPWR _10_/HI _10_/LO sky130_fd_sc_hd__conb_1
Xlogical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_14_
+ _60_/A VGND VGND VPWR VPWR _69_/A sky130_fd_sc_hd__ebufn_4
XFILLER_3_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_2.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_1.mux_l2_in_3_ _10_/HI chanx_right_in[17] mux_top_ipin_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xlogical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
+ logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR top_width_0_height_0__pin_15_lower sky130_fd_sc_hd__ebufn_4
XFILLER_6_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_top_ipin_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_86_ chanx_right_in[4] VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_2
XFILLER_12_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_1.mux_l4_in_0_ mux_top_ipin_1.mux_l3_in_1_/X mux_top_ipin_1.mux_l3_in_0_/X
+ mux_top_ipin_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_69_ _69_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7] sky130_fd_sc_hd__buf_2
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_6.mux_l2_in_3_ _15_/HI chanx_right_in[16] mux_top_ipin_6.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_1.mux_l3_in_1_ mux_top_ipin_1.mux_l2_in_3_/X mux_top_ipin_1.mux_l2_in_2_/X
+ mux_top_ipin_1.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_2.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
Xlogical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
+ logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR top_width_0_height_0__pin_9_lower sky130_fd_sc_hd__ebufn_4
Xmux_top_ipin_1.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[11] mux_top_ipin_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_6.mux_l4_in_0_ mux_top_ipin_6.mux_l3_in_1_/X mux_top_ipin_6.mux_l3_in_0_/X
+ mux_top_ipin_6.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_top_ipin_8.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_85_ chanx_right_in[3] VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_6.mux_l3_in_1_ mux_top_ipin_6.mux_l2_in_3_/X mux_top_ipin_6.mux_l2_in_2_/X
+ mux_top_ipin_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xlogical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_16_
+ _61_/A VGND VGND VPWR VPWR _70_/A sky130_fd_sc_hd__ebufn_4
Xmux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_1.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_2_ sky130_fd_sc_hd__buf_4
XFILLER_5_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_top_ipin_5.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
X_68_ _68_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6] sky130_fd_sc_hd__buf_2
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_6.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[10] mux_top_ipin_6.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_1.mux_l3_in_0_ mux_top_ipin_1.mux_l2_in_1_/X mux_top_ipin_1.mux_l2_in_0_/X
+ mux_top_ipin_1.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xlogical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
+ logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR top_width_0_height_0__pin_3_lower sky130_fd_sc_hd__ebufn_4
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_1.mux_l2_in_1_ chanx_left_in[11] mux_top_ipin_1.mux_l1_in_2_/X mux_top_ipin_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_top_ipin_8.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xlogical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _54_/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
Xmux_top_ipin_1.mux_l1_in_2_ chanx_right_in[5] chanx_left_in[5] mux_top_ipin_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_6.mux_l3_in_0_ mux_top_ipin_6.mux_l2_in_1_/X mux_top_ipin_6.mux_l2_in_0_/X
+ mux_top_ipin_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_84_ chanx_right_in[2] VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_2
XFILLER_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_top_ipin_4.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xlogical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_/CLK logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ sky130_fd_sc_hd__dfxtp_1
X_67_ _67_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5] sky130_fd_sc_hd__buf_2
XFILLER_2_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_6.mux_l2_in_1_ chanx_left_in[10] mux_top_ipin_6.mux_l1_in_2_/X mux_top_ipin_6.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_6.mux_l1_in_2_ chanx_right_in[6] chanx_left_in[6] mux_top_ipin_6.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_1.mux_l2_in_0_ mux_top_ipin_1.mux_l1_in_1_/X mux_top_ipin_1.mux_l1_in_0_/X
+ mux_top_ipin_1.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xlogical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N VGND VGND VPWR VPWR _60_/A sky130_fd_sc_hd__or2b_4
.ends

