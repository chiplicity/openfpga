magic
tech sky130A
magscale 1 2
timestamp 1605173835
<< locali >>
rect 12081 33439 12115 33609
rect 12081 29019 12115 29189
rect 11989 20315 12023 20417
rect 12265 19703 12299 19941
rect 9689 14875 9723 15045
rect 8125 6647 8159 6749
rect 6377 5151 6411 5253
rect 6469 5083 6503 5321
<< viali >>
rect 4813 36873 4847 36907
rect 4629 36669 4663 36703
rect 5273 36533 5307 36567
rect 4997 36329 5031 36363
rect 6561 36329 6595 36363
rect 4813 36193 4847 36227
rect 6377 36193 6411 36227
rect 4721 35785 4755 35819
rect 5825 35785 5859 35819
rect 7297 35785 7331 35819
rect 8401 35785 8435 35819
rect 9873 35717 9907 35751
rect 4537 35581 4571 35615
rect 5641 35581 5675 35615
rect 7113 35581 7147 35615
rect 8217 35581 8251 35615
rect 9689 35581 9723 35615
rect 4445 35513 4479 35547
rect 5089 35445 5123 35479
rect 6193 35445 6227 35479
rect 6653 35445 6687 35479
rect 7665 35445 7699 35479
rect 8033 35445 8067 35479
rect 8861 35445 8895 35479
rect 10241 35445 10275 35479
rect 1593 35241 1627 35275
rect 4261 35241 4295 35275
rect 5641 35241 5675 35275
rect 8309 35241 8343 35275
rect 1409 35105 1443 35139
rect 2513 35105 2547 35139
rect 4077 35105 4111 35139
rect 5457 35105 5491 35139
rect 6929 35105 6963 35139
rect 8125 35105 8159 35139
rect 10057 35105 10091 35139
rect 7021 35037 7055 35071
rect 7205 35037 7239 35071
rect 10149 35037 10183 35071
rect 10241 35037 10275 35071
rect 2697 34969 2731 35003
rect 2053 34901 2087 34935
rect 6561 34901 6595 34935
rect 7757 34901 7791 34935
rect 9689 34901 9723 34935
rect 10701 34901 10735 34935
rect 2145 34697 2179 34731
rect 2513 34697 2547 34731
rect 3249 34697 3283 34731
rect 4353 34697 4387 34731
rect 6285 34697 6319 34731
rect 9781 34697 9815 34731
rect 3709 34629 3743 34663
rect 5457 34629 5491 34663
rect 9045 34629 9079 34663
rect 1593 34561 1627 34595
rect 6653 34561 6687 34595
rect 1409 34493 1443 34527
rect 3065 34493 3099 34527
rect 4077 34493 4111 34527
rect 4169 34493 4203 34527
rect 4721 34493 4755 34527
rect 5273 34493 5307 34527
rect 5825 34493 5859 34527
rect 7021 34493 7055 34527
rect 7481 34493 7515 34527
rect 7665 34493 7699 34527
rect 7932 34493 7966 34527
rect 9873 34493 9907 34527
rect 10129 34493 10163 34527
rect 5181 34357 5215 34391
rect 9321 34357 9355 34391
rect 11253 34357 11287 34391
rect 2881 34153 2915 34187
rect 4261 34153 4295 34187
rect 6009 34153 6043 34187
rect 8769 34153 8803 34187
rect 9873 34153 9907 34187
rect 10241 34153 10275 34187
rect 1685 34085 1719 34119
rect 5917 34085 5951 34119
rect 7634 34085 7668 34119
rect 1409 34017 1443 34051
rect 2697 34017 2731 34051
rect 4077 34017 4111 34051
rect 7389 34017 7423 34051
rect 10793 34017 10827 34051
rect 12357 34017 12391 34051
rect 6101 33949 6135 33983
rect 10885 33949 10919 33983
rect 10977 33949 11011 33983
rect 12449 33949 12483 33983
rect 12541 33949 12575 33983
rect 5549 33881 5583 33915
rect 7205 33881 7239 33915
rect 5457 33813 5491 33847
rect 6929 33813 6963 33847
rect 9413 33813 9447 33847
rect 10425 33813 10459 33847
rect 11989 33813 12023 33847
rect 1593 33609 1627 33643
rect 5917 33609 5951 33643
rect 6561 33609 6595 33643
rect 12081 33609 12115 33643
rect 2421 33541 2455 33575
rect 9321 33541 9355 33575
rect 10885 33541 10919 33575
rect 6193 33473 6227 33507
rect 7297 33473 7331 33507
rect 7481 33473 7515 33507
rect 9229 33473 9263 33507
rect 9873 33473 9907 33507
rect 12449 33541 12483 33575
rect 13093 33473 13127 33507
rect 13461 33473 13495 33507
rect 1409 33405 1443 33439
rect 1961 33405 1995 33439
rect 3341 33405 3375 33439
rect 4169 33405 4203 33439
rect 7205 33405 7239 33439
rect 8861 33405 8895 33439
rect 9689 33405 9723 33439
rect 12081 33405 12115 33439
rect 12173 33405 12207 33439
rect 12817 33405 12851 33439
rect 3709 33337 3743 33371
rect 4436 33337 4470 33371
rect 9781 33337 9815 33371
rect 11069 33337 11103 33371
rect 12909 33337 12943 33371
rect 2789 33269 2823 33303
rect 3985 33269 4019 33303
rect 5549 33269 5583 33303
rect 6837 33269 6871 33303
rect 7849 33269 7883 33303
rect 8309 33269 8343 33303
rect 10425 33269 10459 33303
rect 11805 33269 11839 33303
rect 4261 33065 4295 33099
rect 5273 33065 5307 33099
rect 8769 33065 8803 33099
rect 10149 33065 10183 33099
rect 11621 33065 11655 33099
rect 12081 33065 12115 33099
rect 12541 33065 12575 33099
rect 12909 33065 12943 33099
rect 1685 32997 1719 33031
rect 1409 32929 1443 32963
rect 4077 32929 4111 32963
rect 5365 32929 5399 32963
rect 5632 32929 5666 32963
rect 7297 32929 7331 32963
rect 8125 32929 8159 32963
rect 8217 32929 8251 32963
rect 10508 32929 10542 32963
rect 8309 32861 8343 32895
rect 10241 32861 10275 32895
rect 6745 32793 6779 32827
rect 7757 32793 7791 32827
rect 9137 32793 9171 32827
rect 1593 32521 1627 32555
rect 4169 32521 4203 32555
rect 5181 32521 5215 32555
rect 6193 32521 6227 32555
rect 6653 32521 6687 32555
rect 8585 32521 8619 32555
rect 9781 32521 9815 32555
rect 11437 32521 11471 32555
rect 5089 32453 5123 32487
rect 8217 32453 8251 32487
rect 8769 32453 8803 32487
rect 5641 32385 5675 32419
rect 5733 32385 5767 32419
rect 7757 32385 7791 32419
rect 9321 32385 9355 32419
rect 10977 32385 11011 32419
rect 7113 32317 7147 32351
rect 9137 32317 9171 32351
rect 10793 32317 10827 32351
rect 4721 32249 4755 32283
rect 5549 32249 5583 32283
rect 7665 32249 7699 32283
rect 10149 32249 10183 32283
rect 10701 32249 10735 32283
rect 7205 32181 7239 32215
rect 7573 32181 7607 32215
rect 9229 32181 9263 32215
rect 10333 32181 10367 32215
rect 5365 31977 5399 32011
rect 7757 31977 7791 32011
rect 8585 31977 8619 32011
rect 9505 31977 9539 32011
rect 10701 31977 10735 32011
rect 6644 31909 6678 31943
rect 10057 31909 10091 31943
rect 6377 31841 6411 31875
rect 10149 31841 10183 31875
rect 4905 31773 4939 31807
rect 10333 31773 10367 31807
rect 8033 31637 8067 31671
rect 9045 31637 9079 31671
rect 9689 31637 9723 31671
rect 11161 31637 11195 31671
rect 7665 31433 7699 31467
rect 9229 31433 9263 31467
rect 6469 31365 6503 31399
rect 7113 31365 7147 31399
rect 9137 31365 9171 31399
rect 4353 31297 4387 31331
rect 5365 31297 5399 31331
rect 8217 31297 8251 31331
rect 8769 31297 8803 31331
rect 9689 31297 9723 31331
rect 9873 31297 9907 31331
rect 5181 31229 5215 31263
rect 8125 31229 8159 31263
rect 9597 31229 9631 31263
rect 4721 31161 4755 31195
rect 5273 31161 5307 31195
rect 8033 31161 8067 31195
rect 4813 31093 4847 31127
rect 6101 31093 6135 31127
rect 7481 31093 7515 31127
rect 10241 31093 10275 31127
rect 4905 30889 4939 30923
rect 7757 30889 7791 30923
rect 9321 30889 9355 30923
rect 9965 30889 9999 30923
rect 5457 30753 5491 30787
rect 11612 30753 11646 30787
rect 5549 30685 5583 30719
rect 5641 30685 5675 30719
rect 11345 30685 11379 30719
rect 1869 30549 1903 30583
rect 5089 30549 5123 30583
rect 6929 30549 6963 30583
rect 10885 30549 10919 30583
rect 12725 30549 12759 30583
rect 13001 30549 13035 30583
rect 4721 30277 4755 30311
rect 6653 30277 6687 30311
rect 10793 30277 10827 30311
rect 1685 30209 1719 30243
rect 2421 30209 2455 30243
rect 5825 30209 5859 30243
rect 7297 30209 7331 30243
rect 7389 30209 7423 30243
rect 10701 30209 10735 30243
rect 11437 30209 11471 30243
rect 12265 30209 12299 30243
rect 13093 30209 13127 30243
rect 3341 30141 3375 30175
rect 7205 30141 7239 30175
rect 11253 30141 11287 30175
rect 12817 30141 12851 30175
rect 2145 30073 2179 30107
rect 3249 30073 3283 30107
rect 3608 30073 3642 30107
rect 10333 30073 10367 30107
rect 1777 30005 1811 30039
rect 2237 30005 2271 30039
rect 5089 30005 5123 30039
rect 5549 30005 5583 30039
rect 6837 30005 6871 30039
rect 11161 30005 11195 30039
rect 11897 30005 11931 30039
rect 12449 30005 12483 30039
rect 12909 30005 12943 30039
rect 13461 30005 13495 30039
rect 2145 29801 2179 29835
rect 4169 29801 4203 29835
rect 6285 29801 6319 29835
rect 7021 29801 7055 29835
rect 13737 29801 13771 29835
rect 1685 29733 1719 29767
rect 9934 29733 9968 29767
rect 1409 29665 1443 29699
rect 4537 29665 4571 29699
rect 4629 29665 4663 29699
rect 9689 29665 9723 29699
rect 12624 29665 12658 29699
rect 4813 29597 4847 29631
rect 6377 29597 6411 29631
rect 6469 29597 6503 29631
rect 11437 29597 11471 29631
rect 12357 29597 12391 29631
rect 3433 29529 3467 29563
rect 3801 29461 3835 29495
rect 5917 29461 5951 29495
rect 8217 29461 8251 29495
rect 11069 29461 11103 29495
rect 1685 29257 1719 29291
rect 5089 29257 5123 29291
rect 6377 29257 6411 29291
rect 9505 29257 9539 29291
rect 9965 29257 9999 29291
rect 12449 29257 12483 29291
rect 11437 29189 11471 29223
rect 12081 29189 12115 29223
rect 12173 29189 12207 29223
rect 13829 29189 13863 29223
rect 8585 29121 8619 29155
rect 8769 29121 8803 29155
rect 3249 29053 3283 29087
rect 3709 29053 3743 29087
rect 6009 29053 6043 29087
rect 8033 29053 8067 29087
rect 10057 29053 10091 29087
rect 10313 29053 10347 29087
rect 13093 29121 13127 29155
rect 13461 29121 13495 29155
rect 12817 29053 12851 29087
rect 12909 29053 12943 29087
rect 3617 28985 3651 29019
rect 3976 28985 4010 29019
rect 8493 28985 8527 29019
rect 11805 28985 11839 29019
rect 12081 28985 12115 29019
rect 5549 28917 5583 28951
rect 7665 28917 7699 28951
rect 8125 28917 8159 28951
rect 9229 28917 9263 28951
rect 3709 28713 3743 28747
rect 4353 28713 4387 28747
rect 6837 28713 6871 28747
rect 8033 28713 8067 28747
rect 11069 28713 11103 28747
rect 11989 28713 12023 28747
rect 12449 28713 12483 28747
rect 13001 28713 13035 28747
rect 9505 28645 9539 28679
rect 5713 28577 5747 28611
rect 8401 28577 8435 28611
rect 9945 28577 9979 28611
rect 12357 28577 12391 28611
rect 5457 28509 5491 28543
rect 8493 28509 8527 28543
rect 8677 28509 8711 28543
rect 9045 28509 9079 28543
rect 9689 28509 9723 28543
rect 12541 28509 12575 28543
rect 7941 28441 7975 28475
rect 4721 28373 4755 28407
rect 5273 28373 5307 28407
rect 3617 28169 3651 28203
rect 4721 28169 4755 28203
rect 9045 28169 9079 28203
rect 10793 28169 10827 28203
rect 12081 28169 12115 28203
rect 8861 28101 8895 28135
rect 10701 28101 10735 28135
rect 1593 28033 1627 28067
rect 4077 28033 4111 28067
rect 4169 28033 4203 28067
rect 5825 28033 5859 28067
rect 9597 28033 9631 28067
rect 11345 28033 11379 28067
rect 12449 28033 12483 28067
rect 1409 27965 1443 27999
rect 3525 27965 3559 27999
rect 3985 27965 4019 27999
rect 5641 27965 5675 27999
rect 6837 27965 6871 27999
rect 10057 27965 10091 27999
rect 5089 27897 5123 27931
rect 5549 27897 5583 27931
rect 6653 27897 6687 27931
rect 7082 27897 7116 27931
rect 8585 27897 8619 27931
rect 11161 27897 11195 27931
rect 2237 27829 2271 27863
rect 5181 27829 5215 27863
rect 6193 27829 6227 27863
rect 8217 27829 8251 27863
rect 9413 27829 9447 27863
rect 9505 27829 9539 27863
rect 11253 27829 11287 27863
rect 3709 27625 3743 27659
rect 5273 27625 5307 27659
rect 8677 27625 8711 27659
rect 11069 27625 11103 27659
rect 12081 27625 12115 27659
rect 12449 27625 12483 27659
rect 9689 27557 9723 27591
rect 5825 27489 5859 27523
rect 7288 27489 7322 27523
rect 5917 27421 5951 27455
rect 6009 27421 6043 27455
rect 7021 27421 7055 27455
rect 5457 27285 5491 27319
rect 6929 27285 6963 27319
rect 8401 27285 8435 27319
rect 9045 27285 9079 27319
rect 10241 27285 10275 27319
rect 10701 27285 10735 27319
rect 11437 27285 11471 27319
rect 4997 27081 5031 27115
rect 6653 27081 6687 27115
rect 7021 27081 7055 27115
rect 7205 27081 7239 27115
rect 8217 27081 8251 27115
rect 10609 27081 10643 27115
rect 4905 27013 4939 27047
rect 4537 26945 4571 26979
rect 5457 26945 5491 26979
rect 5549 26945 5583 26979
rect 7757 26945 7791 26979
rect 10517 26945 10551 26979
rect 11253 26945 11287 26979
rect 4169 26877 4203 26911
rect 5365 26877 5399 26911
rect 7573 26877 7607 26911
rect 7665 26809 7699 26843
rect 10977 26809 11011 26843
rect 6009 26741 6043 26775
rect 10149 26741 10183 26775
rect 11069 26741 11103 26775
rect 4997 26537 5031 26571
rect 7573 26537 7607 26571
rect 10425 26537 10459 26571
rect 11989 26537 12023 26571
rect 12449 26537 12483 26571
rect 10793 26469 10827 26503
rect 10885 26401 10919 26435
rect 12357 26401 12391 26435
rect 10333 26333 10367 26367
rect 10977 26333 11011 26367
rect 12541 26333 12575 26367
rect 8953 26265 8987 26299
rect 5549 26197 5583 26231
rect 7297 26197 7331 26231
rect 8585 26197 8619 26231
rect 9321 26197 9355 26231
rect 6193 25993 6227 26027
rect 8493 25993 8527 26027
rect 10425 25993 10459 26027
rect 11437 25993 11471 26027
rect 11989 25993 12023 26027
rect 12633 25993 12667 26027
rect 8401 25857 8435 25891
rect 9321 25857 9355 25891
rect 9505 25857 9539 25891
rect 11069 25857 11103 25891
rect 6377 25789 6411 25823
rect 7021 25789 7055 25823
rect 8677 25789 8711 25823
rect 9965 25789 9999 25823
rect 10793 25789 10827 25823
rect 7941 25721 7975 25755
rect 9229 25721 9263 25755
rect 8861 25653 8895 25687
rect 10241 25653 10275 25687
rect 10885 25653 10919 25687
rect 13001 25653 13035 25687
rect 7849 25449 7883 25483
rect 8309 25449 8343 25483
rect 9689 25449 9723 25483
rect 10057 25449 10091 25483
rect 10701 25449 10735 25483
rect 11069 25449 11103 25483
rect 12633 25449 12667 25483
rect 4353 25381 4387 25415
rect 6193 25381 6227 25415
rect 10149 25381 10183 25415
rect 11498 25381 11532 25415
rect 4077 25313 4111 25347
rect 6101 25313 6135 25347
rect 8217 25313 8251 25347
rect 11253 25313 11287 25347
rect 6285 25245 6319 25279
rect 8401 25245 8435 25279
rect 10333 25245 10367 25279
rect 9229 25177 9263 25211
rect 4905 25109 4939 25143
rect 5733 25109 5767 25143
rect 7665 25109 7699 25143
rect 6193 24905 6227 24939
rect 7573 24905 7607 24939
rect 10793 24905 10827 24939
rect 11529 24905 11563 24939
rect 11897 24905 11931 24939
rect 5917 24837 5951 24871
rect 4721 24769 4755 24803
rect 5365 24769 5399 24803
rect 8217 24769 8251 24803
rect 8585 24769 8619 24803
rect 8953 24769 8987 24803
rect 11161 24769 11195 24803
rect 4353 24701 4387 24735
rect 5181 24701 5215 24735
rect 7481 24701 7515 24735
rect 7941 24701 7975 24735
rect 9137 24701 9171 24735
rect 9404 24701 9438 24735
rect 3985 24633 4019 24667
rect 7113 24633 7147 24667
rect 4813 24565 4847 24599
rect 5273 24565 5307 24599
rect 6653 24565 6687 24599
rect 8033 24565 8067 24599
rect 10517 24565 10551 24599
rect 5825 24361 5859 24395
rect 6837 24361 6871 24395
rect 7297 24361 7331 24395
rect 8769 24361 8803 24395
rect 9137 24361 9171 24395
rect 9689 24361 9723 24395
rect 11253 24361 11287 24395
rect 11621 24361 11655 24395
rect 6285 24293 6319 24327
rect 7656 24293 7690 24327
rect 10057 24293 10091 24327
rect 11713 24293 11747 24327
rect 6193 24225 6227 24259
rect 4813 24157 4847 24191
rect 6377 24157 6411 24191
rect 7389 24157 7423 24191
rect 10149 24157 10183 24191
rect 10333 24157 10367 24191
rect 11805 24157 11839 24191
rect 4445 24021 4479 24055
rect 9413 24021 9447 24055
rect 5917 23817 5951 23851
rect 6285 23817 6319 23851
rect 9045 23817 9079 23851
rect 10517 23817 10551 23851
rect 11345 23817 11379 23851
rect 11989 23817 12023 23851
rect 6469 23749 6503 23783
rect 8217 23749 8251 23783
rect 8493 23749 8527 23783
rect 8861 23749 8895 23783
rect 11713 23749 11747 23783
rect 4905 23681 4939 23715
rect 9505 23681 9539 23715
rect 9689 23681 9723 23715
rect 4261 23613 4295 23647
rect 6653 23613 6687 23647
rect 6837 23613 6871 23647
rect 7093 23613 7127 23647
rect 9413 23613 9447 23647
rect 4721 23545 4755 23579
rect 4813 23545 4847 23579
rect 4353 23477 4387 23511
rect 5549 23477 5583 23511
rect 10057 23477 10091 23511
rect 4445 23273 4479 23307
rect 6653 23273 6687 23307
rect 6929 23273 6963 23307
rect 7481 23273 7515 23307
rect 9137 23273 9171 23307
rect 9873 23273 9907 23307
rect 5540 23205 5574 23239
rect 4997 23137 5031 23171
rect 7849 23137 7883 23171
rect 7941 23137 7975 23171
rect 5273 23069 5307 23103
rect 8033 23069 8067 23103
rect 4813 22933 4847 22967
rect 7389 22933 7423 22967
rect 8493 22933 8527 22967
rect 3433 22729 3467 22763
rect 3801 22729 3835 22763
rect 4169 22729 4203 22763
rect 6837 22729 6871 22763
rect 7941 22729 7975 22763
rect 8401 22729 8435 22763
rect 4261 22593 4295 22627
rect 7481 22593 7515 22627
rect 10241 22593 10275 22627
rect 7205 22525 7239 22559
rect 7297 22525 7331 22559
rect 8585 22525 8619 22559
rect 8861 22525 8895 22559
rect 9965 22525 9999 22559
rect 4506 22457 4540 22491
rect 6653 22457 6687 22491
rect 5641 22389 5675 22423
rect 6193 22389 6227 22423
rect 8217 22389 8251 22423
rect 9781 22389 9815 22423
rect 5457 22185 5491 22219
rect 6653 22185 6687 22219
rect 7573 22185 7607 22219
rect 6101 22117 6135 22151
rect 6745 22117 6779 22151
rect 4333 22049 4367 22083
rect 10497 22049 10531 22083
rect 4077 21981 4111 22015
rect 6929 21981 6963 22015
rect 10241 21981 10275 22015
rect 6285 21913 6319 21947
rect 5733 21845 5767 21879
rect 7941 21845 7975 21879
rect 11621 21845 11655 21879
rect 3801 21641 3835 21675
rect 4813 21641 4847 21675
rect 6285 21641 6319 21675
rect 6469 21641 6503 21675
rect 10333 21641 10367 21675
rect 4721 21573 4755 21607
rect 1593 21505 1627 21539
rect 5365 21505 5399 21539
rect 5917 21505 5951 21539
rect 1409 21437 1443 21471
rect 5273 21437 5307 21471
rect 6653 21437 6687 21471
rect 8493 21437 8527 21471
rect 5181 21369 5215 21403
rect 7113 21369 7147 21403
rect 8401 21369 8435 21403
rect 8738 21369 8772 21403
rect 2237 21301 2271 21335
rect 4169 21301 4203 21335
rect 7481 21301 7515 21335
rect 9873 21301 9907 21335
rect 10701 21301 10735 21335
rect 2697 21097 2731 21131
rect 5181 21097 5215 21131
rect 6561 21097 6595 21131
rect 11069 21097 11103 21131
rect 1685 21029 1719 21063
rect 4905 21029 4939 21063
rect 9956 21029 9990 21063
rect 12142 21029 12176 21063
rect 1409 20961 1443 20995
rect 7757 20961 7791 20995
rect 8585 20961 8619 20995
rect 9137 20961 9171 20995
rect 9689 20961 9723 20995
rect 11897 20961 11931 20995
rect 7849 20893 7883 20927
rect 8033 20893 8067 20927
rect 7021 20825 7055 20859
rect 7389 20757 7423 20791
rect 9505 20757 9539 20791
rect 13277 20757 13311 20791
rect 5917 20553 5951 20587
rect 6653 20553 6687 20587
rect 8585 20553 8619 20587
rect 9045 20553 9079 20587
rect 11161 20485 11195 20519
rect 12449 20485 12483 20519
rect 2605 20417 2639 20451
rect 6929 20417 6963 20451
rect 9413 20417 9447 20451
rect 9781 20417 9815 20451
rect 10425 20417 10459 20451
rect 11805 20417 11839 20451
rect 11989 20417 12023 20451
rect 12265 20417 12299 20451
rect 12909 20417 12943 20451
rect 13001 20417 13035 20451
rect 7196 20349 7230 20383
rect 10241 20349 10275 20383
rect 13461 20349 13495 20383
rect 2513 20281 2547 20315
rect 2850 20281 2884 20315
rect 6285 20281 6319 20315
rect 11989 20281 12023 20315
rect 12817 20281 12851 20315
rect 1685 20213 1719 20247
rect 3985 20213 4019 20247
rect 8309 20213 8343 20247
rect 9873 20213 9907 20247
rect 10333 20213 10367 20247
rect 11437 20213 11471 20247
rect 2421 20009 2455 20043
rect 6101 20009 6135 20043
rect 6929 20009 6963 20043
rect 8125 20009 8159 20043
rect 9137 20009 9171 20043
rect 9965 20009 9999 20043
rect 11437 20009 11471 20043
rect 2881 19941 2915 19975
rect 10057 19941 10091 19975
rect 12081 19941 12115 19975
rect 12265 19941 12299 19975
rect 2789 19873 2823 19907
rect 4905 19873 4939 19907
rect 4997 19873 5031 19907
rect 6469 19873 6503 19907
rect 7297 19873 7331 19907
rect 11529 19873 11563 19907
rect 2973 19805 3007 19839
rect 5181 19805 5215 19839
rect 5641 19805 5675 19839
rect 6561 19805 6595 19839
rect 6653 19805 6687 19839
rect 7389 19805 7423 19839
rect 7573 19805 7607 19839
rect 8217 19805 8251 19839
rect 8309 19805 8343 19839
rect 11621 19805 11655 19839
rect 7757 19737 7791 19771
rect 11069 19737 11103 19771
rect 12449 19873 12483 19907
rect 13001 19873 13035 19907
rect 13093 19805 13127 19839
rect 13185 19805 13219 19839
rect 12633 19737 12667 19771
rect 3893 19669 3927 19703
rect 4537 19669 4571 19703
rect 6009 19669 6043 19703
rect 8769 19669 8803 19703
rect 10517 19669 10551 19703
rect 10885 19669 10919 19703
rect 12265 19669 12299 19703
rect 10057 19465 10091 19499
rect 11529 19465 11563 19499
rect 3801 19397 3835 19431
rect 7389 19397 7423 19431
rect 9965 19397 9999 19431
rect 11069 19397 11103 19431
rect 4261 19329 4295 19363
rect 4353 19329 4387 19363
rect 8033 19329 8067 19363
rect 9045 19329 9079 19363
rect 10609 19329 10643 19363
rect 13001 19329 13035 19363
rect 1409 19261 1443 19295
rect 1685 19261 1719 19295
rect 2513 19261 2547 19295
rect 7205 19261 7239 19295
rect 7757 19261 7791 19295
rect 8953 19261 8987 19295
rect 10425 19261 10459 19295
rect 12817 19261 12851 19295
rect 3341 19193 3375 19227
rect 5273 19193 5307 19227
rect 8861 19193 8895 19227
rect 9505 19193 9539 19227
rect 12909 19193 12943 19227
rect 2881 19125 2915 19159
rect 3709 19125 3743 19159
rect 4169 19125 4203 19159
rect 4813 19125 4847 19159
rect 5365 19125 5399 19159
rect 6101 19125 6135 19159
rect 6653 19125 6687 19159
rect 7849 19125 7883 19159
rect 8493 19125 8527 19159
rect 10517 19125 10551 19159
rect 11805 19125 11839 19159
rect 12173 19125 12207 19159
rect 12449 19125 12483 19159
rect 13461 19125 13495 19159
rect 1593 18921 1627 18955
rect 2513 18921 2547 18955
rect 4077 18921 4111 18955
rect 6009 18921 6043 18955
rect 7113 18921 7147 18955
rect 9229 18921 9263 18955
rect 9689 18921 9723 18955
rect 10149 18921 10183 18955
rect 11253 18921 11287 18955
rect 13001 18921 13035 18955
rect 3801 18853 3835 18887
rect 4445 18853 4479 18887
rect 5549 18853 5583 18887
rect 6101 18853 6135 18887
rect 12725 18853 12759 18887
rect 7205 18785 7239 18819
rect 10057 18785 10091 18819
rect 11621 18785 11655 18819
rect 4537 18717 4571 18751
rect 4629 18717 4663 18751
rect 6285 18717 6319 18751
rect 10241 18717 10275 18751
rect 11713 18717 11747 18751
rect 11805 18717 11839 18751
rect 5641 18649 5675 18683
rect 8493 18649 8527 18683
rect 11069 18649 11103 18683
rect 3249 18581 3283 18615
rect 6745 18581 6779 18615
rect 10701 18581 10735 18615
rect 4537 18377 4571 18411
rect 4813 18377 4847 18411
rect 5641 18377 5675 18411
rect 6009 18377 6043 18411
rect 6653 18377 6687 18411
rect 8493 18377 8527 18411
rect 9045 18377 9079 18411
rect 11437 18377 11471 18411
rect 12081 18377 12115 18411
rect 9321 18309 9355 18343
rect 10885 18241 10919 18275
rect 3157 18173 3191 18207
rect 6837 18173 6871 18207
rect 7093 18173 7127 18207
rect 10149 18173 10183 18207
rect 10793 18173 10827 18207
rect 3065 18105 3099 18139
rect 3424 18105 3458 18139
rect 10701 18105 10735 18139
rect 5365 18037 5399 18071
rect 8217 18037 8251 18071
rect 9781 18037 9815 18071
rect 10333 18037 10367 18071
rect 11713 18037 11747 18071
rect 2421 17833 2455 17867
rect 4353 17833 4387 17867
rect 4629 17833 4663 17867
rect 6377 17833 6411 17867
rect 7849 17833 7883 17867
rect 8493 17833 8527 17867
rect 10885 17833 10919 17867
rect 3801 17765 3835 17799
rect 8401 17765 8435 17799
rect 2789 17697 2823 17731
rect 5253 17697 5287 17731
rect 10793 17697 10827 17731
rect 2881 17629 2915 17663
rect 3065 17629 3099 17663
rect 4997 17629 5031 17663
rect 8585 17629 8619 17663
rect 10977 17629 11011 17663
rect 8033 17561 8067 17595
rect 10425 17561 10459 17595
rect 6837 17493 6871 17527
rect 7297 17493 7331 17527
rect 10057 17493 10091 17527
rect 2513 17289 2547 17323
rect 3709 17289 3743 17323
rect 7389 17289 7423 17323
rect 8493 17289 8527 17323
rect 10977 17289 11011 17323
rect 8769 17221 8803 17255
rect 2789 17153 2823 17187
rect 4261 17153 4295 17187
rect 8125 17153 8159 17187
rect 10609 17153 10643 17187
rect 3249 17085 3283 17119
rect 7757 17085 7791 17119
rect 3617 17017 3651 17051
rect 4077 17017 4111 17051
rect 10425 17017 10459 17051
rect 4169 16949 4203 16983
rect 5089 16949 5123 16983
rect 5457 16949 5491 16983
rect 7573 16949 7607 16983
rect 9781 16949 9815 16983
rect 9965 16949 9999 16983
rect 10333 16949 10367 16983
rect 3801 16745 3835 16779
rect 5089 16745 5123 16779
rect 7021 16745 7055 16779
rect 10057 16745 10091 16779
rect 10793 16745 10827 16779
rect 12357 16745 12391 16779
rect 5457 16609 5491 16643
rect 5641 16609 5675 16643
rect 5908 16609 5942 16643
rect 8217 16609 8251 16643
rect 11233 16609 11267 16643
rect 8309 16541 8343 16575
rect 8401 16541 8435 16575
rect 10977 16541 11011 16575
rect 5273 16473 5307 16507
rect 7389 16473 7423 16507
rect 7849 16405 7883 16439
rect 10425 16405 10459 16439
rect 4997 16201 5031 16235
rect 6009 16201 6043 16235
rect 11345 16201 11379 16235
rect 1593 16065 1627 16099
rect 5549 16065 5583 16099
rect 7021 16065 7055 16099
rect 9229 16065 9263 16099
rect 1409 15997 1443 16031
rect 4905 15997 4939 16031
rect 5457 15997 5491 16031
rect 6653 15929 6687 15963
rect 7266 15929 7300 15963
rect 9045 15929 9079 15963
rect 9474 15929 9508 15963
rect 2237 15861 2271 15895
rect 5365 15861 5399 15895
rect 8401 15861 8435 15895
rect 8769 15861 8803 15895
rect 10609 15861 10643 15895
rect 10977 15861 11011 15895
rect 6561 15657 6595 15691
rect 7941 15657 7975 15691
rect 8125 15657 8159 15691
rect 9229 15657 9263 15691
rect 10333 15657 10367 15691
rect 6929 15521 6963 15555
rect 7021 15453 7055 15487
rect 7113 15453 7147 15487
rect 10425 15453 10459 15487
rect 10517 15453 10551 15487
rect 5457 15385 5491 15419
rect 5089 15317 5123 15351
rect 5733 15317 5767 15351
rect 8585 15317 8619 15351
rect 9965 15317 9999 15351
rect 6653 15113 6687 15147
rect 8125 15113 8159 15147
rect 9137 15113 9171 15147
rect 9965 15113 9999 15147
rect 11069 15113 11103 15147
rect 5917 15045 5951 15079
rect 7113 15045 7147 15079
rect 9689 15045 9723 15079
rect 9781 15045 9815 15079
rect 7665 14977 7699 15011
rect 9505 14977 9539 15011
rect 3157 14909 3191 14943
rect 7481 14909 7515 14943
rect 10517 14977 10551 15011
rect 10333 14909 10367 14943
rect 3065 14841 3099 14875
rect 3402 14841 3436 14875
rect 6285 14841 6319 14875
rect 7573 14841 7607 14875
rect 9689 14841 9723 14875
rect 10425 14841 10459 14875
rect 4537 14773 4571 14807
rect 3157 14569 3191 14603
rect 4997 14569 5031 14603
rect 7205 14569 7239 14603
rect 7665 14569 7699 14603
rect 8033 14569 8067 14603
rect 10057 14569 10091 14603
rect 10333 14501 10367 14535
rect 4905 14433 4939 14467
rect 6285 14433 6319 14467
rect 7573 14433 7607 14467
rect 8125 14433 8159 14467
rect 5089 14365 5123 14399
rect 5549 14365 5583 14399
rect 8217 14365 8251 14399
rect 4537 14297 4571 14331
rect 4445 14229 4479 14263
rect 6101 14229 6135 14263
rect 6653 14229 6687 14263
rect 7389 14229 7423 14263
rect 2697 14025 2731 14059
rect 4537 14025 4571 14059
rect 6469 14025 6503 14059
rect 7389 14025 7423 14059
rect 7757 14025 7791 14059
rect 4997 13957 5031 13991
rect 8125 13957 8159 13991
rect 5549 13889 5583 13923
rect 10149 13889 10183 13923
rect 10793 13889 10827 13923
rect 2789 13821 2823 13855
rect 3056 13821 3090 13855
rect 5457 13821 5491 13855
rect 6009 13821 6043 13855
rect 8401 13821 8435 13855
rect 9413 13821 9447 13855
rect 9781 13821 9815 13855
rect 10701 13821 10735 13855
rect 10609 13753 10643 13787
rect 4169 13685 4203 13719
rect 4905 13685 4939 13719
rect 5365 13685 5399 13719
rect 10241 13685 10275 13719
rect 3709 13481 3743 13515
rect 4445 13481 4479 13515
rect 8401 13481 8435 13515
rect 8953 13481 8987 13515
rect 9413 13481 9447 13515
rect 9689 13481 9723 13515
rect 11253 13481 11287 13515
rect 1685 13413 1719 13447
rect 2973 13413 3007 13447
rect 1409 13345 1443 13379
rect 4793 13345 4827 13379
rect 7012 13345 7046 13379
rect 9137 13345 9171 13379
rect 10057 13345 10091 13379
rect 11621 13345 11655 13379
rect 11713 13345 11747 13379
rect 4537 13277 4571 13311
rect 6745 13277 6779 13311
rect 10149 13277 10183 13311
rect 10333 13277 10367 13311
rect 11805 13277 11839 13311
rect 2237 13141 2271 13175
rect 2881 13141 2915 13175
rect 5917 13141 5951 13175
rect 6653 13141 6687 13175
rect 8125 13141 8159 13175
rect 3157 12937 3191 12971
rect 3525 12937 3559 12971
rect 5089 12937 5123 12971
rect 6285 12937 6319 12971
rect 7849 12937 7883 12971
rect 8217 12937 8251 12971
rect 8401 12937 8435 12971
rect 10609 12937 10643 12971
rect 11161 12937 11195 12971
rect 3617 12869 3651 12903
rect 4629 12869 4663 12903
rect 6653 12869 6687 12903
rect 11713 12869 11747 12903
rect 1961 12801 1995 12835
rect 2697 12801 2731 12835
rect 4169 12801 4203 12835
rect 5641 12801 5675 12835
rect 5825 12801 5859 12835
rect 7481 12801 7515 12835
rect 8953 12801 8987 12835
rect 11253 12801 11287 12835
rect 12081 12801 12115 12835
rect 2421 12733 2455 12767
rect 3985 12733 4019 12767
rect 5549 12733 5583 12767
rect 7297 12733 7331 12767
rect 8585 12733 8619 12767
rect 9220 12733 9254 12767
rect 7205 12665 7239 12699
rect 2053 12597 2087 12631
rect 2513 12597 2547 12631
rect 4077 12597 4111 12631
rect 5181 12597 5215 12631
rect 6837 12597 6871 12631
rect 10333 12597 10367 12631
rect 1593 12393 1627 12427
rect 3709 12393 3743 12427
rect 4445 12393 4479 12427
rect 5181 12393 5215 12427
rect 6653 12393 6687 12427
rect 9045 12393 9079 12427
rect 10241 12393 10275 12427
rect 7082 12325 7116 12359
rect 9321 12325 9355 12359
rect 4537 12257 4571 12291
rect 5825 12257 5859 12291
rect 8677 12257 8711 12291
rect 10793 12257 10827 12291
rect 11060 12257 11094 12291
rect 4721 12189 4755 12223
rect 6837 12189 6871 12223
rect 9965 12121 9999 12155
rect 2145 12053 2179 12087
rect 3249 12053 3283 12087
rect 4077 12053 4111 12087
rect 5641 12053 5675 12087
rect 8217 12053 8251 12087
rect 12173 12053 12207 12087
rect 3157 11849 3191 11883
rect 4629 11849 4663 11883
rect 5733 11849 5767 11883
rect 6929 11849 6963 11883
rect 3065 11781 3099 11815
rect 10793 11781 10827 11815
rect 12173 11781 12207 11815
rect 3709 11713 3743 11747
rect 7481 11713 7515 11747
rect 8493 11713 8527 11747
rect 11253 11713 11287 11747
rect 11437 11713 11471 11747
rect 3525 11645 3559 11679
rect 6285 11645 6319 11679
rect 7389 11645 7423 11679
rect 8585 11645 8619 11679
rect 8852 11645 8886 11679
rect 7297 11577 7331 11611
rect 7941 11577 7975 11611
rect 10701 11577 10735 11611
rect 11161 11577 11195 11611
rect 3617 11509 3651 11543
rect 4261 11509 4295 11543
rect 4905 11509 4939 11543
rect 6653 11509 6687 11543
rect 9965 11509 9999 11543
rect 10333 11509 10367 11543
rect 11897 11509 11931 11543
rect 3249 11305 3283 11339
rect 6653 11305 6687 11339
rect 7297 11305 7331 11339
rect 7757 11305 7791 11339
rect 9505 11305 9539 11339
rect 11253 11305 11287 11339
rect 7021 11237 7055 11271
rect 8401 11237 8435 11271
rect 10885 11237 10919 11271
rect 7665 11169 7699 11203
rect 8677 11169 8711 11203
rect 10057 11169 10091 11203
rect 11621 11169 11655 11203
rect 7941 11101 7975 11135
rect 10149 11101 10183 11135
rect 10241 11101 10275 11135
rect 11713 11101 11747 11135
rect 11897 11101 11931 11135
rect 3893 11033 3927 11067
rect 9689 11033 9723 11067
rect 7665 10761 7699 10795
rect 9321 10761 9355 10795
rect 10149 10761 10183 10795
rect 11345 10693 11379 10727
rect 1593 10625 1627 10659
rect 4353 10625 4387 10659
rect 7941 10625 7975 10659
rect 10793 10625 10827 10659
rect 1409 10557 1443 10591
rect 2145 10557 2179 10591
rect 3709 10557 3743 10591
rect 4261 10557 4295 10591
rect 4169 10489 4203 10523
rect 8208 10489 8242 10523
rect 3801 10421 3835 10455
rect 6837 10421 6871 10455
rect 7389 10421 7423 10455
rect 9689 10421 9723 10455
rect 10517 10421 10551 10455
rect 10609 10421 10643 10455
rect 11621 10421 11655 10455
rect 11989 10421 12023 10455
rect 2421 10217 2455 10251
rect 3893 10217 3927 10251
rect 5825 10217 5859 10251
rect 7481 10217 7515 10251
rect 7941 10217 7975 10251
rect 8585 10217 8619 10251
rect 9781 10217 9815 10251
rect 11529 10217 11563 10251
rect 5733 10149 5767 10183
rect 6929 10149 6963 10183
rect 9045 10149 9079 10183
rect 11897 10149 11931 10183
rect 7849 10081 7883 10115
rect 10149 10081 10183 10115
rect 10241 10081 10275 10115
rect 5273 10013 5307 10047
rect 6009 10013 6043 10047
rect 7389 10013 7423 10047
rect 8125 10013 8159 10047
rect 10333 10013 10367 10047
rect 10885 9945 10919 9979
rect 5365 9877 5399 9911
rect 9413 9877 9447 9911
rect 11253 9877 11287 9911
rect 5917 9673 5951 9707
rect 7849 9673 7883 9707
rect 2329 9605 2363 9639
rect 9873 9605 9907 9639
rect 2789 9537 2823 9571
rect 2881 9537 2915 9571
rect 3893 9537 3927 9571
rect 7481 9537 7515 9571
rect 8493 9537 8527 9571
rect 10149 9537 10183 9571
rect 10517 9537 10551 9571
rect 11253 9537 11287 9571
rect 7205 9469 7239 9503
rect 11161 9469 11195 9503
rect 3801 9401 3835 9435
rect 4138 9401 4172 9435
rect 7297 9401 7331 9435
rect 8401 9401 8435 9435
rect 8738 9401 8772 9435
rect 11069 9401 11103 9435
rect 2237 9333 2271 9367
rect 2697 9333 2731 9367
rect 3433 9333 3467 9367
rect 5273 9333 5307 9367
rect 5641 9333 5675 9367
rect 6561 9333 6595 9367
rect 6837 9333 6871 9367
rect 10701 9333 10735 9367
rect 2421 9129 2455 9163
rect 6929 9129 6963 9163
rect 7757 9129 7791 9163
rect 8309 9129 8343 9163
rect 9505 9129 9539 9163
rect 11621 9129 11655 9163
rect 5334 9061 5368 9095
rect 9965 9061 9999 9095
rect 10508 9061 10542 9095
rect 7665 8993 7699 9027
rect 5089 8925 5123 8959
rect 7941 8925 7975 8959
rect 10241 8925 10275 8959
rect 4905 8789 4939 8823
rect 6469 8789 6503 8823
rect 7297 8789 7331 8823
rect 8677 8789 8711 8823
rect 4169 8585 4203 8619
rect 5089 8585 5123 8619
rect 6653 8585 6687 8619
rect 8493 8585 8527 8619
rect 10793 8585 10827 8619
rect 8217 8517 8251 8551
rect 8861 8517 8895 8551
rect 10425 8517 10459 8551
rect 1593 8449 1627 8483
rect 4721 8449 4755 8483
rect 5641 8449 5675 8483
rect 5825 8449 5859 8483
rect 1409 8381 1443 8415
rect 2789 8381 2823 8415
rect 5549 8381 5583 8415
rect 6193 8381 6227 8415
rect 6837 8381 6871 8415
rect 7093 8381 7127 8415
rect 9045 8381 9079 8415
rect 9301 8381 9335 8415
rect 2697 8313 2731 8347
rect 3034 8313 3068 8347
rect 2237 8245 2271 8279
rect 5181 8245 5215 8279
rect 11161 8245 11195 8279
rect 2237 8041 2271 8075
rect 6101 8041 6135 8075
rect 7757 8041 7791 8075
rect 6009 7973 6043 8007
rect 7205 7905 7239 7939
rect 11428 7905 11462 7939
rect 4629 7837 4663 7871
rect 6193 7837 6227 7871
rect 6837 7837 6871 7871
rect 9045 7837 9079 7871
rect 11161 7837 11195 7871
rect 5273 7769 5307 7803
rect 1685 7701 1719 7735
rect 2881 7701 2915 7735
rect 5641 7701 5675 7735
rect 7389 7701 7423 7735
rect 8125 7701 8159 7735
rect 12541 7701 12575 7735
rect 2145 7497 2179 7531
rect 2605 7497 2639 7531
rect 4537 7497 4571 7531
rect 4905 7497 4939 7531
rect 6101 7497 6135 7531
rect 7205 7497 7239 7531
rect 8677 7497 8711 7531
rect 11253 7497 11287 7531
rect 3341 7429 3375 7463
rect 4997 7429 5031 7463
rect 1593 7361 1627 7395
rect 4169 7361 4203 7395
rect 5457 7361 5491 7395
rect 5549 7361 5583 7395
rect 1409 7293 1443 7327
rect 2697 7293 2731 7327
rect 5365 7293 5399 7327
rect 7297 7293 7331 7327
rect 6653 7225 6687 7259
rect 7564 7225 7598 7259
rect 2881 7157 2915 7191
rect 8953 7157 8987 7191
rect 11621 7157 11655 7191
rect 4905 6953 4939 6987
rect 5733 6953 5767 6987
rect 12357 6953 12391 6987
rect 1409 6817 1443 6851
rect 2697 6817 2731 6851
rect 4997 6817 5031 6851
rect 6101 6817 6135 6851
rect 6929 6817 6963 6851
rect 7665 6817 7699 6851
rect 9045 6817 9079 6851
rect 9689 6817 9723 6851
rect 10977 6817 11011 6851
rect 11233 6817 11267 6851
rect 1593 6749 1627 6783
rect 7757 6749 7791 6783
rect 7849 6749 7883 6783
rect 8125 6749 8159 6783
rect 8677 6749 8711 6783
rect 7297 6681 7331 6715
rect 9413 6681 9447 6715
rect 10241 6681 10275 6715
rect 2421 6613 2455 6647
rect 2881 6613 2915 6647
rect 3341 6613 3375 6647
rect 3893 6613 3927 6647
rect 4353 6613 4387 6647
rect 5181 6613 5215 6647
rect 6285 6613 6319 6647
rect 8125 6613 8159 6647
rect 8309 6613 8343 6647
rect 9873 6613 9907 6647
rect 2053 6409 2087 6443
rect 5181 6409 5215 6443
rect 5549 6409 5583 6443
rect 6837 6409 6871 6443
rect 9045 6409 9079 6443
rect 9781 6409 9815 6443
rect 11621 6409 11655 6443
rect 4721 6341 4755 6375
rect 6285 6341 6319 6375
rect 7297 6273 7331 6307
rect 7481 6273 7515 6307
rect 9965 6273 9999 6307
rect 2145 6205 2179 6239
rect 4537 6205 4571 6239
rect 5641 6205 5675 6239
rect 7205 6205 7239 6239
rect 8401 6205 8435 6239
rect 2390 6137 2424 6171
rect 9413 6137 9447 6171
rect 10210 6137 10244 6171
rect 1685 6069 1719 6103
rect 3525 6069 3559 6103
rect 4077 6069 4111 6103
rect 4353 6069 4387 6103
rect 5825 6069 5859 6103
rect 6653 6069 6687 6103
rect 7849 6069 7883 6103
rect 8309 6069 8343 6103
rect 8585 6069 8619 6103
rect 11345 6069 11379 6103
rect 12081 6069 12115 6103
rect 2421 5865 2455 5899
rect 2789 5865 2823 5899
rect 6653 5865 6687 5899
rect 7849 5865 7883 5899
rect 8309 5865 8343 5899
rect 8953 5865 8987 5899
rect 11069 5865 11103 5899
rect 11437 5865 11471 5899
rect 8217 5797 8251 5831
rect 9956 5797 9990 5831
rect 2881 5729 2915 5763
rect 3893 5729 3927 5763
rect 4344 5729 4378 5763
rect 6193 5729 6227 5763
rect 9689 5729 9723 5763
rect 3065 5661 3099 5695
rect 4077 5661 4111 5695
rect 5825 5661 5859 5695
rect 6745 5661 6779 5695
rect 6929 5661 6963 5695
rect 8401 5661 8435 5695
rect 6285 5593 6319 5627
rect 1869 5525 1903 5559
rect 2237 5525 2271 5559
rect 3525 5525 3559 5559
rect 5457 5525 5491 5559
rect 7297 5525 7331 5559
rect 7757 5525 7791 5559
rect 9505 5525 9539 5559
rect 1961 5321 1995 5355
rect 3065 5321 3099 5355
rect 4629 5321 4663 5355
rect 6193 5321 6227 5355
rect 6469 5321 6503 5355
rect 7941 5321 7975 5355
rect 8401 5321 8435 5355
rect 9781 5321 9815 5355
rect 10517 5321 10551 5355
rect 12081 5321 12115 5355
rect 1777 5253 1811 5287
rect 6377 5253 6411 5287
rect 2421 5185 2455 5219
rect 2605 5185 2639 5219
rect 3985 5185 4019 5219
rect 4169 5185 4203 5219
rect 5733 5185 5767 5219
rect 2329 5117 2363 5151
rect 3433 5117 3467 5151
rect 5457 5117 5491 5151
rect 6377 5117 6411 5151
rect 6561 5253 6595 5287
rect 7389 5185 7423 5219
rect 9045 5185 9079 5219
rect 10149 5185 10183 5219
rect 11253 5185 11287 5219
rect 7205 5117 7239 5151
rect 8769 5117 8803 5151
rect 10977 5117 11011 5151
rect 4997 5049 5031 5083
rect 6469 5049 6503 5083
rect 7297 5049 7331 5083
rect 11069 5049 11103 5083
rect 3525 4981 3559 5015
rect 3893 4981 3927 5015
rect 5089 4981 5123 5015
rect 5549 4981 5583 5015
rect 6837 4981 6871 5015
rect 8309 4981 8343 5015
rect 8861 4981 8895 5015
rect 10609 4981 10643 5015
rect 11621 4981 11655 5015
rect 12449 4981 12483 5015
rect 4353 4777 4387 4811
rect 4721 4777 4755 4811
rect 5733 4777 5767 4811
rect 7573 4777 7607 4811
rect 9045 4777 9079 4811
rect 10057 4777 10091 4811
rect 11069 4777 11103 4811
rect 11253 4777 11287 4811
rect 11621 4777 11655 4811
rect 12449 4777 12483 4811
rect 4813 4709 4847 4743
rect 1409 4641 1443 4675
rect 2697 4641 2731 4675
rect 3617 4641 3651 4675
rect 5457 4641 5491 4675
rect 6193 4641 6227 4675
rect 6460 4641 6494 4675
rect 8401 4641 8435 4675
rect 11713 4641 11747 4675
rect 12817 4641 12851 4675
rect 1593 4573 1627 4607
rect 4905 4573 4939 4607
rect 8309 4573 8343 4607
rect 10149 4573 10183 4607
rect 10241 4573 10275 4607
rect 11805 4573 11839 4607
rect 2881 4505 2915 4539
rect 9689 4505 9723 4539
rect 13001 4505 13035 4539
rect 2513 4437 2547 4471
rect 7941 4437 7975 4471
rect 8585 4437 8619 4471
rect 9505 4437 9539 4471
rect 10701 4437 10735 4471
rect 2053 4233 2087 4267
rect 3893 4233 3927 4267
rect 5273 4233 5307 4267
rect 7941 4233 7975 4267
rect 8953 4233 8987 4267
rect 9781 4233 9815 4267
rect 10057 4233 10091 4267
rect 13461 4233 13495 4267
rect 2329 4165 2363 4199
rect 3709 4165 3743 4199
rect 11253 4165 11287 4199
rect 4353 4097 4387 4131
rect 4537 4097 4571 4131
rect 7389 4097 7423 4131
rect 8493 4097 8527 4131
rect 9413 4097 9447 4131
rect 10609 4097 10643 4131
rect 12909 4097 12943 4131
rect 13001 4097 13035 4131
rect 2145 4029 2179 4063
rect 3433 4029 3467 4063
rect 4261 4029 4295 4063
rect 5457 4029 5491 4063
rect 6009 4029 6043 4063
rect 6837 4029 6871 4063
rect 8309 4029 8343 4063
rect 11805 4029 11839 4063
rect 12173 4029 12207 4063
rect 1685 3961 1719 3995
rect 7757 3961 7791 3995
rect 10425 3961 10459 3995
rect 2697 3893 2731 3927
rect 4997 3893 5031 3927
rect 5641 3893 5675 3927
rect 6377 3893 6411 3927
rect 7021 3893 7055 3927
rect 8401 3893 8435 3927
rect 10517 3893 10551 3927
rect 12449 3893 12483 3927
rect 12817 3893 12851 3927
rect 2421 3689 2455 3723
rect 2789 3689 2823 3723
rect 4077 3689 4111 3723
rect 5089 3689 5123 3723
rect 5549 3689 5583 3723
rect 6837 3689 6871 3723
rect 8033 3689 8067 3723
rect 9137 3689 9171 3723
rect 10149 3689 10183 3723
rect 11161 3689 11195 3723
rect 11713 3689 11747 3723
rect 12081 3689 12115 3723
rect 2329 3621 2363 3655
rect 4445 3621 4479 3655
rect 5825 3621 5859 3655
rect 6929 3621 6963 3655
rect 8493 3621 8527 3655
rect 10609 3621 10643 3655
rect 4537 3553 4571 3587
rect 8401 3553 8435 3587
rect 10517 3553 10551 3587
rect 11529 3553 11563 3587
rect 13277 3553 13311 3587
rect 2881 3485 2915 3519
rect 3065 3485 3099 3519
rect 4721 3485 4755 3519
rect 7021 3485 7055 3519
rect 8677 3485 8711 3519
rect 10057 3485 10091 3519
rect 10793 3485 10827 3519
rect 12173 3485 12207 3519
rect 12265 3485 12299 3519
rect 12725 3485 12759 3519
rect 3525 3417 3559 3451
rect 3893 3417 3927 3451
rect 6469 3417 6503 3451
rect 7573 3417 7607 3451
rect 7941 3417 7975 3451
rect 9505 3417 9539 3451
rect 13461 3417 13495 3451
rect 1961 3349 1995 3383
rect 6285 3349 6319 3383
rect 13093 3349 13127 3383
rect 3341 3145 3375 3179
rect 3709 3145 3743 3179
rect 4077 3145 4111 3179
rect 5549 3145 5583 3179
rect 6193 3145 6227 3179
rect 7665 3145 7699 3179
rect 8033 3145 8067 3179
rect 9597 3145 9631 3179
rect 9965 3145 9999 3179
rect 10241 3145 10275 3179
rect 11805 3145 11839 3179
rect 12449 3145 12483 3179
rect 13461 3145 13495 3179
rect 6469 3077 6503 3111
rect 10425 3077 10459 3111
rect 10977 3009 11011 3043
rect 12173 3009 12207 3043
rect 12909 3009 12943 3043
rect 13001 3009 13035 3043
rect 1961 2941 1995 2975
rect 4169 2941 4203 2975
rect 6837 2941 6871 2975
rect 8217 2941 8251 2975
rect 10885 2941 10919 2975
rect 2228 2873 2262 2907
rect 4414 2873 4448 2907
rect 8462 2873 8496 2907
rect 10793 2873 10827 2907
rect 12817 2873 12851 2907
rect 13829 2873 13863 2907
rect 1869 2805 1903 2839
rect 7021 2805 7055 2839
rect 2421 2601 2455 2635
rect 4077 2601 4111 2635
rect 4445 2601 4479 2635
rect 8125 2601 8159 2635
rect 8493 2601 8527 2635
rect 10057 2601 10091 2635
rect 11069 2601 11103 2635
rect 11437 2601 11471 2635
rect 11897 2601 11931 2635
rect 3525 2533 3559 2567
rect 5549 2533 5583 2567
rect 7665 2533 7699 2567
rect 8585 2533 8619 2567
rect 9229 2533 9263 2567
rect 10425 2533 10459 2567
rect 12173 2533 12207 2567
rect 1409 2465 1443 2499
rect 1961 2465 1995 2499
rect 2789 2465 2823 2499
rect 5181 2465 5215 2499
rect 5641 2465 5675 2499
rect 6469 2465 6503 2499
rect 6929 2465 6963 2499
rect 8033 2465 8067 2499
rect 9597 2465 9631 2499
rect 10517 2465 10551 2499
rect 12633 2465 12667 2499
rect 13185 2465 13219 2499
rect 2329 2397 2363 2431
rect 2881 2397 2915 2431
rect 2973 2397 3007 2431
rect 3893 2397 3927 2431
rect 4537 2397 4571 2431
rect 4629 2397 4663 2431
rect 8677 2397 8711 2431
rect 10701 2397 10735 2431
rect 5825 2329 5859 2363
rect 12817 2329 12851 2363
rect 7113 2261 7147 2295
<< metal1 >>
rect 11146 37680 11152 37732
rect 11204 37720 11210 37732
rect 11790 37720 11796 37732
rect 11204 37692 11796 37720
rect 11204 37680 11210 37692
rect 11790 37680 11796 37692
rect 11848 37680 11854 37732
rect 1104 37562 14812 37584
rect 1104 37510 6315 37562
rect 6367 37510 6379 37562
rect 6431 37510 6443 37562
rect 6495 37510 6507 37562
rect 6559 37510 11648 37562
rect 11700 37510 11712 37562
rect 11764 37510 11776 37562
rect 11828 37510 11840 37562
rect 11892 37510 14812 37562
rect 1104 37488 14812 37510
rect 1104 37018 14812 37040
rect 1104 36966 3648 37018
rect 3700 36966 3712 37018
rect 3764 36966 3776 37018
rect 3828 36966 3840 37018
rect 3892 36966 8982 37018
rect 9034 36966 9046 37018
rect 9098 36966 9110 37018
rect 9162 36966 9174 37018
rect 9226 36966 14315 37018
rect 14367 36966 14379 37018
rect 14431 36966 14443 37018
rect 14495 36966 14507 37018
rect 14559 36966 14812 37018
rect 1104 36944 14812 36966
rect 4522 36864 4528 36916
rect 4580 36904 4586 36916
rect 4801 36907 4859 36913
rect 4801 36904 4813 36907
rect 4580 36876 4813 36904
rect 4580 36864 4586 36876
rect 4801 36873 4813 36876
rect 4847 36873 4859 36907
rect 4801 36867 4859 36873
rect 4617 36703 4675 36709
rect 4617 36669 4629 36703
rect 4663 36700 4675 36703
rect 4663 36672 5304 36700
rect 4663 36669 4675 36672
rect 4617 36663 4675 36669
rect 5276 36573 5304 36672
rect 5261 36567 5319 36573
rect 5261 36533 5273 36567
rect 5307 36564 5319 36567
rect 7926 36564 7932 36576
rect 5307 36536 7932 36564
rect 5307 36533 5319 36536
rect 5261 36527 5319 36533
rect 7926 36524 7932 36536
rect 7984 36524 7990 36576
rect 1104 36474 14812 36496
rect 1104 36422 6315 36474
rect 6367 36422 6379 36474
rect 6431 36422 6443 36474
rect 6495 36422 6507 36474
rect 6559 36422 11648 36474
rect 11700 36422 11712 36474
rect 11764 36422 11776 36474
rect 11828 36422 11840 36474
rect 11892 36422 14812 36474
rect 1104 36400 14812 36422
rect 4982 36360 4988 36372
rect 4943 36332 4988 36360
rect 4982 36320 4988 36332
rect 5040 36320 5046 36372
rect 6178 36320 6184 36372
rect 6236 36360 6242 36372
rect 6549 36363 6607 36369
rect 6549 36360 6561 36363
rect 6236 36332 6561 36360
rect 6236 36320 6242 36332
rect 6549 36329 6561 36332
rect 6595 36329 6607 36363
rect 6549 36323 6607 36329
rect 4801 36227 4859 36233
rect 4801 36193 4813 36227
rect 4847 36224 4859 36227
rect 5074 36224 5080 36236
rect 4847 36196 5080 36224
rect 4847 36193 4859 36196
rect 4801 36187 4859 36193
rect 5074 36184 5080 36196
rect 5132 36184 5138 36236
rect 6365 36227 6423 36233
rect 6365 36193 6377 36227
rect 6411 36224 6423 36227
rect 6730 36224 6736 36236
rect 6411 36196 6736 36224
rect 6411 36193 6423 36196
rect 6365 36187 6423 36193
rect 6730 36184 6736 36196
rect 6788 36184 6794 36236
rect 1104 35930 14812 35952
rect 1104 35878 3648 35930
rect 3700 35878 3712 35930
rect 3764 35878 3776 35930
rect 3828 35878 3840 35930
rect 3892 35878 8982 35930
rect 9034 35878 9046 35930
rect 9098 35878 9110 35930
rect 9162 35878 9174 35930
rect 9226 35878 14315 35930
rect 14367 35878 14379 35930
rect 14431 35878 14443 35930
rect 14495 35878 14507 35930
rect 14559 35878 14812 35930
rect 1104 35856 14812 35878
rect 4709 35819 4767 35825
rect 4709 35785 4721 35819
rect 4755 35816 4767 35819
rect 5350 35816 5356 35828
rect 4755 35788 5356 35816
rect 4755 35785 4767 35788
rect 4709 35779 4767 35785
rect 5350 35776 5356 35788
rect 5408 35776 5414 35828
rect 5718 35776 5724 35828
rect 5776 35816 5782 35828
rect 5813 35819 5871 35825
rect 5813 35816 5825 35819
rect 5776 35788 5825 35816
rect 5776 35776 5782 35788
rect 5813 35785 5825 35788
rect 5859 35785 5871 35819
rect 5813 35779 5871 35785
rect 6914 35776 6920 35828
rect 6972 35816 6978 35828
rect 7285 35819 7343 35825
rect 7285 35816 7297 35819
rect 6972 35788 7297 35816
rect 6972 35776 6978 35788
rect 7285 35785 7297 35788
rect 7331 35785 7343 35819
rect 7285 35779 7343 35785
rect 7742 35776 7748 35828
rect 7800 35816 7806 35828
rect 8389 35819 8447 35825
rect 8389 35816 8401 35819
rect 7800 35788 8401 35816
rect 7800 35776 7806 35788
rect 8389 35785 8401 35788
rect 8435 35785 8447 35819
rect 8389 35779 8447 35785
rect 9858 35748 9864 35760
rect 9819 35720 9864 35748
rect 9858 35708 9864 35720
rect 9916 35708 9922 35760
rect 4525 35615 4583 35621
rect 4525 35581 4537 35615
rect 4571 35612 4583 35615
rect 5629 35615 5687 35621
rect 4571 35584 4605 35612
rect 4571 35581 4583 35584
rect 4525 35575 4583 35581
rect 5629 35581 5641 35615
rect 5675 35612 5687 35615
rect 7101 35615 7159 35621
rect 5675 35584 6224 35612
rect 5675 35581 5687 35584
rect 5629 35575 5687 35581
rect 4433 35547 4491 35553
rect 4433 35513 4445 35547
rect 4479 35544 4491 35547
rect 4540 35544 4568 35575
rect 4982 35544 4988 35556
rect 4479 35516 4988 35544
rect 4479 35513 4491 35516
rect 4433 35507 4491 35513
rect 4982 35504 4988 35516
rect 5040 35504 5046 35556
rect 6196 35488 6224 35584
rect 7101 35581 7113 35615
rect 7147 35612 7159 35615
rect 8205 35615 8263 35621
rect 7147 35584 7696 35612
rect 7147 35581 7159 35584
rect 7101 35575 7159 35581
rect 7668 35488 7696 35584
rect 8205 35581 8217 35615
rect 8251 35612 8263 35615
rect 9677 35615 9735 35621
rect 8251 35584 8892 35612
rect 8251 35581 8263 35584
rect 8205 35575 8263 35581
rect 8864 35488 8892 35584
rect 9677 35581 9689 35615
rect 9723 35612 9735 35615
rect 9723 35584 10088 35612
rect 9723 35581 9735 35584
rect 9677 35575 9735 35581
rect 10060 35488 10088 35584
rect 5074 35476 5080 35488
rect 5035 35448 5080 35476
rect 5074 35436 5080 35448
rect 5132 35436 5138 35488
rect 6178 35476 6184 35488
rect 6139 35448 6184 35476
rect 6178 35436 6184 35448
rect 6236 35436 6242 35488
rect 6641 35479 6699 35485
rect 6641 35445 6653 35479
rect 6687 35476 6699 35479
rect 6730 35476 6736 35488
rect 6687 35448 6736 35476
rect 6687 35445 6699 35448
rect 6641 35439 6699 35445
rect 6730 35436 6736 35448
rect 6788 35436 6794 35488
rect 7650 35476 7656 35488
rect 7611 35448 7656 35476
rect 7650 35436 7656 35448
rect 7708 35436 7714 35488
rect 7834 35436 7840 35488
rect 7892 35476 7898 35488
rect 8021 35479 8079 35485
rect 8021 35476 8033 35479
rect 7892 35448 8033 35476
rect 7892 35436 7898 35448
rect 8021 35445 8033 35448
rect 8067 35445 8079 35479
rect 8846 35476 8852 35488
rect 8807 35448 8852 35476
rect 8021 35439 8079 35445
rect 8846 35436 8852 35448
rect 8904 35436 8910 35488
rect 10042 35436 10048 35488
rect 10100 35476 10106 35488
rect 10229 35479 10287 35485
rect 10229 35476 10241 35479
rect 10100 35448 10241 35476
rect 10100 35436 10106 35448
rect 10229 35445 10241 35448
rect 10275 35445 10287 35479
rect 10229 35439 10287 35445
rect 1104 35386 14812 35408
rect 1104 35334 6315 35386
rect 6367 35334 6379 35386
rect 6431 35334 6443 35386
rect 6495 35334 6507 35386
rect 6559 35334 11648 35386
rect 11700 35334 11712 35386
rect 11764 35334 11776 35386
rect 11828 35334 11840 35386
rect 11892 35334 14812 35386
rect 1104 35312 14812 35334
rect 566 35232 572 35284
rect 624 35272 630 35284
rect 1581 35275 1639 35281
rect 1581 35272 1593 35275
rect 624 35244 1593 35272
rect 624 35232 630 35244
rect 1581 35241 1593 35244
rect 1627 35241 1639 35275
rect 4246 35272 4252 35284
rect 4207 35244 4252 35272
rect 1581 35235 1639 35241
rect 4246 35232 4252 35244
rect 4304 35232 4310 35284
rect 5629 35275 5687 35281
rect 5629 35241 5641 35275
rect 5675 35272 5687 35275
rect 6638 35272 6644 35284
rect 5675 35244 6644 35272
rect 5675 35241 5687 35244
rect 5629 35235 5687 35241
rect 6638 35232 6644 35244
rect 6696 35232 6702 35284
rect 7374 35232 7380 35284
rect 7432 35272 7438 35284
rect 8297 35275 8355 35281
rect 8297 35272 8309 35275
rect 7432 35244 8309 35272
rect 7432 35232 7438 35244
rect 8297 35241 8309 35244
rect 8343 35241 8355 35275
rect 8297 35235 8355 35241
rect 9766 35232 9772 35284
rect 9824 35272 9830 35284
rect 10594 35272 10600 35284
rect 9824 35244 10600 35272
rect 9824 35232 9830 35244
rect 10594 35232 10600 35244
rect 10652 35232 10658 35284
rect 1397 35139 1455 35145
rect 1397 35105 1409 35139
rect 1443 35136 1455 35139
rect 1946 35136 1952 35148
rect 1443 35108 1952 35136
rect 1443 35105 1455 35108
rect 1397 35099 1455 35105
rect 1946 35096 1952 35108
rect 2004 35096 2010 35148
rect 2498 35136 2504 35148
rect 2459 35108 2504 35136
rect 2498 35096 2504 35108
rect 2556 35096 2562 35148
rect 4062 35136 4068 35148
rect 4023 35108 4068 35136
rect 4062 35096 4068 35108
rect 4120 35096 4126 35148
rect 5442 35136 5448 35148
rect 5403 35108 5448 35136
rect 5442 35096 5448 35108
rect 5500 35096 5506 35148
rect 6914 35136 6920 35148
rect 6875 35108 6920 35136
rect 6914 35096 6920 35108
rect 6972 35096 6978 35148
rect 7374 35096 7380 35148
rect 7432 35136 7438 35148
rect 8113 35139 8171 35145
rect 8113 35136 8125 35139
rect 7432 35108 8125 35136
rect 7432 35096 7438 35108
rect 8113 35105 8125 35108
rect 8159 35105 8171 35139
rect 8113 35099 8171 35105
rect 9306 35096 9312 35148
rect 9364 35136 9370 35148
rect 10045 35139 10103 35145
rect 10045 35136 10057 35139
rect 9364 35108 10057 35136
rect 9364 35096 9370 35108
rect 10045 35105 10057 35108
rect 10091 35105 10103 35139
rect 10045 35099 10103 35105
rect 7006 35068 7012 35080
rect 6967 35040 7012 35068
rect 7006 35028 7012 35040
rect 7064 35028 7070 35080
rect 7193 35071 7251 35077
rect 7193 35037 7205 35071
rect 7239 35068 7251 35071
rect 7239 35040 7788 35068
rect 7239 35037 7251 35040
rect 7193 35031 7251 35037
rect 1394 34960 1400 35012
rect 1452 35000 1458 35012
rect 2685 35003 2743 35009
rect 2685 35000 2697 35003
rect 1452 34972 2697 35000
rect 1452 34960 1458 34972
rect 2685 34969 2697 34972
rect 2731 34969 2743 35003
rect 2685 34963 2743 34969
rect 7760 34944 7788 35040
rect 9766 35028 9772 35080
rect 9824 35068 9830 35080
rect 10137 35071 10195 35077
rect 10137 35068 10149 35071
rect 9824 35040 10149 35068
rect 9824 35028 9830 35040
rect 10137 35037 10149 35040
rect 10183 35037 10195 35071
rect 10137 35031 10195 35037
rect 10229 35071 10287 35077
rect 10229 35037 10241 35071
rect 10275 35037 10287 35071
rect 10229 35031 10287 35037
rect 9858 34960 9864 35012
rect 9916 35000 9922 35012
rect 10244 35000 10272 35031
rect 9916 34972 10272 35000
rect 9916 34960 9922 34972
rect 2038 34932 2044 34944
rect 1999 34904 2044 34932
rect 2038 34892 2044 34904
rect 2096 34892 2102 34944
rect 5718 34892 5724 34944
rect 5776 34932 5782 34944
rect 6549 34935 6607 34941
rect 6549 34932 6561 34935
rect 5776 34904 6561 34932
rect 5776 34892 5782 34904
rect 6549 34901 6561 34904
rect 6595 34901 6607 34935
rect 7742 34932 7748 34944
rect 7703 34904 7748 34932
rect 6549 34895 6607 34901
rect 7742 34892 7748 34904
rect 7800 34892 7806 34944
rect 9677 34935 9735 34941
rect 9677 34901 9689 34935
rect 9723 34932 9735 34935
rect 10134 34932 10140 34944
rect 9723 34904 10140 34932
rect 9723 34901 9735 34904
rect 9677 34895 9735 34901
rect 10134 34892 10140 34904
rect 10192 34892 10198 34944
rect 10226 34892 10232 34944
rect 10284 34932 10290 34944
rect 10689 34935 10747 34941
rect 10689 34932 10701 34935
rect 10284 34904 10701 34932
rect 10284 34892 10290 34904
rect 10689 34901 10701 34904
rect 10735 34901 10747 34935
rect 10689 34895 10747 34901
rect 1104 34842 14812 34864
rect 1104 34790 3648 34842
rect 3700 34790 3712 34842
rect 3764 34790 3776 34842
rect 3828 34790 3840 34842
rect 3892 34790 8982 34842
rect 9034 34790 9046 34842
rect 9098 34790 9110 34842
rect 9162 34790 9174 34842
rect 9226 34790 14315 34842
rect 14367 34790 14379 34842
rect 14431 34790 14443 34842
rect 14495 34790 14507 34842
rect 14559 34790 14812 34842
rect 1104 34768 14812 34790
rect 1946 34688 1952 34740
rect 2004 34728 2010 34740
rect 2133 34731 2191 34737
rect 2133 34728 2145 34731
rect 2004 34700 2145 34728
rect 2004 34688 2010 34700
rect 2133 34697 2145 34700
rect 2179 34697 2191 34731
rect 2498 34728 2504 34740
rect 2459 34700 2504 34728
rect 2133 34691 2191 34697
rect 2498 34688 2504 34700
rect 2556 34688 2562 34740
rect 3234 34728 3240 34740
rect 3195 34700 3240 34728
rect 3234 34688 3240 34700
rect 3292 34688 3298 34740
rect 4338 34728 4344 34740
rect 4299 34700 4344 34728
rect 4338 34688 4344 34700
rect 4396 34688 4402 34740
rect 6273 34731 6331 34737
rect 6273 34697 6285 34731
rect 6319 34728 6331 34731
rect 6914 34728 6920 34740
rect 6319 34700 6920 34728
rect 6319 34697 6331 34700
rect 6273 34691 6331 34697
rect 6914 34688 6920 34700
rect 6972 34728 6978 34740
rect 8294 34728 8300 34740
rect 6972 34700 8300 34728
rect 6972 34688 6978 34700
rect 8294 34688 8300 34700
rect 8352 34688 8358 34740
rect 9766 34728 9772 34740
rect 9727 34700 9772 34728
rect 9766 34688 9772 34700
rect 9824 34688 9830 34740
rect 3694 34660 3700 34672
rect 3068 34632 3700 34660
rect 1578 34592 1584 34604
rect 1539 34564 1584 34592
rect 1578 34552 1584 34564
rect 1636 34552 1642 34604
rect 2038 34592 2044 34604
rect 1688 34564 2044 34592
rect 1397 34527 1455 34533
rect 1397 34493 1409 34527
rect 1443 34524 1455 34527
rect 1688 34524 1716 34564
rect 2038 34552 2044 34564
rect 2096 34552 2102 34604
rect 1443 34496 1716 34524
rect 1443 34493 1455 34496
rect 1397 34487 1455 34493
rect 1762 34484 1768 34536
rect 1820 34524 1826 34536
rect 3068 34533 3096 34632
rect 3694 34620 3700 34632
rect 3752 34620 3758 34672
rect 3970 34620 3976 34672
rect 4028 34660 4034 34672
rect 5445 34663 5503 34669
rect 5445 34660 5457 34663
rect 4028 34632 5457 34660
rect 4028 34620 4034 34632
rect 5445 34629 5457 34632
rect 5491 34629 5503 34663
rect 5445 34623 5503 34629
rect 9033 34663 9091 34669
rect 9033 34629 9045 34663
rect 9079 34660 9091 34663
rect 9858 34660 9864 34672
rect 9079 34632 9864 34660
rect 9079 34629 9091 34632
rect 9033 34623 9091 34629
rect 9858 34620 9864 34632
rect 9916 34620 9922 34672
rect 3326 34552 3332 34604
rect 3384 34592 3390 34604
rect 4338 34592 4344 34604
rect 3384 34564 4344 34592
rect 3384 34552 3390 34564
rect 4338 34552 4344 34564
rect 4396 34552 4402 34604
rect 6641 34595 6699 34601
rect 6641 34561 6653 34595
rect 6687 34592 6699 34595
rect 9876 34592 9904 34620
rect 6687 34564 7788 34592
rect 9876 34564 9996 34592
rect 6687 34561 6699 34564
rect 6641 34555 6699 34561
rect 7760 34536 7788 34564
rect 3053 34527 3111 34533
rect 1820 34496 2820 34524
rect 1820 34484 1826 34496
rect 2792 34468 2820 34496
rect 3053 34493 3065 34527
rect 3099 34493 3111 34527
rect 4062 34524 4068 34536
rect 4023 34496 4068 34524
rect 3053 34487 3111 34493
rect 4062 34484 4068 34496
rect 4120 34484 4126 34536
rect 4157 34527 4215 34533
rect 4157 34493 4169 34527
rect 4203 34524 4215 34527
rect 4246 34524 4252 34536
rect 4203 34496 4252 34524
rect 4203 34493 4215 34496
rect 4157 34487 4215 34493
rect 4246 34484 4252 34496
rect 4304 34524 4310 34536
rect 4709 34527 4767 34533
rect 4709 34524 4721 34527
rect 4304 34496 4721 34524
rect 4304 34484 4310 34496
rect 4709 34493 4721 34496
rect 4755 34493 4767 34527
rect 4709 34487 4767 34493
rect 5261 34527 5319 34533
rect 5261 34493 5273 34527
rect 5307 34493 5319 34527
rect 5261 34487 5319 34493
rect 2774 34416 2780 34468
rect 2832 34416 2838 34468
rect 5276 34400 5304 34487
rect 5442 34484 5448 34536
rect 5500 34524 5506 34536
rect 5813 34527 5871 34533
rect 5813 34524 5825 34527
rect 5500 34496 5825 34524
rect 5500 34484 5506 34496
rect 5813 34493 5825 34496
rect 5859 34493 5871 34527
rect 7006 34524 7012 34536
rect 6967 34496 7012 34524
rect 5813 34487 5871 34493
rect 7006 34484 7012 34496
rect 7064 34484 7070 34536
rect 7374 34484 7380 34536
rect 7432 34524 7438 34536
rect 7469 34527 7527 34533
rect 7469 34524 7481 34527
rect 7432 34496 7481 34524
rect 7432 34484 7438 34496
rect 7469 34493 7481 34496
rect 7515 34493 7527 34527
rect 7469 34487 7527 34493
rect 7653 34527 7711 34533
rect 7653 34493 7665 34527
rect 7699 34493 7711 34527
rect 7653 34487 7711 34493
rect 7668 34456 7696 34487
rect 7742 34484 7748 34536
rect 7800 34524 7806 34536
rect 7920 34527 7978 34533
rect 7920 34524 7932 34527
rect 7800 34496 7932 34524
rect 7800 34484 7806 34496
rect 7920 34493 7932 34496
rect 7966 34524 7978 34527
rect 9861 34527 9919 34533
rect 7966 34496 8340 34524
rect 7966 34493 7978 34496
rect 7920 34487 7978 34493
rect 7834 34456 7840 34468
rect 7668 34428 7840 34456
rect 7834 34416 7840 34428
rect 7892 34456 7898 34468
rect 8110 34456 8116 34468
rect 7892 34428 8116 34456
rect 7892 34416 7898 34428
rect 8110 34416 8116 34428
rect 8168 34416 8174 34468
rect 8312 34456 8340 34496
rect 9861 34493 9873 34527
rect 9907 34493 9919 34527
rect 9968 34524 9996 34564
rect 10117 34527 10175 34533
rect 10117 34524 10129 34527
rect 9968 34496 10129 34524
rect 9861 34487 9919 34493
rect 10117 34493 10129 34496
rect 10163 34493 10175 34527
rect 10117 34487 10175 34493
rect 8754 34456 8760 34468
rect 8312 34428 8760 34456
rect 8754 34416 8760 34428
rect 8812 34416 8818 34468
rect 9876 34456 9904 34487
rect 10226 34456 10232 34468
rect 9876 34428 10232 34456
rect 10226 34416 10232 34428
rect 10284 34416 10290 34468
rect 5169 34391 5227 34397
rect 5169 34357 5181 34391
rect 5215 34388 5227 34391
rect 5258 34388 5264 34400
rect 5215 34360 5264 34388
rect 5215 34357 5227 34360
rect 5169 34351 5227 34357
rect 5258 34348 5264 34360
rect 5316 34348 5322 34400
rect 7742 34348 7748 34400
rect 7800 34388 7806 34400
rect 8202 34388 8208 34400
rect 7800 34360 8208 34388
rect 7800 34348 7806 34360
rect 8202 34348 8208 34360
rect 8260 34388 8266 34400
rect 9306 34388 9312 34400
rect 8260 34360 9312 34388
rect 8260 34348 8266 34360
rect 9306 34348 9312 34360
rect 9364 34348 9370 34400
rect 11241 34391 11299 34397
rect 11241 34357 11253 34391
rect 11287 34388 11299 34391
rect 12158 34388 12164 34400
rect 11287 34360 12164 34388
rect 11287 34357 11299 34360
rect 11241 34351 11299 34357
rect 12158 34348 12164 34360
rect 12216 34348 12222 34400
rect 1104 34298 14812 34320
rect 1104 34246 6315 34298
rect 6367 34246 6379 34298
rect 6431 34246 6443 34298
rect 6495 34246 6507 34298
rect 6559 34246 11648 34298
rect 11700 34246 11712 34298
rect 11764 34246 11776 34298
rect 11828 34246 11840 34298
rect 11892 34246 14812 34298
rect 1104 34224 14812 34246
rect 2774 34144 2780 34196
rect 2832 34184 2838 34196
rect 2869 34187 2927 34193
rect 2869 34184 2881 34187
rect 2832 34156 2881 34184
rect 2832 34144 2838 34156
rect 2869 34153 2881 34156
rect 2915 34153 2927 34187
rect 2869 34147 2927 34153
rect 4249 34187 4307 34193
rect 4249 34153 4261 34187
rect 4295 34184 4307 34187
rect 4338 34184 4344 34196
rect 4295 34156 4344 34184
rect 4295 34153 4307 34156
rect 4249 34147 4307 34153
rect 4338 34144 4344 34156
rect 4396 34144 4402 34196
rect 5994 34184 6000 34196
rect 5955 34156 6000 34184
rect 5994 34144 6000 34156
rect 6052 34144 6058 34196
rect 8754 34184 8760 34196
rect 8715 34156 8760 34184
rect 8754 34144 8760 34156
rect 8812 34144 8818 34196
rect 9858 34184 9864 34196
rect 9819 34156 9864 34184
rect 9858 34144 9864 34156
rect 9916 34184 9922 34196
rect 10229 34187 10287 34193
rect 10229 34184 10241 34187
rect 9916 34156 10241 34184
rect 9916 34144 9922 34156
rect 10229 34153 10241 34156
rect 10275 34153 10287 34187
rect 10229 34147 10287 34153
rect 1486 34076 1492 34128
rect 1544 34116 1550 34128
rect 1673 34119 1731 34125
rect 1673 34116 1685 34119
rect 1544 34088 1685 34116
rect 1544 34076 1550 34088
rect 1673 34085 1685 34088
rect 1719 34085 1731 34119
rect 5902 34116 5908 34128
rect 5863 34088 5908 34116
rect 1673 34079 1731 34085
rect 5902 34076 5908 34088
rect 5960 34076 5966 34128
rect 7558 34076 7564 34128
rect 7616 34125 7622 34128
rect 7616 34119 7680 34125
rect 7616 34085 7634 34119
rect 7668 34085 7680 34119
rect 7616 34079 7680 34085
rect 7616 34076 7622 34079
rect 12434 34076 12440 34128
rect 12492 34116 12498 34128
rect 12710 34116 12716 34128
rect 12492 34088 12716 34116
rect 12492 34076 12498 34088
rect 12710 34076 12716 34088
rect 12768 34076 12774 34128
rect 1397 34051 1455 34057
rect 1397 34017 1409 34051
rect 1443 34048 1455 34051
rect 2406 34048 2412 34060
rect 1443 34020 2412 34048
rect 1443 34017 1455 34020
rect 1397 34011 1455 34017
rect 2406 34008 2412 34020
rect 2464 34008 2470 34060
rect 2685 34051 2743 34057
rect 2685 34017 2697 34051
rect 2731 34048 2743 34051
rect 3050 34048 3056 34060
rect 2731 34020 3056 34048
rect 2731 34017 2743 34020
rect 2685 34011 2743 34017
rect 3050 34008 3056 34020
rect 3108 34008 3114 34060
rect 3970 34008 3976 34060
rect 4028 34048 4034 34060
rect 4065 34051 4123 34057
rect 4065 34048 4077 34051
rect 4028 34020 4077 34048
rect 4028 34008 4034 34020
rect 4065 34017 4077 34020
rect 4111 34017 4123 34051
rect 4065 34011 4123 34017
rect 7377 34051 7435 34057
rect 7377 34017 7389 34051
rect 7423 34048 7435 34051
rect 8110 34048 8116 34060
rect 7423 34020 8116 34048
rect 7423 34017 7435 34020
rect 7377 34011 7435 34017
rect 8110 34008 8116 34020
rect 8168 34008 8174 34060
rect 10778 34048 10784 34060
rect 10739 34020 10784 34048
rect 10778 34008 10784 34020
rect 10836 34008 10842 34060
rect 12342 34048 12348 34060
rect 12303 34020 12348 34048
rect 12342 34008 12348 34020
rect 12400 34008 12406 34060
rect 6086 33980 6092 33992
rect 6047 33952 6092 33980
rect 6086 33940 6092 33952
rect 6144 33940 6150 33992
rect 10870 33980 10876 33992
rect 10831 33952 10876 33980
rect 10870 33940 10876 33952
rect 10928 33940 10934 33992
rect 10965 33983 11023 33989
rect 10965 33949 10977 33983
rect 11011 33949 11023 33983
rect 10965 33943 11023 33949
rect 5537 33915 5595 33921
rect 5537 33881 5549 33915
rect 5583 33912 5595 33915
rect 7193 33915 7251 33921
rect 7193 33912 7205 33915
rect 5583 33884 7205 33912
rect 5583 33881 5595 33884
rect 5537 33875 5595 33881
rect 7193 33881 7205 33884
rect 7239 33912 7251 33915
rect 7282 33912 7288 33924
rect 7239 33884 7288 33912
rect 7239 33881 7251 33884
rect 7193 33875 7251 33881
rect 7282 33872 7288 33884
rect 7340 33872 7346 33924
rect 10686 33872 10692 33924
rect 10744 33912 10750 33924
rect 10980 33912 11008 33943
rect 11422 33940 11428 33992
rect 11480 33980 11486 33992
rect 12250 33980 12256 33992
rect 11480 33952 12256 33980
rect 11480 33940 11486 33952
rect 12250 33940 12256 33952
rect 12308 33980 12314 33992
rect 12437 33983 12495 33989
rect 12437 33980 12449 33983
rect 12308 33952 12449 33980
rect 12308 33940 12314 33952
rect 12437 33949 12449 33952
rect 12483 33949 12495 33983
rect 12437 33943 12495 33949
rect 12529 33983 12587 33989
rect 12529 33949 12541 33983
rect 12575 33949 12587 33983
rect 12529 33943 12587 33949
rect 12544 33912 12572 33943
rect 10744 33884 11008 33912
rect 12268 33884 12572 33912
rect 10744 33872 10750 33884
rect 12268 33856 12296 33884
rect 5445 33847 5503 33853
rect 5445 33813 5457 33847
rect 5491 33844 5503 33847
rect 5626 33844 5632 33856
rect 5491 33816 5632 33844
rect 5491 33813 5503 33816
rect 5445 33807 5503 33813
rect 5626 33804 5632 33816
rect 5684 33844 5690 33856
rect 6086 33844 6092 33856
rect 5684 33816 6092 33844
rect 5684 33804 5690 33816
rect 6086 33804 6092 33816
rect 6144 33804 6150 33856
rect 6917 33847 6975 33853
rect 6917 33813 6929 33847
rect 6963 33844 6975 33847
rect 7098 33844 7104 33856
rect 6963 33816 7104 33844
rect 6963 33813 6975 33816
rect 6917 33807 6975 33813
rect 7098 33804 7104 33816
rect 7156 33804 7162 33856
rect 9398 33844 9404 33856
rect 9359 33816 9404 33844
rect 9398 33804 9404 33816
rect 9456 33804 9462 33856
rect 9674 33804 9680 33856
rect 9732 33844 9738 33856
rect 10413 33847 10471 33853
rect 10413 33844 10425 33847
rect 9732 33816 10425 33844
rect 9732 33804 9738 33816
rect 10413 33813 10425 33816
rect 10459 33813 10471 33847
rect 10413 33807 10471 33813
rect 10778 33804 10784 33856
rect 10836 33844 10842 33856
rect 11977 33847 12035 33853
rect 11977 33844 11989 33847
rect 10836 33816 11989 33844
rect 10836 33804 10842 33816
rect 11977 33813 11989 33816
rect 12023 33813 12035 33847
rect 11977 33807 12035 33813
rect 12250 33804 12256 33856
rect 12308 33804 12314 33856
rect 1104 33754 14812 33776
rect 1104 33702 3648 33754
rect 3700 33702 3712 33754
rect 3764 33702 3776 33754
rect 3828 33702 3840 33754
rect 3892 33702 8982 33754
rect 9034 33702 9046 33754
rect 9098 33702 9110 33754
rect 9162 33702 9174 33754
rect 9226 33702 14315 33754
rect 14367 33702 14379 33754
rect 14431 33702 14443 33754
rect 14495 33702 14507 33754
rect 14559 33702 14812 33754
rect 1104 33680 14812 33702
rect 934 33600 940 33652
rect 992 33640 998 33652
rect 1581 33643 1639 33649
rect 1581 33640 1593 33643
rect 992 33612 1593 33640
rect 992 33600 998 33612
rect 1581 33609 1593 33612
rect 1627 33609 1639 33643
rect 1581 33603 1639 33609
rect 5905 33643 5963 33649
rect 5905 33609 5917 33643
rect 5951 33640 5963 33643
rect 5994 33640 6000 33652
rect 5951 33612 6000 33640
rect 5951 33609 5963 33612
rect 5905 33603 5963 33609
rect 5994 33600 6000 33612
rect 6052 33600 6058 33652
rect 6546 33640 6552 33652
rect 6507 33612 6552 33640
rect 6546 33600 6552 33612
rect 6604 33600 6610 33652
rect 12069 33643 12127 33649
rect 12069 33609 12081 33643
rect 12115 33640 12127 33643
rect 12115 33612 12848 33640
rect 12115 33609 12127 33612
rect 12069 33603 12127 33609
rect 2406 33572 2412 33584
rect 2367 33544 2412 33572
rect 2406 33532 2412 33544
rect 2464 33532 2470 33584
rect 7098 33532 7104 33584
rect 7156 33572 7162 33584
rect 9306 33572 9312 33584
rect 7156 33544 7512 33572
rect 9267 33544 9312 33572
rect 7156 33532 7162 33544
rect 5902 33464 5908 33516
rect 5960 33504 5966 33516
rect 6181 33507 6239 33513
rect 6181 33504 6193 33507
rect 5960 33476 6193 33504
rect 5960 33464 5966 33476
rect 6181 33473 6193 33476
rect 6227 33473 6239 33507
rect 7282 33504 7288 33516
rect 7243 33476 7288 33504
rect 6181 33467 6239 33473
rect 7282 33464 7288 33476
rect 7340 33464 7346 33516
rect 7484 33513 7512 33544
rect 9306 33532 9312 33544
rect 9364 33532 9370 33584
rect 10870 33572 10876 33584
rect 10783 33544 10876 33572
rect 10870 33532 10876 33544
rect 10928 33572 10934 33584
rect 12437 33575 12495 33581
rect 12437 33572 12449 33575
rect 10928 33544 12449 33572
rect 10928 33532 10934 33544
rect 12437 33541 12449 33544
rect 12483 33541 12495 33575
rect 12437 33535 12495 33541
rect 7469 33507 7527 33513
rect 7469 33473 7481 33507
rect 7515 33473 7527 33507
rect 7469 33467 7527 33473
rect 9217 33507 9275 33513
rect 9217 33473 9229 33507
rect 9263 33504 9275 33507
rect 9766 33504 9772 33516
rect 9263 33476 9772 33504
rect 9263 33473 9275 33476
rect 9217 33467 9275 33473
rect 9766 33464 9772 33476
rect 9824 33504 9830 33516
rect 9861 33507 9919 33513
rect 9861 33504 9873 33507
rect 9824 33476 9873 33504
rect 9824 33464 9830 33476
rect 9861 33473 9873 33476
rect 9907 33473 9919 33507
rect 9861 33467 9919 33473
rect 1397 33439 1455 33445
rect 1397 33405 1409 33439
rect 1443 33436 1455 33439
rect 1946 33436 1952 33448
rect 1443 33408 1952 33436
rect 1443 33405 1455 33408
rect 1397 33399 1455 33405
rect 1946 33396 1952 33408
rect 2004 33396 2010 33448
rect 3329 33439 3387 33445
rect 3329 33405 3341 33439
rect 3375 33436 3387 33439
rect 4157 33439 4215 33445
rect 4157 33436 4169 33439
rect 3375 33408 4169 33436
rect 3375 33405 3387 33408
rect 3329 33399 3387 33405
rect 4157 33405 4169 33408
rect 4203 33436 4215 33439
rect 5350 33436 5356 33448
rect 4203 33408 5356 33436
rect 4203 33405 4215 33408
rect 4157 33399 4215 33405
rect 5350 33396 5356 33408
rect 5408 33396 5414 33448
rect 6546 33396 6552 33448
rect 6604 33436 6610 33448
rect 7190 33436 7196 33448
rect 6604 33408 7196 33436
rect 6604 33396 6610 33408
rect 7190 33396 7196 33408
rect 7248 33396 7254 33448
rect 8849 33439 8907 33445
rect 8849 33405 8861 33439
rect 8895 33436 8907 33439
rect 9674 33436 9680 33448
rect 8895 33408 9680 33436
rect 8895 33405 8907 33408
rect 8849 33399 8907 33405
rect 9674 33396 9680 33408
rect 9732 33396 9738 33448
rect 11238 33396 11244 33448
rect 11296 33436 11302 33448
rect 12820 33445 12848 33612
rect 12894 33464 12900 33516
rect 12952 33504 12958 33516
rect 13081 33507 13139 33513
rect 13081 33504 13093 33507
rect 12952 33476 13093 33504
rect 12952 33464 12958 33476
rect 13081 33473 13093 33476
rect 13127 33504 13139 33507
rect 13449 33507 13507 33513
rect 13449 33504 13461 33507
rect 13127 33476 13461 33504
rect 13127 33473 13139 33476
rect 13081 33467 13139 33473
rect 13449 33473 13461 33476
rect 13495 33473 13507 33507
rect 13449 33467 13507 33473
rect 12069 33439 12127 33445
rect 12069 33436 12081 33439
rect 11296 33408 12081 33436
rect 11296 33396 11302 33408
rect 12069 33405 12081 33408
rect 12115 33436 12127 33439
rect 12161 33439 12219 33445
rect 12161 33436 12173 33439
rect 12115 33408 12173 33436
rect 12115 33405 12127 33408
rect 12069 33399 12127 33405
rect 12161 33405 12173 33408
rect 12207 33405 12219 33439
rect 12161 33399 12219 33405
rect 12805 33439 12863 33445
rect 12805 33405 12817 33439
rect 12851 33405 12863 33439
rect 12805 33399 12863 33405
rect 3697 33371 3755 33377
rect 3697 33337 3709 33371
rect 3743 33368 3755 33371
rect 4424 33371 4482 33377
rect 4424 33368 4436 33371
rect 3743 33340 4436 33368
rect 3743 33337 3755 33340
rect 3697 33331 3755 33337
rect 4424 33337 4436 33340
rect 4470 33368 4482 33371
rect 4706 33368 4712 33380
rect 4470 33340 4712 33368
rect 4470 33337 4482 33340
rect 4424 33331 4482 33337
rect 4706 33328 4712 33340
rect 4764 33328 4770 33380
rect 9398 33328 9404 33380
rect 9456 33368 9462 33380
rect 9769 33371 9827 33377
rect 9769 33368 9781 33371
rect 9456 33340 9781 33368
rect 9456 33328 9462 33340
rect 9769 33337 9781 33340
rect 9815 33337 9827 33371
rect 9769 33331 9827 33337
rect 11057 33371 11115 33377
rect 11057 33337 11069 33371
rect 11103 33368 11115 33371
rect 12342 33368 12348 33380
rect 11103 33340 12348 33368
rect 11103 33337 11115 33340
rect 11057 33331 11115 33337
rect 12342 33328 12348 33340
rect 12400 33328 12406 33380
rect 12710 33328 12716 33380
rect 12768 33368 12774 33380
rect 12897 33371 12955 33377
rect 12897 33368 12909 33371
rect 12768 33340 12909 33368
rect 12768 33328 12774 33340
rect 12897 33337 12909 33340
rect 12943 33368 12955 33371
rect 13170 33368 13176 33380
rect 12943 33340 13176 33368
rect 12943 33337 12955 33340
rect 12897 33331 12955 33337
rect 13170 33328 13176 33340
rect 13228 33328 13234 33380
rect 2777 33303 2835 33309
rect 2777 33269 2789 33303
rect 2823 33300 2835 33303
rect 3050 33300 3056 33312
rect 2823 33272 3056 33300
rect 2823 33269 2835 33272
rect 2777 33263 2835 33269
rect 3050 33260 3056 33272
rect 3108 33260 3114 33312
rect 3970 33300 3976 33312
rect 3931 33272 3976 33300
rect 3970 33260 3976 33272
rect 4028 33260 4034 33312
rect 5537 33303 5595 33309
rect 5537 33269 5549 33303
rect 5583 33300 5595 33303
rect 5626 33300 5632 33312
rect 5583 33272 5632 33300
rect 5583 33269 5595 33272
rect 5537 33263 5595 33269
rect 5626 33260 5632 33272
rect 5684 33260 5690 33312
rect 6822 33300 6828 33312
rect 6783 33272 6828 33300
rect 6822 33260 6828 33272
rect 6880 33260 6886 33312
rect 7282 33260 7288 33312
rect 7340 33300 7346 33312
rect 7558 33300 7564 33312
rect 7340 33272 7564 33300
rect 7340 33260 7346 33272
rect 7558 33260 7564 33272
rect 7616 33300 7622 33312
rect 7837 33303 7895 33309
rect 7837 33300 7849 33303
rect 7616 33272 7849 33300
rect 7616 33260 7622 33272
rect 7837 33269 7849 33272
rect 7883 33269 7895 33303
rect 7837 33263 7895 33269
rect 8110 33260 8116 33312
rect 8168 33300 8174 33312
rect 8297 33303 8355 33309
rect 8297 33300 8309 33303
rect 8168 33272 8309 33300
rect 8168 33260 8174 33272
rect 8297 33269 8309 33272
rect 8343 33300 8355 33303
rect 9582 33300 9588 33312
rect 8343 33272 9588 33300
rect 8343 33269 8355 33272
rect 8297 33263 8355 33269
rect 9582 33260 9588 33272
rect 9640 33260 9646 33312
rect 9858 33260 9864 33312
rect 9916 33300 9922 33312
rect 10413 33303 10471 33309
rect 10413 33300 10425 33303
rect 9916 33272 10425 33300
rect 9916 33260 9922 33272
rect 10413 33269 10425 33272
rect 10459 33300 10471 33303
rect 10686 33300 10692 33312
rect 10459 33272 10692 33300
rect 10459 33269 10471 33272
rect 10413 33263 10471 33269
rect 10686 33260 10692 33272
rect 10744 33300 10750 33312
rect 10870 33300 10876 33312
rect 10744 33272 10876 33300
rect 10744 33260 10750 33272
rect 10870 33260 10876 33272
rect 10928 33260 10934 33312
rect 11422 33260 11428 33312
rect 11480 33300 11486 33312
rect 11793 33303 11851 33309
rect 11793 33300 11805 33303
rect 11480 33272 11805 33300
rect 11480 33260 11486 33272
rect 11793 33269 11805 33272
rect 11839 33269 11851 33303
rect 11793 33263 11851 33269
rect 1104 33210 14812 33232
rect 1104 33158 6315 33210
rect 6367 33158 6379 33210
rect 6431 33158 6443 33210
rect 6495 33158 6507 33210
rect 6559 33158 11648 33210
rect 11700 33158 11712 33210
rect 11764 33158 11776 33210
rect 11828 33158 11840 33210
rect 11892 33158 14812 33210
rect 1104 33136 14812 33158
rect 4154 33056 4160 33108
rect 4212 33096 4218 33108
rect 4249 33099 4307 33105
rect 4249 33096 4261 33099
rect 4212 33068 4261 33096
rect 4212 33056 4218 33068
rect 4249 33065 4261 33068
rect 4295 33065 4307 33099
rect 4249 33059 4307 33065
rect 5261 33099 5319 33105
rect 5261 33065 5273 33099
rect 5307 33096 5319 33099
rect 5534 33096 5540 33108
rect 5307 33068 5540 33096
rect 5307 33065 5319 33068
rect 5261 33059 5319 33065
rect 5534 33056 5540 33068
rect 5592 33096 5598 33108
rect 6822 33096 6828 33108
rect 5592 33068 6828 33096
rect 5592 33056 5598 33068
rect 6822 33056 6828 33068
rect 6880 33056 6886 33108
rect 7558 33056 7564 33108
rect 7616 33096 7622 33108
rect 8757 33099 8815 33105
rect 8757 33096 8769 33099
rect 7616 33068 8769 33096
rect 7616 33056 7622 33068
rect 8757 33065 8769 33068
rect 8803 33096 8815 33099
rect 9306 33096 9312 33108
rect 8803 33068 9312 33096
rect 8803 33065 8815 33068
rect 8757 33059 8815 33065
rect 9306 33056 9312 33068
rect 9364 33056 9370 33108
rect 10137 33099 10195 33105
rect 10137 33065 10149 33099
rect 10183 33096 10195 33099
rect 10778 33096 10784 33108
rect 10183 33068 10784 33096
rect 10183 33065 10195 33068
rect 10137 33059 10195 33065
rect 10778 33056 10784 33068
rect 10836 33056 10842 33108
rect 10870 33056 10876 33108
rect 10928 33096 10934 33108
rect 11609 33099 11667 33105
rect 11609 33096 11621 33099
rect 10928 33068 11621 33096
rect 10928 33056 10934 33068
rect 11609 33065 11621 33068
rect 11655 33065 11667 33099
rect 11609 33059 11667 33065
rect 12069 33099 12127 33105
rect 12069 33065 12081 33099
rect 12115 33096 12127 33099
rect 12342 33096 12348 33108
rect 12115 33068 12348 33096
rect 12115 33065 12127 33068
rect 12069 33059 12127 33065
rect 12342 33056 12348 33068
rect 12400 33056 12406 33108
rect 12529 33099 12587 33105
rect 12529 33065 12541 33099
rect 12575 33096 12587 33099
rect 12710 33096 12716 33108
rect 12575 33068 12716 33096
rect 12575 33065 12587 33068
rect 12529 33059 12587 33065
rect 12710 33056 12716 33068
rect 12768 33056 12774 33108
rect 12894 33096 12900 33108
rect 12855 33068 12900 33096
rect 12894 33056 12900 33068
rect 12952 33056 12958 33108
rect 1670 33028 1676 33040
rect 1631 33000 1676 33028
rect 1670 32988 1676 33000
rect 1728 32988 1734 33040
rect 1394 32960 1400 32972
rect 1355 32932 1400 32960
rect 1394 32920 1400 32932
rect 1452 32920 1458 32972
rect 4065 32963 4123 32969
rect 4065 32929 4077 32963
rect 4111 32960 4123 32963
rect 4154 32960 4160 32972
rect 4111 32932 4160 32960
rect 4111 32929 4123 32932
rect 4065 32923 4123 32929
rect 4154 32920 4160 32932
rect 4212 32920 4218 32972
rect 5350 32960 5356 32972
rect 5311 32932 5356 32960
rect 5350 32920 5356 32932
rect 5408 32920 5414 32972
rect 5626 32969 5632 32972
rect 5620 32960 5632 32969
rect 5539 32932 5632 32960
rect 5620 32923 5632 32932
rect 5684 32960 5690 32972
rect 6178 32960 6184 32972
rect 5684 32932 6184 32960
rect 5626 32920 5632 32923
rect 5684 32920 5690 32932
rect 6178 32920 6184 32932
rect 6236 32920 6242 32972
rect 7285 32963 7343 32969
rect 7285 32929 7297 32963
rect 7331 32960 7343 32963
rect 7742 32960 7748 32972
rect 7331 32932 7748 32960
rect 7331 32929 7343 32932
rect 7285 32923 7343 32929
rect 7742 32920 7748 32932
rect 7800 32920 7806 32972
rect 8110 32960 8116 32972
rect 8071 32932 8116 32960
rect 8110 32920 8116 32932
rect 8168 32920 8174 32972
rect 8202 32920 8208 32972
rect 8260 32960 8266 32972
rect 8260 32932 8305 32960
rect 8260 32920 8266 32932
rect 9674 32920 9680 32972
rect 9732 32920 9738 32972
rect 10502 32969 10508 32972
rect 10496 32960 10508 32969
rect 10463 32932 10508 32960
rect 10496 32923 10508 32932
rect 10502 32920 10508 32923
rect 10560 32920 10566 32972
rect 12250 32920 12256 32972
rect 12308 32960 12314 32972
rect 12912 32960 12940 33056
rect 12308 32932 12940 32960
rect 12308 32920 12314 32932
rect 8297 32895 8355 32901
rect 8297 32892 8309 32895
rect 7116 32864 8309 32892
rect 7116 32836 7144 32864
rect 8297 32861 8309 32864
rect 8343 32861 8355 32895
rect 9692 32892 9720 32920
rect 10226 32892 10232 32904
rect 9692 32864 10232 32892
rect 8297 32855 8355 32861
rect 10226 32852 10232 32864
rect 10284 32852 10290 32904
rect 12710 32852 12716 32904
rect 12768 32892 12774 32904
rect 14642 32892 14648 32904
rect 12768 32864 14648 32892
rect 12768 32852 12774 32864
rect 14642 32852 14648 32864
rect 14700 32852 14706 32904
rect 6638 32784 6644 32836
rect 6696 32824 6702 32836
rect 6733 32827 6791 32833
rect 6733 32824 6745 32827
rect 6696 32796 6745 32824
rect 6696 32784 6702 32796
rect 6733 32793 6745 32796
rect 6779 32824 6791 32827
rect 7098 32824 7104 32836
rect 6779 32796 7104 32824
rect 6779 32793 6791 32796
rect 6733 32787 6791 32793
rect 7098 32784 7104 32796
rect 7156 32784 7162 32836
rect 7745 32827 7803 32833
rect 7745 32793 7757 32827
rect 7791 32824 7803 32827
rect 8846 32824 8852 32836
rect 7791 32796 8852 32824
rect 7791 32793 7803 32796
rect 7745 32787 7803 32793
rect 8846 32784 8852 32796
rect 8904 32824 8910 32836
rect 9125 32827 9183 32833
rect 9125 32824 9137 32827
rect 8904 32796 9137 32824
rect 8904 32784 8910 32796
rect 9125 32793 9137 32796
rect 9171 32793 9183 32827
rect 9125 32787 9183 32793
rect 10244 32756 10272 32852
rect 11514 32756 11520 32768
rect 10244 32728 11520 32756
rect 11514 32716 11520 32728
rect 11572 32716 11578 32768
rect 1104 32666 14812 32688
rect 1104 32614 3648 32666
rect 3700 32614 3712 32666
rect 3764 32614 3776 32666
rect 3828 32614 3840 32666
rect 3892 32614 8982 32666
rect 9034 32614 9046 32666
rect 9098 32614 9110 32666
rect 9162 32614 9174 32666
rect 9226 32614 14315 32666
rect 14367 32614 14379 32666
rect 14431 32614 14443 32666
rect 14495 32614 14507 32666
rect 14559 32614 14812 32666
rect 1104 32592 14812 32614
rect 1394 32512 1400 32564
rect 1452 32552 1458 32564
rect 1581 32555 1639 32561
rect 1581 32552 1593 32555
rect 1452 32524 1593 32552
rect 1452 32512 1458 32524
rect 1581 32521 1593 32524
rect 1627 32521 1639 32555
rect 4154 32552 4160 32564
rect 4115 32524 4160 32552
rect 1581 32515 1639 32521
rect 4154 32512 4160 32524
rect 4212 32512 4218 32564
rect 5166 32552 5172 32564
rect 5127 32524 5172 32552
rect 5166 32512 5172 32524
rect 5224 32512 5230 32564
rect 6178 32552 6184 32564
rect 6139 32524 6184 32552
rect 6178 32512 6184 32524
rect 6236 32512 6242 32564
rect 6638 32552 6644 32564
rect 6599 32524 6644 32552
rect 6638 32512 6644 32524
rect 6696 32512 6702 32564
rect 8110 32512 8116 32564
rect 8168 32552 8174 32564
rect 8570 32552 8576 32564
rect 8168 32524 8576 32552
rect 8168 32512 8174 32524
rect 8570 32512 8576 32524
rect 8628 32512 8634 32564
rect 9674 32512 9680 32564
rect 9732 32552 9738 32564
rect 9769 32555 9827 32561
rect 9769 32552 9781 32555
rect 9732 32524 9781 32552
rect 9732 32512 9738 32524
rect 9769 32521 9781 32524
rect 9815 32521 9827 32555
rect 9769 32515 9827 32521
rect 11425 32555 11483 32561
rect 11425 32521 11437 32555
rect 11471 32552 11483 32555
rect 12250 32552 12256 32564
rect 11471 32524 12256 32552
rect 11471 32521 11483 32524
rect 11425 32515 11483 32521
rect 5077 32487 5135 32493
rect 5077 32453 5089 32487
rect 5123 32484 5135 32487
rect 6656 32484 6684 32512
rect 8202 32484 8208 32496
rect 5123 32456 5764 32484
rect 6656 32456 7788 32484
rect 8163 32456 8208 32484
rect 5123 32453 5135 32456
rect 5077 32447 5135 32453
rect 5534 32376 5540 32428
rect 5592 32416 5598 32428
rect 5736 32425 5764 32456
rect 5629 32419 5687 32425
rect 5629 32416 5641 32419
rect 5592 32388 5641 32416
rect 5592 32376 5598 32388
rect 5629 32385 5641 32388
rect 5675 32385 5687 32419
rect 5629 32379 5687 32385
rect 5721 32419 5779 32425
rect 5721 32385 5733 32419
rect 5767 32416 5779 32419
rect 7282 32416 7288 32428
rect 5767 32388 7288 32416
rect 5767 32385 5779 32388
rect 5721 32379 5779 32385
rect 7282 32376 7288 32388
rect 7340 32376 7346 32428
rect 7760 32425 7788 32456
rect 8202 32444 8208 32456
rect 8260 32444 8266 32496
rect 8294 32444 8300 32496
rect 8352 32484 8358 32496
rect 8757 32487 8815 32493
rect 8757 32484 8769 32487
rect 8352 32456 8769 32484
rect 8352 32444 8358 32456
rect 8757 32453 8769 32456
rect 8803 32453 8815 32487
rect 8757 32447 8815 32453
rect 7745 32419 7803 32425
rect 7745 32385 7757 32419
rect 7791 32385 7803 32419
rect 9306 32416 9312 32428
rect 9267 32388 9312 32416
rect 7745 32379 7803 32385
rect 9306 32376 9312 32388
rect 9364 32376 9370 32428
rect 5258 32308 5264 32360
rect 5316 32348 5322 32360
rect 7101 32351 7159 32357
rect 7101 32348 7113 32351
rect 5316 32320 7113 32348
rect 5316 32308 5322 32320
rect 7101 32317 7113 32320
rect 7147 32348 7159 32351
rect 7147 32320 7512 32348
rect 7147 32317 7159 32320
rect 7101 32311 7159 32317
rect 4709 32283 4767 32289
rect 4709 32249 4721 32283
rect 4755 32280 4767 32283
rect 5537 32283 5595 32289
rect 5537 32280 5549 32283
rect 4755 32252 5549 32280
rect 4755 32249 4767 32252
rect 4709 32243 4767 32249
rect 5537 32249 5549 32252
rect 5583 32280 5595 32283
rect 5583 32252 7236 32280
rect 5583 32249 5595 32252
rect 5537 32243 5595 32249
rect 7208 32221 7236 32252
rect 7484 32224 7512 32320
rect 8846 32308 8852 32360
rect 8904 32348 8910 32360
rect 9125 32351 9183 32357
rect 9125 32348 9137 32351
rect 8904 32320 9137 32348
rect 8904 32308 8910 32320
rect 9125 32317 9137 32320
rect 9171 32317 9183 32351
rect 9784 32348 9812 32515
rect 10502 32376 10508 32428
rect 10560 32416 10566 32428
rect 10965 32419 11023 32425
rect 10965 32416 10977 32419
rect 10560 32388 10977 32416
rect 10560 32376 10566 32388
rect 10965 32385 10977 32388
rect 11011 32416 11023 32419
rect 11440 32416 11468 32515
rect 12250 32512 12256 32524
rect 12308 32512 12314 32564
rect 11011 32388 11468 32416
rect 11011 32385 11023 32388
rect 10965 32379 11023 32385
rect 10781 32351 10839 32357
rect 10781 32348 10793 32351
rect 9784 32320 10793 32348
rect 9125 32311 9183 32317
rect 10781 32317 10793 32320
rect 10827 32317 10839 32351
rect 10781 32311 10839 32317
rect 7653 32283 7711 32289
rect 7653 32249 7665 32283
rect 7699 32280 7711 32283
rect 7742 32280 7748 32292
rect 7699 32252 7748 32280
rect 7699 32249 7711 32252
rect 7653 32243 7711 32249
rect 7742 32240 7748 32252
rect 7800 32240 7806 32292
rect 9674 32240 9680 32292
rect 9732 32280 9738 32292
rect 10137 32283 10195 32289
rect 10137 32280 10149 32283
rect 9732 32252 10149 32280
rect 9732 32240 9738 32252
rect 10137 32249 10149 32252
rect 10183 32280 10195 32283
rect 10689 32283 10747 32289
rect 10689 32280 10701 32283
rect 10183 32252 10701 32280
rect 10183 32249 10195 32252
rect 10137 32243 10195 32249
rect 10689 32249 10701 32252
rect 10735 32249 10747 32283
rect 10689 32243 10747 32249
rect 7193 32215 7251 32221
rect 7193 32181 7205 32215
rect 7239 32181 7251 32215
rect 7193 32175 7251 32181
rect 7466 32172 7472 32224
rect 7524 32212 7530 32224
rect 7561 32215 7619 32221
rect 7561 32212 7573 32215
rect 7524 32184 7573 32212
rect 7524 32172 7530 32184
rect 7561 32181 7573 32184
rect 7607 32181 7619 32215
rect 7561 32175 7619 32181
rect 8846 32172 8852 32224
rect 8904 32212 8910 32224
rect 9217 32215 9275 32221
rect 9217 32212 9229 32215
rect 8904 32184 9229 32212
rect 8904 32172 8910 32184
rect 9217 32181 9229 32184
rect 9263 32181 9275 32215
rect 10318 32212 10324 32224
rect 10279 32184 10324 32212
rect 9217 32175 9275 32181
rect 10318 32172 10324 32184
rect 10376 32172 10382 32224
rect 1104 32122 14812 32144
rect 1104 32070 6315 32122
rect 6367 32070 6379 32122
rect 6431 32070 6443 32122
rect 6495 32070 6507 32122
rect 6559 32070 11648 32122
rect 11700 32070 11712 32122
rect 11764 32070 11776 32122
rect 11828 32070 11840 32122
rect 11892 32070 14812 32122
rect 1104 32048 14812 32070
rect 5350 32008 5356 32020
rect 5311 31980 5356 32008
rect 5350 31968 5356 31980
rect 5408 32008 5414 32020
rect 6178 32008 6184 32020
rect 5408 31980 6184 32008
rect 5408 31968 5414 31980
rect 6178 31968 6184 31980
rect 6236 31968 6242 32020
rect 7282 31968 7288 32020
rect 7340 32008 7346 32020
rect 7745 32011 7803 32017
rect 7745 32008 7757 32011
rect 7340 31980 7757 32008
rect 7340 31968 7346 31980
rect 7745 31977 7757 31980
rect 7791 31977 7803 32011
rect 8570 32008 8576 32020
rect 8531 31980 8576 32008
rect 7745 31971 7803 31977
rect 8570 31968 8576 31980
rect 8628 31968 8634 32020
rect 9490 32008 9496 32020
rect 9403 31980 9496 32008
rect 9490 31968 9496 31980
rect 9548 32008 9554 32020
rect 10318 32008 10324 32020
rect 9548 31980 10324 32008
rect 9548 31968 9554 31980
rect 10318 31968 10324 31980
rect 10376 31968 10382 32020
rect 10502 31968 10508 32020
rect 10560 32008 10566 32020
rect 10689 32011 10747 32017
rect 10689 32008 10701 32011
rect 10560 31980 10701 32008
rect 10560 31968 10566 31980
rect 10689 31977 10701 31980
rect 10735 31977 10747 32011
rect 10689 31971 10747 31977
rect 6638 31949 6644 31952
rect 6632 31940 6644 31949
rect 6599 31912 6644 31940
rect 6632 31903 6644 31912
rect 6696 31940 6702 31952
rect 6914 31940 6920 31952
rect 6696 31912 6920 31940
rect 6638 31900 6644 31903
rect 6696 31900 6702 31912
rect 6914 31900 6920 31912
rect 6972 31900 6978 31952
rect 10045 31943 10103 31949
rect 10045 31909 10057 31943
rect 10091 31940 10103 31943
rect 10226 31940 10232 31952
rect 10091 31912 10232 31940
rect 10091 31909 10103 31912
rect 10045 31903 10103 31909
rect 10226 31900 10232 31912
rect 10284 31900 10290 31952
rect 6178 31832 6184 31884
rect 6236 31872 6242 31884
rect 6365 31875 6423 31881
rect 6365 31872 6377 31875
rect 6236 31844 6377 31872
rect 6236 31832 6242 31844
rect 6365 31841 6377 31844
rect 6411 31841 6423 31875
rect 10134 31872 10140 31884
rect 10095 31844 10140 31872
rect 6365 31835 6423 31841
rect 10134 31832 10140 31844
rect 10192 31832 10198 31884
rect 4890 31804 4896 31816
rect 4851 31776 4896 31804
rect 4890 31764 4896 31776
rect 4948 31764 4954 31816
rect 10318 31804 10324 31816
rect 10231 31776 10324 31804
rect 10318 31764 10324 31776
rect 10376 31804 10382 31816
rect 10520 31804 10548 31968
rect 10376 31776 10548 31804
rect 10376 31764 10382 31776
rect 7006 31628 7012 31680
rect 7064 31668 7070 31680
rect 8018 31668 8024 31680
rect 7064 31640 8024 31668
rect 7064 31628 7070 31640
rect 8018 31628 8024 31640
rect 8076 31628 8082 31680
rect 8846 31628 8852 31680
rect 8904 31668 8910 31680
rect 9033 31671 9091 31677
rect 9033 31668 9045 31671
rect 8904 31640 9045 31668
rect 8904 31628 8910 31640
rect 9033 31637 9045 31640
rect 9079 31637 9091 31671
rect 9033 31631 9091 31637
rect 9582 31628 9588 31680
rect 9640 31668 9646 31680
rect 9677 31671 9735 31677
rect 9677 31668 9689 31671
rect 9640 31640 9689 31668
rect 9640 31628 9646 31640
rect 9677 31637 9689 31640
rect 9723 31637 9735 31671
rect 9677 31631 9735 31637
rect 11149 31671 11207 31677
rect 11149 31637 11161 31671
rect 11195 31668 11207 31671
rect 11514 31668 11520 31680
rect 11195 31640 11520 31668
rect 11195 31637 11207 31640
rect 11149 31631 11207 31637
rect 11514 31628 11520 31640
rect 11572 31628 11578 31680
rect 1104 31578 14812 31600
rect 1104 31526 3648 31578
rect 3700 31526 3712 31578
rect 3764 31526 3776 31578
rect 3828 31526 3840 31578
rect 3892 31526 8982 31578
rect 9034 31526 9046 31578
rect 9098 31526 9110 31578
rect 9162 31526 9174 31578
rect 9226 31526 14315 31578
rect 14367 31526 14379 31578
rect 14431 31526 14443 31578
rect 14495 31526 14507 31578
rect 14559 31526 14812 31578
rect 1104 31504 14812 31526
rect 7653 31467 7711 31473
rect 7653 31433 7665 31467
rect 7699 31464 7711 31467
rect 8846 31464 8852 31476
rect 7699 31436 8852 31464
rect 7699 31433 7711 31436
rect 7653 31427 7711 31433
rect 8846 31424 8852 31436
rect 8904 31424 8910 31476
rect 9217 31467 9275 31473
rect 9217 31433 9229 31467
rect 9263 31464 9275 31467
rect 9398 31464 9404 31476
rect 9263 31436 9404 31464
rect 9263 31433 9275 31436
rect 9217 31427 9275 31433
rect 9398 31424 9404 31436
rect 9456 31424 9462 31476
rect 10318 31464 10324 31476
rect 9508 31436 10324 31464
rect 6457 31399 6515 31405
rect 6457 31365 6469 31399
rect 6503 31396 6515 31399
rect 6914 31396 6920 31408
rect 6503 31368 6920 31396
rect 6503 31365 6515 31368
rect 6457 31359 6515 31365
rect 6914 31356 6920 31368
rect 6972 31396 6978 31408
rect 7101 31399 7159 31405
rect 7101 31396 7113 31399
rect 6972 31368 7113 31396
rect 6972 31356 6978 31368
rect 7101 31365 7113 31368
rect 7147 31365 7159 31399
rect 7101 31359 7159 31365
rect 9125 31399 9183 31405
rect 9125 31365 9137 31399
rect 9171 31396 9183 31399
rect 9508 31396 9536 31436
rect 10318 31424 10324 31436
rect 10376 31424 10382 31476
rect 9171 31368 9536 31396
rect 9171 31365 9183 31368
rect 9125 31359 9183 31365
rect 9582 31356 9588 31408
rect 9640 31356 9646 31408
rect 4154 31288 4160 31340
rect 4212 31328 4218 31340
rect 4341 31331 4399 31337
rect 4341 31328 4353 31331
rect 4212 31300 4353 31328
rect 4212 31288 4218 31300
rect 4341 31297 4353 31300
rect 4387 31328 4399 31331
rect 5350 31328 5356 31340
rect 4387 31300 5356 31328
rect 4387 31297 4399 31300
rect 4341 31291 4399 31297
rect 5350 31288 5356 31300
rect 5408 31288 5414 31340
rect 8018 31288 8024 31340
rect 8076 31328 8082 31340
rect 8205 31331 8263 31337
rect 8205 31328 8217 31331
rect 8076 31300 8217 31328
rect 8076 31288 8082 31300
rect 8205 31297 8217 31300
rect 8251 31297 8263 31331
rect 8205 31291 8263 31297
rect 8757 31331 8815 31337
rect 8757 31297 8769 31331
rect 8803 31328 8815 31331
rect 9600 31328 9628 31356
rect 9677 31331 9735 31337
rect 9677 31328 9689 31331
rect 8803 31300 9689 31328
rect 8803 31297 8815 31300
rect 8757 31291 8815 31297
rect 9677 31297 9689 31300
rect 9723 31297 9735 31331
rect 9858 31328 9864 31340
rect 9819 31300 9864 31328
rect 9677 31291 9735 31297
rect 9858 31288 9864 31300
rect 9916 31288 9922 31340
rect 4890 31220 4896 31272
rect 4948 31260 4954 31272
rect 5169 31263 5227 31269
rect 5169 31260 5181 31263
rect 4948 31232 5181 31260
rect 4948 31220 4954 31232
rect 5169 31229 5181 31232
rect 5215 31229 5227 31263
rect 8110 31260 8116 31272
rect 8023 31232 8116 31260
rect 5169 31223 5227 31229
rect 8110 31220 8116 31232
rect 8168 31220 8174 31272
rect 9490 31220 9496 31272
rect 9548 31260 9554 31272
rect 9585 31263 9643 31269
rect 9585 31260 9597 31263
rect 9548 31232 9597 31260
rect 9548 31220 9554 31232
rect 9585 31229 9597 31232
rect 9631 31229 9643 31263
rect 9585 31223 9643 31229
rect 4709 31195 4767 31201
rect 4709 31161 4721 31195
rect 4755 31192 4767 31195
rect 5258 31192 5264 31204
rect 4755 31164 5264 31192
rect 4755 31161 4767 31164
rect 4709 31155 4767 31161
rect 5258 31152 5264 31164
rect 5316 31152 5322 31204
rect 7650 31192 7656 31204
rect 7484 31164 7656 31192
rect 4798 31124 4804 31136
rect 4759 31096 4804 31124
rect 4798 31084 4804 31096
rect 4856 31084 4862 31136
rect 6089 31127 6147 31133
rect 6089 31093 6101 31127
rect 6135 31124 6147 31127
rect 6178 31124 6184 31136
rect 6135 31096 6184 31124
rect 6135 31093 6147 31096
rect 6089 31087 6147 31093
rect 6178 31084 6184 31096
rect 6236 31084 6242 31136
rect 7098 31084 7104 31136
rect 7156 31124 7162 31136
rect 7484 31133 7512 31164
rect 7650 31152 7656 31164
rect 7708 31192 7714 31204
rect 8021 31195 8079 31201
rect 8021 31192 8033 31195
rect 7708 31164 8033 31192
rect 7708 31152 7714 31164
rect 8021 31161 8033 31164
rect 8067 31161 8079 31195
rect 8128 31192 8156 31220
rect 8128 31164 9628 31192
rect 8021 31155 8079 31161
rect 9600 31136 9628 31164
rect 9674 31152 9680 31204
rect 9732 31192 9738 31204
rect 9950 31192 9956 31204
rect 9732 31164 9956 31192
rect 9732 31152 9738 31164
rect 9950 31152 9956 31164
rect 10008 31152 10014 31204
rect 7469 31127 7527 31133
rect 7469 31124 7481 31127
rect 7156 31096 7481 31124
rect 7156 31084 7162 31096
rect 7469 31093 7481 31096
rect 7515 31093 7527 31127
rect 7469 31087 7527 31093
rect 9582 31084 9588 31136
rect 9640 31084 9646 31136
rect 10226 31124 10232 31136
rect 10187 31096 10232 31124
rect 10226 31084 10232 31096
rect 10284 31084 10290 31136
rect 1104 31034 14812 31056
rect 1104 30982 6315 31034
rect 6367 30982 6379 31034
rect 6431 30982 6443 31034
rect 6495 30982 6507 31034
rect 6559 30982 11648 31034
rect 11700 30982 11712 31034
rect 11764 30982 11776 31034
rect 11828 30982 11840 31034
rect 11892 30982 14812 31034
rect 1104 30960 14812 30982
rect 4890 30920 4896 30932
rect 4851 30892 4896 30920
rect 4890 30880 4896 30892
rect 4948 30880 4954 30932
rect 7745 30923 7803 30929
rect 7745 30889 7757 30923
rect 7791 30920 7803 30923
rect 8110 30920 8116 30932
rect 7791 30892 8116 30920
rect 7791 30889 7803 30892
rect 7745 30883 7803 30889
rect 8110 30880 8116 30892
rect 8168 30880 8174 30932
rect 9306 30920 9312 30932
rect 9267 30892 9312 30920
rect 9306 30880 9312 30892
rect 9364 30880 9370 30932
rect 9953 30923 10011 30929
rect 9953 30889 9965 30923
rect 9999 30920 10011 30923
rect 10134 30920 10140 30932
rect 9999 30892 10140 30920
rect 9999 30889 10011 30892
rect 9953 30883 10011 30889
rect 10134 30880 10140 30892
rect 10192 30880 10198 30932
rect 7466 30812 7472 30864
rect 7524 30852 7530 30864
rect 8018 30852 8024 30864
rect 7524 30824 8024 30852
rect 7524 30812 7530 30824
rect 8018 30812 8024 30824
rect 8076 30812 8082 30864
rect 5074 30744 5080 30796
rect 5132 30784 5138 30796
rect 5442 30784 5448 30796
rect 5132 30756 5448 30784
rect 5132 30744 5138 30756
rect 5442 30744 5448 30756
rect 5500 30744 5506 30796
rect 11600 30787 11658 30793
rect 11600 30753 11612 30787
rect 11646 30784 11658 30787
rect 11974 30784 11980 30796
rect 11646 30756 11980 30784
rect 11646 30753 11658 30756
rect 11600 30747 11658 30753
rect 11974 30744 11980 30756
rect 12032 30744 12038 30796
rect 5534 30716 5540 30728
rect 5495 30688 5540 30716
rect 5534 30676 5540 30688
rect 5592 30676 5598 30728
rect 5629 30719 5687 30725
rect 5629 30685 5641 30719
rect 5675 30685 5687 30719
rect 5629 30679 5687 30685
rect 11333 30719 11391 30725
rect 11333 30685 11345 30719
rect 11379 30685 11391 30719
rect 11333 30679 11391 30685
rect 5350 30608 5356 30660
rect 5408 30648 5414 30660
rect 5644 30648 5672 30679
rect 5408 30620 5672 30648
rect 5408 30608 5414 30620
rect 1857 30583 1915 30589
rect 1857 30549 1869 30583
rect 1903 30580 1915 30583
rect 2222 30580 2228 30592
rect 1903 30552 2228 30580
rect 1903 30549 1915 30552
rect 1857 30543 1915 30549
rect 2222 30540 2228 30552
rect 2280 30540 2286 30592
rect 5077 30583 5135 30589
rect 5077 30549 5089 30583
rect 5123 30580 5135 30583
rect 6917 30583 6975 30589
rect 6917 30580 6929 30583
rect 5123 30552 6929 30580
rect 5123 30549 5135 30552
rect 5077 30543 5135 30549
rect 6917 30549 6929 30552
rect 6963 30580 6975 30583
rect 7282 30580 7288 30592
rect 6963 30552 7288 30580
rect 6963 30549 6975 30552
rect 6917 30543 6975 30549
rect 7282 30540 7288 30552
rect 7340 30540 7346 30592
rect 10502 30540 10508 30592
rect 10560 30580 10566 30592
rect 10778 30580 10784 30592
rect 10560 30552 10784 30580
rect 10560 30540 10566 30552
rect 10778 30540 10784 30552
rect 10836 30540 10842 30592
rect 10873 30583 10931 30589
rect 10873 30549 10885 30583
rect 10919 30580 10931 30583
rect 11238 30580 11244 30592
rect 10919 30552 11244 30580
rect 10919 30549 10931 30552
rect 10873 30543 10931 30549
rect 11238 30540 11244 30552
rect 11296 30540 11302 30592
rect 11348 30580 11376 30679
rect 11514 30580 11520 30592
rect 11348 30552 11520 30580
rect 11514 30540 11520 30552
rect 11572 30540 11578 30592
rect 12434 30540 12440 30592
rect 12492 30580 12498 30592
rect 12713 30583 12771 30589
rect 12713 30580 12725 30583
rect 12492 30552 12725 30580
rect 12492 30540 12498 30552
rect 12713 30549 12725 30552
rect 12759 30549 12771 30583
rect 12713 30543 12771 30549
rect 12894 30540 12900 30592
rect 12952 30580 12958 30592
rect 12989 30583 13047 30589
rect 12989 30580 13001 30583
rect 12952 30552 13001 30580
rect 12952 30540 12958 30552
rect 12989 30549 13001 30552
rect 13035 30549 13047 30583
rect 12989 30543 13047 30549
rect 1104 30490 14812 30512
rect 1104 30438 3648 30490
rect 3700 30438 3712 30490
rect 3764 30438 3776 30490
rect 3828 30438 3840 30490
rect 3892 30438 8982 30490
rect 9034 30438 9046 30490
rect 9098 30438 9110 30490
rect 9162 30438 9174 30490
rect 9226 30438 14315 30490
rect 14367 30438 14379 30490
rect 14431 30438 14443 30490
rect 14495 30438 14507 30490
rect 14559 30438 14812 30490
rect 1104 30416 14812 30438
rect 10318 30336 10324 30388
rect 10376 30376 10382 30388
rect 10686 30376 10692 30388
rect 10376 30348 10692 30376
rect 10376 30336 10382 30348
rect 10686 30336 10692 30348
rect 10744 30336 10750 30388
rect 4706 30308 4712 30320
rect 4667 30280 4712 30308
rect 4706 30268 4712 30280
rect 4764 30268 4770 30320
rect 4798 30268 4804 30320
rect 4856 30308 4862 30320
rect 6641 30311 6699 30317
rect 6641 30308 6653 30311
rect 4856 30280 6653 30308
rect 4856 30268 4862 30280
rect 6641 30277 6653 30280
rect 6687 30308 6699 30311
rect 10778 30308 10784 30320
rect 6687 30280 7420 30308
rect 10739 30280 10784 30308
rect 6687 30277 6699 30280
rect 6641 30271 6699 30277
rect 1673 30243 1731 30249
rect 1673 30209 1685 30243
rect 1719 30240 1731 30243
rect 2406 30240 2412 30252
rect 1719 30212 2412 30240
rect 1719 30209 1731 30212
rect 1673 30203 1731 30209
rect 2406 30200 2412 30212
rect 2464 30200 2470 30252
rect 5534 30200 5540 30252
rect 5592 30240 5598 30252
rect 5813 30243 5871 30249
rect 5813 30240 5825 30243
rect 5592 30212 5825 30240
rect 5592 30200 5598 30212
rect 5813 30209 5825 30212
rect 5859 30209 5871 30243
rect 7282 30240 7288 30252
rect 7243 30212 7288 30240
rect 5813 30203 5871 30209
rect 7282 30200 7288 30212
rect 7340 30200 7346 30252
rect 7392 30249 7420 30280
rect 10778 30268 10784 30280
rect 10836 30268 10842 30320
rect 12434 30308 12440 30320
rect 11440 30280 12440 30308
rect 7377 30243 7435 30249
rect 7377 30209 7389 30243
rect 7423 30209 7435 30243
rect 10686 30240 10692 30252
rect 10599 30212 10692 30240
rect 7377 30203 7435 30209
rect 10686 30200 10692 30212
rect 10744 30240 10750 30252
rect 11440 30249 11468 30280
rect 12434 30268 12440 30280
rect 12492 30268 12498 30320
rect 11425 30243 11483 30249
rect 11425 30240 11437 30243
rect 10744 30212 11437 30240
rect 10744 30200 10750 30212
rect 11425 30209 11437 30212
rect 11471 30209 11483 30243
rect 11425 30203 11483 30209
rect 12253 30243 12311 30249
rect 12253 30209 12265 30243
rect 12299 30240 12311 30243
rect 13081 30243 13139 30249
rect 13081 30240 13093 30243
rect 12299 30212 13093 30240
rect 12299 30209 12311 30212
rect 12253 30203 12311 30209
rect 13081 30209 13093 30212
rect 13127 30240 13139 30243
rect 13722 30240 13728 30252
rect 13127 30212 13728 30240
rect 13127 30209 13139 30212
rect 13081 30203 13139 30209
rect 13722 30200 13728 30212
rect 13780 30200 13786 30252
rect 3326 30172 3332 30184
rect 3287 30144 3332 30172
rect 3326 30132 3332 30144
rect 3384 30132 3390 30184
rect 7190 30172 7196 30184
rect 7151 30144 7196 30172
rect 7190 30132 7196 30144
rect 7248 30132 7254 30184
rect 11238 30172 11244 30184
rect 11199 30144 11244 30172
rect 11238 30132 11244 30144
rect 11296 30132 11302 30184
rect 12805 30175 12863 30181
rect 12805 30141 12817 30175
rect 12851 30172 12863 30175
rect 12894 30172 12900 30184
rect 12851 30144 12900 30172
rect 12851 30141 12863 30144
rect 12805 30135 12863 30141
rect 12894 30132 12900 30144
rect 12952 30132 12958 30184
rect 2130 30104 2136 30116
rect 2091 30076 2136 30104
rect 2130 30064 2136 30076
rect 2188 30064 2194 30116
rect 3237 30107 3295 30113
rect 3237 30073 3249 30107
rect 3283 30104 3295 30107
rect 3596 30107 3654 30113
rect 3596 30104 3608 30107
rect 3283 30076 3608 30104
rect 3283 30073 3295 30076
rect 3237 30067 3295 30073
rect 3596 30073 3608 30076
rect 3642 30104 3654 30107
rect 4798 30104 4804 30116
rect 3642 30076 4804 30104
rect 3642 30073 3654 30076
rect 3596 30067 3654 30073
rect 4798 30064 4804 30076
rect 4856 30064 4862 30116
rect 10321 30107 10379 30113
rect 10321 30073 10333 30107
rect 10367 30104 10379 30107
rect 10367 30076 11192 30104
rect 10367 30073 10379 30076
rect 10321 30067 10379 30073
rect 11164 30048 11192 30076
rect 1762 30036 1768 30048
rect 1723 30008 1768 30036
rect 1762 29996 1768 30008
rect 1820 29996 1826 30048
rect 2222 30036 2228 30048
rect 2183 30008 2228 30036
rect 2222 29996 2228 30008
rect 2280 29996 2286 30048
rect 4522 29996 4528 30048
rect 4580 30036 4586 30048
rect 5074 30036 5080 30048
rect 4580 30008 5080 30036
rect 4580 29996 4586 30008
rect 5074 29996 5080 30008
rect 5132 29996 5138 30048
rect 5537 30039 5595 30045
rect 5537 30005 5549 30039
rect 5583 30036 5595 30039
rect 5626 30036 5632 30048
rect 5583 30008 5632 30036
rect 5583 30005 5595 30008
rect 5537 29999 5595 30005
rect 5626 29996 5632 30008
rect 5684 29996 5690 30048
rect 6822 30036 6828 30048
rect 6783 30008 6828 30036
rect 6822 29996 6828 30008
rect 6880 29996 6886 30048
rect 11146 30036 11152 30048
rect 11107 30008 11152 30036
rect 11146 29996 11152 30008
rect 11204 29996 11210 30048
rect 11885 30039 11943 30045
rect 11885 30005 11897 30039
rect 11931 30036 11943 30039
rect 11974 30036 11980 30048
rect 11931 30008 11980 30036
rect 11931 30005 11943 30008
rect 11885 29999 11943 30005
rect 11974 29996 11980 30008
rect 12032 29996 12038 30048
rect 12437 30039 12495 30045
rect 12437 30005 12449 30039
rect 12483 30036 12495 30039
rect 12526 30036 12532 30048
rect 12483 30008 12532 30036
rect 12483 30005 12495 30008
rect 12437 29999 12495 30005
rect 12526 29996 12532 30008
rect 12584 29996 12590 30048
rect 12894 30036 12900 30048
rect 12855 30008 12900 30036
rect 12894 29996 12900 30008
rect 12952 30036 12958 30048
rect 13449 30039 13507 30045
rect 13449 30036 13461 30039
rect 12952 30008 13461 30036
rect 12952 29996 12958 30008
rect 13449 30005 13461 30008
rect 13495 30005 13507 30039
rect 13449 29999 13507 30005
rect 1104 29946 14812 29968
rect 1104 29894 6315 29946
rect 6367 29894 6379 29946
rect 6431 29894 6443 29946
rect 6495 29894 6507 29946
rect 6559 29894 11648 29946
rect 11700 29894 11712 29946
rect 11764 29894 11776 29946
rect 11828 29894 11840 29946
rect 11892 29894 14812 29946
rect 1104 29872 14812 29894
rect 2130 29832 2136 29844
rect 2091 29804 2136 29832
rect 2130 29792 2136 29804
rect 2188 29792 2194 29844
rect 4154 29832 4160 29844
rect 4115 29804 4160 29832
rect 4154 29792 4160 29804
rect 4212 29792 4218 29844
rect 6273 29835 6331 29841
rect 6273 29801 6285 29835
rect 6319 29832 6331 29835
rect 6638 29832 6644 29844
rect 6319 29804 6644 29832
rect 6319 29801 6331 29804
rect 6273 29795 6331 29801
rect 6638 29792 6644 29804
rect 6696 29792 6702 29844
rect 7009 29835 7067 29841
rect 7009 29801 7021 29835
rect 7055 29832 7067 29835
rect 7190 29832 7196 29844
rect 7055 29804 7196 29832
rect 7055 29801 7067 29804
rect 7009 29795 7067 29801
rect 7190 29792 7196 29804
rect 7248 29792 7254 29844
rect 13722 29832 13728 29844
rect 13683 29804 13728 29832
rect 13722 29792 13728 29804
rect 13780 29792 13786 29844
rect 1670 29764 1676 29776
rect 1631 29736 1676 29764
rect 1670 29724 1676 29736
rect 1728 29724 1734 29776
rect 9306 29724 9312 29776
rect 9364 29764 9370 29776
rect 9922 29767 9980 29773
rect 9922 29764 9934 29767
rect 9364 29736 9934 29764
rect 9364 29724 9370 29736
rect 9922 29733 9934 29736
rect 9968 29733 9980 29767
rect 9922 29727 9980 29733
rect 1397 29699 1455 29705
rect 1397 29665 1409 29699
rect 1443 29696 1455 29699
rect 1762 29696 1768 29708
rect 1443 29668 1768 29696
rect 1443 29665 1455 29668
rect 1397 29659 1455 29665
rect 1762 29656 1768 29668
rect 1820 29656 1826 29708
rect 4525 29699 4583 29705
rect 4525 29665 4537 29699
rect 4571 29665 4583 29699
rect 4525 29659 4583 29665
rect 4617 29699 4675 29705
rect 4617 29665 4629 29699
rect 4663 29696 4675 29699
rect 4982 29696 4988 29708
rect 4663 29668 4988 29696
rect 4663 29665 4675 29668
rect 4617 29659 4675 29665
rect 3326 29520 3332 29572
rect 3384 29560 3390 29572
rect 3421 29563 3479 29569
rect 3421 29560 3433 29563
rect 3384 29532 3433 29560
rect 3384 29520 3390 29532
rect 3421 29529 3433 29532
rect 3467 29560 3479 29563
rect 4246 29560 4252 29572
rect 3467 29532 4252 29560
rect 3467 29529 3479 29532
rect 3421 29523 3479 29529
rect 4246 29520 4252 29532
rect 4304 29520 4310 29572
rect 3510 29452 3516 29504
rect 3568 29492 3574 29504
rect 3789 29495 3847 29501
rect 3789 29492 3801 29495
rect 3568 29464 3801 29492
rect 3568 29452 3574 29464
rect 3789 29461 3801 29464
rect 3835 29492 3847 29495
rect 4540 29492 4568 29659
rect 4982 29656 4988 29668
rect 5040 29656 5046 29708
rect 9677 29699 9735 29705
rect 9677 29665 9689 29699
rect 9723 29696 9735 29699
rect 10226 29696 10232 29708
rect 9723 29668 10232 29696
rect 9723 29665 9735 29668
rect 9677 29659 9735 29665
rect 10226 29656 10232 29668
rect 10284 29696 10290 29708
rect 10284 29668 11468 29696
rect 10284 29656 10290 29668
rect 4798 29628 4804 29640
rect 4759 29600 4804 29628
rect 4798 29588 4804 29600
rect 4856 29588 4862 29640
rect 5994 29588 6000 29640
rect 6052 29628 6058 29640
rect 6365 29631 6423 29637
rect 6365 29628 6377 29631
rect 6052 29600 6377 29628
rect 6052 29588 6058 29600
rect 6365 29597 6377 29600
rect 6411 29597 6423 29631
rect 6365 29591 6423 29597
rect 6454 29588 6460 29640
rect 6512 29628 6518 29640
rect 11440 29637 11468 29668
rect 12434 29656 12440 29708
rect 12492 29696 12498 29708
rect 12612 29699 12670 29705
rect 12612 29696 12624 29699
rect 12492 29668 12624 29696
rect 12492 29656 12498 29668
rect 12612 29665 12624 29668
rect 12658 29696 12670 29699
rect 12986 29696 12992 29708
rect 12658 29668 12992 29696
rect 12658 29665 12670 29668
rect 12612 29659 12670 29665
rect 12986 29656 12992 29668
rect 13044 29656 13050 29708
rect 11425 29631 11483 29637
rect 6512 29600 6557 29628
rect 6512 29588 6518 29600
rect 11425 29597 11437 29631
rect 11471 29628 11483 29631
rect 11514 29628 11520 29640
rect 11471 29600 11520 29628
rect 11471 29597 11483 29600
rect 11425 29591 11483 29597
rect 11514 29588 11520 29600
rect 11572 29628 11578 29640
rect 12342 29628 12348 29640
rect 11572 29600 12348 29628
rect 11572 29588 11578 29600
rect 12342 29588 12348 29600
rect 12400 29588 12406 29640
rect 5902 29492 5908 29504
rect 3835 29464 4568 29492
rect 5863 29464 5908 29492
rect 3835 29461 3847 29464
rect 3789 29455 3847 29461
rect 5902 29452 5908 29464
rect 5960 29452 5966 29504
rect 8205 29495 8263 29501
rect 8205 29461 8217 29495
rect 8251 29492 8263 29495
rect 8570 29492 8576 29504
rect 8251 29464 8576 29492
rect 8251 29461 8263 29464
rect 8205 29455 8263 29461
rect 8570 29452 8576 29464
rect 8628 29452 8634 29504
rect 9950 29452 9956 29504
rect 10008 29492 10014 29504
rect 11057 29495 11115 29501
rect 11057 29492 11069 29495
rect 10008 29464 11069 29492
rect 10008 29452 10014 29464
rect 11057 29461 11069 29464
rect 11103 29461 11115 29495
rect 11057 29455 11115 29461
rect 1104 29402 14812 29424
rect 1104 29350 3648 29402
rect 3700 29350 3712 29402
rect 3764 29350 3776 29402
rect 3828 29350 3840 29402
rect 3892 29350 8982 29402
rect 9034 29350 9046 29402
rect 9098 29350 9110 29402
rect 9162 29350 9174 29402
rect 9226 29350 14315 29402
rect 14367 29350 14379 29402
rect 14431 29350 14443 29402
rect 14495 29350 14507 29402
rect 14559 29350 14812 29402
rect 1104 29328 14812 29350
rect 1673 29291 1731 29297
rect 1673 29257 1685 29291
rect 1719 29288 1731 29291
rect 1762 29288 1768 29300
rect 1719 29260 1768 29288
rect 1719 29257 1731 29260
rect 1673 29251 1731 29257
rect 1762 29248 1768 29260
rect 1820 29248 1826 29300
rect 4798 29248 4804 29300
rect 4856 29288 4862 29300
rect 5077 29291 5135 29297
rect 5077 29288 5089 29291
rect 4856 29260 5089 29288
rect 4856 29248 4862 29260
rect 5077 29257 5089 29260
rect 5123 29257 5135 29291
rect 5077 29251 5135 29257
rect 6365 29291 6423 29297
rect 6365 29257 6377 29291
rect 6411 29288 6423 29291
rect 6638 29288 6644 29300
rect 6411 29260 6644 29288
rect 6411 29257 6423 29260
rect 6365 29251 6423 29257
rect 6638 29248 6644 29260
rect 6696 29248 6702 29300
rect 9306 29248 9312 29300
rect 9364 29288 9370 29300
rect 9493 29291 9551 29297
rect 9493 29288 9505 29291
rect 9364 29260 9505 29288
rect 9364 29248 9370 29260
rect 9493 29257 9505 29260
rect 9539 29257 9551 29291
rect 9493 29251 9551 29257
rect 9950 29248 9956 29300
rect 10008 29288 10014 29300
rect 10008 29260 10053 29288
rect 10008 29248 10014 29260
rect 10962 29248 10968 29300
rect 11020 29288 11026 29300
rect 11020 29260 11100 29288
rect 11020 29248 11026 29260
rect 8570 29152 8576 29164
rect 8531 29124 8576 29152
rect 8570 29112 8576 29124
rect 8628 29112 8634 29164
rect 8757 29155 8815 29161
rect 8757 29121 8769 29155
rect 8803 29152 8815 29155
rect 9582 29152 9588 29164
rect 8803 29124 9588 29152
rect 8803 29121 8815 29124
rect 8757 29115 8815 29121
rect 3237 29087 3295 29093
rect 3237 29053 3249 29087
rect 3283 29084 3295 29087
rect 3418 29084 3424 29096
rect 3283 29056 3424 29084
rect 3283 29053 3295 29056
rect 3237 29047 3295 29053
rect 3418 29044 3424 29056
rect 3476 29084 3482 29096
rect 3697 29087 3755 29093
rect 3697 29084 3709 29087
rect 3476 29056 3709 29084
rect 3476 29044 3482 29056
rect 3697 29053 3709 29056
rect 3743 29053 3755 29087
rect 5994 29084 6000 29096
rect 5955 29056 6000 29084
rect 3697 29047 3755 29053
rect 5994 29044 6000 29056
rect 6052 29044 6058 29096
rect 8021 29087 8079 29093
rect 8021 29053 8033 29087
rect 8067 29084 8079 29087
rect 8294 29084 8300 29096
rect 8067 29056 8300 29084
rect 8067 29053 8079 29056
rect 8021 29047 8079 29053
rect 8294 29044 8300 29056
rect 8352 29084 8358 29096
rect 8772 29084 8800 29115
rect 9582 29112 9588 29124
rect 9640 29112 9646 29164
rect 9968 29152 9996 29248
rect 9968 29124 10180 29152
rect 10045 29087 10103 29093
rect 10045 29084 10057 29087
rect 8352 29056 8800 29084
rect 9692 29056 10057 29084
rect 8352 29044 8358 29056
rect 3605 29019 3663 29025
rect 3605 28985 3617 29019
rect 3651 29016 3663 29019
rect 3964 29019 4022 29025
rect 3964 29016 3976 29019
rect 3651 28988 3976 29016
rect 3651 28985 3663 28988
rect 3605 28979 3663 28985
rect 3964 28985 3976 28988
rect 4010 29016 4022 29019
rect 4062 29016 4068 29028
rect 4010 28988 4068 29016
rect 4010 28985 4022 28988
rect 3964 28979 4022 28985
rect 4062 28976 4068 28988
rect 4120 28976 4126 29028
rect 5166 28976 5172 29028
rect 5224 28976 5230 29028
rect 6454 29016 6460 29028
rect 5552 28988 6460 29016
rect 4614 28908 4620 28960
rect 4672 28948 4678 28960
rect 5184 28948 5212 28976
rect 4672 28920 5212 28948
rect 4672 28908 4678 28920
rect 5258 28908 5264 28960
rect 5316 28948 5322 28960
rect 5552 28957 5580 28988
rect 6454 28976 6460 28988
rect 6512 28976 6518 29028
rect 8481 29019 8539 29025
rect 8481 29016 8493 29019
rect 7668 28988 8493 29016
rect 7668 28960 7696 28988
rect 8481 28985 8493 28988
rect 8527 28985 8539 29019
rect 8481 28979 8539 28985
rect 9692 28960 9720 29056
rect 10045 29053 10057 29056
rect 10091 29053 10103 29087
rect 10152 29084 10180 29124
rect 10301 29087 10359 29093
rect 10301 29084 10313 29087
rect 10152 29056 10313 29084
rect 10045 29047 10103 29053
rect 10301 29053 10313 29056
rect 10347 29053 10359 29087
rect 11072 29084 11100 29260
rect 11238 29248 11244 29300
rect 11296 29288 11302 29300
rect 12437 29291 12495 29297
rect 12437 29288 12449 29291
rect 11296 29260 12449 29288
rect 11296 29248 11302 29260
rect 12437 29257 12449 29260
rect 12483 29257 12495 29291
rect 12437 29251 12495 29257
rect 11425 29223 11483 29229
rect 11425 29189 11437 29223
rect 11471 29189 11483 29223
rect 11425 29183 11483 29189
rect 11238 29112 11244 29164
rect 11296 29152 11302 29164
rect 11440 29152 11468 29183
rect 11882 29180 11888 29232
rect 11940 29220 11946 29232
rect 12069 29223 12127 29229
rect 12069 29220 12081 29223
rect 11940 29192 12081 29220
rect 11940 29180 11946 29192
rect 12069 29189 12081 29192
rect 12115 29220 12127 29223
rect 12161 29223 12219 29229
rect 12161 29220 12173 29223
rect 12115 29192 12173 29220
rect 12115 29189 12127 29192
rect 12069 29183 12127 29189
rect 12161 29189 12173 29192
rect 12207 29189 12219 29223
rect 12161 29183 12219 29189
rect 12342 29180 12348 29232
rect 12400 29220 12406 29232
rect 13817 29223 13875 29229
rect 13817 29220 13829 29223
rect 12400 29192 13829 29220
rect 12400 29180 12406 29192
rect 13817 29189 13829 29192
rect 13863 29189 13875 29223
rect 13817 29183 13875 29189
rect 11296 29124 11468 29152
rect 11296 29112 11302 29124
rect 11974 29112 11980 29164
rect 12032 29152 12038 29164
rect 13081 29155 13139 29161
rect 13081 29152 13093 29155
rect 12032 29124 13093 29152
rect 12032 29112 12038 29124
rect 13081 29121 13093 29124
rect 13127 29152 13139 29155
rect 13449 29155 13507 29161
rect 13449 29152 13461 29155
rect 13127 29124 13461 29152
rect 13127 29121 13139 29124
rect 13081 29115 13139 29121
rect 13449 29121 13461 29124
rect 13495 29121 13507 29155
rect 13449 29115 13507 29121
rect 12805 29087 12863 29093
rect 12805 29084 12817 29087
rect 10301 29047 10359 29053
rect 10980 29056 11100 29084
rect 12176 29056 12817 29084
rect 10980 28960 11008 29056
rect 12176 29028 12204 29056
rect 12805 29053 12817 29056
rect 12851 29053 12863 29087
rect 12805 29047 12863 29053
rect 12897 29087 12955 29093
rect 12897 29053 12909 29087
rect 12943 29084 12955 29087
rect 14182 29084 14188 29096
rect 12943 29056 14188 29084
rect 12943 29053 12955 29056
rect 12897 29047 12955 29053
rect 11514 28976 11520 29028
rect 11572 29016 11578 29028
rect 11793 29019 11851 29025
rect 11793 29016 11805 29019
rect 11572 28988 11805 29016
rect 11572 28976 11578 28988
rect 11793 28985 11805 28988
rect 11839 29016 11851 29019
rect 12069 29019 12127 29025
rect 11839 28988 12020 29016
rect 11839 28985 11851 28988
rect 11793 28979 11851 28985
rect 5537 28951 5595 28957
rect 5537 28948 5549 28951
rect 5316 28920 5549 28948
rect 5316 28908 5322 28920
rect 5537 28917 5549 28920
rect 5583 28917 5595 28951
rect 7650 28948 7656 28960
rect 7611 28920 7656 28948
rect 5537 28911 5595 28917
rect 7650 28908 7656 28920
rect 7708 28908 7714 28960
rect 8110 28948 8116 28960
rect 8071 28920 8116 28948
rect 8110 28908 8116 28920
rect 8168 28908 8174 28960
rect 9217 28951 9275 28957
rect 9217 28917 9229 28951
rect 9263 28948 9275 28951
rect 9674 28948 9680 28960
rect 9263 28920 9680 28948
rect 9263 28917 9275 28920
rect 9217 28911 9275 28917
rect 9674 28908 9680 28920
rect 9732 28908 9738 28960
rect 10962 28908 10968 28960
rect 11020 28908 11026 28960
rect 11992 28948 12020 28988
rect 12069 28985 12081 29019
rect 12115 29016 12127 29019
rect 12158 29016 12164 29028
rect 12115 28988 12164 29016
rect 12115 28985 12127 28988
rect 12069 28979 12127 28985
rect 12158 28976 12164 28988
rect 12216 28976 12222 29028
rect 12912 29016 12940 29047
rect 14182 29044 14188 29056
rect 14240 29044 14246 29096
rect 12268 28988 12940 29016
rect 12268 28948 12296 28988
rect 11992 28920 12296 28948
rect 1104 28858 14812 28880
rect 1104 28806 6315 28858
rect 6367 28806 6379 28858
rect 6431 28806 6443 28858
rect 6495 28806 6507 28858
rect 6559 28806 11648 28858
rect 11700 28806 11712 28858
rect 11764 28806 11776 28858
rect 11828 28806 11840 28858
rect 11892 28806 14812 28858
rect 1104 28784 14812 28806
rect 3694 28744 3700 28756
rect 3655 28716 3700 28744
rect 3694 28704 3700 28716
rect 3752 28744 3758 28756
rect 4062 28744 4068 28756
rect 3752 28716 4068 28744
rect 3752 28704 3758 28716
rect 4062 28704 4068 28716
rect 4120 28704 4126 28756
rect 4341 28747 4399 28753
rect 4341 28713 4353 28747
rect 4387 28744 4399 28747
rect 4798 28744 4804 28756
rect 4387 28716 4804 28744
rect 4387 28713 4399 28716
rect 4341 28707 4399 28713
rect 4798 28704 4804 28716
rect 4856 28704 4862 28756
rect 5534 28704 5540 28756
rect 5592 28744 5598 28756
rect 6825 28747 6883 28753
rect 6825 28744 6837 28747
rect 5592 28716 6837 28744
rect 5592 28704 5598 28716
rect 6825 28713 6837 28716
rect 6871 28713 6883 28747
rect 6825 28707 6883 28713
rect 7650 28704 7656 28756
rect 7708 28744 7714 28756
rect 8021 28747 8079 28753
rect 8021 28744 8033 28747
rect 7708 28716 8033 28744
rect 7708 28704 7714 28716
rect 8021 28713 8033 28716
rect 8067 28713 8079 28747
rect 8021 28707 8079 28713
rect 9582 28704 9588 28756
rect 9640 28744 9646 28756
rect 11057 28747 11115 28753
rect 11057 28744 11069 28747
rect 9640 28716 11069 28744
rect 9640 28704 9646 28716
rect 11057 28713 11069 28716
rect 11103 28713 11115 28747
rect 11057 28707 11115 28713
rect 11146 28704 11152 28756
rect 11204 28744 11210 28756
rect 11977 28747 12035 28753
rect 11977 28744 11989 28747
rect 11204 28716 11989 28744
rect 11204 28704 11210 28716
rect 11977 28713 11989 28716
rect 12023 28713 12035 28747
rect 11977 28707 12035 28713
rect 12066 28704 12072 28756
rect 12124 28744 12130 28756
rect 12437 28747 12495 28753
rect 12437 28744 12449 28747
rect 12124 28716 12449 28744
rect 12124 28704 12130 28716
rect 12437 28713 12449 28716
rect 12483 28713 12495 28747
rect 12986 28744 12992 28756
rect 12947 28716 12992 28744
rect 12437 28707 12495 28713
rect 12986 28704 12992 28716
rect 13044 28704 13050 28756
rect 9493 28679 9551 28685
rect 9493 28645 9505 28679
rect 9539 28676 9551 28679
rect 9674 28676 9680 28688
rect 9539 28648 9680 28676
rect 9539 28645 9551 28648
rect 9493 28639 9551 28645
rect 9674 28636 9680 28648
rect 9732 28676 9738 28688
rect 10226 28676 10232 28688
rect 9732 28648 10232 28676
rect 9732 28636 9738 28648
rect 10226 28636 10232 28648
rect 10284 28636 10290 28688
rect 5258 28568 5264 28620
rect 5316 28608 5322 28620
rect 5701 28611 5759 28617
rect 5701 28608 5713 28611
rect 5316 28580 5713 28608
rect 5316 28568 5322 28580
rect 5701 28577 5713 28580
rect 5747 28577 5759 28611
rect 8386 28608 8392 28620
rect 8347 28580 8392 28608
rect 5701 28571 5759 28577
rect 8386 28568 8392 28580
rect 8444 28568 8450 28620
rect 9933 28611 9991 28617
rect 9933 28608 9945 28611
rect 9416 28580 9945 28608
rect 9416 28552 9444 28580
rect 9933 28577 9945 28580
rect 9979 28577 9991 28611
rect 12342 28608 12348 28620
rect 12303 28580 12348 28608
rect 9933 28571 9991 28577
rect 12342 28568 12348 28580
rect 12400 28568 12406 28620
rect 5445 28543 5503 28549
rect 5445 28509 5457 28543
rect 5491 28509 5503 28543
rect 8478 28540 8484 28552
rect 8439 28512 8484 28540
rect 5445 28503 5503 28509
rect 5460 28416 5488 28503
rect 8478 28500 8484 28512
rect 8536 28500 8542 28552
rect 8665 28543 8723 28549
rect 8665 28509 8677 28543
rect 8711 28540 8723 28543
rect 9033 28543 9091 28549
rect 9033 28540 9045 28543
rect 8711 28512 9045 28540
rect 8711 28509 8723 28512
rect 8665 28503 8723 28509
rect 9033 28509 9045 28512
rect 9079 28540 9091 28543
rect 9398 28540 9404 28552
rect 9079 28512 9404 28540
rect 9079 28509 9091 28512
rect 9033 28503 9091 28509
rect 7929 28475 7987 28481
rect 7929 28441 7941 28475
rect 7975 28472 7987 28475
rect 8680 28472 8708 28503
rect 9398 28500 9404 28512
rect 9456 28500 9462 28552
rect 9674 28540 9680 28552
rect 9635 28512 9680 28540
rect 9674 28500 9680 28512
rect 9732 28500 9738 28552
rect 11974 28500 11980 28552
rect 12032 28540 12038 28552
rect 12434 28540 12440 28552
rect 12032 28512 12440 28540
rect 12032 28500 12038 28512
rect 12434 28500 12440 28512
rect 12492 28540 12498 28552
rect 12529 28543 12587 28549
rect 12529 28540 12541 28543
rect 12492 28512 12541 28540
rect 12492 28500 12498 28512
rect 12529 28509 12541 28512
rect 12575 28509 12587 28543
rect 12529 28503 12587 28509
rect 7975 28444 8708 28472
rect 7975 28441 7987 28444
rect 7929 28435 7987 28441
rect 4709 28407 4767 28413
rect 4709 28373 4721 28407
rect 4755 28404 4767 28407
rect 4982 28404 4988 28416
rect 4755 28376 4988 28404
rect 4755 28373 4767 28376
rect 4709 28367 4767 28373
rect 4982 28364 4988 28376
rect 5040 28364 5046 28416
rect 5258 28404 5264 28416
rect 5219 28376 5264 28404
rect 5258 28364 5264 28376
rect 5316 28364 5322 28416
rect 5442 28404 5448 28416
rect 5355 28376 5448 28404
rect 5442 28364 5448 28376
rect 5500 28404 5506 28416
rect 6178 28404 6184 28416
rect 5500 28376 6184 28404
rect 5500 28364 5506 28376
rect 6178 28364 6184 28376
rect 6236 28404 6242 28416
rect 6822 28404 6828 28416
rect 6236 28376 6828 28404
rect 6236 28364 6242 28376
rect 6822 28364 6828 28376
rect 6880 28364 6886 28416
rect 1104 28314 14812 28336
rect 1104 28262 3648 28314
rect 3700 28262 3712 28314
rect 3764 28262 3776 28314
rect 3828 28262 3840 28314
rect 3892 28262 8982 28314
rect 9034 28262 9046 28314
rect 9098 28262 9110 28314
rect 9162 28262 9174 28314
rect 9226 28262 14315 28314
rect 14367 28262 14379 28314
rect 14431 28262 14443 28314
rect 14495 28262 14507 28314
rect 14559 28262 14812 28314
rect 1104 28240 14812 28262
rect 3510 28160 3516 28212
rect 3568 28200 3574 28212
rect 3605 28203 3663 28209
rect 3605 28200 3617 28203
rect 3568 28172 3617 28200
rect 3568 28160 3574 28172
rect 3605 28169 3617 28172
rect 3651 28169 3663 28203
rect 3605 28163 3663 28169
rect 4246 28160 4252 28212
rect 4304 28200 4310 28212
rect 4709 28203 4767 28209
rect 4709 28200 4721 28203
rect 4304 28172 4721 28200
rect 4304 28160 4310 28172
rect 4709 28169 4721 28172
rect 4755 28200 4767 28203
rect 5442 28200 5448 28212
rect 4755 28172 5448 28200
rect 4755 28169 4767 28172
rect 4709 28163 4767 28169
rect 5442 28160 5448 28172
rect 5500 28160 5506 28212
rect 5994 28160 6000 28212
rect 6052 28200 6058 28212
rect 6178 28200 6184 28212
rect 6052 28172 6184 28200
rect 6052 28160 6058 28172
rect 6178 28160 6184 28172
rect 6236 28160 6242 28212
rect 8570 28160 8576 28212
rect 8628 28200 8634 28212
rect 9033 28203 9091 28209
rect 9033 28200 9045 28203
rect 8628 28172 9045 28200
rect 8628 28160 8634 28172
rect 9033 28169 9045 28172
rect 9079 28169 9091 28203
rect 10778 28200 10784 28212
rect 10739 28172 10784 28200
rect 9033 28163 9091 28169
rect 10778 28160 10784 28172
rect 10836 28160 10842 28212
rect 12066 28200 12072 28212
rect 12027 28172 12072 28200
rect 12066 28160 12072 28172
rect 12124 28160 12130 28212
rect 8846 28132 8852 28144
rect 8807 28104 8852 28132
rect 8846 28092 8852 28104
rect 8904 28092 8910 28144
rect 10686 28132 10692 28144
rect 10647 28104 10692 28132
rect 10686 28092 10692 28104
rect 10744 28132 10750 28144
rect 10744 28104 11376 28132
rect 10744 28092 10750 28104
rect 1578 28064 1584 28076
rect 1539 28036 1584 28064
rect 1578 28024 1584 28036
rect 1636 28024 1642 28076
rect 4062 28064 4068 28076
rect 4023 28036 4068 28064
rect 4062 28024 4068 28036
rect 4120 28024 4126 28076
rect 4154 28024 4160 28076
rect 4212 28064 4218 28076
rect 4212 28036 4257 28064
rect 4212 28024 4218 28036
rect 5258 28024 5264 28076
rect 5316 28064 5322 28076
rect 5813 28067 5871 28073
rect 5813 28064 5825 28067
rect 5316 28036 5825 28064
rect 5316 28024 5322 28036
rect 5813 28033 5825 28036
rect 5859 28064 5871 28067
rect 5994 28064 6000 28076
rect 5859 28036 6000 28064
rect 5859 28033 5871 28036
rect 5813 28027 5871 28033
rect 5994 28024 6000 28036
rect 6052 28024 6058 28076
rect 11348 28073 11376 28104
rect 9585 28067 9643 28073
rect 9585 28033 9597 28067
rect 9631 28064 9643 28067
rect 11333 28067 11391 28073
rect 9631 28036 9665 28064
rect 9631 28033 9643 28036
rect 9585 28027 9643 28033
rect 11333 28033 11345 28067
rect 11379 28033 11391 28067
rect 11333 28027 11391 28033
rect 1397 27999 1455 28005
rect 1397 27965 1409 27999
rect 1443 27996 1455 27999
rect 3513 27999 3571 28005
rect 1443 27968 2268 27996
rect 1443 27965 1455 27968
rect 1397 27959 1455 27965
rect 2240 27872 2268 27968
rect 3513 27965 3525 27999
rect 3559 27996 3571 27999
rect 3973 27999 4031 28005
rect 3973 27996 3985 27999
rect 3559 27968 3985 27996
rect 3559 27965 3571 27968
rect 3513 27959 3571 27965
rect 3973 27965 3985 27968
rect 4019 27996 4031 27999
rect 4614 27996 4620 28008
rect 4019 27968 4620 27996
rect 4019 27965 4031 27968
rect 3973 27959 4031 27965
rect 4614 27956 4620 27968
rect 4672 27956 4678 28008
rect 5629 27999 5687 28005
rect 5629 27996 5641 27999
rect 5092 27968 5641 27996
rect 5092 27940 5120 27968
rect 5629 27965 5641 27968
rect 5675 27996 5687 27999
rect 5718 27996 5724 28008
rect 5675 27968 5724 27996
rect 5675 27965 5687 27968
rect 5629 27959 5687 27965
rect 5718 27956 5724 27968
rect 5776 27956 5782 28008
rect 6822 27996 6828 28008
rect 6783 27968 6828 27996
rect 6822 27956 6828 27968
rect 6880 27956 6886 28008
rect 9398 27956 9404 28008
rect 9456 27996 9462 28008
rect 9600 27996 9628 28027
rect 12066 28024 12072 28076
rect 12124 28064 12130 28076
rect 12342 28064 12348 28076
rect 12124 28036 12348 28064
rect 12124 28024 12130 28036
rect 12342 28024 12348 28036
rect 12400 28064 12406 28076
rect 12437 28067 12495 28073
rect 12437 28064 12449 28067
rect 12400 28036 12449 28064
rect 12400 28024 12406 28036
rect 12437 28033 12449 28036
rect 12483 28033 12495 28067
rect 12437 28027 12495 28033
rect 10045 27999 10103 28005
rect 10045 27996 10057 27999
rect 9456 27968 10057 27996
rect 9456 27956 9462 27968
rect 10045 27965 10057 27968
rect 10091 27965 10103 27999
rect 10045 27959 10103 27965
rect 5074 27928 5080 27940
rect 5035 27900 5080 27928
rect 5074 27888 5080 27900
rect 5132 27888 5138 27940
rect 5534 27928 5540 27940
rect 5495 27900 5540 27928
rect 5534 27888 5540 27900
rect 5592 27888 5598 27940
rect 6641 27931 6699 27937
rect 6641 27897 6653 27931
rect 6687 27928 6699 27931
rect 7006 27928 7012 27940
rect 6687 27900 7012 27928
rect 6687 27897 6699 27900
rect 6641 27891 6699 27897
rect 7006 27888 7012 27900
rect 7064 27937 7070 27940
rect 7064 27931 7128 27937
rect 7064 27897 7082 27931
rect 7116 27897 7128 27931
rect 7064 27891 7128 27897
rect 7064 27888 7070 27891
rect 8478 27888 8484 27940
rect 8536 27928 8542 27940
rect 8573 27931 8631 27937
rect 8573 27928 8585 27931
rect 8536 27900 8585 27928
rect 8536 27888 8542 27900
rect 8573 27897 8585 27900
rect 8619 27928 8631 27931
rect 9582 27928 9588 27940
rect 8619 27900 9588 27928
rect 8619 27897 8631 27900
rect 8573 27891 8631 27897
rect 9582 27888 9588 27900
rect 9640 27888 9646 27940
rect 11149 27931 11207 27937
rect 11149 27897 11161 27931
rect 11195 27928 11207 27931
rect 11422 27928 11428 27940
rect 11195 27900 11428 27928
rect 11195 27897 11207 27900
rect 11149 27891 11207 27897
rect 11422 27888 11428 27900
rect 11480 27888 11486 27940
rect 2222 27860 2228 27872
rect 2183 27832 2228 27860
rect 2222 27820 2228 27832
rect 2280 27820 2286 27872
rect 5166 27860 5172 27872
rect 5127 27832 5172 27860
rect 5166 27820 5172 27832
rect 5224 27820 5230 27872
rect 5994 27820 6000 27872
rect 6052 27860 6058 27872
rect 6181 27863 6239 27869
rect 6181 27860 6193 27863
rect 6052 27832 6193 27860
rect 6052 27820 6058 27832
rect 6181 27829 6193 27832
rect 6227 27860 6239 27863
rect 8205 27863 8263 27869
rect 8205 27860 8217 27863
rect 6227 27832 8217 27860
rect 6227 27829 6239 27832
rect 6181 27823 6239 27829
rect 8205 27829 8217 27832
rect 8251 27829 8263 27863
rect 8205 27823 8263 27829
rect 8846 27820 8852 27872
rect 8904 27860 8910 27872
rect 9306 27860 9312 27872
rect 8904 27832 9312 27860
rect 8904 27820 8910 27832
rect 9306 27820 9312 27832
rect 9364 27860 9370 27872
rect 9401 27863 9459 27869
rect 9401 27860 9413 27863
rect 9364 27832 9413 27860
rect 9364 27820 9370 27832
rect 9401 27829 9413 27832
rect 9447 27829 9459 27863
rect 9401 27823 9459 27829
rect 9490 27820 9496 27872
rect 9548 27860 9554 27872
rect 11238 27860 11244 27872
rect 9548 27832 9593 27860
rect 11199 27832 11244 27860
rect 9548 27820 9554 27832
rect 11238 27820 11244 27832
rect 11296 27820 11302 27872
rect 1104 27770 14812 27792
rect 1104 27718 6315 27770
rect 6367 27718 6379 27770
rect 6431 27718 6443 27770
rect 6495 27718 6507 27770
rect 6559 27718 11648 27770
rect 11700 27718 11712 27770
rect 11764 27718 11776 27770
rect 11828 27718 11840 27770
rect 11892 27718 14812 27770
rect 1104 27696 14812 27718
rect 3697 27659 3755 27665
rect 3697 27625 3709 27659
rect 3743 27656 3755 27659
rect 4062 27656 4068 27668
rect 3743 27628 4068 27656
rect 3743 27625 3755 27628
rect 3697 27619 3755 27625
rect 4062 27616 4068 27628
rect 4120 27616 4126 27668
rect 4706 27616 4712 27668
rect 4764 27656 4770 27668
rect 5261 27659 5319 27665
rect 5261 27656 5273 27659
rect 4764 27628 5273 27656
rect 4764 27616 4770 27628
rect 5261 27625 5273 27628
rect 5307 27656 5319 27659
rect 5534 27656 5540 27668
rect 5307 27628 5540 27656
rect 5307 27625 5319 27628
rect 5261 27619 5319 27625
rect 5534 27616 5540 27628
rect 5592 27616 5598 27668
rect 8386 27616 8392 27668
rect 8444 27656 8450 27668
rect 8665 27659 8723 27665
rect 8665 27656 8677 27659
rect 8444 27628 8677 27656
rect 8444 27616 8450 27628
rect 8665 27625 8677 27628
rect 8711 27625 8723 27659
rect 8665 27619 8723 27625
rect 11057 27659 11115 27665
rect 11057 27625 11069 27659
rect 11103 27656 11115 27659
rect 11238 27656 11244 27668
rect 11103 27628 11244 27656
rect 11103 27625 11115 27628
rect 11057 27619 11115 27625
rect 3050 27548 3056 27600
rect 3108 27588 3114 27600
rect 3326 27588 3332 27600
rect 3108 27560 3332 27588
rect 3108 27548 3114 27560
rect 3326 27548 3332 27560
rect 3384 27548 3390 27600
rect 8680 27588 8708 27619
rect 11238 27616 11244 27628
rect 11296 27616 11302 27668
rect 12066 27656 12072 27668
rect 12027 27628 12072 27656
rect 12066 27616 12072 27628
rect 12124 27616 12130 27668
rect 12434 27656 12440 27668
rect 12395 27628 12440 27656
rect 12434 27616 12440 27628
rect 12492 27616 12498 27668
rect 9677 27591 9735 27597
rect 9677 27588 9689 27591
rect 8680 27560 9689 27588
rect 9677 27557 9689 27560
rect 9723 27557 9735 27591
rect 9677 27551 9735 27557
rect 5810 27520 5816 27532
rect 5771 27492 5816 27520
rect 5810 27480 5816 27492
rect 5868 27480 5874 27532
rect 6638 27480 6644 27532
rect 6696 27520 6702 27532
rect 7276 27523 7334 27529
rect 7276 27520 7288 27523
rect 6696 27492 7288 27520
rect 6696 27480 6702 27492
rect 7276 27489 7288 27492
rect 7322 27520 7334 27523
rect 8202 27520 8208 27532
rect 7322 27492 8208 27520
rect 7322 27489 7334 27492
rect 7276 27483 7334 27489
rect 8202 27480 8208 27492
rect 8260 27480 8266 27532
rect 5534 27412 5540 27464
rect 5592 27452 5598 27464
rect 5905 27455 5963 27461
rect 5905 27452 5917 27455
rect 5592 27424 5917 27452
rect 5592 27412 5598 27424
rect 5905 27421 5917 27424
rect 5951 27421 5963 27455
rect 5905 27415 5963 27421
rect 5994 27412 6000 27464
rect 6052 27452 6058 27464
rect 6052 27424 6097 27452
rect 6052 27412 6058 27424
rect 6822 27412 6828 27464
rect 6880 27452 6886 27464
rect 7009 27455 7067 27461
rect 7009 27452 7021 27455
rect 6880 27424 7021 27452
rect 6880 27412 6886 27424
rect 7009 27421 7021 27424
rect 7055 27421 7067 27455
rect 7009 27415 7067 27421
rect 5350 27276 5356 27328
rect 5408 27316 5414 27328
rect 5445 27319 5503 27325
rect 5445 27316 5457 27319
rect 5408 27288 5457 27316
rect 5408 27276 5414 27288
rect 5445 27285 5457 27288
rect 5491 27285 5503 27319
rect 5445 27279 5503 27285
rect 6917 27319 6975 27325
rect 6917 27285 6929 27319
rect 6963 27316 6975 27319
rect 7024 27316 7052 27415
rect 8202 27316 8208 27328
rect 6963 27288 8208 27316
rect 6963 27285 6975 27288
rect 6917 27279 6975 27285
rect 8202 27276 8208 27288
rect 8260 27276 8266 27328
rect 8386 27316 8392 27328
rect 8347 27288 8392 27316
rect 8386 27276 8392 27288
rect 8444 27276 8450 27328
rect 8662 27276 8668 27328
rect 8720 27316 8726 27328
rect 9033 27319 9091 27325
rect 9033 27316 9045 27319
rect 8720 27288 9045 27316
rect 8720 27276 8726 27288
rect 9033 27285 9045 27288
rect 9079 27316 9091 27319
rect 9490 27316 9496 27328
rect 9079 27288 9496 27316
rect 9079 27285 9091 27288
rect 9033 27279 9091 27285
rect 9490 27276 9496 27288
rect 9548 27276 9554 27328
rect 10226 27316 10232 27328
rect 10187 27288 10232 27316
rect 10226 27276 10232 27288
rect 10284 27276 10290 27328
rect 10686 27316 10692 27328
rect 10647 27288 10692 27316
rect 10686 27276 10692 27288
rect 10744 27276 10750 27328
rect 11422 27316 11428 27328
rect 11383 27288 11428 27316
rect 11422 27276 11428 27288
rect 11480 27276 11486 27328
rect 1104 27226 14812 27248
rect 1104 27174 3648 27226
rect 3700 27174 3712 27226
rect 3764 27174 3776 27226
rect 3828 27174 3840 27226
rect 3892 27174 8982 27226
rect 9034 27174 9046 27226
rect 9098 27174 9110 27226
rect 9162 27174 9174 27226
rect 9226 27174 14315 27226
rect 14367 27174 14379 27226
rect 14431 27174 14443 27226
rect 14495 27174 14507 27226
rect 14559 27174 14812 27226
rect 1104 27152 14812 27174
rect 4982 27112 4988 27124
rect 4943 27084 4988 27112
rect 4982 27072 4988 27084
rect 5040 27072 5046 27124
rect 6638 27112 6644 27124
rect 6599 27084 6644 27112
rect 6638 27072 6644 27084
rect 6696 27072 6702 27124
rect 7006 27112 7012 27124
rect 6967 27084 7012 27112
rect 7006 27072 7012 27084
rect 7064 27072 7070 27124
rect 7190 27112 7196 27124
rect 7151 27084 7196 27112
rect 7190 27072 7196 27084
rect 7248 27072 7254 27124
rect 8202 27112 8208 27124
rect 8163 27084 8208 27112
rect 8202 27072 8208 27084
rect 8260 27072 8266 27124
rect 10597 27115 10655 27121
rect 10597 27081 10609 27115
rect 10643 27112 10655 27115
rect 11238 27112 11244 27124
rect 10643 27084 11244 27112
rect 10643 27081 10655 27084
rect 10597 27075 10655 27081
rect 11238 27072 11244 27084
rect 11296 27072 11302 27124
rect 12802 27072 12808 27124
rect 12860 27112 12866 27124
rect 12860 27084 12940 27112
rect 12860 27072 12866 27084
rect 4893 27047 4951 27053
rect 4893 27013 4905 27047
rect 4939 27044 4951 27047
rect 5994 27044 6000 27056
rect 4939 27016 6000 27044
rect 4939 27013 4951 27016
rect 4893 27007 4951 27013
rect 5994 27004 6000 27016
rect 6052 27004 6058 27056
rect 4525 26979 4583 26985
rect 4525 26945 4537 26979
rect 4571 26976 4583 26979
rect 5166 26976 5172 26988
rect 4571 26948 5172 26976
rect 4571 26945 4583 26948
rect 4525 26939 4583 26945
rect 5166 26936 5172 26948
rect 5224 26976 5230 26988
rect 5445 26979 5503 26985
rect 5445 26976 5457 26979
rect 5224 26948 5457 26976
rect 5224 26936 5230 26948
rect 5445 26945 5457 26948
rect 5491 26945 5503 26979
rect 5445 26939 5503 26945
rect 5537 26979 5595 26985
rect 5537 26945 5549 26979
rect 5583 26945 5595 26979
rect 7024 26976 7052 27072
rect 7745 26979 7803 26985
rect 7745 26976 7757 26979
rect 7024 26948 7757 26976
rect 5537 26939 5595 26945
rect 7745 26945 7757 26948
rect 7791 26976 7803 26979
rect 8386 26976 8392 26988
rect 7791 26948 8392 26976
rect 7791 26945 7803 26948
rect 7745 26939 7803 26945
rect 4157 26911 4215 26917
rect 4157 26877 4169 26911
rect 4203 26908 4215 26911
rect 5350 26908 5356 26920
rect 4203 26880 5356 26908
rect 4203 26877 4215 26880
rect 4157 26871 4215 26877
rect 5350 26868 5356 26880
rect 5408 26868 5414 26920
rect 5552 26908 5580 26939
rect 8386 26936 8392 26948
rect 8444 26936 8450 26988
rect 10505 26979 10563 26985
rect 10505 26945 10517 26979
rect 10551 26976 10563 26979
rect 11241 26979 11299 26985
rect 11241 26976 11253 26979
rect 10551 26948 11253 26976
rect 10551 26945 10563 26948
rect 10505 26939 10563 26945
rect 11241 26945 11253 26948
rect 11287 26976 11299 26979
rect 12434 26976 12440 26988
rect 11287 26948 12440 26976
rect 11287 26945 11299 26948
rect 11241 26939 11299 26945
rect 12434 26936 12440 26948
rect 12492 26936 12498 26988
rect 12912 26920 12940 27084
rect 7558 26908 7564 26920
rect 5460 26880 5580 26908
rect 7471 26880 7564 26908
rect 4982 26800 4988 26852
rect 5040 26840 5046 26852
rect 5460 26840 5488 26880
rect 7558 26868 7564 26880
rect 7616 26908 7622 26920
rect 8110 26908 8116 26920
rect 7616 26880 8116 26908
rect 7616 26868 7622 26880
rect 8110 26868 8116 26880
rect 8168 26868 8174 26920
rect 12894 26868 12900 26920
rect 12952 26868 12958 26920
rect 5040 26812 5488 26840
rect 5040 26800 5046 26812
rect 7282 26800 7288 26852
rect 7340 26840 7346 26852
rect 7653 26843 7711 26849
rect 7653 26840 7665 26843
rect 7340 26812 7665 26840
rect 7340 26800 7346 26812
rect 7653 26809 7665 26812
rect 7699 26809 7711 26843
rect 10965 26843 11023 26849
rect 10965 26840 10977 26843
rect 7653 26803 7711 26809
rect 10152 26812 10977 26840
rect 10152 26784 10180 26812
rect 10965 26809 10977 26812
rect 11011 26809 11023 26843
rect 10965 26803 11023 26809
rect 5534 26732 5540 26784
rect 5592 26772 5598 26784
rect 5997 26775 6055 26781
rect 5997 26772 6009 26775
rect 5592 26744 6009 26772
rect 5592 26732 5598 26744
rect 5997 26741 6009 26744
rect 6043 26741 6055 26775
rect 10134 26772 10140 26784
rect 10095 26744 10140 26772
rect 5997 26735 6055 26741
rect 10134 26732 10140 26744
rect 10192 26732 10198 26784
rect 10686 26732 10692 26784
rect 10744 26772 10750 26784
rect 11057 26775 11115 26781
rect 11057 26772 11069 26775
rect 10744 26744 11069 26772
rect 10744 26732 10750 26744
rect 11057 26741 11069 26744
rect 11103 26741 11115 26775
rect 11057 26735 11115 26741
rect 1104 26682 14812 26704
rect 1104 26630 6315 26682
rect 6367 26630 6379 26682
rect 6431 26630 6443 26682
rect 6495 26630 6507 26682
rect 6559 26630 11648 26682
rect 11700 26630 11712 26682
rect 11764 26630 11776 26682
rect 11828 26630 11840 26682
rect 11892 26630 14812 26682
rect 1104 26608 14812 26630
rect 4062 26528 4068 26580
rect 4120 26568 4126 26580
rect 4982 26568 4988 26580
rect 4120 26540 4988 26568
rect 4120 26528 4126 26540
rect 4982 26528 4988 26540
rect 5040 26528 5046 26580
rect 7558 26568 7564 26580
rect 7519 26540 7564 26568
rect 7558 26528 7564 26540
rect 7616 26528 7622 26580
rect 10134 26528 10140 26580
rect 10192 26568 10198 26580
rect 10413 26571 10471 26577
rect 10413 26568 10425 26571
rect 10192 26540 10425 26568
rect 10192 26528 10198 26540
rect 10413 26537 10425 26540
rect 10459 26537 10471 26571
rect 10413 26531 10471 26537
rect 11422 26528 11428 26580
rect 11480 26568 11486 26580
rect 11977 26571 12035 26577
rect 11977 26568 11989 26571
rect 11480 26540 11989 26568
rect 11480 26528 11486 26540
rect 11977 26537 11989 26540
rect 12023 26537 12035 26571
rect 11977 26531 12035 26537
rect 12437 26571 12495 26577
rect 12437 26537 12449 26571
rect 12483 26568 12495 26571
rect 12986 26568 12992 26580
rect 12483 26540 12992 26568
rect 12483 26537 12495 26540
rect 12437 26531 12495 26537
rect 12986 26528 12992 26540
rect 13044 26528 13050 26580
rect 10318 26460 10324 26512
rect 10376 26500 10382 26512
rect 10778 26500 10784 26512
rect 10376 26472 10784 26500
rect 10376 26460 10382 26472
rect 10778 26460 10784 26472
rect 10836 26460 10842 26512
rect 10410 26392 10416 26444
rect 10468 26432 10474 26444
rect 10873 26435 10931 26441
rect 10873 26432 10885 26435
rect 10468 26404 10885 26432
rect 10468 26392 10474 26404
rect 10873 26401 10885 26404
rect 10919 26401 10931 26435
rect 10873 26395 10931 26401
rect 11146 26392 11152 26444
rect 11204 26432 11210 26444
rect 11974 26432 11980 26444
rect 11204 26404 11980 26432
rect 11204 26392 11210 26404
rect 11974 26392 11980 26404
rect 12032 26432 12038 26444
rect 12345 26435 12403 26441
rect 12345 26432 12357 26435
rect 12032 26404 12357 26432
rect 12032 26392 12038 26404
rect 12345 26401 12357 26404
rect 12391 26401 12403 26435
rect 12345 26395 12403 26401
rect 10321 26367 10379 26373
rect 10321 26333 10333 26367
rect 10367 26364 10379 26367
rect 10965 26367 11023 26373
rect 10965 26364 10977 26367
rect 10367 26336 10977 26364
rect 10367 26333 10379 26336
rect 10321 26327 10379 26333
rect 10965 26333 10977 26336
rect 11011 26364 11023 26367
rect 11054 26364 11060 26376
rect 11011 26336 11060 26364
rect 11011 26333 11023 26336
rect 10965 26327 11023 26333
rect 11054 26324 11060 26336
rect 11112 26324 11118 26376
rect 12434 26324 12440 26376
rect 12492 26364 12498 26376
rect 12529 26367 12587 26373
rect 12529 26364 12541 26367
rect 12492 26336 12541 26364
rect 12492 26324 12498 26336
rect 12529 26333 12541 26336
rect 12575 26333 12587 26367
rect 12529 26327 12587 26333
rect 8941 26299 8999 26305
rect 8941 26265 8953 26299
rect 8987 26296 8999 26299
rect 9398 26296 9404 26308
rect 8987 26268 9404 26296
rect 8987 26265 8999 26268
rect 8941 26259 8999 26265
rect 9398 26256 9404 26268
rect 9456 26256 9462 26308
rect 5537 26231 5595 26237
rect 5537 26197 5549 26231
rect 5583 26228 5595 26231
rect 5810 26228 5816 26240
rect 5583 26200 5816 26228
rect 5583 26197 5595 26200
rect 5537 26191 5595 26197
rect 5810 26188 5816 26200
rect 5868 26228 5874 26240
rect 7006 26228 7012 26240
rect 5868 26200 7012 26228
rect 5868 26188 5874 26200
rect 7006 26188 7012 26200
rect 7064 26188 7070 26240
rect 7282 26228 7288 26240
rect 7243 26200 7288 26228
rect 7282 26188 7288 26200
rect 7340 26188 7346 26240
rect 8570 26228 8576 26240
rect 8531 26200 8576 26228
rect 8570 26188 8576 26200
rect 8628 26188 8634 26240
rect 9309 26231 9367 26237
rect 9309 26197 9321 26231
rect 9355 26228 9367 26231
rect 9582 26228 9588 26240
rect 9355 26200 9588 26228
rect 9355 26197 9367 26200
rect 9309 26191 9367 26197
rect 9582 26188 9588 26200
rect 9640 26188 9646 26240
rect 1104 26138 14812 26160
rect 1104 26086 3648 26138
rect 3700 26086 3712 26138
rect 3764 26086 3776 26138
rect 3828 26086 3840 26138
rect 3892 26086 8982 26138
rect 9034 26086 9046 26138
rect 9098 26086 9110 26138
rect 9162 26086 9174 26138
rect 9226 26086 14315 26138
rect 14367 26086 14379 26138
rect 14431 26086 14443 26138
rect 14495 26086 14507 26138
rect 14559 26086 14812 26138
rect 1104 26064 14812 26086
rect 6181 26027 6239 26033
rect 6181 25993 6193 26027
rect 6227 26024 6239 26027
rect 6822 26024 6828 26036
rect 6227 25996 6828 26024
rect 6227 25993 6239 25996
rect 6181 25987 6239 25993
rect 6822 25984 6828 25996
rect 6880 25984 6886 26036
rect 8481 26027 8539 26033
rect 8481 25993 8493 26027
rect 8527 26024 8539 26027
rect 10226 26024 10232 26036
rect 8527 25996 10232 26024
rect 8527 25993 8539 25996
rect 8481 25987 8539 25993
rect 10226 25984 10232 25996
rect 10284 25984 10290 26036
rect 10413 26027 10471 26033
rect 10413 25993 10425 26027
rect 10459 26024 10471 26027
rect 10686 26024 10692 26036
rect 10459 25996 10692 26024
rect 10459 25993 10471 25996
rect 10413 25987 10471 25993
rect 10686 25984 10692 25996
rect 10744 25984 10750 26036
rect 10778 25984 10784 26036
rect 10836 26024 10842 26036
rect 11425 26027 11483 26033
rect 11425 26024 11437 26027
rect 10836 25996 11437 26024
rect 10836 25984 10842 25996
rect 11425 25993 11437 25996
rect 11471 25993 11483 26027
rect 11974 26024 11980 26036
rect 11935 25996 11980 26024
rect 11425 25987 11483 25993
rect 11974 25984 11980 25996
rect 12032 25984 12038 26036
rect 12434 25984 12440 26036
rect 12492 26024 12498 26036
rect 12621 26027 12679 26033
rect 12621 26024 12633 26027
rect 12492 25996 12633 26024
rect 12492 25984 12498 25996
rect 12621 25993 12633 25996
rect 12667 25993 12679 26027
rect 12621 25987 12679 25993
rect 10962 25916 10968 25968
rect 11020 25956 11026 25968
rect 11146 25956 11152 25968
rect 11020 25928 11152 25956
rect 11020 25916 11026 25928
rect 11146 25916 11152 25928
rect 11204 25916 11210 25968
rect 8389 25891 8447 25897
rect 8389 25857 8401 25891
rect 8435 25888 8447 25891
rect 9306 25888 9312 25900
rect 8435 25860 9312 25888
rect 8435 25857 8447 25860
rect 8389 25851 8447 25857
rect 9306 25848 9312 25860
rect 9364 25848 9370 25900
rect 9398 25848 9404 25900
rect 9456 25888 9462 25900
rect 9493 25891 9551 25897
rect 9493 25888 9505 25891
rect 9456 25860 9505 25888
rect 9456 25848 9462 25860
rect 9493 25857 9505 25860
rect 9539 25888 9551 25891
rect 9766 25888 9772 25900
rect 9539 25860 9772 25888
rect 9539 25857 9551 25860
rect 9493 25851 9551 25857
rect 9766 25848 9772 25860
rect 9824 25848 9830 25900
rect 11054 25888 11060 25900
rect 11015 25860 11060 25888
rect 11054 25848 11060 25860
rect 11112 25848 11118 25900
rect 5626 25780 5632 25832
rect 5684 25820 5690 25832
rect 6365 25823 6423 25829
rect 6365 25820 6377 25823
rect 5684 25792 6377 25820
rect 5684 25780 5690 25792
rect 6365 25789 6377 25792
rect 6411 25820 6423 25823
rect 7009 25823 7067 25829
rect 7009 25820 7021 25823
rect 6411 25792 7021 25820
rect 6411 25789 6423 25792
rect 6365 25783 6423 25789
rect 7009 25789 7021 25792
rect 7055 25789 7067 25823
rect 7009 25783 7067 25789
rect 8570 25780 8576 25832
rect 8628 25820 8634 25832
rect 8665 25823 8723 25829
rect 8665 25820 8677 25823
rect 8628 25792 8677 25820
rect 8628 25780 8634 25792
rect 8665 25789 8677 25792
rect 8711 25789 8723 25823
rect 8665 25783 8723 25789
rect 9953 25823 10011 25829
rect 9953 25789 9965 25823
rect 9999 25820 10011 25823
rect 10410 25820 10416 25832
rect 9999 25792 10416 25820
rect 9999 25789 10011 25792
rect 9953 25783 10011 25789
rect 10410 25780 10416 25792
rect 10468 25780 10474 25832
rect 10502 25780 10508 25832
rect 10560 25820 10566 25832
rect 10781 25823 10839 25829
rect 10781 25820 10793 25823
rect 10560 25792 10793 25820
rect 10560 25780 10566 25792
rect 10781 25789 10793 25792
rect 10827 25789 10839 25823
rect 10781 25783 10839 25789
rect 7929 25755 7987 25761
rect 7929 25721 7941 25755
rect 7975 25752 7987 25755
rect 9217 25755 9275 25761
rect 7975 25724 8892 25752
rect 7975 25721 7987 25724
rect 7929 25715 7987 25721
rect 8864 25696 8892 25724
rect 9217 25721 9229 25755
rect 9263 25752 9275 25755
rect 9582 25752 9588 25764
rect 9263 25724 9588 25752
rect 9263 25721 9275 25724
rect 9217 25715 9275 25721
rect 9582 25712 9588 25724
rect 9640 25712 9646 25764
rect 10594 25712 10600 25764
rect 10652 25752 10658 25764
rect 10962 25752 10968 25764
rect 10652 25724 10968 25752
rect 10652 25712 10658 25724
rect 10962 25712 10968 25724
rect 11020 25712 11026 25764
rect 5994 25644 6000 25696
rect 6052 25684 6058 25696
rect 6178 25684 6184 25696
rect 6052 25656 6184 25684
rect 6052 25644 6058 25656
rect 6178 25644 6184 25656
rect 6236 25644 6242 25696
rect 8846 25684 8852 25696
rect 8807 25656 8852 25684
rect 8846 25644 8852 25656
rect 8904 25644 8910 25696
rect 9950 25644 9956 25696
rect 10008 25684 10014 25696
rect 10229 25687 10287 25693
rect 10229 25684 10241 25687
rect 10008 25656 10241 25684
rect 10008 25644 10014 25656
rect 10229 25653 10241 25656
rect 10275 25684 10287 25687
rect 10873 25687 10931 25693
rect 10873 25684 10885 25687
rect 10275 25656 10885 25684
rect 10275 25653 10287 25656
rect 10229 25647 10287 25653
rect 10873 25653 10885 25656
rect 10919 25653 10931 25687
rect 10873 25647 10931 25653
rect 11238 25644 11244 25696
rect 11296 25684 11302 25696
rect 12986 25684 12992 25696
rect 11296 25656 12992 25684
rect 11296 25644 11302 25656
rect 12986 25644 12992 25656
rect 13044 25644 13050 25696
rect 1104 25594 14812 25616
rect 1104 25542 6315 25594
rect 6367 25542 6379 25594
rect 6431 25542 6443 25594
rect 6495 25542 6507 25594
rect 6559 25542 11648 25594
rect 11700 25542 11712 25594
rect 11764 25542 11776 25594
rect 11828 25542 11840 25594
rect 11892 25542 14812 25594
rect 1104 25520 14812 25542
rect 7282 25440 7288 25492
rect 7340 25480 7346 25492
rect 7837 25483 7895 25489
rect 7837 25480 7849 25483
rect 7340 25452 7849 25480
rect 7340 25440 7346 25452
rect 7837 25449 7849 25452
rect 7883 25449 7895 25483
rect 7837 25443 7895 25449
rect 8297 25483 8355 25489
rect 8297 25449 8309 25483
rect 8343 25480 8355 25483
rect 8846 25480 8852 25492
rect 8343 25452 8852 25480
rect 8343 25449 8355 25452
rect 8297 25443 8355 25449
rect 8846 25440 8852 25452
rect 8904 25440 8910 25492
rect 9306 25440 9312 25492
rect 9364 25480 9370 25492
rect 9677 25483 9735 25489
rect 9677 25480 9689 25483
rect 9364 25452 9689 25480
rect 9364 25440 9370 25452
rect 9677 25449 9689 25452
rect 9723 25449 9735 25483
rect 9677 25443 9735 25449
rect 10045 25483 10103 25489
rect 10045 25449 10057 25483
rect 10091 25480 10103 25483
rect 10502 25480 10508 25492
rect 10091 25452 10508 25480
rect 10091 25449 10103 25452
rect 10045 25443 10103 25449
rect 10502 25440 10508 25452
rect 10560 25480 10566 25492
rect 10689 25483 10747 25489
rect 10689 25480 10701 25483
rect 10560 25452 10701 25480
rect 10560 25440 10566 25452
rect 10689 25449 10701 25452
rect 10735 25449 10747 25483
rect 11054 25480 11060 25492
rect 11015 25452 11060 25480
rect 10689 25443 10747 25449
rect 11054 25440 11060 25452
rect 11112 25440 11118 25492
rect 12434 25440 12440 25492
rect 12492 25480 12498 25492
rect 12621 25483 12679 25489
rect 12621 25480 12633 25483
rect 12492 25452 12633 25480
rect 12492 25440 12498 25452
rect 12621 25449 12633 25452
rect 12667 25449 12679 25483
rect 12621 25443 12679 25449
rect 4338 25412 4344 25424
rect 4299 25384 4344 25412
rect 4338 25372 4344 25384
rect 4396 25372 4402 25424
rect 6178 25412 6184 25424
rect 6139 25384 6184 25412
rect 6178 25372 6184 25384
rect 6236 25372 6242 25424
rect 9950 25372 9956 25424
rect 10008 25412 10014 25424
rect 10137 25415 10195 25421
rect 10137 25412 10149 25415
rect 10008 25384 10149 25412
rect 10008 25372 10014 25384
rect 10137 25381 10149 25384
rect 10183 25381 10195 25415
rect 11072 25412 11100 25440
rect 11422 25412 11428 25424
rect 11072 25384 11428 25412
rect 10137 25375 10195 25381
rect 11422 25372 11428 25384
rect 11480 25421 11486 25424
rect 11480 25415 11544 25421
rect 11480 25381 11498 25415
rect 11532 25381 11544 25415
rect 11480 25375 11544 25381
rect 11480 25372 11486 25375
rect 4062 25344 4068 25356
rect 4023 25316 4068 25344
rect 4062 25304 4068 25316
rect 4120 25304 4126 25356
rect 6089 25347 6147 25353
rect 6089 25313 6101 25347
rect 6135 25344 6147 25347
rect 6822 25344 6828 25356
rect 6135 25316 6828 25344
rect 6135 25313 6147 25316
rect 6089 25307 6147 25313
rect 6822 25304 6828 25316
rect 6880 25304 6886 25356
rect 7558 25304 7564 25356
rect 7616 25344 7622 25356
rect 8205 25347 8263 25353
rect 8205 25344 8217 25347
rect 7616 25316 8217 25344
rect 7616 25304 7622 25316
rect 8205 25313 8217 25316
rect 8251 25313 8263 25347
rect 8205 25307 8263 25313
rect 10226 25304 10232 25356
rect 10284 25344 10290 25356
rect 11241 25347 11299 25353
rect 11241 25344 11253 25347
rect 10284 25316 11253 25344
rect 10284 25304 10290 25316
rect 11241 25313 11253 25316
rect 11287 25344 11299 25347
rect 11882 25344 11888 25356
rect 11287 25316 11888 25344
rect 11287 25313 11299 25316
rect 11241 25307 11299 25313
rect 11882 25304 11888 25316
rect 11940 25304 11946 25356
rect 6270 25276 6276 25288
rect 6231 25248 6276 25276
rect 6270 25236 6276 25248
rect 6328 25236 6334 25288
rect 8294 25236 8300 25288
rect 8352 25276 8358 25288
rect 8389 25279 8447 25285
rect 8389 25276 8401 25279
rect 8352 25248 8401 25276
rect 8352 25236 8358 25248
rect 8389 25245 8401 25248
rect 8435 25245 8447 25279
rect 10318 25276 10324 25288
rect 10279 25248 10324 25276
rect 8389 25239 8447 25245
rect 10318 25236 10324 25248
rect 10376 25236 10382 25288
rect 9217 25211 9275 25217
rect 9217 25177 9229 25211
rect 9263 25208 9275 25211
rect 10336 25208 10364 25236
rect 9263 25180 10364 25208
rect 9263 25177 9275 25180
rect 9217 25171 9275 25177
rect 4893 25143 4951 25149
rect 4893 25109 4905 25143
rect 4939 25140 4951 25143
rect 5258 25140 5264 25152
rect 4939 25112 5264 25140
rect 4939 25109 4951 25112
rect 4893 25103 4951 25109
rect 5258 25100 5264 25112
rect 5316 25100 5322 25152
rect 5534 25100 5540 25152
rect 5592 25140 5598 25152
rect 5721 25143 5779 25149
rect 5721 25140 5733 25143
rect 5592 25112 5733 25140
rect 5592 25100 5598 25112
rect 5721 25109 5733 25112
rect 5767 25109 5779 25143
rect 7650 25140 7656 25152
rect 7611 25112 7656 25140
rect 5721 25103 5779 25109
rect 7650 25100 7656 25112
rect 7708 25100 7714 25152
rect 1104 25050 14812 25072
rect 1104 24998 3648 25050
rect 3700 24998 3712 25050
rect 3764 24998 3776 25050
rect 3828 24998 3840 25050
rect 3892 24998 8982 25050
rect 9034 24998 9046 25050
rect 9098 24998 9110 25050
rect 9162 24998 9174 25050
rect 9226 24998 14315 25050
rect 14367 24998 14379 25050
rect 14431 24998 14443 25050
rect 14495 24998 14507 25050
rect 14559 24998 14812 25050
rect 1104 24976 14812 24998
rect 6178 24936 6184 24948
rect 6139 24908 6184 24936
rect 6178 24896 6184 24908
rect 6236 24896 6242 24948
rect 7558 24936 7564 24948
rect 7519 24908 7564 24936
rect 7558 24896 7564 24908
rect 7616 24896 7622 24948
rect 9766 24936 9772 24948
rect 8312 24908 9772 24936
rect 5905 24871 5963 24877
rect 5905 24837 5917 24871
rect 5951 24868 5963 24871
rect 6270 24868 6276 24880
rect 5951 24840 6276 24868
rect 5951 24837 5963 24840
rect 5905 24831 5963 24837
rect 6270 24828 6276 24840
rect 6328 24868 6334 24880
rect 6730 24868 6736 24880
rect 6328 24840 6736 24868
rect 6328 24828 6334 24840
rect 6730 24828 6736 24840
rect 6788 24828 6794 24880
rect 7650 24828 7656 24880
rect 7708 24868 7714 24880
rect 8312 24868 8340 24908
rect 9766 24896 9772 24908
rect 9824 24896 9830 24948
rect 10502 24896 10508 24948
rect 10560 24936 10566 24948
rect 10686 24936 10692 24948
rect 10560 24908 10692 24936
rect 10560 24896 10566 24908
rect 10686 24896 10692 24908
rect 10744 24936 10750 24948
rect 10781 24939 10839 24945
rect 10781 24936 10793 24939
rect 10744 24908 10793 24936
rect 10744 24896 10750 24908
rect 10781 24905 10793 24908
rect 10827 24905 10839 24939
rect 10781 24899 10839 24905
rect 11422 24896 11428 24948
rect 11480 24936 11486 24948
rect 11517 24939 11575 24945
rect 11517 24936 11529 24939
rect 11480 24908 11529 24936
rect 11480 24896 11486 24908
rect 11517 24905 11529 24908
rect 11563 24905 11575 24939
rect 11882 24936 11888 24948
rect 11843 24908 11888 24936
rect 11517 24899 11575 24905
rect 11882 24896 11888 24908
rect 11940 24896 11946 24948
rect 7708 24840 8340 24868
rect 7708 24828 7714 24840
rect 4709 24803 4767 24809
rect 4709 24769 4721 24803
rect 4755 24800 4767 24803
rect 5350 24800 5356 24812
rect 4755 24772 5356 24800
rect 4755 24769 4767 24772
rect 4709 24763 4767 24769
rect 5350 24760 5356 24772
rect 5408 24760 5414 24812
rect 8220 24809 8248 24840
rect 8205 24803 8263 24809
rect 8205 24769 8217 24803
rect 8251 24769 8263 24803
rect 8205 24763 8263 24769
rect 8294 24760 8300 24812
rect 8352 24800 8358 24812
rect 8573 24803 8631 24809
rect 8573 24800 8585 24803
rect 8352 24772 8585 24800
rect 8352 24760 8358 24772
rect 8573 24769 8585 24772
rect 8619 24769 8631 24803
rect 8573 24763 8631 24769
rect 8754 24760 8760 24812
rect 8812 24800 8818 24812
rect 8941 24803 8999 24809
rect 8941 24800 8953 24803
rect 8812 24772 8953 24800
rect 8812 24760 8818 24772
rect 8941 24769 8953 24772
rect 8987 24769 8999 24803
rect 8941 24763 8999 24769
rect 4341 24735 4399 24741
rect 4341 24701 4353 24735
rect 4387 24732 4399 24735
rect 5169 24735 5227 24741
rect 5169 24732 5181 24735
rect 4387 24704 5181 24732
rect 4387 24701 4399 24704
rect 4341 24695 4399 24701
rect 5169 24701 5181 24704
rect 5215 24732 5227 24735
rect 5442 24732 5448 24744
rect 5215 24704 5448 24732
rect 5215 24701 5227 24704
rect 5169 24695 5227 24701
rect 5442 24692 5448 24704
rect 5500 24692 5506 24744
rect 7469 24735 7527 24741
rect 7469 24701 7481 24735
rect 7515 24732 7527 24735
rect 7926 24732 7932 24744
rect 7515 24704 7932 24732
rect 7515 24701 7527 24704
rect 7469 24695 7527 24701
rect 7926 24692 7932 24704
rect 7984 24692 7990 24744
rect 3973 24667 4031 24673
rect 3973 24633 3985 24667
rect 4019 24664 4031 24667
rect 4062 24664 4068 24676
rect 4019 24636 4068 24664
rect 4019 24633 4031 24636
rect 3973 24627 4031 24633
rect 4062 24624 4068 24636
rect 4120 24664 4126 24676
rect 7101 24667 7159 24673
rect 4120 24636 4844 24664
rect 4120 24624 4126 24636
rect 4816 24605 4844 24636
rect 7101 24633 7113 24667
rect 7147 24664 7159 24667
rect 8956 24664 8984 24763
rect 10318 24760 10324 24812
rect 10376 24800 10382 24812
rect 11149 24803 11207 24809
rect 11149 24800 11161 24803
rect 10376 24772 11161 24800
rect 10376 24760 10382 24772
rect 11149 24769 11161 24772
rect 11195 24769 11207 24803
rect 11149 24763 11207 24769
rect 9122 24732 9128 24744
rect 9083 24704 9128 24732
rect 9122 24692 9128 24704
rect 9180 24692 9186 24744
rect 9214 24692 9220 24744
rect 9272 24732 9278 24744
rect 9392 24735 9450 24741
rect 9392 24732 9404 24735
rect 9272 24704 9404 24732
rect 9272 24692 9278 24704
rect 9392 24701 9404 24704
rect 9438 24732 9450 24735
rect 10336 24732 10364 24760
rect 9438 24704 10364 24732
rect 9438 24701 9450 24704
rect 9392 24695 9450 24701
rect 9306 24664 9312 24676
rect 7147 24636 8064 24664
rect 8956 24636 9312 24664
rect 7147 24633 7159 24636
rect 7101 24627 7159 24633
rect 8036 24608 8064 24636
rect 9306 24624 9312 24636
rect 9364 24624 9370 24676
rect 4801 24599 4859 24605
rect 4801 24565 4813 24599
rect 4847 24565 4859 24599
rect 5258 24596 5264 24608
rect 5219 24568 5264 24596
rect 4801 24559 4859 24565
rect 5258 24556 5264 24568
rect 5316 24556 5322 24608
rect 6641 24599 6699 24605
rect 6641 24565 6653 24599
rect 6687 24596 6699 24599
rect 6822 24596 6828 24608
rect 6687 24568 6828 24596
rect 6687 24565 6699 24568
rect 6641 24559 6699 24565
rect 6822 24556 6828 24568
rect 6880 24556 6886 24608
rect 8018 24556 8024 24608
rect 8076 24596 8082 24608
rect 8076 24568 8121 24596
rect 8076 24556 8082 24568
rect 9766 24556 9772 24608
rect 9824 24596 9830 24608
rect 10505 24599 10563 24605
rect 10505 24596 10517 24599
rect 9824 24568 10517 24596
rect 9824 24556 9830 24568
rect 10505 24565 10517 24568
rect 10551 24565 10563 24599
rect 10505 24559 10563 24565
rect 1104 24506 14812 24528
rect 1104 24454 6315 24506
rect 6367 24454 6379 24506
rect 6431 24454 6443 24506
rect 6495 24454 6507 24506
rect 6559 24454 11648 24506
rect 11700 24454 11712 24506
rect 11764 24454 11776 24506
rect 11828 24454 11840 24506
rect 11892 24454 14812 24506
rect 1104 24432 14812 24454
rect 5813 24395 5871 24401
rect 5813 24361 5825 24395
rect 5859 24392 5871 24395
rect 6178 24392 6184 24404
rect 5859 24364 6184 24392
rect 5859 24361 5871 24364
rect 5813 24355 5871 24361
rect 6178 24352 6184 24364
rect 6236 24352 6242 24404
rect 6730 24352 6736 24404
rect 6788 24392 6794 24404
rect 6825 24395 6883 24401
rect 6825 24392 6837 24395
rect 6788 24364 6837 24392
rect 6788 24352 6794 24364
rect 6825 24361 6837 24364
rect 6871 24361 6883 24395
rect 6825 24355 6883 24361
rect 7285 24395 7343 24401
rect 7285 24361 7297 24395
rect 7331 24392 7343 24395
rect 7558 24392 7564 24404
rect 7331 24364 7564 24392
rect 7331 24361 7343 24364
rect 7285 24355 7343 24361
rect 7558 24352 7564 24364
rect 7616 24352 7622 24404
rect 8757 24395 8815 24401
rect 8757 24361 8769 24395
rect 8803 24392 8815 24395
rect 9125 24395 9183 24401
rect 9125 24392 9137 24395
rect 8803 24364 9137 24392
rect 8803 24361 8815 24364
rect 8757 24355 8815 24361
rect 9125 24361 9137 24364
rect 9171 24392 9183 24395
rect 9214 24392 9220 24404
rect 9171 24364 9220 24392
rect 9171 24361 9183 24364
rect 9125 24355 9183 24361
rect 9214 24352 9220 24364
rect 9272 24352 9278 24404
rect 9674 24392 9680 24404
rect 9635 24364 9680 24392
rect 9674 24352 9680 24364
rect 9732 24352 9738 24404
rect 11238 24392 11244 24404
rect 11199 24364 11244 24392
rect 11238 24352 11244 24364
rect 11296 24352 11302 24404
rect 11609 24395 11667 24401
rect 11609 24361 11621 24395
rect 11655 24392 11667 24395
rect 12250 24392 12256 24404
rect 11655 24364 12256 24392
rect 11655 24361 11667 24364
rect 11609 24355 11667 24361
rect 12250 24352 12256 24364
rect 12308 24352 12314 24404
rect 6270 24324 6276 24336
rect 6183 24296 6276 24324
rect 6270 24284 6276 24296
rect 6328 24324 6334 24336
rect 6914 24324 6920 24336
rect 6328 24296 6920 24324
rect 6328 24284 6334 24296
rect 6914 24284 6920 24296
rect 6972 24284 6978 24336
rect 7466 24284 7472 24336
rect 7524 24324 7530 24336
rect 7644 24327 7702 24333
rect 7644 24324 7656 24327
rect 7524 24296 7656 24324
rect 7524 24284 7530 24296
rect 7644 24293 7656 24296
rect 7690 24293 7702 24327
rect 7644 24287 7702 24293
rect 10045 24327 10103 24333
rect 10045 24293 10057 24327
rect 10091 24324 10103 24327
rect 10778 24324 10784 24336
rect 10091 24296 10784 24324
rect 10091 24293 10103 24296
rect 10045 24287 10103 24293
rect 10778 24284 10784 24296
rect 10836 24284 10842 24336
rect 11422 24284 11428 24336
rect 11480 24324 11486 24336
rect 11701 24327 11759 24333
rect 11701 24324 11713 24327
rect 11480 24296 11713 24324
rect 11480 24284 11486 24296
rect 11701 24293 11713 24296
rect 11747 24293 11759 24327
rect 11701 24287 11759 24293
rect 6086 24216 6092 24268
rect 6144 24256 6150 24268
rect 6181 24259 6239 24265
rect 6181 24256 6193 24259
rect 6144 24228 6193 24256
rect 6144 24216 6150 24228
rect 6181 24225 6193 24228
rect 6227 24225 6239 24259
rect 10410 24256 10416 24268
rect 6181 24219 6239 24225
rect 10152 24228 10416 24256
rect 4798 24188 4804 24200
rect 4759 24160 4804 24188
rect 4798 24148 4804 24160
rect 4856 24148 4862 24200
rect 5534 24148 5540 24200
rect 5592 24188 5598 24200
rect 6365 24191 6423 24197
rect 6365 24188 6377 24191
rect 5592 24160 6377 24188
rect 5592 24148 5598 24160
rect 6365 24157 6377 24160
rect 6411 24157 6423 24191
rect 6365 24151 6423 24157
rect 7377 24191 7435 24197
rect 7377 24157 7389 24191
rect 7423 24157 7435 24191
rect 7377 24151 7435 24157
rect 4430 24052 4436 24064
rect 4391 24024 4436 24052
rect 4430 24012 4436 24024
rect 4488 24012 4494 24064
rect 7190 24012 7196 24064
rect 7248 24052 7254 24064
rect 7392 24052 7420 24151
rect 9950 24148 9956 24200
rect 10008 24188 10014 24200
rect 10152 24197 10180 24228
rect 10410 24216 10416 24228
rect 10468 24216 10474 24268
rect 10137 24191 10195 24197
rect 10137 24188 10149 24191
rect 10008 24160 10149 24188
rect 10008 24148 10014 24160
rect 10137 24157 10149 24160
rect 10183 24157 10195 24191
rect 10318 24188 10324 24200
rect 10279 24160 10324 24188
rect 10137 24151 10195 24157
rect 10318 24148 10324 24160
rect 10376 24148 10382 24200
rect 11514 24148 11520 24200
rect 11572 24188 11578 24200
rect 11793 24191 11851 24197
rect 11793 24188 11805 24191
rect 11572 24160 11805 24188
rect 11572 24148 11578 24160
rect 11793 24157 11805 24160
rect 11839 24157 11851 24191
rect 11793 24151 11851 24157
rect 9122 24080 9128 24132
rect 9180 24080 9186 24132
rect 8386 24052 8392 24064
rect 7248 24024 8392 24052
rect 7248 24012 7254 24024
rect 8386 24012 8392 24024
rect 8444 24052 8450 24064
rect 9140 24052 9168 24080
rect 9401 24055 9459 24061
rect 9401 24052 9413 24055
rect 8444 24024 9413 24052
rect 8444 24012 8450 24024
rect 9401 24021 9413 24024
rect 9447 24021 9459 24055
rect 9401 24015 9459 24021
rect 1104 23962 14812 23984
rect 1104 23910 3648 23962
rect 3700 23910 3712 23962
rect 3764 23910 3776 23962
rect 3828 23910 3840 23962
rect 3892 23910 8982 23962
rect 9034 23910 9046 23962
rect 9098 23910 9110 23962
rect 9162 23910 9174 23962
rect 9226 23910 14315 23962
rect 14367 23910 14379 23962
rect 14431 23910 14443 23962
rect 14495 23910 14507 23962
rect 14559 23910 14812 23962
rect 1104 23888 14812 23910
rect 5810 23808 5816 23860
rect 5868 23848 5874 23860
rect 5905 23851 5963 23857
rect 5905 23848 5917 23851
rect 5868 23820 5917 23848
rect 5868 23808 5874 23820
rect 5905 23817 5917 23820
rect 5951 23848 5963 23851
rect 6086 23848 6092 23860
rect 5951 23820 6092 23848
rect 5951 23817 5963 23820
rect 5905 23811 5963 23817
rect 6086 23808 6092 23820
rect 6144 23808 6150 23860
rect 6270 23848 6276 23860
rect 6231 23820 6276 23848
rect 6270 23808 6276 23820
rect 6328 23808 6334 23860
rect 7466 23808 7472 23860
rect 7524 23848 7530 23860
rect 7524 23820 7788 23848
rect 7524 23808 7530 23820
rect 5626 23740 5632 23792
rect 5684 23780 5690 23792
rect 6457 23783 6515 23789
rect 6457 23780 6469 23783
rect 5684 23752 6469 23780
rect 5684 23740 5690 23752
rect 6457 23749 6469 23752
rect 6503 23749 6515 23783
rect 6457 23743 6515 23749
rect 6730 23740 6736 23792
rect 6788 23740 6794 23792
rect 7760 23780 7788 23820
rect 8018 23808 8024 23860
rect 8076 23848 8082 23860
rect 9033 23851 9091 23857
rect 9033 23848 9045 23851
rect 8076 23820 9045 23848
rect 8076 23808 8082 23820
rect 9033 23817 9045 23820
rect 9079 23817 9091 23851
rect 9033 23811 9091 23817
rect 10502 23808 10508 23860
rect 10560 23848 10566 23860
rect 10778 23848 10784 23860
rect 10560 23820 10784 23848
rect 10560 23808 10566 23820
rect 10778 23808 10784 23820
rect 10836 23808 10842 23860
rect 11146 23808 11152 23860
rect 11204 23848 11210 23860
rect 11333 23851 11391 23857
rect 11333 23848 11345 23851
rect 11204 23820 11345 23848
rect 11204 23808 11210 23820
rect 11333 23817 11345 23820
rect 11379 23848 11391 23851
rect 11422 23848 11428 23860
rect 11379 23820 11428 23848
rect 11379 23817 11391 23820
rect 11333 23811 11391 23817
rect 11422 23808 11428 23820
rect 11480 23808 11486 23860
rect 11514 23808 11520 23860
rect 11572 23848 11578 23860
rect 11977 23851 12035 23857
rect 11977 23848 11989 23851
rect 11572 23820 11989 23848
rect 11572 23808 11578 23820
rect 11977 23817 11989 23820
rect 12023 23817 12035 23851
rect 11977 23811 12035 23817
rect 8205 23783 8263 23789
rect 8205 23780 8217 23783
rect 7760 23752 8217 23780
rect 8205 23749 8217 23752
rect 8251 23780 8263 23783
rect 8481 23783 8539 23789
rect 8481 23780 8493 23783
rect 8251 23752 8493 23780
rect 8251 23749 8263 23752
rect 8205 23743 8263 23749
rect 8481 23749 8493 23752
rect 8527 23749 8539 23783
rect 8846 23780 8852 23792
rect 8807 23752 8852 23780
rect 8481 23743 8539 23749
rect 8846 23740 8852 23752
rect 8904 23780 8910 23792
rect 11701 23783 11759 23789
rect 11701 23780 11713 23783
rect 8904 23752 9536 23780
rect 8904 23740 8910 23752
rect 4430 23672 4436 23724
rect 4488 23712 4494 23724
rect 4893 23715 4951 23721
rect 4893 23712 4905 23715
rect 4488 23684 4905 23712
rect 4488 23672 4494 23684
rect 4893 23681 4905 23684
rect 4939 23681 4951 23715
rect 4893 23675 4951 23681
rect 5718 23672 5724 23724
rect 5776 23712 5782 23724
rect 6086 23712 6092 23724
rect 5776 23684 6092 23712
rect 5776 23672 5782 23684
rect 6086 23672 6092 23684
rect 6144 23672 6150 23724
rect 6748 23712 6776 23740
rect 9508 23721 9536 23752
rect 11440 23752 11713 23780
rect 11440 23724 11468 23752
rect 11701 23749 11713 23752
rect 11747 23780 11759 23783
rect 12250 23780 12256 23792
rect 11747 23752 12256 23780
rect 11747 23749 11759 23752
rect 11701 23743 11759 23749
rect 12250 23740 12256 23752
rect 12308 23740 12314 23792
rect 9493 23715 9551 23721
rect 6748 23684 6960 23712
rect 4249 23647 4307 23653
rect 4249 23613 4261 23647
rect 4295 23644 4307 23647
rect 6641 23647 6699 23653
rect 4295 23616 4844 23644
rect 4295 23613 4307 23616
rect 4249 23607 4307 23613
rect 4706 23576 4712 23588
rect 4667 23548 4712 23576
rect 4706 23536 4712 23548
rect 4764 23536 4770 23588
rect 4816 23585 4844 23616
rect 6641 23613 6653 23647
rect 6687 23613 6699 23647
rect 6641 23607 6699 23613
rect 6825 23647 6883 23653
rect 6825 23613 6837 23647
rect 6871 23613 6883 23647
rect 6932 23644 6960 23684
rect 9493 23681 9505 23715
rect 9539 23681 9551 23715
rect 9493 23675 9551 23681
rect 9677 23715 9735 23721
rect 9677 23681 9689 23715
rect 9723 23712 9735 23715
rect 9858 23712 9864 23724
rect 9723 23684 9864 23712
rect 9723 23681 9735 23684
rect 9677 23675 9735 23681
rect 9858 23672 9864 23684
rect 9916 23712 9922 23724
rect 10318 23712 10324 23724
rect 9916 23684 10324 23712
rect 9916 23672 9922 23684
rect 10318 23672 10324 23684
rect 10376 23672 10382 23724
rect 10778 23672 10784 23724
rect 10836 23712 10842 23724
rect 11054 23712 11060 23724
rect 10836 23684 11060 23712
rect 10836 23672 10842 23684
rect 11054 23672 11060 23684
rect 11112 23672 11118 23724
rect 11422 23672 11428 23724
rect 11480 23672 11486 23724
rect 7081 23647 7139 23653
rect 7081 23644 7093 23647
rect 6932 23616 7093 23644
rect 6825 23607 6883 23613
rect 7081 23613 7093 23616
rect 7127 23613 7139 23647
rect 9398 23644 9404 23656
rect 9359 23616 9404 23644
rect 7081 23607 7139 23613
rect 4801 23579 4859 23585
rect 4801 23545 4813 23579
rect 4847 23576 4859 23579
rect 5074 23576 5080 23588
rect 4847 23548 5080 23576
rect 4847 23545 4859 23548
rect 4801 23539 4859 23545
rect 5074 23536 5080 23548
rect 5132 23576 5138 23588
rect 5442 23576 5448 23588
rect 5132 23548 5448 23576
rect 5132 23536 5138 23548
rect 5442 23536 5448 23548
rect 5500 23536 5506 23588
rect 5718 23536 5724 23588
rect 5776 23576 5782 23588
rect 6546 23576 6552 23588
rect 5776 23548 6552 23576
rect 5776 23536 5782 23548
rect 6546 23536 6552 23548
rect 6604 23536 6610 23588
rect 4338 23508 4344 23520
rect 4299 23480 4344 23508
rect 4338 23468 4344 23480
rect 4396 23468 4402 23520
rect 5534 23508 5540 23520
rect 5495 23480 5540 23508
rect 5534 23468 5540 23480
rect 5592 23468 5598 23520
rect 6656 23508 6684 23607
rect 6840 23576 6868 23607
rect 9398 23604 9404 23616
rect 9456 23604 9462 23656
rect 7190 23576 7196 23588
rect 6840 23548 7196 23576
rect 7190 23536 7196 23548
rect 7248 23536 7254 23588
rect 7558 23508 7564 23520
rect 6656 23480 7564 23508
rect 7558 23468 7564 23480
rect 7616 23468 7622 23520
rect 9950 23468 9956 23520
rect 10008 23508 10014 23520
rect 10045 23511 10103 23517
rect 10045 23508 10057 23511
rect 10008 23480 10057 23508
rect 10008 23468 10014 23480
rect 10045 23477 10057 23480
rect 10091 23477 10103 23511
rect 10045 23471 10103 23477
rect 1104 23418 14812 23440
rect 1104 23366 6315 23418
rect 6367 23366 6379 23418
rect 6431 23366 6443 23418
rect 6495 23366 6507 23418
rect 6559 23366 11648 23418
rect 11700 23366 11712 23418
rect 11764 23366 11776 23418
rect 11828 23366 11840 23418
rect 11892 23366 14812 23418
rect 1104 23344 14812 23366
rect 4433 23307 4491 23313
rect 4433 23273 4445 23307
rect 4479 23304 4491 23307
rect 4706 23304 4712 23316
rect 4479 23276 4712 23304
rect 4479 23273 4491 23276
rect 4433 23267 4491 23273
rect 4706 23264 4712 23276
rect 4764 23264 4770 23316
rect 6638 23304 6644 23316
rect 6599 23276 6644 23304
rect 6638 23264 6644 23276
rect 6696 23264 6702 23316
rect 6914 23304 6920 23316
rect 6875 23276 6920 23304
rect 6914 23264 6920 23276
rect 6972 23264 6978 23316
rect 7466 23304 7472 23316
rect 7427 23276 7472 23304
rect 7466 23264 7472 23276
rect 7524 23264 7530 23316
rect 9125 23307 9183 23313
rect 9125 23273 9137 23307
rect 9171 23304 9183 23307
rect 9398 23304 9404 23316
rect 9171 23276 9404 23304
rect 9171 23273 9183 23276
rect 9125 23267 9183 23273
rect 9398 23264 9404 23276
rect 9456 23264 9462 23316
rect 9858 23304 9864 23316
rect 9819 23276 9864 23304
rect 9858 23264 9864 23276
rect 9916 23264 9922 23316
rect 5534 23245 5540 23248
rect 5528 23236 5540 23245
rect 5495 23208 5540 23236
rect 5528 23199 5540 23208
rect 5534 23196 5540 23199
rect 5592 23196 5598 23248
rect 5626 23196 5632 23248
rect 5684 23196 5690 23248
rect 4062 23128 4068 23180
rect 4120 23168 4126 23180
rect 4985 23171 5043 23177
rect 4985 23168 4997 23171
rect 4120 23140 4997 23168
rect 4120 23128 4126 23140
rect 4985 23137 4997 23140
rect 5031 23168 5043 23171
rect 5644 23168 5672 23196
rect 7834 23168 7840 23180
rect 5031 23140 5672 23168
rect 7795 23140 7840 23168
rect 5031 23137 5043 23140
rect 4985 23131 5043 23137
rect 7834 23128 7840 23140
rect 7892 23128 7898 23180
rect 7929 23171 7987 23177
rect 7929 23137 7941 23171
rect 7975 23168 7987 23171
rect 8202 23168 8208 23180
rect 7975 23140 8208 23168
rect 7975 23137 7987 23140
rect 7929 23131 7987 23137
rect 8202 23128 8208 23140
rect 8260 23128 8266 23180
rect 5261 23103 5319 23109
rect 5261 23100 5273 23103
rect 4816 23072 5273 23100
rect 4246 22924 4252 22976
rect 4304 22964 4310 22976
rect 4816 22973 4844 23072
rect 5261 23069 5273 23072
rect 5307 23069 5319 23103
rect 5261 23063 5319 23069
rect 6638 23060 6644 23112
rect 6696 23100 6702 23112
rect 8018 23100 8024 23112
rect 6696 23072 8024 23100
rect 6696 23060 6702 23072
rect 8018 23060 8024 23072
rect 8076 23060 8082 23112
rect 4801 22967 4859 22973
rect 4801 22964 4813 22967
rect 4304 22936 4813 22964
rect 4304 22924 4310 22936
rect 4801 22933 4813 22936
rect 4847 22933 4859 22967
rect 4801 22927 4859 22933
rect 7377 22967 7435 22973
rect 7377 22933 7389 22967
rect 7423 22964 7435 22967
rect 7466 22964 7472 22976
rect 7423 22936 7472 22964
rect 7423 22933 7435 22936
rect 7377 22927 7435 22933
rect 7466 22924 7472 22936
rect 7524 22924 7530 22976
rect 8386 22924 8392 22976
rect 8444 22964 8450 22976
rect 8481 22967 8539 22973
rect 8481 22964 8493 22967
rect 8444 22936 8493 22964
rect 8444 22924 8450 22936
rect 8481 22933 8493 22936
rect 8527 22933 8539 22967
rect 8481 22927 8539 22933
rect 1104 22874 14812 22896
rect 1104 22822 3648 22874
rect 3700 22822 3712 22874
rect 3764 22822 3776 22874
rect 3828 22822 3840 22874
rect 3892 22822 8982 22874
rect 9034 22822 9046 22874
rect 9098 22822 9110 22874
rect 9162 22822 9174 22874
rect 9226 22822 14315 22874
rect 14367 22822 14379 22874
rect 14431 22822 14443 22874
rect 14495 22822 14507 22874
rect 14559 22822 14812 22874
rect 1104 22800 14812 22822
rect 3418 22760 3424 22772
rect 3379 22732 3424 22760
rect 3418 22720 3424 22732
rect 3476 22720 3482 22772
rect 3789 22763 3847 22769
rect 3789 22729 3801 22763
rect 3835 22760 3847 22763
rect 4062 22760 4068 22772
rect 3835 22732 4068 22760
rect 3835 22729 3847 22732
rect 3789 22723 3847 22729
rect 4062 22720 4068 22732
rect 4120 22720 4126 22772
rect 4157 22763 4215 22769
rect 4157 22729 4169 22763
rect 4203 22760 4215 22763
rect 4430 22760 4436 22772
rect 4203 22732 4436 22760
rect 4203 22729 4215 22732
rect 4157 22723 4215 22729
rect 4430 22720 4436 22732
rect 4488 22720 4494 22772
rect 6822 22760 6828 22772
rect 6783 22732 6828 22760
rect 6822 22720 6828 22732
rect 6880 22720 6886 22772
rect 7929 22763 7987 22769
rect 7929 22729 7941 22763
rect 7975 22760 7987 22763
rect 8018 22760 8024 22772
rect 7975 22732 8024 22760
rect 7975 22729 7987 22732
rect 7929 22723 7987 22729
rect 8018 22720 8024 22732
rect 8076 22720 8082 22772
rect 8389 22763 8447 22769
rect 8389 22729 8401 22763
rect 8435 22760 8447 22763
rect 8478 22760 8484 22772
rect 8435 22732 8484 22760
rect 8435 22729 8447 22732
rect 8389 22723 8447 22729
rect 8478 22720 8484 22732
rect 8536 22720 8542 22772
rect 3436 22624 3464 22720
rect 4062 22624 4068 22636
rect 3436 22596 4068 22624
rect 4062 22584 4068 22596
rect 4120 22624 4126 22636
rect 4246 22624 4252 22636
rect 4120 22596 4252 22624
rect 4120 22584 4126 22596
rect 4246 22584 4252 22596
rect 4304 22584 4310 22636
rect 7469 22627 7527 22633
rect 7469 22593 7481 22627
rect 7515 22593 7527 22627
rect 8496 22624 8524 22720
rect 10229 22627 10287 22633
rect 10229 22624 10241 22627
rect 8496 22596 10241 22624
rect 7469 22587 7527 22593
rect 6914 22516 6920 22568
rect 6972 22556 6978 22568
rect 7193 22559 7251 22565
rect 7193 22556 7205 22559
rect 6972 22528 7205 22556
rect 6972 22516 6978 22528
rect 7193 22525 7205 22528
rect 7239 22525 7251 22559
rect 7193 22519 7251 22525
rect 7282 22516 7288 22568
rect 7340 22556 7346 22568
rect 7340 22528 7385 22556
rect 7340 22516 7346 22528
rect 4430 22448 4436 22500
rect 4488 22497 4494 22500
rect 4488 22491 4552 22497
rect 4488 22457 4506 22491
rect 4540 22457 4552 22491
rect 6638 22488 6644 22500
rect 6551 22460 6644 22488
rect 4488 22451 4552 22457
rect 4488 22448 4494 22451
rect 6638 22448 6644 22460
rect 6696 22488 6702 22500
rect 7300 22488 7328 22516
rect 6696 22460 7328 22488
rect 6696 22448 6702 22460
rect 5534 22380 5540 22432
rect 5592 22420 5598 22432
rect 5629 22423 5687 22429
rect 5629 22420 5641 22423
rect 5592 22392 5641 22420
rect 5592 22380 5598 22392
rect 5629 22389 5641 22392
rect 5675 22420 5687 22423
rect 5718 22420 5724 22432
rect 5675 22392 5724 22420
rect 5675 22389 5687 22392
rect 5629 22383 5687 22389
rect 5718 22380 5724 22392
rect 5776 22420 5782 22432
rect 6181 22423 6239 22429
rect 6181 22420 6193 22423
rect 5776 22392 6193 22420
rect 5776 22380 5782 22392
rect 6181 22389 6193 22392
rect 6227 22420 6239 22423
rect 6914 22420 6920 22432
rect 6227 22392 6920 22420
rect 6227 22389 6239 22392
rect 6181 22383 6239 22389
rect 6914 22380 6920 22392
rect 6972 22420 6978 22432
rect 7484 22420 7512 22587
rect 7558 22516 7564 22568
rect 7616 22556 7622 22568
rect 9968 22565 9996 22596
rect 10229 22593 10241 22596
rect 10275 22593 10287 22627
rect 10229 22587 10287 22593
rect 8573 22559 8631 22565
rect 8573 22556 8585 22559
rect 7616 22528 8585 22556
rect 7616 22516 7622 22528
rect 8573 22525 8585 22528
rect 8619 22556 8631 22559
rect 8849 22559 8907 22565
rect 8849 22556 8861 22559
rect 8619 22528 8861 22556
rect 8619 22525 8631 22528
rect 8573 22519 8631 22525
rect 8849 22525 8861 22528
rect 8895 22525 8907 22559
rect 8849 22519 8907 22525
rect 9953 22559 10011 22565
rect 9953 22525 9965 22559
rect 9999 22525 10011 22559
rect 9953 22519 10011 22525
rect 8202 22420 8208 22432
rect 6972 22392 7512 22420
rect 8163 22392 8208 22420
rect 6972 22380 6978 22392
rect 8202 22380 8208 22392
rect 8260 22380 8266 22432
rect 9769 22423 9827 22429
rect 9769 22389 9781 22423
rect 9815 22420 9827 22423
rect 10226 22420 10232 22432
rect 9815 22392 10232 22420
rect 9815 22389 9827 22392
rect 9769 22383 9827 22389
rect 10226 22380 10232 22392
rect 10284 22380 10290 22432
rect 1104 22330 14812 22352
rect 1104 22278 6315 22330
rect 6367 22278 6379 22330
rect 6431 22278 6443 22330
rect 6495 22278 6507 22330
rect 6559 22278 11648 22330
rect 11700 22278 11712 22330
rect 11764 22278 11776 22330
rect 11828 22278 11840 22330
rect 11892 22278 14812 22330
rect 1104 22256 14812 22278
rect 4430 22176 4436 22228
rect 4488 22216 4494 22228
rect 5445 22219 5503 22225
rect 5445 22216 5457 22219
rect 4488 22188 5457 22216
rect 4488 22176 4494 22188
rect 5445 22185 5457 22188
rect 5491 22185 5503 22219
rect 5445 22179 5503 22185
rect 5994 22176 6000 22228
rect 6052 22216 6058 22228
rect 6641 22219 6699 22225
rect 6641 22216 6653 22219
rect 6052 22188 6653 22216
rect 6052 22176 6058 22188
rect 6288 22160 6316 22188
rect 6641 22185 6653 22188
rect 6687 22185 6699 22219
rect 7558 22216 7564 22228
rect 7471 22188 7564 22216
rect 6641 22179 6699 22185
rect 7558 22176 7564 22188
rect 7616 22216 7622 22228
rect 7834 22216 7840 22228
rect 7616 22188 7840 22216
rect 7616 22176 7622 22188
rect 7834 22176 7840 22188
rect 7892 22176 7898 22228
rect 4062 22108 4068 22160
rect 4120 22148 4126 22160
rect 6089 22151 6147 22157
rect 6089 22148 6101 22151
rect 4120 22120 6101 22148
rect 4120 22108 4126 22120
rect 5920 22092 5948 22120
rect 6089 22117 6101 22120
rect 6135 22117 6147 22151
rect 6089 22111 6147 22117
rect 6270 22108 6276 22160
rect 6328 22108 6334 22160
rect 6733 22151 6791 22157
rect 6733 22117 6745 22151
rect 6779 22148 6791 22151
rect 7098 22148 7104 22160
rect 6779 22120 7104 22148
rect 6779 22117 6791 22120
rect 6733 22111 6791 22117
rect 7098 22108 7104 22120
rect 7156 22108 7162 22160
rect 4154 22040 4160 22092
rect 4212 22080 4218 22092
rect 4321 22083 4379 22089
rect 4321 22080 4333 22083
rect 4212 22052 4333 22080
rect 4212 22040 4218 22052
rect 4321 22049 4333 22052
rect 4367 22049 4379 22083
rect 4321 22043 4379 22049
rect 5902 22040 5908 22092
rect 5960 22040 5966 22092
rect 10318 22040 10324 22092
rect 10376 22080 10382 22092
rect 10485 22083 10543 22089
rect 10485 22080 10497 22083
rect 10376 22052 10497 22080
rect 10376 22040 10382 22052
rect 10485 22049 10497 22052
rect 10531 22049 10543 22083
rect 10485 22043 10543 22049
rect 4062 22012 4068 22024
rect 4023 21984 4068 22012
rect 4062 21972 4068 21984
rect 4120 21972 4126 22024
rect 6914 22012 6920 22024
rect 6875 21984 6920 22012
rect 6914 21972 6920 21984
rect 6972 21972 6978 22024
rect 10226 22012 10232 22024
rect 10187 21984 10232 22012
rect 10226 21972 10232 21984
rect 10284 21972 10290 22024
rect 6273 21947 6331 21953
rect 6273 21913 6285 21947
rect 6319 21944 6331 21947
rect 7558 21944 7564 21956
rect 6319 21916 7564 21944
rect 6319 21913 6331 21916
rect 6273 21907 6331 21913
rect 7558 21904 7564 21916
rect 7616 21904 7622 21956
rect 5718 21876 5724 21888
rect 5679 21848 5724 21876
rect 5718 21836 5724 21848
rect 5776 21836 5782 21888
rect 7929 21879 7987 21885
rect 7929 21845 7941 21879
rect 7975 21876 7987 21879
rect 8478 21876 8484 21888
rect 7975 21848 8484 21876
rect 7975 21845 7987 21848
rect 7929 21839 7987 21845
rect 8478 21836 8484 21848
rect 8536 21836 8542 21888
rect 9950 21836 9956 21888
rect 10008 21876 10014 21888
rect 11609 21879 11667 21885
rect 11609 21876 11621 21879
rect 10008 21848 11621 21876
rect 10008 21836 10014 21848
rect 11609 21845 11621 21848
rect 11655 21845 11667 21879
rect 11609 21839 11667 21845
rect 1104 21786 14812 21808
rect 1104 21734 3648 21786
rect 3700 21734 3712 21786
rect 3764 21734 3776 21786
rect 3828 21734 3840 21786
rect 3892 21734 8982 21786
rect 9034 21734 9046 21786
rect 9098 21734 9110 21786
rect 9162 21734 9174 21786
rect 9226 21734 14315 21786
rect 14367 21734 14379 21786
rect 14431 21734 14443 21786
rect 14495 21734 14507 21786
rect 14559 21734 14812 21786
rect 1104 21712 14812 21734
rect 3789 21675 3847 21681
rect 3789 21641 3801 21675
rect 3835 21672 3847 21675
rect 4062 21672 4068 21684
rect 3835 21644 4068 21672
rect 3835 21641 3847 21644
rect 3789 21635 3847 21641
rect 4062 21632 4068 21644
rect 4120 21632 4126 21684
rect 4798 21672 4804 21684
rect 4759 21644 4804 21672
rect 4798 21632 4804 21644
rect 4856 21632 4862 21684
rect 4982 21672 4988 21684
rect 4895 21644 4988 21672
rect 4709 21607 4767 21613
rect 4709 21573 4721 21607
rect 4755 21604 4767 21607
rect 4908 21604 4936 21644
rect 4982 21632 4988 21644
rect 5040 21672 5046 21684
rect 5166 21672 5172 21684
rect 5040 21644 5172 21672
rect 5040 21632 5046 21644
rect 5166 21632 5172 21644
rect 5224 21632 5230 21684
rect 5534 21632 5540 21684
rect 5592 21672 5598 21684
rect 6270 21672 6276 21684
rect 5592 21644 6276 21672
rect 5592 21632 5598 21644
rect 6270 21632 6276 21644
rect 6328 21632 6334 21684
rect 6457 21675 6515 21681
rect 6457 21641 6469 21675
rect 6503 21672 6515 21675
rect 7466 21672 7472 21684
rect 6503 21644 7472 21672
rect 6503 21641 6515 21644
rect 6457 21635 6515 21641
rect 7466 21632 7472 21644
rect 7524 21632 7530 21684
rect 10318 21672 10324 21684
rect 10279 21644 10324 21672
rect 10318 21632 10324 21644
rect 10376 21632 10382 21684
rect 4755 21576 4936 21604
rect 4755 21573 4767 21576
rect 4709 21567 4767 21573
rect 1578 21536 1584 21548
rect 1539 21508 1584 21536
rect 1578 21496 1584 21508
rect 1636 21496 1642 21548
rect 5166 21496 5172 21548
rect 5224 21496 5230 21548
rect 5350 21536 5356 21548
rect 5311 21508 5356 21536
rect 5350 21496 5356 21508
rect 5408 21536 5414 21548
rect 5718 21536 5724 21548
rect 5408 21508 5724 21536
rect 5408 21496 5414 21508
rect 5718 21496 5724 21508
rect 5776 21536 5782 21548
rect 5905 21539 5963 21545
rect 5905 21536 5917 21539
rect 5776 21508 5917 21536
rect 5776 21496 5782 21508
rect 5905 21505 5917 21508
rect 5951 21505 5963 21539
rect 5905 21499 5963 21505
rect 1397 21471 1455 21477
rect 1397 21437 1409 21471
rect 1443 21468 1455 21471
rect 1443 21440 2268 21468
rect 1443 21437 1455 21440
rect 1397 21431 1455 21437
rect 2240 21341 2268 21440
rect 4338 21428 4344 21480
rect 4396 21468 4402 21480
rect 5184 21468 5212 21496
rect 5261 21471 5319 21477
rect 5261 21468 5273 21471
rect 4396 21440 5273 21468
rect 4396 21428 4402 21440
rect 5261 21437 5273 21440
rect 5307 21437 5319 21471
rect 5261 21431 5319 21437
rect 6641 21471 6699 21477
rect 6641 21437 6653 21471
rect 6687 21468 6699 21471
rect 6730 21468 6736 21480
rect 6687 21440 6736 21468
rect 6687 21437 6699 21440
rect 6641 21431 6699 21437
rect 6730 21428 6736 21440
rect 6788 21428 6794 21480
rect 8478 21468 8484 21480
rect 8439 21440 8484 21468
rect 8478 21428 8484 21440
rect 8536 21428 8542 21480
rect 4982 21360 4988 21412
rect 5040 21400 5046 21412
rect 5169 21403 5227 21409
rect 5169 21400 5181 21403
rect 5040 21372 5181 21400
rect 5040 21360 5046 21372
rect 5169 21369 5181 21372
rect 5215 21400 5227 21403
rect 5718 21400 5724 21412
rect 5215 21372 5724 21400
rect 5215 21369 5227 21372
rect 5169 21363 5227 21369
rect 5718 21360 5724 21372
rect 5776 21360 5782 21412
rect 7098 21400 7104 21412
rect 7011 21372 7104 21400
rect 7098 21360 7104 21372
rect 7156 21400 7162 21412
rect 7558 21400 7564 21412
rect 7156 21372 7564 21400
rect 7156 21360 7162 21372
rect 7558 21360 7564 21372
rect 7616 21360 7622 21412
rect 8389 21403 8447 21409
rect 8389 21369 8401 21403
rect 8435 21400 8447 21403
rect 8726 21403 8784 21409
rect 8726 21400 8738 21403
rect 8435 21372 8738 21400
rect 8435 21369 8447 21372
rect 8389 21363 8447 21369
rect 8726 21369 8738 21372
rect 8772 21400 8784 21403
rect 8846 21400 8852 21412
rect 8772 21372 8852 21400
rect 8772 21369 8784 21372
rect 8726 21363 8784 21369
rect 8846 21360 8852 21372
rect 8904 21360 8910 21412
rect 2225 21335 2283 21341
rect 2225 21301 2237 21335
rect 2271 21332 2283 21335
rect 2406 21332 2412 21344
rect 2271 21304 2412 21332
rect 2271 21301 2283 21304
rect 2225 21295 2283 21301
rect 2406 21292 2412 21304
rect 2464 21292 2470 21344
rect 4154 21332 4160 21344
rect 4115 21304 4160 21332
rect 4154 21292 4160 21304
rect 4212 21292 4218 21344
rect 7466 21332 7472 21344
rect 7427 21304 7472 21332
rect 7466 21292 7472 21304
rect 7524 21292 7530 21344
rect 9398 21292 9404 21344
rect 9456 21332 9462 21344
rect 9861 21335 9919 21341
rect 9861 21332 9873 21335
rect 9456 21304 9873 21332
rect 9456 21292 9462 21304
rect 9861 21301 9873 21304
rect 9907 21301 9919 21335
rect 9861 21295 9919 21301
rect 10226 21292 10232 21344
rect 10284 21332 10290 21344
rect 10689 21335 10747 21341
rect 10689 21332 10701 21335
rect 10284 21304 10701 21332
rect 10284 21292 10290 21304
rect 10689 21301 10701 21304
rect 10735 21332 10747 21335
rect 11974 21332 11980 21344
rect 10735 21304 11980 21332
rect 10735 21301 10747 21304
rect 10689 21295 10747 21301
rect 11974 21292 11980 21304
rect 12032 21292 12038 21344
rect 1104 21242 14812 21264
rect 1104 21190 6315 21242
rect 6367 21190 6379 21242
rect 6431 21190 6443 21242
rect 6495 21190 6507 21242
rect 6559 21190 11648 21242
rect 11700 21190 11712 21242
rect 11764 21190 11776 21242
rect 11828 21190 11840 21242
rect 11892 21190 14812 21242
rect 1104 21168 14812 21190
rect 2590 21088 2596 21140
rect 2648 21128 2654 21140
rect 2685 21131 2743 21137
rect 2685 21128 2697 21131
rect 2648 21100 2697 21128
rect 2648 21088 2654 21100
rect 2685 21097 2697 21100
rect 2731 21128 2743 21131
rect 4062 21128 4068 21140
rect 2731 21100 4068 21128
rect 2731 21097 2743 21100
rect 2685 21091 2743 21097
rect 4062 21088 4068 21100
rect 4120 21088 4126 21140
rect 5166 21128 5172 21140
rect 5127 21100 5172 21128
rect 5166 21088 5172 21100
rect 5224 21088 5230 21140
rect 6549 21131 6607 21137
rect 6549 21097 6561 21131
rect 6595 21128 6607 21131
rect 6730 21128 6736 21140
rect 6595 21100 6736 21128
rect 6595 21097 6607 21100
rect 6549 21091 6607 21097
rect 6730 21088 6736 21100
rect 6788 21088 6794 21140
rect 8846 21088 8852 21140
rect 8904 21128 8910 21140
rect 11057 21131 11115 21137
rect 11057 21128 11069 21131
rect 8904 21100 11069 21128
rect 8904 21088 8910 21100
rect 11057 21097 11069 21100
rect 11103 21128 11115 21131
rect 11238 21128 11244 21140
rect 11103 21100 11244 21128
rect 11103 21097 11115 21100
rect 11057 21091 11115 21097
rect 11238 21088 11244 21100
rect 11296 21088 11302 21140
rect 1670 21060 1676 21072
rect 1631 21032 1676 21060
rect 1670 21020 1676 21032
rect 1728 21020 1734 21072
rect 4893 21063 4951 21069
rect 4893 21029 4905 21063
rect 4939 21060 4951 21063
rect 5350 21060 5356 21072
rect 4939 21032 5356 21060
rect 4939 21029 4951 21032
rect 4893 21023 4951 21029
rect 5350 21020 5356 21032
rect 5408 21020 5414 21072
rect 5442 21020 5448 21072
rect 5500 21060 5506 21072
rect 8754 21060 8760 21072
rect 5500 21032 8760 21060
rect 5500 21020 5506 21032
rect 8754 21020 8760 21032
rect 8812 21020 8818 21072
rect 9950 21069 9956 21072
rect 9944 21060 9956 21069
rect 9911 21032 9956 21060
rect 9944 21023 9956 21032
rect 9950 21020 9956 21023
rect 10008 21020 10014 21072
rect 12066 21020 12072 21072
rect 12124 21069 12130 21072
rect 12124 21063 12188 21069
rect 12124 21029 12142 21063
rect 12176 21029 12188 21063
rect 12124 21023 12188 21029
rect 12124 21020 12130 21023
rect 1397 20995 1455 21001
rect 1397 20961 1409 20995
rect 1443 20992 1455 20995
rect 1443 20964 1716 20992
rect 1443 20961 1455 20964
rect 1397 20955 1455 20961
rect 1688 20936 1716 20964
rect 3970 20952 3976 21004
rect 4028 20992 4034 21004
rect 7098 20992 7104 21004
rect 4028 20964 7104 20992
rect 4028 20952 4034 20964
rect 7098 20952 7104 20964
rect 7156 20952 7162 21004
rect 7466 20952 7472 21004
rect 7524 20992 7530 21004
rect 7745 20995 7803 21001
rect 7745 20992 7757 20995
rect 7524 20964 7757 20992
rect 7524 20952 7530 20964
rect 7745 20961 7757 20964
rect 7791 20992 7803 20995
rect 8202 20992 8208 21004
rect 7791 20964 8208 20992
rect 7791 20961 7803 20964
rect 7745 20955 7803 20961
rect 8202 20952 8208 20964
rect 8260 20952 8266 21004
rect 8478 20952 8484 21004
rect 8536 20992 8542 21004
rect 8573 20995 8631 21001
rect 8573 20992 8585 20995
rect 8536 20964 8585 20992
rect 8536 20952 8542 20964
rect 8573 20961 8585 20964
rect 8619 20992 8631 20995
rect 9125 20995 9183 21001
rect 9125 20992 9137 20995
rect 8619 20964 9137 20992
rect 8619 20961 8631 20964
rect 8573 20955 8631 20961
rect 9125 20961 9137 20964
rect 9171 20992 9183 20995
rect 9677 20995 9735 21001
rect 9677 20992 9689 20995
rect 9171 20964 9689 20992
rect 9171 20961 9183 20964
rect 9125 20955 9183 20961
rect 9677 20961 9689 20964
rect 9723 20992 9735 20995
rect 10226 20992 10232 21004
rect 9723 20964 10232 20992
rect 9723 20961 9735 20964
rect 9677 20955 9735 20961
rect 10226 20952 10232 20964
rect 10284 20952 10290 21004
rect 11885 20995 11943 21001
rect 11885 20961 11897 20995
rect 11931 20992 11943 20995
rect 11974 20992 11980 21004
rect 11931 20964 11980 20992
rect 11931 20961 11943 20964
rect 11885 20955 11943 20961
rect 11974 20952 11980 20964
rect 12032 20952 12038 21004
rect 1670 20884 1676 20936
rect 1728 20884 1734 20936
rect 6914 20884 6920 20936
rect 6972 20924 6978 20936
rect 7650 20924 7656 20936
rect 6972 20896 7656 20924
rect 6972 20884 6978 20896
rect 7650 20884 7656 20896
rect 7708 20924 7714 20936
rect 7837 20927 7895 20933
rect 7837 20924 7849 20927
rect 7708 20896 7849 20924
rect 7708 20884 7714 20896
rect 7837 20893 7849 20896
rect 7883 20893 7895 20927
rect 8018 20924 8024 20936
rect 7979 20896 8024 20924
rect 7837 20887 7895 20893
rect 8018 20884 8024 20896
rect 8076 20884 8082 20936
rect 7009 20859 7067 20865
rect 7009 20825 7021 20859
rect 7055 20856 7067 20859
rect 8036 20856 8064 20884
rect 7055 20828 8064 20856
rect 7055 20825 7067 20828
rect 7009 20819 7067 20825
rect 7374 20788 7380 20800
rect 7335 20760 7380 20788
rect 7374 20748 7380 20760
rect 7432 20748 7438 20800
rect 9493 20791 9551 20797
rect 9493 20757 9505 20791
rect 9539 20788 9551 20791
rect 9582 20788 9588 20800
rect 9539 20760 9588 20788
rect 9539 20757 9551 20760
rect 9493 20751 9551 20757
rect 9582 20748 9588 20760
rect 9640 20748 9646 20800
rect 12526 20748 12532 20800
rect 12584 20788 12590 20800
rect 13265 20791 13323 20797
rect 13265 20788 13277 20791
rect 12584 20760 13277 20788
rect 12584 20748 12590 20760
rect 13265 20757 13277 20760
rect 13311 20757 13323 20791
rect 13265 20751 13323 20757
rect 1104 20698 14812 20720
rect 1104 20646 3648 20698
rect 3700 20646 3712 20698
rect 3764 20646 3776 20698
rect 3828 20646 3840 20698
rect 3892 20646 8982 20698
rect 9034 20646 9046 20698
rect 9098 20646 9110 20698
rect 9162 20646 9174 20698
rect 9226 20646 14315 20698
rect 14367 20646 14379 20698
rect 14431 20646 14443 20698
rect 14495 20646 14507 20698
rect 14559 20646 14812 20698
rect 1104 20624 14812 20646
rect 5902 20584 5908 20596
rect 5863 20556 5908 20584
rect 5902 20544 5908 20556
rect 5960 20544 5966 20596
rect 6641 20587 6699 20593
rect 6641 20553 6653 20587
rect 6687 20584 6699 20587
rect 6822 20584 6828 20596
rect 6687 20556 6828 20584
rect 6687 20553 6699 20556
rect 6641 20547 6699 20553
rect 6822 20544 6828 20556
rect 6880 20544 6886 20596
rect 8294 20544 8300 20596
rect 8352 20584 8358 20596
rect 8573 20587 8631 20593
rect 8573 20584 8585 20587
rect 8352 20556 8585 20584
rect 8352 20544 8358 20556
rect 8573 20553 8585 20556
rect 8619 20553 8631 20587
rect 8573 20547 8631 20553
rect 9033 20587 9091 20593
rect 9033 20553 9045 20587
rect 9079 20584 9091 20587
rect 9398 20584 9404 20596
rect 9079 20556 9404 20584
rect 9079 20553 9091 20556
rect 9033 20547 9091 20553
rect 2590 20448 2596 20460
rect 2551 20420 2596 20448
rect 2590 20408 2596 20420
rect 2648 20408 2654 20460
rect 5920 20448 5948 20544
rect 8018 20476 8024 20528
rect 8076 20516 8082 20528
rect 9048 20516 9076 20547
rect 9398 20544 9404 20556
rect 9456 20544 9462 20596
rect 9766 20544 9772 20596
rect 9824 20584 9830 20596
rect 10226 20584 10232 20596
rect 9824 20556 10232 20584
rect 9824 20544 9830 20556
rect 10226 20544 10232 20556
rect 10284 20544 10290 20596
rect 8076 20488 9076 20516
rect 11149 20519 11207 20525
rect 8076 20476 8082 20488
rect 11149 20485 11161 20519
rect 11195 20516 11207 20519
rect 12434 20516 12440 20528
rect 11195 20488 12440 20516
rect 11195 20485 11207 20488
rect 11149 20479 11207 20485
rect 12434 20476 12440 20488
rect 12492 20516 12498 20528
rect 12492 20488 12585 20516
rect 12492 20476 12498 20488
rect 6917 20451 6975 20457
rect 6917 20448 6929 20451
rect 5920 20420 6929 20448
rect 6917 20417 6929 20420
rect 6963 20417 6975 20451
rect 6917 20411 6975 20417
rect 5534 20340 5540 20392
rect 5592 20380 5598 20392
rect 5902 20380 5908 20392
rect 5592 20352 5908 20380
rect 5592 20340 5598 20352
rect 5902 20340 5908 20352
rect 5960 20340 5966 20392
rect 6086 20340 6092 20392
rect 6144 20380 6150 20392
rect 6822 20380 6828 20392
rect 6144 20352 6828 20380
rect 6144 20340 6150 20352
rect 6822 20340 6828 20352
rect 6880 20340 6886 20392
rect 7184 20383 7242 20389
rect 7184 20349 7196 20383
rect 7230 20380 7242 20383
rect 8036 20380 8064 20476
rect 9401 20451 9459 20457
rect 9401 20417 9413 20451
rect 9447 20448 9459 20451
rect 9769 20451 9827 20457
rect 9769 20448 9781 20451
rect 9447 20420 9781 20448
rect 9447 20417 9459 20420
rect 9401 20411 9459 20417
rect 9769 20417 9781 20420
rect 9815 20448 9827 20451
rect 9950 20448 9956 20460
rect 9815 20420 9956 20448
rect 9815 20417 9827 20420
rect 9769 20411 9827 20417
rect 9950 20408 9956 20420
rect 10008 20448 10014 20460
rect 10413 20451 10471 20457
rect 10413 20448 10425 20451
rect 10008 20420 10425 20448
rect 10008 20408 10014 20420
rect 10413 20417 10425 20420
rect 10459 20417 10471 20451
rect 10413 20411 10471 20417
rect 10870 20408 10876 20460
rect 10928 20448 10934 20460
rect 11793 20451 11851 20457
rect 11793 20448 11805 20451
rect 10928 20420 11805 20448
rect 10928 20408 10934 20420
rect 11793 20417 11805 20420
rect 11839 20448 11851 20451
rect 11977 20451 12035 20457
rect 11977 20448 11989 20451
rect 11839 20420 11989 20448
rect 11839 20417 11851 20420
rect 11793 20411 11851 20417
rect 11977 20417 11989 20420
rect 12023 20417 12035 20451
rect 12250 20448 12256 20460
rect 12163 20420 12256 20448
rect 11977 20411 12035 20417
rect 12250 20408 12256 20420
rect 12308 20448 12314 20460
rect 12894 20448 12900 20460
rect 12308 20420 12900 20448
rect 12308 20408 12314 20420
rect 12894 20408 12900 20420
rect 12952 20408 12958 20460
rect 12989 20451 13047 20457
rect 12989 20417 13001 20451
rect 13035 20417 13047 20451
rect 12989 20411 13047 20417
rect 9858 20380 9864 20392
rect 7230 20352 8064 20380
rect 9784 20352 9864 20380
rect 7230 20349 7242 20352
rect 7184 20343 7242 20349
rect 9784 20324 9812 20352
rect 9858 20340 9864 20352
rect 9916 20340 9922 20392
rect 10226 20380 10232 20392
rect 10187 20352 10232 20380
rect 10226 20340 10232 20352
rect 10284 20340 10290 20392
rect 12066 20380 12072 20392
rect 11440 20352 12072 20380
rect 2501 20315 2559 20321
rect 2501 20281 2513 20315
rect 2547 20312 2559 20315
rect 2838 20315 2896 20321
rect 2838 20312 2850 20315
rect 2547 20284 2850 20312
rect 2547 20281 2559 20284
rect 2501 20275 2559 20281
rect 2838 20281 2850 20284
rect 2884 20312 2896 20315
rect 3510 20312 3516 20324
rect 2884 20284 3516 20312
rect 2884 20281 2896 20284
rect 2838 20275 2896 20281
rect 3510 20272 3516 20284
rect 3568 20272 3574 20324
rect 6273 20315 6331 20321
rect 6273 20281 6285 20315
rect 6319 20312 6331 20315
rect 6319 20284 7144 20312
rect 6319 20281 6331 20284
rect 6273 20275 6331 20281
rect 1670 20244 1676 20256
rect 1631 20216 1676 20244
rect 1670 20204 1676 20216
rect 1728 20204 1734 20256
rect 2958 20204 2964 20256
rect 3016 20244 3022 20256
rect 3973 20247 4031 20253
rect 3973 20244 3985 20247
rect 3016 20216 3985 20244
rect 3016 20204 3022 20216
rect 3973 20213 3985 20216
rect 4019 20244 4031 20247
rect 4154 20244 4160 20256
rect 4019 20216 4160 20244
rect 4019 20213 4031 20216
rect 3973 20207 4031 20213
rect 4154 20204 4160 20216
rect 4212 20204 4218 20256
rect 7116 20244 7144 20284
rect 9766 20272 9772 20324
rect 9824 20272 9830 20324
rect 7282 20244 7288 20256
rect 7116 20216 7288 20244
rect 7282 20204 7288 20216
rect 7340 20204 7346 20256
rect 8294 20244 8300 20256
rect 8255 20216 8300 20244
rect 8294 20204 8300 20216
rect 8352 20204 8358 20256
rect 9674 20204 9680 20256
rect 9732 20244 9738 20256
rect 9861 20247 9919 20253
rect 9861 20244 9873 20247
rect 9732 20216 9873 20244
rect 9732 20204 9738 20216
rect 9861 20213 9873 20216
rect 9907 20213 9919 20247
rect 9861 20207 9919 20213
rect 10318 20204 10324 20256
rect 10376 20244 10382 20256
rect 10376 20216 10421 20244
rect 10376 20204 10382 20216
rect 11330 20204 11336 20256
rect 11388 20244 11394 20256
rect 11440 20253 11468 20352
rect 12066 20340 12072 20352
rect 12124 20380 12130 20392
rect 13004 20380 13032 20411
rect 13170 20380 13176 20392
rect 12124 20352 13176 20380
rect 12124 20340 12130 20352
rect 13170 20340 13176 20352
rect 13228 20380 13234 20392
rect 13449 20383 13507 20389
rect 13449 20380 13461 20383
rect 13228 20352 13461 20380
rect 13228 20340 13234 20352
rect 13449 20349 13461 20352
rect 13495 20349 13507 20383
rect 13449 20343 13507 20349
rect 11977 20315 12035 20321
rect 11977 20281 11989 20315
rect 12023 20312 12035 20315
rect 12805 20315 12863 20321
rect 12805 20312 12817 20315
rect 12023 20284 12817 20312
rect 12023 20281 12035 20284
rect 11977 20275 12035 20281
rect 12805 20281 12817 20284
rect 12851 20281 12863 20315
rect 12805 20275 12863 20281
rect 11425 20247 11483 20253
rect 11425 20244 11437 20247
rect 11388 20216 11437 20244
rect 11388 20204 11394 20216
rect 11425 20213 11437 20216
rect 11471 20213 11483 20247
rect 11425 20207 11483 20213
rect 1104 20154 14812 20176
rect 1104 20102 6315 20154
rect 6367 20102 6379 20154
rect 6431 20102 6443 20154
rect 6495 20102 6507 20154
rect 6559 20102 11648 20154
rect 11700 20102 11712 20154
rect 11764 20102 11776 20154
rect 11828 20102 11840 20154
rect 11892 20102 14812 20154
rect 1104 20080 14812 20102
rect 2406 20040 2412 20052
rect 2367 20012 2412 20040
rect 2406 20000 2412 20012
rect 2464 20000 2470 20052
rect 6086 20040 6092 20052
rect 6047 20012 6092 20040
rect 6086 20000 6092 20012
rect 6144 20000 6150 20052
rect 6917 20043 6975 20049
rect 6917 20040 6929 20043
rect 6564 20012 6929 20040
rect 2866 19972 2872 19984
rect 2827 19944 2872 19972
rect 2866 19932 2872 19944
rect 2924 19932 2930 19984
rect 2774 19864 2780 19916
rect 2832 19904 2838 19916
rect 2832 19876 2877 19904
rect 2832 19864 2838 19876
rect 4798 19864 4804 19916
rect 4856 19904 4862 19916
rect 4893 19907 4951 19913
rect 4893 19904 4905 19907
rect 4856 19876 4905 19904
rect 4856 19864 4862 19876
rect 4893 19873 4905 19876
rect 4939 19873 4951 19907
rect 4893 19867 4951 19873
rect 4985 19907 5043 19913
rect 4985 19873 4997 19907
rect 5031 19904 5043 19907
rect 5258 19904 5264 19916
rect 5031 19876 5264 19904
rect 5031 19873 5043 19876
rect 4985 19867 5043 19873
rect 5258 19864 5264 19876
rect 5316 19864 5322 19916
rect 5534 19864 5540 19916
rect 5592 19904 5598 19916
rect 6454 19904 6460 19916
rect 5592 19876 6460 19904
rect 5592 19864 5598 19876
rect 6454 19864 6460 19876
rect 6512 19864 6518 19916
rect 2958 19836 2964 19848
rect 2919 19808 2964 19836
rect 2958 19796 2964 19808
rect 3016 19796 3022 19848
rect 5166 19836 5172 19848
rect 5127 19808 5172 19836
rect 5166 19796 5172 19808
rect 5224 19796 5230 19848
rect 6564 19845 6592 20012
rect 6917 20009 6929 20012
rect 6963 20009 6975 20043
rect 6917 20003 6975 20009
rect 7374 20000 7380 20052
rect 7432 20040 7438 20052
rect 7834 20040 7840 20052
rect 7432 20012 7840 20040
rect 7432 20000 7438 20012
rect 7834 20000 7840 20012
rect 7892 20040 7898 20052
rect 8113 20043 8171 20049
rect 8113 20040 8125 20043
rect 7892 20012 8125 20040
rect 7892 20000 7898 20012
rect 8113 20009 8125 20012
rect 8159 20009 8171 20043
rect 8113 20003 8171 20009
rect 8846 20000 8852 20052
rect 8904 20040 8910 20052
rect 9125 20043 9183 20049
rect 9125 20040 9137 20043
rect 8904 20012 9137 20040
rect 8904 20000 8910 20012
rect 9125 20009 9137 20012
rect 9171 20009 9183 20043
rect 9125 20003 9183 20009
rect 9953 20043 10011 20049
rect 9953 20009 9965 20043
rect 9999 20040 10011 20043
rect 10318 20040 10324 20052
rect 9999 20012 10324 20040
rect 9999 20009 10011 20012
rect 9953 20003 10011 20009
rect 10318 20000 10324 20012
rect 10376 20000 10382 20052
rect 11425 20043 11483 20049
rect 11425 20009 11437 20043
rect 11471 20040 11483 20043
rect 12434 20040 12440 20052
rect 11471 20012 12440 20040
rect 11471 20009 11483 20012
rect 11425 20003 11483 20009
rect 12434 20000 12440 20012
rect 12492 20000 12498 20052
rect 10045 19975 10103 19981
rect 10045 19941 10057 19975
rect 10091 19972 10103 19975
rect 10870 19972 10876 19984
rect 10091 19944 10876 19972
rect 10091 19941 10103 19944
rect 10045 19935 10103 19941
rect 10870 19932 10876 19944
rect 10928 19932 10934 19984
rect 11882 19932 11888 19984
rect 11940 19972 11946 19984
rect 12069 19975 12127 19981
rect 12069 19972 12081 19975
rect 11940 19944 12081 19972
rect 11940 19932 11946 19944
rect 12069 19941 12081 19944
rect 12115 19941 12127 19975
rect 12069 19935 12127 19941
rect 12158 19932 12164 19984
rect 12216 19972 12222 19984
rect 12253 19975 12311 19981
rect 12253 19972 12265 19975
rect 12216 19944 12265 19972
rect 12216 19932 12222 19944
rect 12253 19941 12265 19944
rect 12299 19941 12311 19975
rect 12253 19935 12311 19941
rect 7282 19904 7288 19916
rect 7243 19876 7288 19904
rect 7282 19864 7288 19876
rect 7340 19864 7346 19916
rect 11517 19907 11575 19913
rect 11517 19904 11529 19907
rect 7576 19876 8340 19904
rect 5629 19839 5687 19845
rect 5629 19805 5641 19839
rect 5675 19836 5687 19839
rect 6549 19839 6607 19845
rect 6549 19836 6561 19839
rect 5675 19808 6561 19836
rect 5675 19805 5687 19808
rect 5629 19799 5687 19805
rect 6549 19805 6561 19808
rect 6595 19805 6607 19839
rect 6549 19799 6607 19805
rect 6641 19839 6699 19845
rect 6641 19805 6653 19839
rect 6687 19805 6699 19839
rect 6641 19799 6699 19805
rect 7377 19839 7435 19845
rect 7377 19805 7389 19839
rect 7423 19836 7435 19839
rect 7466 19836 7472 19848
rect 7423 19808 7472 19836
rect 7423 19805 7435 19808
rect 7377 19799 7435 19805
rect 6086 19728 6092 19780
rect 6144 19768 6150 19780
rect 6656 19768 6684 19799
rect 7466 19796 7472 19808
rect 7524 19796 7530 19848
rect 7576 19845 7604 19876
rect 8312 19848 8340 19876
rect 11440 19876 11529 19904
rect 7561 19839 7619 19845
rect 7561 19805 7573 19839
rect 7607 19805 7619 19839
rect 8202 19836 8208 19848
rect 8163 19808 8208 19836
rect 7561 19799 7619 19805
rect 8202 19796 8208 19808
rect 8260 19796 8266 19848
rect 8294 19796 8300 19848
rect 8352 19836 8358 19848
rect 8352 19808 8397 19836
rect 8352 19796 8358 19808
rect 9950 19796 9956 19848
rect 10008 19836 10014 19848
rect 10502 19836 10508 19848
rect 10008 19808 10508 19836
rect 10008 19796 10014 19808
rect 10502 19796 10508 19808
rect 10560 19796 10566 19848
rect 6144 19740 6684 19768
rect 6144 19728 6150 19740
rect 7006 19728 7012 19780
rect 7064 19768 7070 19780
rect 7745 19771 7803 19777
rect 7745 19768 7757 19771
rect 7064 19740 7757 19768
rect 7064 19728 7070 19740
rect 7745 19737 7757 19740
rect 7791 19737 7803 19771
rect 7745 19731 7803 19737
rect 10226 19728 10232 19780
rect 10284 19768 10290 19780
rect 11057 19771 11115 19777
rect 11057 19768 11069 19771
rect 10284 19740 11069 19768
rect 10284 19728 10290 19740
rect 11057 19737 11069 19740
rect 11103 19737 11115 19771
rect 11440 19768 11468 19876
rect 11517 19873 11529 19876
rect 11563 19873 11575 19907
rect 11517 19867 11575 19873
rect 11790 19864 11796 19916
rect 11848 19904 11854 19916
rect 12437 19907 12495 19913
rect 12437 19904 12449 19907
rect 11848 19876 12449 19904
rect 11848 19864 11854 19876
rect 12437 19873 12449 19876
rect 12483 19873 12495 19907
rect 12437 19867 12495 19873
rect 11606 19836 11612 19848
rect 11567 19808 11612 19836
rect 11606 19796 11612 19808
rect 11664 19836 11670 19848
rect 12342 19836 12348 19848
rect 11664 19808 12348 19836
rect 11664 19796 11670 19808
rect 12342 19796 12348 19808
rect 12400 19796 12406 19848
rect 12452 19836 12480 19867
rect 12618 19864 12624 19916
rect 12676 19904 12682 19916
rect 12986 19904 12992 19916
rect 12676 19876 12992 19904
rect 12676 19864 12682 19876
rect 12986 19864 12992 19876
rect 13044 19864 13050 19916
rect 12526 19836 12532 19848
rect 12452 19808 12532 19836
rect 12526 19796 12532 19808
rect 12584 19796 12590 19848
rect 13078 19836 13084 19848
rect 13039 19808 13084 19836
rect 13078 19796 13084 19808
rect 13136 19796 13142 19848
rect 13170 19796 13176 19848
rect 13228 19836 13234 19848
rect 13228 19808 13273 19836
rect 13228 19796 13234 19808
rect 11514 19768 11520 19780
rect 11440 19740 11520 19768
rect 11057 19731 11115 19737
rect 11514 19728 11520 19740
rect 11572 19768 11578 19780
rect 12621 19771 12679 19777
rect 12621 19768 12633 19771
rect 11572 19740 12633 19768
rect 11572 19728 11578 19740
rect 12621 19737 12633 19740
rect 12667 19737 12679 19771
rect 12621 19731 12679 19737
rect 3881 19703 3939 19709
rect 3881 19669 3893 19703
rect 3927 19700 3939 19703
rect 4246 19700 4252 19712
rect 3927 19672 4252 19700
rect 3927 19669 3939 19672
rect 3881 19663 3939 19669
rect 4246 19660 4252 19672
rect 4304 19700 4310 19712
rect 4525 19703 4583 19709
rect 4525 19700 4537 19703
rect 4304 19672 4537 19700
rect 4304 19660 4310 19672
rect 4525 19669 4537 19672
rect 4571 19669 4583 19703
rect 4525 19663 4583 19669
rect 5997 19703 6055 19709
rect 5997 19669 6009 19703
rect 6043 19700 6055 19703
rect 7466 19700 7472 19712
rect 6043 19672 7472 19700
rect 6043 19669 6055 19672
rect 5997 19663 6055 19669
rect 7466 19660 7472 19672
rect 7524 19660 7530 19712
rect 8754 19700 8760 19712
rect 8715 19672 8760 19700
rect 8754 19660 8760 19672
rect 8812 19660 8818 19712
rect 10502 19700 10508 19712
rect 10463 19672 10508 19700
rect 10502 19660 10508 19672
rect 10560 19660 10566 19712
rect 10870 19700 10876 19712
rect 10831 19672 10876 19700
rect 10870 19660 10876 19672
rect 10928 19660 10934 19712
rect 12158 19660 12164 19712
rect 12216 19700 12222 19712
rect 12253 19703 12311 19709
rect 12253 19700 12265 19703
rect 12216 19672 12265 19700
rect 12216 19660 12222 19672
rect 12253 19669 12265 19672
rect 12299 19669 12311 19703
rect 12253 19663 12311 19669
rect 1104 19610 14812 19632
rect 1104 19558 3648 19610
rect 3700 19558 3712 19610
rect 3764 19558 3776 19610
rect 3828 19558 3840 19610
rect 3892 19558 8982 19610
rect 9034 19558 9046 19610
rect 9098 19558 9110 19610
rect 9162 19558 9174 19610
rect 9226 19558 14315 19610
rect 14367 19558 14379 19610
rect 14431 19558 14443 19610
rect 14495 19558 14507 19610
rect 14559 19558 14812 19610
rect 1104 19536 14812 19558
rect 10045 19499 10103 19505
rect 10045 19465 10057 19499
rect 10091 19496 10103 19499
rect 10318 19496 10324 19508
rect 10091 19468 10324 19496
rect 10091 19465 10103 19468
rect 10045 19459 10103 19465
rect 10318 19456 10324 19468
rect 10376 19456 10382 19508
rect 11514 19496 11520 19508
rect 11475 19468 11520 19496
rect 11514 19456 11520 19468
rect 11572 19456 11578 19508
rect 2774 19388 2780 19440
rect 2832 19428 2838 19440
rect 3789 19431 3847 19437
rect 3789 19428 3801 19431
rect 2832 19400 3801 19428
rect 2832 19388 2838 19400
rect 3789 19397 3801 19400
rect 3835 19397 3847 19431
rect 3789 19391 3847 19397
rect 7377 19431 7435 19437
rect 7377 19397 7389 19431
rect 7423 19428 7435 19431
rect 8202 19428 8208 19440
rect 7423 19400 8208 19428
rect 7423 19397 7435 19400
rect 7377 19391 7435 19397
rect 8202 19388 8208 19400
rect 8260 19388 8266 19440
rect 9953 19431 10011 19437
rect 9953 19397 9965 19431
rect 9999 19428 10011 19431
rect 10410 19428 10416 19440
rect 9999 19400 10416 19428
rect 9999 19397 10011 19400
rect 9953 19391 10011 19397
rect 10410 19388 10416 19400
rect 10468 19428 10474 19440
rect 11057 19431 11115 19437
rect 11057 19428 11069 19431
rect 10468 19400 11069 19428
rect 10468 19388 10474 19400
rect 2958 19360 2964 19372
rect 2700 19332 2964 19360
rect 1394 19292 1400 19304
rect 1355 19264 1400 19292
rect 1394 19252 1400 19264
rect 1452 19252 1458 19304
rect 1670 19292 1676 19304
rect 1631 19264 1676 19292
rect 1670 19252 1676 19264
rect 1728 19252 1734 19304
rect 2501 19295 2559 19301
rect 2501 19261 2513 19295
rect 2547 19292 2559 19295
rect 2700 19292 2728 19332
rect 2958 19320 2964 19332
rect 3016 19320 3022 19372
rect 4246 19360 4252 19372
rect 4207 19332 4252 19360
rect 4246 19320 4252 19332
rect 4304 19320 4310 19372
rect 4341 19363 4399 19369
rect 4341 19329 4353 19363
rect 4387 19329 4399 19363
rect 8018 19360 8024 19372
rect 7979 19332 8024 19360
rect 4341 19323 4399 19329
rect 2547 19264 2728 19292
rect 2547 19261 2559 19264
rect 2501 19255 2559 19261
rect 3510 19252 3516 19304
rect 3568 19292 3574 19304
rect 4356 19292 4384 19323
rect 8018 19320 8024 19332
rect 8076 19320 8082 19372
rect 8846 19320 8852 19372
rect 8904 19360 8910 19372
rect 10612 19369 10640 19400
rect 11057 19397 11069 19400
rect 11103 19428 11115 19431
rect 11606 19428 11612 19440
rect 11103 19400 11612 19428
rect 11103 19397 11115 19400
rect 11057 19391 11115 19397
rect 11606 19388 11612 19400
rect 11664 19388 11670 19440
rect 9033 19363 9091 19369
rect 9033 19360 9045 19363
rect 8904 19332 9045 19360
rect 8904 19320 8910 19332
rect 9033 19329 9045 19332
rect 9079 19329 9091 19363
rect 9033 19323 9091 19329
rect 10597 19363 10655 19369
rect 10597 19329 10609 19363
rect 10643 19329 10655 19363
rect 10597 19323 10655 19329
rect 12526 19320 12532 19372
rect 12584 19360 12590 19372
rect 12986 19360 12992 19372
rect 12584 19332 12848 19360
rect 12947 19332 12992 19360
rect 12584 19320 12590 19332
rect 7190 19292 7196 19304
rect 3568 19264 4384 19292
rect 7151 19264 7196 19292
rect 3568 19252 3574 19264
rect 7190 19252 7196 19264
rect 7248 19292 7254 19304
rect 7745 19295 7803 19301
rect 7745 19292 7757 19295
rect 7248 19264 7757 19292
rect 7248 19252 7254 19264
rect 7745 19261 7757 19264
rect 7791 19292 7803 19295
rect 7926 19292 7932 19304
rect 7791 19264 7932 19292
rect 7791 19261 7803 19264
rect 7745 19255 7803 19261
rect 7926 19252 7932 19264
rect 7984 19252 7990 19304
rect 8754 19252 8760 19304
rect 8812 19292 8818 19304
rect 8941 19295 8999 19301
rect 8941 19292 8953 19295
rect 8812 19264 8953 19292
rect 8812 19252 8818 19264
rect 8941 19261 8953 19264
rect 8987 19261 8999 19295
rect 10410 19292 10416 19304
rect 10323 19264 10416 19292
rect 8941 19255 8999 19261
rect 10410 19252 10416 19264
rect 10468 19292 10474 19304
rect 10870 19292 10876 19304
rect 10468 19264 10876 19292
rect 10468 19252 10474 19264
rect 10870 19252 10876 19264
rect 10928 19252 10934 19304
rect 12820 19301 12848 19332
rect 12986 19320 12992 19332
rect 13044 19320 13050 19372
rect 12805 19295 12863 19301
rect 12805 19261 12817 19295
rect 12851 19261 12863 19295
rect 12805 19255 12863 19261
rect 3329 19227 3387 19233
rect 3329 19193 3341 19227
rect 3375 19224 3387 19227
rect 5258 19224 5264 19236
rect 3375 19196 4200 19224
rect 5219 19196 5264 19224
rect 3375 19193 3387 19196
rect 3329 19187 3387 19193
rect 4172 19168 4200 19196
rect 5258 19184 5264 19196
rect 5316 19184 5322 19236
rect 8846 19224 8852 19236
rect 8807 19196 8852 19224
rect 8846 19184 8852 19196
rect 8904 19224 8910 19236
rect 9493 19227 9551 19233
rect 9493 19224 9505 19227
rect 8904 19196 9505 19224
rect 8904 19184 8910 19196
rect 9493 19193 9505 19196
rect 9539 19193 9551 19227
rect 12897 19227 12955 19233
rect 12897 19224 12909 19227
rect 9493 19187 9551 19193
rect 12176 19196 12909 19224
rect 2866 19156 2872 19168
rect 2827 19128 2872 19156
rect 2866 19116 2872 19128
rect 2924 19116 2930 19168
rect 3697 19159 3755 19165
rect 3697 19125 3709 19159
rect 3743 19156 3755 19159
rect 3970 19156 3976 19168
rect 3743 19128 3976 19156
rect 3743 19125 3755 19128
rect 3697 19119 3755 19125
rect 3970 19116 3976 19128
rect 4028 19116 4034 19168
rect 4154 19156 4160 19168
rect 4115 19128 4160 19156
rect 4154 19116 4160 19128
rect 4212 19116 4218 19168
rect 4798 19156 4804 19168
rect 4759 19128 4804 19156
rect 4798 19116 4804 19128
rect 4856 19116 4862 19168
rect 5350 19156 5356 19168
rect 5311 19128 5356 19156
rect 5350 19116 5356 19128
rect 5408 19116 5414 19168
rect 6086 19156 6092 19168
rect 6047 19128 6092 19156
rect 6086 19116 6092 19128
rect 6144 19116 6150 19168
rect 6641 19159 6699 19165
rect 6641 19125 6653 19159
rect 6687 19156 6699 19159
rect 6822 19156 6828 19168
rect 6687 19128 6828 19156
rect 6687 19125 6699 19128
rect 6641 19119 6699 19125
rect 6822 19116 6828 19128
rect 6880 19156 6886 19168
rect 7837 19159 7895 19165
rect 7837 19156 7849 19159
rect 6880 19128 7849 19156
rect 6880 19116 6886 19128
rect 7837 19125 7849 19128
rect 7883 19156 7895 19159
rect 8110 19156 8116 19168
rect 7883 19128 8116 19156
rect 7883 19125 7895 19128
rect 7837 19119 7895 19125
rect 8110 19116 8116 19128
rect 8168 19116 8174 19168
rect 8478 19156 8484 19168
rect 8439 19128 8484 19156
rect 8478 19116 8484 19128
rect 8536 19116 8542 19168
rect 10502 19156 10508 19168
rect 10463 19128 10508 19156
rect 10502 19116 10508 19128
rect 10560 19116 10566 19168
rect 11330 19116 11336 19168
rect 11388 19156 11394 19168
rect 11514 19156 11520 19168
rect 11388 19128 11520 19156
rect 11388 19116 11394 19128
rect 11514 19116 11520 19128
rect 11572 19156 11578 19168
rect 11793 19159 11851 19165
rect 11793 19156 11805 19159
rect 11572 19128 11805 19156
rect 11572 19116 11578 19128
rect 11793 19125 11805 19128
rect 11839 19125 11851 19159
rect 11793 19119 11851 19125
rect 11974 19116 11980 19168
rect 12032 19156 12038 19168
rect 12176 19165 12204 19196
rect 12897 19193 12909 19196
rect 12943 19193 12955 19227
rect 12897 19187 12955 19193
rect 12161 19159 12219 19165
rect 12161 19156 12173 19159
rect 12032 19128 12173 19156
rect 12032 19116 12038 19128
rect 12161 19125 12173 19128
rect 12207 19125 12219 19159
rect 12161 19119 12219 19125
rect 12434 19116 12440 19168
rect 12492 19156 12498 19168
rect 12492 19128 12537 19156
rect 12492 19116 12498 19128
rect 12618 19116 12624 19168
rect 12676 19156 12682 19168
rect 13449 19159 13507 19165
rect 13449 19156 13461 19159
rect 12676 19128 13461 19156
rect 12676 19116 12682 19128
rect 13449 19125 13461 19128
rect 13495 19125 13507 19159
rect 13449 19119 13507 19125
rect 1104 19066 14812 19088
rect 1104 19014 6315 19066
rect 6367 19014 6379 19066
rect 6431 19014 6443 19066
rect 6495 19014 6507 19066
rect 6559 19014 11648 19066
rect 11700 19014 11712 19066
rect 11764 19014 11776 19066
rect 11828 19014 11840 19066
rect 11892 19014 14812 19066
rect 1104 18992 14812 19014
rect 1394 18912 1400 18964
rect 1452 18952 1458 18964
rect 1581 18955 1639 18961
rect 1581 18952 1593 18955
rect 1452 18924 1593 18952
rect 1452 18912 1458 18924
rect 1581 18921 1593 18924
rect 1627 18921 1639 18955
rect 1581 18915 1639 18921
rect 2501 18955 2559 18961
rect 2501 18921 2513 18955
rect 2547 18952 2559 18955
rect 2774 18952 2780 18964
rect 2547 18924 2780 18952
rect 2547 18921 2559 18924
rect 2501 18915 2559 18921
rect 2774 18912 2780 18924
rect 2832 18912 2838 18964
rect 2866 18912 2872 18964
rect 2924 18952 2930 18964
rect 4065 18955 4123 18961
rect 4065 18952 4077 18955
rect 2924 18924 4077 18952
rect 2924 18912 2930 18924
rect 4065 18921 4077 18924
rect 4111 18921 4123 18955
rect 4065 18915 4123 18921
rect 5350 18912 5356 18964
rect 5408 18952 5414 18964
rect 5994 18952 6000 18964
rect 5408 18924 6000 18952
rect 5408 18912 5414 18924
rect 5994 18912 6000 18924
rect 6052 18912 6058 18964
rect 7101 18955 7159 18961
rect 7101 18921 7113 18955
rect 7147 18952 7159 18955
rect 8018 18952 8024 18964
rect 7147 18924 8024 18952
rect 7147 18921 7159 18924
rect 7101 18915 7159 18921
rect 8018 18912 8024 18924
rect 8076 18912 8082 18964
rect 8202 18912 8208 18964
rect 8260 18952 8266 18964
rect 9217 18955 9275 18961
rect 9217 18952 9229 18955
rect 8260 18924 9229 18952
rect 8260 18912 8266 18924
rect 9217 18921 9229 18924
rect 9263 18921 9275 18955
rect 9674 18952 9680 18964
rect 9635 18924 9680 18952
rect 9217 18915 9275 18921
rect 9674 18912 9680 18924
rect 9732 18912 9738 18964
rect 10134 18952 10140 18964
rect 10047 18924 10140 18952
rect 10134 18912 10140 18924
rect 10192 18952 10198 18964
rect 11241 18955 11299 18961
rect 11241 18952 11253 18955
rect 10192 18924 11253 18952
rect 10192 18912 10198 18924
rect 11241 18921 11253 18924
rect 11287 18921 11299 18955
rect 12986 18952 12992 18964
rect 12947 18924 12992 18952
rect 11241 18915 11299 18921
rect 12986 18912 12992 18924
rect 13044 18912 13050 18964
rect 3510 18844 3516 18896
rect 3568 18884 3574 18896
rect 3789 18887 3847 18893
rect 3789 18884 3801 18887
rect 3568 18856 3801 18884
rect 3568 18844 3574 18856
rect 3789 18853 3801 18856
rect 3835 18853 3847 18887
rect 3789 18847 3847 18853
rect 4433 18887 4491 18893
rect 4433 18853 4445 18887
rect 4479 18884 4491 18887
rect 4614 18884 4620 18896
rect 4479 18856 4620 18884
rect 4479 18853 4491 18856
rect 4433 18847 4491 18853
rect 3804 18816 3832 18847
rect 4614 18844 4620 18856
rect 4672 18844 4678 18896
rect 5534 18884 5540 18896
rect 5495 18856 5540 18884
rect 5534 18844 5540 18856
rect 5592 18844 5598 18896
rect 5626 18844 5632 18896
rect 5684 18884 5690 18896
rect 6089 18887 6147 18893
rect 6089 18884 6101 18887
rect 5684 18856 6101 18884
rect 5684 18844 5690 18856
rect 6089 18853 6101 18856
rect 6135 18853 6147 18887
rect 6089 18847 6147 18853
rect 10226 18844 10232 18896
rect 10284 18884 10290 18896
rect 10686 18884 10692 18896
rect 10284 18856 10692 18884
rect 10284 18844 10290 18856
rect 10686 18844 10692 18856
rect 10744 18844 10750 18896
rect 12066 18884 12072 18896
rect 11624 18856 12072 18884
rect 7193 18819 7251 18825
rect 3804 18788 4660 18816
rect 4338 18708 4344 18760
rect 4396 18748 4402 18760
rect 4632 18757 4660 18788
rect 7193 18785 7205 18819
rect 7239 18816 7251 18819
rect 7374 18816 7380 18828
rect 7239 18788 7380 18816
rect 7239 18785 7251 18788
rect 7193 18779 7251 18785
rect 7374 18776 7380 18788
rect 7432 18776 7438 18828
rect 9858 18776 9864 18828
rect 9916 18816 9922 18828
rect 10042 18816 10048 18828
rect 9916 18788 10048 18816
rect 9916 18776 9922 18788
rect 10042 18776 10048 18788
rect 10100 18776 10106 18828
rect 10594 18776 10600 18828
rect 10652 18816 10658 18828
rect 10870 18816 10876 18828
rect 10652 18788 10876 18816
rect 10652 18776 10658 18788
rect 10870 18776 10876 18788
rect 10928 18776 10934 18828
rect 11330 18776 11336 18828
rect 11388 18816 11394 18828
rect 11624 18825 11652 18856
rect 12066 18844 12072 18856
rect 12124 18844 12130 18896
rect 12713 18887 12771 18893
rect 12713 18853 12725 18887
rect 12759 18884 12771 18887
rect 13078 18884 13084 18896
rect 12759 18856 13084 18884
rect 12759 18853 12771 18856
rect 12713 18847 12771 18853
rect 13078 18844 13084 18856
rect 13136 18844 13142 18896
rect 11609 18819 11667 18825
rect 11609 18816 11621 18819
rect 11388 18788 11621 18816
rect 11388 18776 11394 18788
rect 11609 18785 11621 18788
rect 11655 18785 11667 18819
rect 11609 18779 11667 18785
rect 4525 18751 4583 18757
rect 4525 18748 4537 18751
rect 4396 18720 4537 18748
rect 4396 18708 4402 18720
rect 4525 18717 4537 18720
rect 4571 18717 4583 18751
rect 4525 18711 4583 18717
rect 4617 18751 4675 18757
rect 4617 18717 4629 18751
rect 4663 18748 4675 18751
rect 4706 18748 4712 18760
rect 4663 18720 4712 18748
rect 4663 18717 4675 18720
rect 4617 18711 4675 18717
rect 4706 18708 4712 18720
rect 4764 18708 4770 18760
rect 6273 18751 6331 18757
rect 6273 18717 6285 18751
rect 6319 18748 6331 18751
rect 6822 18748 6828 18760
rect 6319 18720 6828 18748
rect 6319 18717 6331 18720
rect 6273 18711 6331 18717
rect 6822 18708 6828 18720
rect 6880 18708 6886 18760
rect 9306 18708 9312 18760
rect 9364 18748 9370 18760
rect 10229 18751 10287 18757
rect 10229 18748 10241 18751
rect 9364 18720 10241 18748
rect 9364 18708 9370 18720
rect 10229 18717 10241 18720
rect 10275 18717 10287 18751
rect 11698 18748 11704 18760
rect 11659 18720 11704 18748
rect 10229 18711 10287 18717
rect 11698 18708 11704 18720
rect 11756 18708 11762 18760
rect 11793 18751 11851 18757
rect 11793 18717 11805 18751
rect 11839 18748 11851 18751
rect 12066 18748 12072 18760
rect 11839 18720 12072 18748
rect 11839 18717 11851 18720
rect 11793 18711 11851 18717
rect 4154 18640 4160 18692
rect 4212 18680 4218 18692
rect 5629 18683 5687 18689
rect 5629 18680 5641 18683
rect 4212 18652 5641 18680
rect 4212 18640 4218 18652
rect 5629 18649 5641 18652
rect 5675 18649 5687 18683
rect 5629 18643 5687 18649
rect 8386 18640 8392 18692
rect 8444 18680 8450 18692
rect 8481 18683 8539 18689
rect 8481 18680 8493 18683
rect 8444 18652 8493 18680
rect 8444 18640 8450 18652
rect 8481 18649 8493 18652
rect 8527 18649 8539 18683
rect 8481 18643 8539 18649
rect 10594 18640 10600 18692
rect 10652 18680 10658 18692
rect 11057 18683 11115 18689
rect 11057 18680 11069 18683
rect 10652 18652 11069 18680
rect 10652 18640 10658 18652
rect 11057 18649 11069 18652
rect 11103 18649 11115 18683
rect 11057 18643 11115 18649
rect 11238 18640 11244 18692
rect 11296 18680 11302 18692
rect 11808 18680 11836 18711
rect 12066 18708 12072 18720
rect 12124 18748 12130 18760
rect 12986 18748 12992 18760
rect 12124 18720 12992 18748
rect 12124 18708 12130 18720
rect 12986 18708 12992 18720
rect 13044 18708 13050 18760
rect 11296 18652 11836 18680
rect 11296 18640 11302 18652
rect 3234 18612 3240 18624
rect 3195 18584 3240 18612
rect 3234 18572 3240 18584
rect 3292 18572 3298 18624
rect 6730 18612 6736 18624
rect 6691 18584 6736 18612
rect 6730 18572 6736 18584
rect 6788 18572 6794 18624
rect 10686 18612 10692 18624
rect 10647 18584 10692 18612
rect 10686 18572 10692 18584
rect 10744 18572 10750 18624
rect 1104 18522 14812 18544
rect 1104 18470 3648 18522
rect 3700 18470 3712 18522
rect 3764 18470 3776 18522
rect 3828 18470 3840 18522
rect 3892 18470 8982 18522
rect 9034 18470 9046 18522
rect 9098 18470 9110 18522
rect 9162 18470 9174 18522
rect 9226 18470 14315 18522
rect 14367 18470 14379 18522
rect 14431 18470 14443 18522
rect 14495 18470 14507 18522
rect 14559 18470 14812 18522
rect 1104 18448 14812 18470
rect 4525 18411 4583 18417
rect 4525 18377 4537 18411
rect 4571 18408 4583 18411
rect 4706 18408 4712 18420
rect 4571 18380 4712 18408
rect 4571 18377 4583 18380
rect 4525 18371 4583 18377
rect 4706 18368 4712 18380
rect 4764 18408 4770 18420
rect 4801 18411 4859 18417
rect 4801 18408 4813 18411
rect 4764 18380 4813 18408
rect 4764 18368 4770 18380
rect 4801 18377 4813 18380
rect 4847 18377 4859 18411
rect 5626 18408 5632 18420
rect 5587 18380 5632 18408
rect 4801 18371 4859 18377
rect 5626 18368 5632 18380
rect 5684 18368 5690 18420
rect 5994 18408 6000 18420
rect 5955 18380 6000 18408
rect 5994 18368 6000 18380
rect 6052 18368 6058 18420
rect 6641 18411 6699 18417
rect 6641 18377 6653 18411
rect 6687 18408 6699 18411
rect 6730 18408 6736 18420
rect 6687 18380 6736 18408
rect 6687 18377 6699 18380
rect 6641 18371 6699 18377
rect 6730 18368 6736 18380
rect 6788 18408 6794 18420
rect 8294 18408 8300 18420
rect 6788 18380 8300 18408
rect 6788 18368 6794 18380
rect 6840 18272 6868 18380
rect 8294 18368 8300 18380
rect 8352 18408 8358 18420
rect 8481 18411 8539 18417
rect 8481 18408 8493 18411
rect 8352 18380 8493 18408
rect 8352 18368 8358 18380
rect 8481 18377 8493 18380
rect 8527 18377 8539 18411
rect 8481 18371 8539 18377
rect 9033 18411 9091 18417
rect 9033 18377 9045 18411
rect 9079 18408 9091 18411
rect 10134 18408 10140 18420
rect 9079 18380 10140 18408
rect 9079 18377 9091 18380
rect 9033 18371 9091 18377
rect 10134 18368 10140 18380
rect 10192 18368 10198 18420
rect 11425 18411 11483 18417
rect 11425 18377 11437 18411
rect 11471 18408 11483 18411
rect 11698 18408 11704 18420
rect 11471 18380 11704 18408
rect 11471 18377 11483 18380
rect 11425 18371 11483 18377
rect 11698 18368 11704 18380
rect 11756 18368 11762 18420
rect 12066 18408 12072 18420
rect 12027 18380 12072 18408
rect 12066 18368 12072 18380
rect 12124 18368 12130 18420
rect 8018 18300 8024 18352
rect 8076 18340 8082 18352
rect 8570 18340 8576 18352
rect 8076 18312 8576 18340
rect 8076 18300 8082 18312
rect 8570 18300 8576 18312
rect 8628 18340 8634 18352
rect 9306 18340 9312 18352
rect 8628 18312 9312 18340
rect 8628 18300 8634 18312
rect 9306 18300 9312 18312
rect 9364 18300 9370 18352
rect 6840 18244 6960 18272
rect 3145 18207 3203 18213
rect 3145 18173 3157 18207
rect 3191 18204 3203 18207
rect 3234 18204 3240 18216
rect 3191 18176 3240 18204
rect 3191 18173 3203 18176
rect 3145 18167 3203 18173
rect 3234 18164 3240 18176
rect 3292 18204 3298 18216
rect 3292 18176 4108 18204
rect 3292 18164 3298 18176
rect 4080 18148 4108 18176
rect 6730 18164 6736 18216
rect 6788 18204 6794 18216
rect 6825 18207 6883 18213
rect 6825 18204 6837 18207
rect 6788 18176 6837 18204
rect 6788 18164 6794 18176
rect 6825 18173 6837 18176
rect 6871 18173 6883 18207
rect 6932 18204 6960 18244
rect 10594 18232 10600 18284
rect 10652 18272 10658 18284
rect 10873 18275 10931 18281
rect 10873 18272 10885 18275
rect 10652 18244 10885 18272
rect 10652 18232 10658 18244
rect 10873 18241 10885 18244
rect 10919 18241 10931 18275
rect 10873 18235 10931 18241
rect 7081 18207 7139 18213
rect 7081 18204 7093 18207
rect 6932 18176 7093 18204
rect 6825 18167 6883 18173
rect 7081 18173 7093 18176
rect 7127 18173 7139 18207
rect 7081 18167 7139 18173
rect 9766 18164 9772 18216
rect 9824 18204 9830 18216
rect 10137 18207 10195 18213
rect 10137 18204 10149 18207
rect 9824 18176 10149 18204
rect 9824 18164 9830 18176
rect 10137 18173 10149 18176
rect 10183 18204 10195 18207
rect 10318 18204 10324 18216
rect 10183 18176 10324 18204
rect 10183 18173 10195 18176
rect 10137 18167 10195 18173
rect 10318 18164 10324 18176
rect 10376 18204 10382 18216
rect 10781 18207 10839 18213
rect 10781 18204 10793 18207
rect 10376 18176 10793 18204
rect 10376 18164 10382 18176
rect 10781 18173 10793 18176
rect 10827 18173 10839 18207
rect 10781 18167 10839 18173
rect 3053 18139 3111 18145
rect 3053 18105 3065 18139
rect 3099 18136 3111 18139
rect 3412 18139 3470 18145
rect 3412 18136 3424 18139
rect 3099 18108 3424 18136
rect 3099 18105 3111 18108
rect 3053 18099 3111 18105
rect 3412 18105 3424 18108
rect 3458 18136 3470 18139
rect 3458 18108 3832 18136
rect 3458 18105 3470 18108
rect 3412 18099 3470 18105
rect 3804 18080 3832 18108
rect 4062 18096 4068 18148
rect 4120 18096 4126 18148
rect 10226 18096 10232 18148
rect 10284 18136 10290 18148
rect 10686 18136 10692 18148
rect 10284 18108 10692 18136
rect 10284 18096 10290 18108
rect 10686 18096 10692 18108
rect 10744 18096 10750 18148
rect 3786 18028 3792 18080
rect 3844 18068 3850 18080
rect 3970 18068 3976 18080
rect 3844 18040 3976 18068
rect 3844 18028 3850 18040
rect 3970 18028 3976 18040
rect 4028 18068 4034 18080
rect 5166 18068 5172 18080
rect 4028 18040 5172 18068
rect 4028 18028 4034 18040
rect 5166 18028 5172 18040
rect 5224 18068 5230 18080
rect 5353 18071 5411 18077
rect 5353 18068 5365 18071
rect 5224 18040 5365 18068
rect 5224 18028 5230 18040
rect 5353 18037 5365 18040
rect 5399 18068 5411 18071
rect 5534 18068 5540 18080
rect 5399 18040 5540 18068
rect 5399 18037 5411 18040
rect 5353 18031 5411 18037
rect 5534 18028 5540 18040
rect 5592 18028 5598 18080
rect 6086 18028 6092 18080
rect 6144 18068 6150 18080
rect 8205 18071 8263 18077
rect 8205 18068 8217 18071
rect 6144 18040 8217 18068
rect 6144 18028 6150 18040
rect 8205 18037 8217 18040
rect 8251 18037 8263 18071
rect 8205 18031 8263 18037
rect 9769 18071 9827 18077
rect 9769 18037 9781 18071
rect 9815 18068 9827 18071
rect 9858 18068 9864 18080
rect 9815 18040 9864 18068
rect 9815 18037 9827 18040
rect 9769 18031 9827 18037
rect 9858 18028 9864 18040
rect 9916 18028 9922 18080
rect 10318 18068 10324 18080
rect 10279 18040 10324 18068
rect 10318 18028 10324 18040
rect 10376 18028 10382 18080
rect 11330 18028 11336 18080
rect 11388 18068 11394 18080
rect 11701 18071 11759 18077
rect 11701 18068 11713 18071
rect 11388 18040 11713 18068
rect 11388 18028 11394 18040
rect 11701 18037 11713 18040
rect 11747 18037 11759 18071
rect 11701 18031 11759 18037
rect 1104 17978 14812 18000
rect 1104 17926 6315 17978
rect 6367 17926 6379 17978
rect 6431 17926 6443 17978
rect 6495 17926 6507 17978
rect 6559 17926 11648 17978
rect 11700 17926 11712 17978
rect 11764 17926 11776 17978
rect 11828 17926 11840 17978
rect 11892 17926 14812 17978
rect 1104 17904 14812 17926
rect 2409 17867 2467 17873
rect 2409 17833 2421 17867
rect 2455 17864 2467 17867
rect 4338 17864 4344 17876
rect 2455 17836 4344 17864
rect 2455 17833 2467 17836
rect 2409 17827 2467 17833
rect 4338 17824 4344 17836
rect 4396 17824 4402 17876
rect 4614 17864 4620 17876
rect 4575 17836 4620 17864
rect 4614 17824 4620 17836
rect 4672 17824 4678 17876
rect 5534 17824 5540 17876
rect 5592 17864 5598 17876
rect 6365 17867 6423 17873
rect 6365 17864 6377 17867
rect 5592 17836 6377 17864
rect 5592 17824 5598 17836
rect 6365 17833 6377 17836
rect 6411 17864 6423 17867
rect 6822 17864 6828 17876
rect 6411 17836 6828 17864
rect 6411 17833 6423 17836
rect 6365 17827 6423 17833
rect 6822 17824 6828 17836
rect 6880 17824 6886 17876
rect 7834 17864 7840 17876
rect 7795 17836 7840 17864
rect 7834 17824 7840 17836
rect 7892 17824 7898 17876
rect 8478 17864 8484 17876
rect 8439 17836 8484 17864
rect 8478 17824 8484 17836
rect 8536 17824 8542 17876
rect 10318 17824 10324 17876
rect 10376 17864 10382 17876
rect 10778 17864 10784 17876
rect 10376 17836 10784 17864
rect 10376 17824 10382 17836
rect 10778 17824 10784 17836
rect 10836 17864 10842 17876
rect 10873 17867 10931 17873
rect 10873 17864 10885 17867
rect 10836 17836 10885 17864
rect 10836 17824 10842 17836
rect 10873 17833 10885 17836
rect 10919 17833 10931 17867
rect 10873 17827 10931 17833
rect 3786 17796 3792 17808
rect 3747 17768 3792 17796
rect 3786 17756 3792 17768
rect 3844 17756 3850 17808
rect 8386 17796 8392 17808
rect 8347 17768 8392 17796
rect 8386 17756 8392 17768
rect 8444 17756 8450 17808
rect 2774 17688 2780 17740
rect 2832 17728 2838 17740
rect 2832 17700 2877 17728
rect 2832 17688 2838 17700
rect 2866 17660 2872 17672
rect 2827 17632 2872 17660
rect 2866 17620 2872 17632
rect 2924 17620 2930 17672
rect 3053 17663 3111 17669
rect 3053 17629 3065 17663
rect 3099 17660 3111 17663
rect 3804 17660 3832 17756
rect 5074 17688 5080 17740
rect 5132 17728 5138 17740
rect 5241 17731 5299 17737
rect 5241 17728 5253 17731
rect 5132 17700 5253 17728
rect 5132 17688 5138 17700
rect 5241 17697 5253 17700
rect 5287 17697 5299 17731
rect 5241 17691 5299 17697
rect 10781 17731 10839 17737
rect 10781 17697 10793 17731
rect 10827 17728 10839 17731
rect 10870 17728 10876 17740
rect 10827 17700 10876 17728
rect 10827 17697 10839 17700
rect 10781 17691 10839 17697
rect 10870 17688 10876 17700
rect 10928 17688 10934 17740
rect 3099 17632 3832 17660
rect 3099 17629 3111 17632
rect 3053 17623 3111 17629
rect 4062 17620 4068 17672
rect 4120 17660 4126 17672
rect 4982 17660 4988 17672
rect 4120 17632 4988 17660
rect 4120 17620 4126 17632
rect 4982 17620 4988 17632
rect 5040 17620 5046 17672
rect 8570 17660 8576 17672
rect 8531 17632 8576 17660
rect 8570 17620 8576 17632
rect 8628 17620 8634 17672
rect 10318 17620 10324 17672
rect 10376 17660 10382 17672
rect 10965 17663 11023 17669
rect 10965 17660 10977 17663
rect 10376 17632 10977 17660
rect 10376 17620 10382 17632
rect 10965 17629 10977 17632
rect 11011 17660 11023 17663
rect 11514 17660 11520 17672
rect 11011 17632 11520 17660
rect 11011 17629 11023 17632
rect 10965 17623 11023 17629
rect 11514 17620 11520 17632
rect 11572 17620 11578 17672
rect 7466 17552 7472 17604
rect 7524 17592 7530 17604
rect 8021 17595 8079 17601
rect 8021 17592 8033 17595
rect 7524 17564 8033 17592
rect 7524 17552 7530 17564
rect 8021 17561 8033 17564
rect 8067 17561 8079 17595
rect 10410 17592 10416 17604
rect 10371 17564 10416 17592
rect 8021 17555 8079 17561
rect 10410 17552 10416 17564
rect 10468 17552 10474 17604
rect 4982 17484 4988 17536
rect 5040 17524 5046 17536
rect 6730 17524 6736 17536
rect 5040 17496 6736 17524
rect 5040 17484 5046 17496
rect 6730 17484 6736 17496
rect 6788 17524 6794 17536
rect 6825 17527 6883 17533
rect 6825 17524 6837 17527
rect 6788 17496 6837 17524
rect 6788 17484 6794 17496
rect 6825 17493 6837 17496
rect 6871 17493 6883 17527
rect 6825 17487 6883 17493
rect 7285 17527 7343 17533
rect 7285 17493 7297 17527
rect 7331 17524 7343 17527
rect 7374 17524 7380 17536
rect 7331 17496 7380 17524
rect 7331 17493 7343 17496
rect 7285 17487 7343 17493
rect 7374 17484 7380 17496
rect 7432 17484 7438 17536
rect 10045 17527 10103 17533
rect 10045 17493 10057 17527
rect 10091 17524 10103 17527
rect 10594 17524 10600 17536
rect 10091 17496 10600 17524
rect 10091 17493 10103 17496
rect 10045 17487 10103 17493
rect 10594 17484 10600 17496
rect 10652 17484 10658 17536
rect 1104 17434 14812 17456
rect 1104 17382 3648 17434
rect 3700 17382 3712 17434
rect 3764 17382 3776 17434
rect 3828 17382 3840 17434
rect 3892 17382 8982 17434
rect 9034 17382 9046 17434
rect 9098 17382 9110 17434
rect 9162 17382 9174 17434
rect 9226 17382 14315 17434
rect 14367 17382 14379 17434
rect 14431 17382 14443 17434
rect 14495 17382 14507 17434
rect 14559 17382 14812 17434
rect 1104 17360 14812 17382
rect 2501 17323 2559 17329
rect 2501 17289 2513 17323
rect 2547 17320 2559 17323
rect 2774 17320 2780 17332
rect 2547 17292 2780 17320
rect 2547 17289 2559 17292
rect 2501 17283 2559 17289
rect 2774 17280 2780 17292
rect 2832 17280 2838 17332
rect 3697 17323 3755 17329
rect 3697 17289 3709 17323
rect 3743 17320 3755 17323
rect 4614 17320 4620 17332
rect 3743 17292 4620 17320
rect 3743 17289 3755 17292
rect 3697 17283 3755 17289
rect 4614 17280 4620 17292
rect 4672 17280 4678 17332
rect 7282 17280 7288 17332
rect 7340 17320 7346 17332
rect 7377 17323 7435 17329
rect 7377 17320 7389 17323
rect 7340 17292 7389 17320
rect 7340 17280 7346 17292
rect 7377 17289 7389 17292
rect 7423 17289 7435 17323
rect 8478 17320 8484 17332
rect 8439 17292 8484 17320
rect 7377 17283 7435 17289
rect 5626 17212 5632 17264
rect 5684 17252 5690 17264
rect 5810 17252 5816 17264
rect 5684 17224 5816 17252
rect 5684 17212 5690 17224
rect 5810 17212 5816 17224
rect 5868 17212 5874 17264
rect 2777 17187 2835 17193
rect 2777 17153 2789 17187
rect 2823 17184 2835 17187
rect 3970 17184 3976 17196
rect 2823 17156 3976 17184
rect 2823 17153 2835 17156
rect 2777 17147 2835 17153
rect 3970 17144 3976 17156
rect 4028 17184 4034 17196
rect 4249 17187 4307 17193
rect 4249 17184 4261 17187
rect 4028 17156 4261 17184
rect 4028 17144 4034 17156
rect 4249 17153 4261 17156
rect 4295 17153 4307 17187
rect 4249 17147 4307 17153
rect 2866 17076 2872 17128
rect 2924 17116 2930 17128
rect 3237 17119 3295 17125
rect 3237 17116 3249 17119
rect 2924 17088 3249 17116
rect 2924 17076 2930 17088
rect 3237 17085 3249 17088
rect 3283 17116 3295 17119
rect 4154 17116 4160 17128
rect 3283 17088 4160 17116
rect 3283 17085 3295 17088
rect 3237 17079 3295 17085
rect 4154 17076 4160 17088
rect 4212 17076 4218 17128
rect 7392 17116 7420 17283
rect 8478 17280 8484 17292
rect 8536 17280 8542 17332
rect 10870 17280 10876 17332
rect 10928 17320 10934 17332
rect 10965 17323 11023 17329
rect 10965 17320 10977 17323
rect 10928 17292 10977 17320
rect 10928 17280 10934 17292
rect 10965 17289 10977 17292
rect 11011 17320 11023 17323
rect 12342 17320 12348 17332
rect 11011 17292 12348 17320
rect 11011 17289 11023 17292
rect 10965 17283 11023 17289
rect 12342 17280 12348 17292
rect 12400 17280 12406 17332
rect 8386 17212 8392 17264
rect 8444 17252 8450 17264
rect 8757 17255 8815 17261
rect 8757 17252 8769 17255
rect 8444 17224 8769 17252
rect 8444 17212 8450 17224
rect 8757 17221 8769 17224
rect 8803 17221 8815 17255
rect 8757 17215 8815 17221
rect 8113 17187 8171 17193
rect 8113 17153 8125 17187
rect 8159 17184 8171 17187
rect 8570 17184 8576 17196
rect 8159 17156 8576 17184
rect 8159 17153 8171 17156
rect 8113 17147 8171 17153
rect 8570 17144 8576 17156
rect 8628 17144 8634 17196
rect 10594 17184 10600 17196
rect 10555 17156 10600 17184
rect 10594 17144 10600 17156
rect 10652 17144 10658 17196
rect 7745 17119 7803 17125
rect 7745 17116 7757 17119
rect 7392 17088 7757 17116
rect 7745 17085 7757 17088
rect 7791 17085 7803 17119
rect 7745 17079 7803 17085
rect 3605 17051 3663 17057
rect 3605 17017 3617 17051
rect 3651 17048 3663 17051
rect 4065 17051 4123 17057
rect 4065 17048 4077 17051
rect 3651 17020 4077 17048
rect 3651 17017 3663 17020
rect 3605 17011 3663 17017
rect 4065 17017 4077 17020
rect 4111 17048 4123 17051
rect 4246 17048 4252 17060
rect 4111 17020 4252 17048
rect 4111 17017 4123 17020
rect 4065 17011 4123 17017
rect 4246 17008 4252 17020
rect 4304 17008 4310 17060
rect 4982 17008 4988 17060
rect 5040 17048 5046 17060
rect 10413 17051 10471 17057
rect 10413 17048 10425 17051
rect 5040 17020 5488 17048
rect 5040 17008 5046 17020
rect 3970 16940 3976 16992
rect 4028 16980 4034 16992
rect 4157 16983 4215 16989
rect 4157 16980 4169 16983
rect 4028 16952 4169 16980
rect 4028 16940 4034 16952
rect 4157 16949 4169 16952
rect 4203 16949 4215 16983
rect 5074 16980 5080 16992
rect 5035 16952 5080 16980
rect 4157 16943 4215 16949
rect 5074 16940 5080 16952
rect 5132 16940 5138 16992
rect 5460 16989 5488 17020
rect 9784 17020 10425 17048
rect 5445 16983 5503 16989
rect 5445 16949 5457 16983
rect 5491 16980 5503 16983
rect 5718 16980 5724 16992
rect 5491 16952 5724 16980
rect 5491 16949 5503 16952
rect 5445 16943 5503 16949
rect 5718 16940 5724 16952
rect 5776 16940 5782 16992
rect 7558 16980 7564 16992
rect 7519 16952 7564 16980
rect 7558 16940 7564 16952
rect 7616 16940 7622 16992
rect 9674 16940 9680 16992
rect 9732 16980 9738 16992
rect 9784 16989 9812 17020
rect 10413 17017 10425 17020
rect 10459 17017 10471 17051
rect 10413 17011 10471 17017
rect 9769 16983 9827 16989
rect 9769 16980 9781 16983
rect 9732 16952 9781 16980
rect 9732 16940 9738 16952
rect 9769 16949 9781 16952
rect 9815 16949 9827 16983
rect 9950 16980 9956 16992
rect 9911 16952 9956 16980
rect 9769 16943 9827 16949
rect 9950 16940 9956 16952
rect 10008 16940 10014 16992
rect 10042 16940 10048 16992
rect 10100 16980 10106 16992
rect 10321 16983 10379 16989
rect 10321 16980 10333 16983
rect 10100 16952 10333 16980
rect 10100 16940 10106 16952
rect 10321 16949 10333 16952
rect 10367 16949 10379 16983
rect 10321 16943 10379 16949
rect 1104 16890 14812 16912
rect 1104 16838 6315 16890
rect 6367 16838 6379 16890
rect 6431 16838 6443 16890
rect 6495 16838 6507 16890
rect 6559 16838 11648 16890
rect 11700 16838 11712 16890
rect 11764 16838 11776 16890
rect 11828 16838 11840 16890
rect 11892 16838 14812 16890
rect 1104 16816 14812 16838
rect 3789 16779 3847 16785
rect 3789 16745 3801 16779
rect 3835 16776 3847 16779
rect 3970 16776 3976 16788
rect 3835 16748 3976 16776
rect 3835 16745 3847 16748
rect 3789 16739 3847 16745
rect 3970 16736 3976 16748
rect 4028 16736 4034 16788
rect 5074 16776 5080 16788
rect 4987 16748 5080 16776
rect 5074 16736 5080 16748
rect 5132 16776 5138 16788
rect 7009 16779 7067 16785
rect 7009 16776 7021 16779
rect 5132 16748 7021 16776
rect 5132 16736 5138 16748
rect 7009 16745 7021 16748
rect 7055 16745 7067 16779
rect 10042 16776 10048 16788
rect 10003 16748 10048 16776
rect 7009 16739 7067 16745
rect 10042 16736 10048 16748
rect 10100 16736 10106 16788
rect 10778 16776 10784 16788
rect 10739 16748 10784 16776
rect 10778 16736 10784 16748
rect 10836 16736 10842 16788
rect 12345 16779 12403 16785
rect 12345 16745 12357 16779
rect 12391 16745 12403 16779
rect 12345 16739 12403 16745
rect 6086 16708 6092 16720
rect 5920 16680 6092 16708
rect 5920 16652 5948 16680
rect 6086 16668 6092 16680
rect 6144 16668 6150 16720
rect 10318 16668 10324 16720
rect 10376 16708 10382 16720
rect 12360 16708 12388 16739
rect 12434 16736 12440 16788
rect 12492 16776 12498 16788
rect 12618 16776 12624 16788
rect 12492 16748 12624 16776
rect 12492 16736 12498 16748
rect 12618 16736 12624 16748
rect 12676 16736 12682 16788
rect 10376 16680 12388 16708
rect 10376 16668 10382 16680
rect 5442 16640 5448 16652
rect 5403 16612 5448 16640
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 5629 16643 5687 16649
rect 5629 16609 5641 16643
rect 5675 16640 5687 16643
rect 5718 16640 5724 16652
rect 5675 16612 5724 16640
rect 5675 16609 5687 16612
rect 5629 16603 5687 16609
rect 5261 16507 5319 16513
rect 5261 16473 5273 16507
rect 5307 16504 5319 16507
rect 5644 16504 5672 16603
rect 5718 16600 5724 16612
rect 5776 16600 5782 16652
rect 5902 16649 5908 16652
rect 5896 16640 5908 16649
rect 5863 16612 5908 16640
rect 5896 16603 5908 16612
rect 5902 16600 5908 16603
rect 5960 16600 5966 16652
rect 7650 16600 7656 16652
rect 7708 16640 7714 16652
rect 8202 16640 8208 16652
rect 7708 16612 8064 16640
rect 8163 16612 8208 16640
rect 7708 16600 7714 16612
rect 8036 16572 8064 16612
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 10594 16600 10600 16652
rect 10652 16640 10658 16652
rect 11221 16643 11279 16649
rect 11221 16640 11233 16643
rect 10652 16612 11233 16640
rect 10652 16600 10658 16612
rect 11221 16609 11233 16612
rect 11267 16609 11279 16643
rect 11221 16603 11279 16609
rect 8294 16572 8300 16584
rect 8036 16544 8300 16572
rect 8294 16532 8300 16544
rect 8352 16532 8358 16584
rect 8386 16532 8392 16584
rect 8444 16572 8450 16584
rect 10965 16575 11023 16581
rect 8444 16544 8489 16572
rect 8444 16532 8450 16544
rect 10965 16541 10977 16575
rect 11011 16541 11023 16575
rect 10965 16535 11023 16541
rect 5307 16476 5672 16504
rect 5307 16473 5319 16476
rect 5261 16467 5319 16473
rect 7006 16464 7012 16516
rect 7064 16504 7070 16516
rect 7377 16507 7435 16513
rect 7377 16504 7389 16507
rect 7064 16476 7389 16504
rect 7064 16464 7070 16476
rect 7377 16473 7389 16476
rect 7423 16504 7435 16507
rect 9306 16504 9312 16516
rect 7423 16476 9312 16504
rect 7423 16473 7435 16476
rect 7377 16467 7435 16473
rect 9306 16464 9312 16476
rect 9364 16464 9370 16516
rect 7834 16436 7840 16448
rect 7795 16408 7840 16436
rect 7834 16396 7840 16408
rect 7892 16396 7898 16448
rect 10318 16396 10324 16448
rect 10376 16436 10382 16448
rect 10413 16439 10471 16445
rect 10413 16436 10425 16439
rect 10376 16408 10425 16436
rect 10376 16396 10382 16408
rect 10413 16405 10425 16408
rect 10459 16405 10471 16439
rect 10980 16436 11008 16535
rect 11330 16436 11336 16448
rect 10980 16408 11336 16436
rect 10413 16399 10471 16405
rect 11330 16396 11336 16408
rect 11388 16396 11394 16448
rect 1104 16346 14812 16368
rect 1104 16294 3648 16346
rect 3700 16294 3712 16346
rect 3764 16294 3776 16346
rect 3828 16294 3840 16346
rect 3892 16294 8982 16346
rect 9034 16294 9046 16346
rect 9098 16294 9110 16346
rect 9162 16294 9174 16346
rect 9226 16294 14315 16346
rect 14367 16294 14379 16346
rect 14431 16294 14443 16346
rect 14495 16294 14507 16346
rect 14559 16294 14812 16346
rect 1104 16272 14812 16294
rect 4154 16192 4160 16244
rect 4212 16232 4218 16244
rect 4985 16235 5043 16241
rect 4985 16232 4997 16235
rect 4212 16204 4997 16232
rect 4212 16192 4218 16204
rect 4985 16201 4997 16204
rect 5031 16201 5043 16235
rect 4985 16195 5043 16201
rect 5902 16192 5908 16244
rect 5960 16232 5966 16244
rect 5997 16235 6055 16241
rect 5997 16232 6009 16235
rect 5960 16204 6009 16232
rect 5960 16192 5966 16204
rect 5997 16201 6009 16204
rect 6043 16201 6055 16235
rect 11330 16232 11336 16244
rect 11291 16204 11336 16232
rect 5997 16195 6055 16201
rect 11330 16192 11336 16204
rect 11388 16192 11394 16244
rect 1578 16096 1584 16108
rect 1539 16068 1584 16096
rect 1578 16056 1584 16068
rect 1636 16056 1642 16108
rect 5074 16056 5080 16108
rect 5132 16096 5138 16108
rect 5537 16099 5595 16105
rect 5537 16096 5549 16099
rect 5132 16068 5549 16096
rect 5132 16056 5138 16068
rect 5537 16065 5549 16068
rect 5583 16065 5595 16099
rect 7006 16096 7012 16108
rect 6967 16068 7012 16096
rect 5537 16059 5595 16065
rect 7006 16056 7012 16068
rect 7064 16056 7070 16108
rect 9214 16096 9220 16108
rect 9175 16068 9220 16096
rect 9214 16056 9220 16068
rect 9272 16056 9278 16108
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 4893 16031 4951 16037
rect 1443 16000 2268 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 2240 15904 2268 16000
rect 4893 15997 4905 16031
rect 4939 16028 4951 16031
rect 5445 16031 5503 16037
rect 5445 16028 5457 16031
rect 4939 16000 5457 16028
rect 4939 15997 4951 16000
rect 4893 15991 4951 15997
rect 5445 15997 5457 16000
rect 5491 16028 5503 16031
rect 9306 16028 9312 16040
rect 5491 16000 9312 16028
rect 5491 15997 5503 16000
rect 5445 15991 5503 15997
rect 9306 15988 9312 16000
rect 9364 15988 9370 16040
rect 6641 15963 6699 15969
rect 6641 15929 6653 15963
rect 6687 15960 6699 15963
rect 7254 15963 7312 15969
rect 7254 15960 7266 15963
rect 6687 15932 7266 15960
rect 6687 15929 6699 15932
rect 6641 15923 6699 15929
rect 7254 15929 7266 15932
rect 7300 15960 7312 15963
rect 7650 15960 7656 15972
rect 7300 15932 7656 15960
rect 7300 15929 7312 15932
rect 7254 15923 7312 15929
rect 7650 15920 7656 15932
rect 7708 15920 7714 15972
rect 9033 15963 9091 15969
rect 9033 15960 9045 15963
rect 8404 15932 9045 15960
rect 2222 15892 2228 15904
rect 2183 15864 2228 15892
rect 2222 15852 2228 15864
rect 2280 15852 2286 15904
rect 5074 15852 5080 15904
rect 5132 15892 5138 15904
rect 5353 15895 5411 15901
rect 5353 15892 5365 15895
rect 5132 15864 5365 15892
rect 5132 15852 5138 15864
rect 5353 15861 5365 15864
rect 5399 15861 5411 15895
rect 5353 15855 5411 15861
rect 7098 15852 7104 15904
rect 7156 15892 7162 15904
rect 8404 15901 8432 15932
rect 9033 15929 9045 15932
rect 9079 15960 9091 15963
rect 9462 15963 9520 15969
rect 9462 15960 9474 15963
rect 9079 15932 9474 15960
rect 9079 15929 9091 15932
rect 9033 15923 9091 15929
rect 9462 15929 9474 15932
rect 9508 15929 9520 15963
rect 9462 15923 9520 15929
rect 8389 15895 8447 15901
rect 8389 15892 8401 15895
rect 7156 15864 8401 15892
rect 7156 15852 7162 15864
rect 8389 15861 8401 15864
rect 8435 15861 8447 15895
rect 8389 15855 8447 15861
rect 8757 15895 8815 15901
rect 8757 15861 8769 15895
rect 8803 15892 8815 15895
rect 8846 15892 8852 15904
rect 8803 15864 8852 15892
rect 8803 15861 8815 15864
rect 8757 15855 8815 15861
rect 8846 15852 8852 15864
rect 8904 15852 8910 15904
rect 10594 15892 10600 15904
rect 10555 15864 10600 15892
rect 10594 15852 10600 15864
rect 10652 15892 10658 15904
rect 10965 15895 11023 15901
rect 10965 15892 10977 15895
rect 10652 15864 10977 15892
rect 10652 15852 10658 15864
rect 10965 15861 10977 15864
rect 11011 15861 11023 15895
rect 10965 15855 11023 15861
rect 1104 15802 14812 15824
rect 1104 15750 6315 15802
rect 6367 15750 6379 15802
rect 6431 15750 6443 15802
rect 6495 15750 6507 15802
rect 6559 15750 11648 15802
rect 11700 15750 11712 15802
rect 11764 15750 11776 15802
rect 11828 15750 11840 15802
rect 11892 15750 14812 15802
rect 1104 15728 14812 15750
rect 5534 15648 5540 15700
rect 5592 15688 5598 15700
rect 6549 15691 6607 15697
rect 6549 15688 6561 15691
rect 5592 15660 6561 15688
rect 5592 15648 5598 15660
rect 6549 15657 6561 15660
rect 6595 15657 6607 15691
rect 6549 15651 6607 15657
rect 7929 15691 7987 15697
rect 7929 15657 7941 15691
rect 7975 15688 7987 15691
rect 8113 15691 8171 15697
rect 8113 15688 8125 15691
rect 7975 15660 8125 15688
rect 7975 15657 7987 15660
rect 7929 15651 7987 15657
rect 8113 15657 8125 15660
rect 8159 15688 8171 15691
rect 8202 15688 8208 15700
rect 8159 15660 8208 15688
rect 8159 15657 8171 15660
rect 8113 15651 8171 15657
rect 8202 15648 8208 15660
rect 8260 15648 8266 15700
rect 9214 15688 9220 15700
rect 9175 15660 9220 15688
rect 9214 15648 9220 15660
rect 9272 15648 9278 15700
rect 9950 15648 9956 15700
rect 10008 15688 10014 15700
rect 10321 15691 10379 15697
rect 10321 15688 10333 15691
rect 10008 15660 10333 15688
rect 10008 15648 10014 15660
rect 10321 15657 10333 15660
rect 10367 15688 10379 15691
rect 11054 15688 11060 15700
rect 10367 15660 11060 15688
rect 10367 15657 10379 15660
rect 10321 15651 10379 15657
rect 11054 15648 11060 15660
rect 11112 15648 11118 15700
rect 6914 15552 6920 15564
rect 6875 15524 6920 15552
rect 6914 15512 6920 15524
rect 6972 15512 6978 15564
rect 7006 15484 7012 15496
rect 6967 15456 7012 15484
rect 7006 15444 7012 15456
rect 7064 15444 7070 15496
rect 7098 15444 7104 15496
rect 7156 15484 7162 15496
rect 7156 15456 7249 15484
rect 7156 15444 7162 15456
rect 9950 15444 9956 15496
rect 10008 15484 10014 15496
rect 10413 15487 10471 15493
rect 10413 15484 10425 15487
rect 10008 15456 10425 15484
rect 10008 15444 10014 15456
rect 10413 15453 10425 15456
rect 10459 15453 10471 15487
rect 10413 15447 10471 15453
rect 10505 15487 10563 15493
rect 10505 15453 10517 15487
rect 10551 15453 10563 15487
rect 10505 15447 10563 15453
rect 5442 15416 5448 15428
rect 5355 15388 5448 15416
rect 5442 15376 5448 15388
rect 5500 15416 5506 15428
rect 5810 15416 5816 15428
rect 5500 15388 5816 15416
rect 5500 15376 5506 15388
rect 5810 15376 5816 15388
rect 5868 15376 5874 15428
rect 6822 15376 6828 15428
rect 6880 15416 6886 15428
rect 7116 15416 7144 15444
rect 6880 15388 7144 15416
rect 6880 15376 6886 15388
rect 10318 15376 10324 15428
rect 10376 15416 10382 15428
rect 10520 15416 10548 15447
rect 10376 15388 10548 15416
rect 10376 15376 10382 15388
rect 5074 15348 5080 15360
rect 5035 15320 5080 15348
rect 5074 15308 5080 15320
rect 5132 15308 5138 15360
rect 5534 15308 5540 15360
rect 5592 15348 5598 15360
rect 5718 15348 5724 15360
rect 5592 15320 5724 15348
rect 5592 15308 5598 15320
rect 5718 15308 5724 15320
rect 5776 15308 5782 15360
rect 8202 15308 8208 15360
rect 8260 15348 8266 15360
rect 8386 15348 8392 15360
rect 8260 15320 8392 15348
rect 8260 15308 8266 15320
rect 8386 15308 8392 15320
rect 8444 15348 8450 15360
rect 8573 15351 8631 15357
rect 8573 15348 8585 15351
rect 8444 15320 8585 15348
rect 8444 15308 8450 15320
rect 8573 15317 8585 15320
rect 8619 15317 8631 15351
rect 8573 15311 8631 15317
rect 9953 15351 10011 15357
rect 9953 15317 9965 15351
rect 9999 15348 10011 15351
rect 10502 15348 10508 15360
rect 9999 15320 10508 15348
rect 9999 15317 10011 15320
rect 9953 15311 10011 15317
rect 10502 15308 10508 15320
rect 10560 15308 10566 15360
rect 1104 15258 14812 15280
rect 1104 15206 3648 15258
rect 3700 15206 3712 15258
rect 3764 15206 3776 15258
rect 3828 15206 3840 15258
rect 3892 15206 8982 15258
rect 9034 15206 9046 15258
rect 9098 15206 9110 15258
rect 9162 15206 9174 15258
rect 9226 15206 14315 15258
rect 14367 15206 14379 15258
rect 14431 15206 14443 15258
rect 14495 15206 14507 15258
rect 14559 15206 14812 15258
rect 1104 15184 14812 15206
rect 6641 15147 6699 15153
rect 6641 15113 6653 15147
rect 6687 15144 6699 15147
rect 6822 15144 6828 15156
rect 6687 15116 6828 15144
rect 6687 15113 6699 15116
rect 6641 15107 6699 15113
rect 6822 15104 6828 15116
rect 6880 15104 6886 15156
rect 7834 15104 7840 15156
rect 7892 15144 7898 15156
rect 8113 15147 8171 15153
rect 8113 15144 8125 15147
rect 7892 15116 8125 15144
rect 7892 15104 7898 15116
rect 8113 15113 8125 15116
rect 8159 15113 8171 15147
rect 8113 15107 8171 15113
rect 9125 15147 9183 15153
rect 9125 15113 9137 15147
rect 9171 15144 9183 15147
rect 9950 15144 9956 15156
rect 9171 15116 9956 15144
rect 9171 15113 9183 15116
rect 9125 15107 9183 15113
rect 9950 15104 9956 15116
rect 10008 15104 10014 15156
rect 11054 15144 11060 15156
rect 11015 15116 11060 15144
rect 11054 15104 11060 15116
rect 11112 15104 11118 15156
rect 5905 15079 5963 15085
rect 5905 15045 5917 15079
rect 5951 15076 5963 15079
rect 6914 15076 6920 15088
rect 5951 15048 6920 15076
rect 5951 15045 5963 15048
rect 5905 15039 5963 15045
rect 6914 15036 6920 15048
rect 6972 15076 6978 15088
rect 7101 15079 7159 15085
rect 7101 15076 7113 15079
rect 6972 15048 7113 15076
rect 6972 15036 6978 15048
rect 7101 15045 7113 15048
rect 7147 15045 7159 15079
rect 7101 15039 7159 15045
rect 9398 15036 9404 15088
rect 9456 15076 9462 15088
rect 9677 15079 9735 15085
rect 9677 15076 9689 15079
rect 9456 15048 9689 15076
rect 9456 15036 9462 15048
rect 9677 15045 9689 15048
rect 9723 15076 9735 15079
rect 9769 15079 9827 15085
rect 9769 15076 9781 15079
rect 9723 15048 9781 15076
rect 9723 15045 9735 15048
rect 9677 15039 9735 15045
rect 9769 15045 9781 15048
rect 9815 15045 9827 15079
rect 9769 15039 9827 15045
rect 7190 14968 7196 15020
rect 7248 15008 7254 15020
rect 7650 15008 7656 15020
rect 7248 14980 7656 15008
rect 7248 14968 7254 14980
rect 7650 14968 7656 14980
rect 7708 14968 7714 15020
rect 9493 15011 9551 15017
rect 9493 14977 9505 15011
rect 9539 15008 9551 15011
rect 10505 15011 10563 15017
rect 10505 15008 10517 15011
rect 9539 14980 10517 15008
rect 9539 14977 9551 14980
rect 9493 14971 9551 14977
rect 10505 14977 10517 14980
rect 10551 15008 10563 15011
rect 10594 15008 10600 15020
rect 10551 14980 10600 15008
rect 10551 14977 10563 14980
rect 10505 14971 10563 14977
rect 10594 14968 10600 14980
rect 10652 14968 10658 15020
rect 3142 14940 3148 14952
rect 3103 14912 3148 14940
rect 3142 14900 3148 14912
rect 3200 14940 3206 14952
rect 5534 14940 5540 14952
rect 3200 14912 5540 14940
rect 3200 14900 3206 14912
rect 5534 14900 5540 14912
rect 5592 14900 5598 14952
rect 7469 14943 7527 14949
rect 7469 14909 7481 14943
rect 7515 14940 7527 14943
rect 7834 14940 7840 14952
rect 7515 14912 7840 14940
rect 7515 14909 7527 14912
rect 7469 14903 7527 14909
rect 7834 14900 7840 14912
rect 7892 14900 7898 14952
rect 10134 14900 10140 14952
rect 10192 14940 10198 14952
rect 10321 14943 10379 14949
rect 10321 14940 10333 14943
rect 10192 14912 10333 14940
rect 10192 14900 10198 14912
rect 10321 14909 10333 14912
rect 10367 14909 10379 14943
rect 10321 14903 10379 14909
rect 3053 14875 3111 14881
rect 3053 14841 3065 14875
rect 3099 14872 3111 14875
rect 3390 14875 3448 14881
rect 3390 14872 3402 14875
rect 3099 14844 3402 14872
rect 3099 14841 3111 14844
rect 3053 14835 3111 14841
rect 3390 14841 3402 14844
rect 3436 14872 3448 14875
rect 3970 14872 3976 14884
rect 3436 14844 3976 14872
rect 3436 14841 3448 14844
rect 3390 14835 3448 14841
rect 3970 14832 3976 14844
rect 4028 14832 4034 14884
rect 6273 14875 6331 14881
rect 6273 14841 6285 14875
rect 6319 14872 6331 14875
rect 7561 14875 7619 14881
rect 7561 14872 7573 14875
rect 6319 14844 7573 14872
rect 6319 14841 6331 14844
rect 6273 14835 6331 14841
rect 7561 14841 7573 14844
rect 7607 14872 7619 14875
rect 7650 14872 7656 14884
rect 7607 14844 7656 14872
rect 7607 14841 7619 14844
rect 7561 14835 7619 14841
rect 7650 14832 7656 14844
rect 7708 14832 7714 14884
rect 9677 14875 9735 14881
rect 9677 14841 9689 14875
rect 9723 14872 9735 14875
rect 10413 14875 10471 14881
rect 10413 14872 10425 14875
rect 9723 14844 10425 14872
rect 9723 14841 9735 14844
rect 9677 14835 9735 14841
rect 10413 14841 10425 14844
rect 10459 14841 10471 14875
rect 10413 14835 10471 14841
rect 4525 14807 4583 14813
rect 4525 14773 4537 14807
rect 4571 14804 4583 14807
rect 4614 14804 4620 14816
rect 4571 14776 4620 14804
rect 4571 14773 4583 14776
rect 4525 14767 4583 14773
rect 4614 14764 4620 14776
rect 4672 14764 4678 14816
rect 1104 14714 14812 14736
rect 1104 14662 6315 14714
rect 6367 14662 6379 14714
rect 6431 14662 6443 14714
rect 6495 14662 6507 14714
rect 6559 14662 11648 14714
rect 11700 14662 11712 14714
rect 11764 14662 11776 14714
rect 11828 14662 11840 14714
rect 11892 14662 14812 14714
rect 1104 14640 14812 14662
rect 3142 14600 3148 14612
rect 3103 14572 3148 14600
rect 3142 14560 3148 14572
rect 3200 14560 3206 14612
rect 4522 14560 4528 14612
rect 4580 14600 4586 14612
rect 4985 14603 5043 14609
rect 4985 14600 4997 14603
rect 4580 14572 4997 14600
rect 4580 14560 4586 14572
rect 4985 14569 4997 14572
rect 5031 14600 5043 14603
rect 5350 14600 5356 14612
rect 5031 14572 5356 14600
rect 5031 14569 5043 14572
rect 4985 14563 5043 14569
rect 5350 14560 5356 14572
rect 5408 14560 5414 14612
rect 7190 14600 7196 14612
rect 7151 14572 7196 14600
rect 7190 14560 7196 14572
rect 7248 14560 7254 14612
rect 7650 14600 7656 14612
rect 7611 14572 7656 14600
rect 7650 14560 7656 14572
rect 7708 14560 7714 14612
rect 7926 14560 7932 14612
rect 7984 14600 7990 14612
rect 8021 14603 8079 14609
rect 8021 14600 8033 14603
rect 7984 14572 8033 14600
rect 7984 14560 7990 14572
rect 8021 14569 8033 14572
rect 8067 14569 8079 14603
rect 8021 14563 8079 14569
rect 9674 14560 9680 14612
rect 9732 14600 9738 14612
rect 9950 14600 9956 14612
rect 9732 14572 9956 14600
rect 9732 14560 9738 14572
rect 9950 14560 9956 14572
rect 10008 14560 10014 14612
rect 10045 14603 10103 14609
rect 10045 14569 10057 14603
rect 10091 14600 10103 14603
rect 10134 14600 10140 14612
rect 10091 14572 10140 14600
rect 10091 14569 10103 14572
rect 10045 14563 10103 14569
rect 10134 14560 10140 14572
rect 10192 14600 10198 14612
rect 10502 14600 10508 14612
rect 10192 14572 10508 14600
rect 10192 14560 10198 14572
rect 10502 14560 10508 14572
rect 10560 14560 10566 14612
rect 10318 14532 10324 14544
rect 10279 14504 10324 14532
rect 10318 14492 10324 14504
rect 10376 14492 10382 14544
rect 4890 14464 4896 14476
rect 4851 14436 4896 14464
rect 4890 14424 4896 14436
rect 4948 14424 4954 14476
rect 6273 14467 6331 14473
rect 6273 14433 6285 14467
rect 6319 14464 6331 14467
rect 7558 14464 7564 14476
rect 6319 14436 7564 14464
rect 6319 14433 6331 14436
rect 6273 14427 6331 14433
rect 7558 14424 7564 14436
rect 7616 14424 7622 14476
rect 8110 14464 8116 14476
rect 8071 14436 8116 14464
rect 8110 14424 8116 14436
rect 8168 14424 8174 14476
rect 5077 14399 5135 14405
rect 5077 14396 5089 14399
rect 4724 14368 5089 14396
rect 4062 14288 4068 14340
rect 4120 14328 4126 14340
rect 4525 14331 4583 14337
rect 4525 14328 4537 14331
rect 4120 14300 4537 14328
rect 4120 14288 4126 14300
rect 4525 14297 4537 14300
rect 4571 14297 4583 14331
rect 4525 14291 4583 14297
rect 4724 14272 4752 14368
rect 5077 14365 5089 14368
rect 5123 14396 5135 14399
rect 5534 14396 5540 14408
rect 5123 14368 5540 14396
rect 5123 14365 5135 14368
rect 5077 14359 5135 14365
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 8202 14356 8208 14408
rect 8260 14396 8266 14408
rect 8260 14368 8305 14396
rect 8260 14356 8266 14368
rect 3326 14220 3332 14272
rect 3384 14260 3390 14272
rect 4433 14263 4491 14269
rect 4433 14260 4445 14263
rect 3384 14232 4445 14260
rect 3384 14220 3390 14232
rect 4433 14229 4445 14232
rect 4479 14260 4491 14263
rect 4706 14260 4712 14272
rect 4479 14232 4712 14260
rect 4479 14229 4491 14232
rect 4433 14223 4491 14229
rect 4706 14220 4712 14232
rect 4764 14220 4770 14272
rect 5810 14220 5816 14272
rect 5868 14260 5874 14272
rect 6089 14263 6147 14269
rect 6089 14260 6101 14263
rect 5868 14232 6101 14260
rect 5868 14220 5874 14232
rect 6089 14229 6101 14232
rect 6135 14229 6147 14263
rect 6089 14223 6147 14229
rect 6641 14263 6699 14269
rect 6641 14229 6653 14263
rect 6687 14260 6699 14263
rect 6822 14260 6828 14272
rect 6687 14232 6828 14260
rect 6687 14229 6699 14232
rect 6641 14223 6699 14229
rect 6822 14220 6828 14232
rect 6880 14220 6886 14272
rect 7377 14263 7435 14269
rect 7377 14229 7389 14263
rect 7423 14260 7435 14263
rect 8294 14260 8300 14272
rect 7423 14232 8300 14260
rect 7423 14229 7435 14232
rect 7377 14223 7435 14229
rect 8294 14220 8300 14232
rect 8352 14220 8358 14272
rect 1104 14170 14812 14192
rect 1104 14118 3648 14170
rect 3700 14118 3712 14170
rect 3764 14118 3776 14170
rect 3828 14118 3840 14170
rect 3892 14118 8982 14170
rect 9034 14118 9046 14170
rect 9098 14118 9110 14170
rect 9162 14118 9174 14170
rect 9226 14118 14315 14170
rect 14367 14118 14379 14170
rect 14431 14118 14443 14170
rect 14495 14118 14507 14170
rect 14559 14118 14812 14170
rect 1104 14096 14812 14118
rect 2685 14059 2743 14065
rect 2685 14025 2697 14059
rect 2731 14056 2743 14059
rect 3418 14056 3424 14068
rect 2731 14028 3424 14056
rect 2731 14025 2743 14028
rect 2685 14019 2743 14025
rect 3418 14016 3424 14028
rect 3476 14016 3482 14068
rect 4522 14056 4528 14068
rect 4483 14028 4528 14056
rect 4522 14016 4528 14028
rect 4580 14016 4586 14068
rect 6457 14059 6515 14065
rect 6457 14025 6469 14059
rect 6503 14056 6515 14059
rect 7377 14059 7435 14065
rect 7377 14056 7389 14059
rect 6503 14028 7389 14056
rect 6503 14025 6515 14028
rect 6457 14019 6515 14025
rect 7377 14025 7389 14028
rect 7423 14056 7435 14059
rect 7558 14056 7564 14068
rect 7423 14028 7564 14056
rect 7423 14025 7435 14028
rect 7377 14019 7435 14025
rect 7558 14016 7564 14028
rect 7616 14016 7622 14068
rect 7745 14059 7803 14065
rect 7745 14025 7757 14059
rect 7791 14056 7803 14059
rect 7926 14056 7932 14068
rect 7791 14028 7932 14056
rect 7791 14025 7803 14028
rect 7745 14019 7803 14025
rect 7926 14016 7932 14028
rect 7984 14056 7990 14068
rect 8754 14056 8760 14068
rect 7984 14028 8760 14056
rect 7984 14016 7990 14028
rect 8754 14016 8760 14028
rect 8812 14016 8818 14068
rect 4154 13948 4160 14000
rect 4212 13988 4218 14000
rect 4985 13991 5043 13997
rect 4985 13988 4997 13991
rect 4212 13960 4997 13988
rect 4212 13948 4218 13960
rect 4985 13957 4997 13960
rect 5031 13957 5043 13991
rect 8110 13988 8116 14000
rect 8071 13960 8116 13988
rect 4985 13951 5043 13957
rect 8110 13948 8116 13960
rect 8168 13948 8174 14000
rect 5534 13920 5540 13932
rect 5495 13892 5540 13920
rect 5534 13880 5540 13892
rect 5592 13880 5598 13932
rect 9674 13880 9680 13932
rect 9732 13920 9738 13932
rect 10137 13923 10195 13929
rect 10137 13920 10149 13923
rect 9732 13892 10149 13920
rect 9732 13880 9738 13892
rect 10137 13889 10149 13892
rect 10183 13920 10195 13923
rect 10781 13923 10839 13929
rect 10781 13920 10793 13923
rect 10183 13892 10793 13920
rect 10183 13889 10195 13892
rect 10137 13883 10195 13889
rect 10781 13889 10793 13892
rect 10827 13889 10839 13923
rect 10781 13883 10839 13889
rect 2774 13812 2780 13864
rect 2832 13852 2838 13864
rect 3044 13855 3102 13861
rect 2832 13824 2877 13852
rect 2832 13812 2838 13824
rect 3044 13821 3056 13855
rect 3090 13852 3102 13855
rect 3326 13852 3332 13864
rect 3090 13824 3332 13852
rect 3090 13821 3102 13824
rect 3044 13815 3102 13821
rect 3326 13812 3332 13824
rect 3384 13812 3390 13864
rect 5258 13812 5264 13864
rect 5316 13852 5322 13864
rect 5442 13852 5448 13864
rect 5316 13824 5448 13852
rect 5316 13812 5322 13824
rect 5442 13812 5448 13824
rect 5500 13852 5506 13864
rect 5997 13855 6055 13861
rect 5997 13852 6009 13855
rect 5500 13824 6009 13852
rect 5500 13812 5506 13824
rect 5997 13821 6009 13824
rect 6043 13821 6055 13855
rect 5997 13815 6055 13821
rect 8202 13812 8208 13864
rect 8260 13852 8266 13864
rect 8389 13855 8447 13861
rect 8389 13852 8401 13855
rect 8260 13824 8401 13852
rect 8260 13812 8266 13824
rect 8389 13821 8401 13824
rect 8435 13821 8447 13855
rect 8389 13815 8447 13821
rect 9401 13855 9459 13861
rect 9401 13821 9413 13855
rect 9447 13852 9459 13855
rect 9769 13855 9827 13861
rect 9447 13824 9628 13852
rect 9447 13821 9459 13824
rect 9401 13815 9459 13821
rect 5166 13744 5172 13796
rect 5224 13784 5230 13796
rect 5534 13784 5540 13796
rect 5224 13756 5540 13784
rect 5224 13744 5230 13756
rect 5534 13744 5540 13756
rect 5592 13744 5598 13796
rect 9600 13784 9628 13824
rect 9769 13821 9781 13855
rect 9815 13852 9827 13855
rect 10689 13855 10747 13861
rect 10689 13852 10701 13855
rect 9815 13824 10701 13852
rect 9815 13821 9827 13824
rect 9769 13815 9827 13821
rect 10689 13821 10701 13824
rect 10735 13852 10747 13855
rect 11054 13852 11060 13864
rect 10735 13824 11060 13852
rect 10735 13821 10747 13824
rect 10689 13815 10747 13821
rect 11054 13812 11060 13824
rect 11112 13812 11118 13864
rect 10597 13787 10655 13793
rect 10597 13784 10609 13787
rect 9600 13756 10609 13784
rect 10597 13753 10609 13756
rect 10643 13784 10655 13787
rect 11238 13784 11244 13796
rect 10643 13756 11244 13784
rect 10643 13753 10655 13756
rect 10597 13747 10655 13753
rect 11238 13744 11244 13756
rect 11296 13744 11302 13796
rect 3970 13676 3976 13728
rect 4028 13716 4034 13728
rect 4157 13719 4215 13725
rect 4157 13716 4169 13719
rect 4028 13688 4169 13716
rect 4028 13676 4034 13688
rect 4157 13685 4169 13688
rect 4203 13685 4215 13719
rect 4157 13679 4215 13685
rect 4798 13676 4804 13728
rect 4856 13716 4862 13728
rect 4893 13719 4951 13725
rect 4893 13716 4905 13719
rect 4856 13688 4905 13716
rect 4856 13676 4862 13688
rect 4893 13685 4905 13688
rect 4939 13716 4951 13719
rect 5353 13719 5411 13725
rect 5353 13716 5365 13719
rect 4939 13688 5365 13716
rect 4939 13685 4951 13688
rect 4893 13679 4951 13685
rect 5353 13685 5365 13688
rect 5399 13716 5411 13719
rect 5442 13716 5448 13728
rect 5399 13688 5448 13716
rect 5399 13685 5411 13688
rect 5353 13679 5411 13685
rect 5442 13676 5448 13688
rect 5500 13676 5506 13728
rect 10134 13676 10140 13728
rect 10192 13716 10198 13728
rect 10229 13719 10287 13725
rect 10229 13716 10241 13719
rect 10192 13688 10241 13716
rect 10192 13676 10198 13688
rect 10229 13685 10241 13688
rect 10275 13685 10287 13719
rect 10229 13679 10287 13685
rect 1104 13626 14812 13648
rect 1104 13574 6315 13626
rect 6367 13574 6379 13626
rect 6431 13574 6443 13626
rect 6495 13574 6507 13626
rect 6559 13574 11648 13626
rect 11700 13574 11712 13626
rect 11764 13574 11776 13626
rect 11828 13574 11840 13626
rect 11892 13574 14812 13626
rect 1104 13552 14812 13574
rect 3697 13515 3755 13521
rect 3697 13481 3709 13515
rect 3743 13512 3755 13515
rect 4062 13512 4068 13524
rect 3743 13484 4068 13512
rect 3743 13481 3755 13484
rect 3697 13475 3755 13481
rect 4062 13472 4068 13484
rect 4120 13472 4126 13524
rect 4433 13515 4491 13521
rect 4433 13481 4445 13515
rect 4479 13512 4491 13515
rect 4890 13512 4896 13524
rect 4479 13484 4896 13512
rect 4479 13481 4491 13484
rect 4433 13475 4491 13481
rect 1670 13444 1676 13456
rect 1631 13416 1676 13444
rect 1670 13404 1676 13416
rect 1728 13404 1734 13456
rect 2961 13447 3019 13453
rect 2961 13413 2973 13447
rect 3007 13444 3019 13447
rect 4448 13444 4476 13475
rect 4890 13472 4896 13484
rect 4948 13472 4954 13524
rect 8294 13472 8300 13524
rect 8352 13512 8358 13524
rect 8389 13515 8447 13521
rect 8389 13512 8401 13515
rect 8352 13484 8401 13512
rect 8352 13472 8358 13484
rect 8389 13481 8401 13484
rect 8435 13481 8447 13515
rect 8389 13475 8447 13481
rect 6730 13444 6736 13456
rect 3007 13416 4476 13444
rect 6656 13416 6736 13444
rect 3007 13413 3019 13416
rect 2961 13407 3019 13413
rect 1394 13376 1400 13388
rect 1355 13348 1400 13376
rect 1394 13336 1400 13348
rect 1452 13336 1458 13388
rect 4614 13336 4620 13388
rect 4672 13376 4678 13388
rect 4781 13379 4839 13385
rect 4781 13376 4793 13379
rect 4672 13348 4793 13376
rect 4672 13336 4678 13348
rect 4781 13345 4793 13348
rect 4827 13345 4839 13379
rect 4781 13339 4839 13345
rect 4525 13311 4583 13317
rect 4525 13277 4537 13311
rect 4571 13277 4583 13311
rect 4525 13271 4583 13277
rect 2222 13172 2228 13184
rect 2183 13144 2228 13172
rect 2222 13132 2228 13144
rect 2280 13132 2286 13184
rect 2774 13132 2780 13184
rect 2832 13172 2838 13184
rect 2869 13175 2927 13181
rect 2869 13172 2881 13175
rect 2832 13144 2881 13172
rect 2832 13132 2838 13144
rect 2869 13141 2881 13144
rect 2915 13172 2927 13175
rect 3142 13172 3148 13184
rect 2915 13144 3148 13172
rect 2915 13141 2927 13144
rect 2869 13135 2927 13141
rect 3142 13132 3148 13144
rect 3200 13172 3206 13184
rect 4540 13172 4568 13271
rect 6656 13240 6684 13416
rect 6730 13404 6736 13416
rect 6788 13404 6794 13456
rect 7000 13379 7058 13385
rect 7000 13345 7012 13379
rect 7046 13376 7058 13379
rect 7834 13376 7840 13388
rect 7046 13348 7840 13376
rect 7046 13345 7058 13348
rect 7000 13339 7058 13345
rect 7834 13336 7840 13348
rect 7892 13336 7898 13388
rect 8404 13376 8432 13475
rect 8846 13472 8852 13524
rect 8904 13512 8910 13524
rect 8941 13515 8999 13521
rect 8941 13512 8953 13515
rect 8904 13484 8953 13512
rect 8904 13472 8910 13484
rect 8941 13481 8953 13484
rect 8987 13512 8999 13515
rect 9306 13512 9312 13524
rect 8987 13484 9312 13512
rect 8987 13481 8999 13484
rect 8941 13475 8999 13481
rect 9306 13472 9312 13484
rect 9364 13512 9370 13524
rect 9401 13515 9459 13521
rect 9401 13512 9413 13515
rect 9364 13484 9413 13512
rect 9364 13472 9370 13484
rect 9401 13481 9413 13484
rect 9447 13481 9459 13515
rect 9674 13512 9680 13524
rect 9635 13484 9680 13512
rect 9401 13475 9459 13481
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 11238 13512 11244 13524
rect 11199 13484 11244 13512
rect 11238 13472 11244 13484
rect 11296 13472 11302 13524
rect 8570 13376 8576 13388
rect 8404 13348 8576 13376
rect 8570 13336 8576 13348
rect 8628 13376 8634 13388
rect 9125 13379 9183 13385
rect 9125 13376 9137 13379
rect 8628 13348 9137 13376
rect 8628 13336 8634 13348
rect 9125 13345 9137 13348
rect 9171 13345 9183 13379
rect 10042 13376 10048 13388
rect 10003 13348 10048 13376
rect 9125 13339 9183 13345
rect 10042 13336 10048 13348
rect 10100 13336 10106 13388
rect 11606 13376 11612 13388
rect 11567 13348 11612 13376
rect 11606 13336 11612 13348
rect 11664 13336 11670 13388
rect 11698 13336 11704 13388
rect 11756 13376 11762 13388
rect 12250 13376 12256 13388
rect 11756 13348 12256 13376
rect 11756 13336 11762 13348
rect 12250 13336 12256 13348
rect 12308 13336 12314 13388
rect 6733 13311 6791 13317
rect 6733 13277 6745 13311
rect 6779 13277 6791 13311
rect 10134 13308 10140 13320
rect 10095 13280 10140 13308
rect 6733 13271 6791 13277
rect 6104 13212 6684 13240
rect 6104 13184 6132 13212
rect 5166 13172 5172 13184
rect 3200 13144 5172 13172
rect 3200 13132 3206 13144
rect 5166 13132 5172 13144
rect 5224 13132 5230 13184
rect 5902 13172 5908 13184
rect 5863 13144 5908 13172
rect 5902 13132 5908 13144
rect 5960 13132 5966 13184
rect 6086 13132 6092 13184
rect 6144 13132 6150 13184
rect 6641 13175 6699 13181
rect 6641 13141 6653 13175
rect 6687 13172 6699 13175
rect 6748 13172 6776 13271
rect 10134 13268 10140 13280
rect 10192 13268 10198 13320
rect 10318 13308 10324 13320
rect 10279 13280 10324 13308
rect 10318 13268 10324 13280
rect 10376 13268 10382 13320
rect 11790 13308 11796 13320
rect 11751 13280 11796 13308
rect 11790 13268 11796 13280
rect 11848 13268 11854 13320
rect 8386 13240 8392 13252
rect 7944 13212 8392 13240
rect 7650 13172 7656 13184
rect 6687 13144 7656 13172
rect 6687 13141 6699 13144
rect 6641 13135 6699 13141
rect 7650 13132 7656 13144
rect 7708 13172 7714 13184
rect 7944 13172 7972 13212
rect 8386 13200 8392 13212
rect 8444 13200 8450 13252
rect 8110 13172 8116 13184
rect 7708 13144 7972 13172
rect 8071 13144 8116 13172
rect 7708 13132 7714 13144
rect 8110 13132 8116 13144
rect 8168 13132 8174 13184
rect 1104 13082 14812 13104
rect 1104 13030 3648 13082
rect 3700 13030 3712 13082
rect 3764 13030 3776 13082
rect 3828 13030 3840 13082
rect 3892 13030 8982 13082
rect 9034 13030 9046 13082
rect 9098 13030 9110 13082
rect 9162 13030 9174 13082
rect 9226 13030 14315 13082
rect 14367 13030 14379 13082
rect 14431 13030 14443 13082
rect 14495 13030 14507 13082
rect 14559 13030 14812 13082
rect 1104 13008 14812 13030
rect 3142 12968 3148 12980
rect 3103 12940 3148 12968
rect 3142 12928 3148 12940
rect 3200 12928 3206 12980
rect 3234 12928 3240 12980
rect 3292 12968 3298 12980
rect 3513 12971 3571 12977
rect 3513 12968 3525 12971
rect 3292 12940 3525 12968
rect 3292 12928 3298 12940
rect 3513 12937 3525 12940
rect 3559 12968 3571 12971
rect 3970 12968 3976 12980
rect 3559 12940 3976 12968
rect 3559 12937 3571 12940
rect 3513 12931 3571 12937
rect 3970 12928 3976 12940
rect 4028 12928 4034 12980
rect 5077 12971 5135 12977
rect 5077 12937 5089 12971
rect 5123 12968 5135 12971
rect 5258 12968 5264 12980
rect 5123 12940 5264 12968
rect 5123 12937 5135 12940
rect 5077 12931 5135 12937
rect 5258 12928 5264 12940
rect 5316 12928 5322 12980
rect 6273 12971 6331 12977
rect 6273 12937 6285 12971
rect 6319 12968 6331 12971
rect 7834 12968 7840 12980
rect 6319 12940 7840 12968
rect 6319 12937 6331 12940
rect 6273 12931 6331 12937
rect 3605 12903 3663 12909
rect 3605 12869 3617 12903
rect 3651 12869 3663 12903
rect 3605 12863 3663 12869
rect 1949 12835 2007 12841
rect 1949 12801 1961 12835
rect 1995 12832 2007 12835
rect 2682 12832 2688 12844
rect 1995 12804 2688 12832
rect 1995 12801 2007 12804
rect 1949 12795 2007 12801
rect 2682 12792 2688 12804
rect 2740 12792 2746 12844
rect 2222 12724 2228 12776
rect 2280 12764 2286 12776
rect 2409 12767 2467 12773
rect 2409 12764 2421 12767
rect 2280 12736 2421 12764
rect 2280 12724 2286 12736
rect 2409 12733 2421 12736
rect 2455 12764 2467 12767
rect 3620 12764 3648 12863
rect 3988 12832 4016 12928
rect 4614 12900 4620 12912
rect 4575 12872 4620 12900
rect 4614 12860 4620 12872
rect 4672 12860 4678 12912
rect 4157 12835 4215 12841
rect 4157 12832 4169 12835
rect 3988 12804 4169 12832
rect 4157 12801 4169 12804
rect 4203 12801 4215 12835
rect 5276 12832 5304 12928
rect 5629 12835 5687 12841
rect 5629 12832 5641 12835
rect 5276 12804 5641 12832
rect 4157 12795 4215 12801
rect 5629 12801 5641 12804
rect 5675 12801 5687 12835
rect 5629 12795 5687 12801
rect 5813 12835 5871 12841
rect 5813 12801 5825 12835
rect 5859 12832 5871 12835
rect 5902 12832 5908 12844
rect 5859 12804 5908 12832
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 5902 12792 5908 12804
rect 5960 12832 5966 12844
rect 6288 12832 6316 12931
rect 7834 12928 7840 12940
rect 7892 12928 7898 12980
rect 8110 12928 8116 12980
rect 8168 12968 8174 12980
rect 8205 12971 8263 12977
rect 8205 12968 8217 12971
rect 8168 12940 8217 12968
rect 8168 12928 8174 12940
rect 8205 12937 8217 12940
rect 8251 12937 8263 12971
rect 8386 12968 8392 12980
rect 8347 12940 8392 12968
rect 8205 12931 8263 12937
rect 8386 12928 8392 12940
rect 8444 12928 8450 12980
rect 10134 12928 10140 12980
rect 10192 12968 10198 12980
rect 10594 12968 10600 12980
rect 10192 12940 10600 12968
rect 10192 12928 10198 12940
rect 10594 12928 10600 12940
rect 10652 12928 10658 12980
rect 11149 12971 11207 12977
rect 11149 12937 11161 12971
rect 11195 12968 11207 12971
rect 11330 12968 11336 12980
rect 11195 12940 11336 12968
rect 11195 12937 11207 12940
rect 11149 12931 11207 12937
rect 11330 12928 11336 12940
rect 11388 12968 11394 12980
rect 11790 12968 11796 12980
rect 11388 12940 11796 12968
rect 11388 12928 11394 12940
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 6641 12903 6699 12909
rect 6641 12869 6653 12903
rect 6687 12900 6699 12903
rect 7098 12900 7104 12912
rect 6687 12872 7104 12900
rect 6687 12869 6699 12872
rect 6641 12863 6699 12869
rect 7098 12860 7104 12872
rect 7156 12860 7162 12912
rect 5960 12804 6316 12832
rect 7469 12835 7527 12841
rect 5960 12792 5966 12804
rect 7469 12801 7481 12835
rect 7515 12832 7527 12835
rect 7650 12832 7656 12844
rect 7515 12804 7656 12832
rect 7515 12801 7527 12804
rect 7469 12795 7527 12801
rect 7650 12792 7656 12804
rect 7708 12832 7714 12844
rect 8128 12832 8156 12928
rect 11698 12900 11704 12912
rect 11659 12872 11704 12900
rect 11698 12860 11704 12872
rect 11756 12860 11762 12912
rect 7708 12804 8156 12832
rect 7708 12792 7714 12804
rect 8478 12792 8484 12844
rect 8536 12832 8542 12844
rect 8846 12832 8852 12844
rect 8536 12804 8852 12832
rect 8536 12792 8542 12804
rect 8846 12792 8852 12804
rect 8904 12832 8910 12844
rect 8941 12835 8999 12841
rect 8941 12832 8953 12835
rect 8904 12804 8953 12832
rect 8904 12792 8910 12804
rect 8941 12801 8953 12804
rect 8987 12801 8999 12835
rect 8941 12795 8999 12801
rect 11241 12835 11299 12841
rect 11241 12801 11253 12835
rect 11287 12832 11299 12835
rect 11606 12832 11612 12844
rect 11287 12804 11612 12832
rect 11287 12801 11299 12804
rect 11241 12795 11299 12801
rect 11606 12792 11612 12804
rect 11664 12832 11670 12844
rect 12069 12835 12127 12841
rect 12069 12832 12081 12835
rect 11664 12804 12081 12832
rect 11664 12792 11670 12804
rect 12069 12801 12081 12804
rect 12115 12801 12127 12835
rect 12069 12795 12127 12801
rect 2455 12736 3648 12764
rect 3973 12767 4031 12773
rect 2455 12733 2467 12736
rect 2409 12727 2467 12733
rect 3973 12733 3985 12767
rect 4019 12764 4031 12767
rect 4062 12764 4068 12776
rect 4019 12736 4068 12764
rect 4019 12733 4031 12736
rect 3973 12727 4031 12733
rect 4062 12724 4068 12736
rect 4120 12724 4126 12776
rect 4798 12724 4804 12776
rect 4856 12764 4862 12776
rect 5534 12764 5540 12776
rect 4856 12736 5540 12764
rect 4856 12724 4862 12736
rect 5534 12724 5540 12736
rect 5592 12764 5598 12776
rect 6730 12764 6736 12776
rect 5592 12736 6736 12764
rect 5592 12724 5598 12736
rect 6730 12724 6736 12736
rect 6788 12724 6794 12776
rect 6822 12724 6828 12776
rect 6880 12764 6886 12776
rect 7285 12767 7343 12773
rect 7285 12764 7297 12767
rect 6880 12736 7297 12764
rect 6880 12724 6886 12736
rect 7285 12733 7297 12736
rect 7331 12733 7343 12767
rect 8570 12764 8576 12776
rect 8531 12736 8576 12764
rect 7285 12727 7343 12733
rect 8570 12724 8576 12736
rect 8628 12724 8634 12776
rect 9030 12724 9036 12776
rect 9088 12764 9094 12776
rect 9208 12767 9266 12773
rect 9208 12764 9220 12767
rect 9088 12736 9220 12764
rect 9088 12724 9094 12736
rect 9208 12733 9220 12736
rect 9254 12764 9266 12767
rect 9582 12764 9588 12776
rect 9254 12736 9588 12764
rect 9254 12733 9266 12736
rect 9208 12727 9266 12733
rect 9582 12724 9588 12736
rect 9640 12724 9646 12776
rect 7098 12656 7104 12708
rect 7156 12696 7162 12708
rect 7193 12699 7251 12705
rect 7193 12696 7205 12699
rect 7156 12668 7205 12696
rect 7156 12656 7162 12668
rect 7193 12665 7205 12668
rect 7239 12665 7251 12699
rect 7193 12659 7251 12665
rect 8662 12656 8668 12708
rect 8720 12696 8726 12708
rect 8846 12696 8852 12708
rect 8720 12668 8852 12696
rect 8720 12656 8726 12668
rect 8846 12656 8852 12668
rect 8904 12656 8910 12708
rect 2038 12628 2044 12640
rect 1999 12600 2044 12628
rect 2038 12588 2044 12600
rect 2096 12588 2102 12640
rect 2498 12588 2504 12640
rect 2556 12628 2562 12640
rect 4062 12628 4068 12640
rect 2556 12600 2601 12628
rect 4023 12600 4068 12628
rect 2556 12588 2562 12600
rect 4062 12588 4068 12600
rect 4120 12588 4126 12640
rect 5169 12631 5227 12637
rect 5169 12597 5181 12631
rect 5215 12628 5227 12631
rect 5534 12628 5540 12640
rect 5215 12600 5540 12628
rect 5215 12597 5227 12600
rect 5169 12591 5227 12597
rect 5534 12588 5540 12600
rect 5592 12588 5598 12640
rect 5718 12588 5724 12640
rect 5776 12628 5782 12640
rect 6825 12631 6883 12637
rect 6825 12628 6837 12631
rect 5776 12600 6837 12628
rect 5776 12588 5782 12600
rect 6825 12597 6837 12600
rect 6871 12597 6883 12631
rect 6825 12591 6883 12597
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 10318 12628 10324 12640
rect 9732 12600 10324 12628
rect 9732 12588 9738 12600
rect 10318 12588 10324 12600
rect 10376 12588 10382 12640
rect 1104 12538 14812 12560
rect 1104 12486 6315 12538
rect 6367 12486 6379 12538
rect 6431 12486 6443 12538
rect 6495 12486 6507 12538
rect 6559 12486 11648 12538
rect 11700 12486 11712 12538
rect 11764 12486 11776 12538
rect 11828 12486 11840 12538
rect 11892 12486 14812 12538
rect 1104 12464 14812 12486
rect 1394 12384 1400 12436
rect 1452 12424 1458 12436
rect 1581 12427 1639 12433
rect 1581 12424 1593 12427
rect 1452 12396 1593 12424
rect 1452 12384 1458 12396
rect 1581 12393 1593 12396
rect 1627 12393 1639 12427
rect 1581 12387 1639 12393
rect 3697 12427 3755 12433
rect 3697 12393 3709 12427
rect 3743 12424 3755 12427
rect 4062 12424 4068 12436
rect 3743 12396 4068 12424
rect 3743 12393 3755 12396
rect 3697 12387 3755 12393
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 4246 12384 4252 12436
rect 4304 12424 4310 12436
rect 4433 12427 4491 12433
rect 4433 12424 4445 12427
rect 4304 12396 4445 12424
rect 4304 12384 4310 12396
rect 4433 12393 4445 12396
rect 4479 12424 4491 12427
rect 4522 12424 4528 12436
rect 4479 12396 4528 12424
rect 4479 12393 4491 12396
rect 4433 12387 4491 12393
rect 4522 12384 4528 12396
rect 4580 12384 4586 12436
rect 4798 12384 4804 12436
rect 4856 12424 4862 12436
rect 5169 12427 5227 12433
rect 5169 12424 5181 12427
rect 4856 12396 5181 12424
rect 4856 12384 4862 12396
rect 5169 12393 5181 12396
rect 5215 12393 5227 12427
rect 5169 12387 5227 12393
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 6641 12427 6699 12433
rect 6641 12424 6653 12427
rect 5592 12396 6653 12424
rect 5592 12384 5598 12396
rect 6641 12393 6653 12396
rect 6687 12424 6699 12427
rect 6822 12424 6828 12436
rect 6687 12396 6828 12424
rect 6687 12393 6699 12396
rect 6641 12387 6699 12393
rect 6822 12384 6828 12396
rect 6880 12384 6886 12436
rect 9030 12424 9036 12436
rect 8991 12396 9036 12424
rect 9030 12384 9036 12396
rect 9088 12384 9094 12436
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 10229 12427 10287 12433
rect 10229 12424 10241 12427
rect 10100 12396 10241 12424
rect 10100 12384 10106 12396
rect 10229 12393 10241 12396
rect 10275 12393 10287 12427
rect 10229 12387 10287 12393
rect 2958 12316 2964 12368
rect 3016 12356 3022 12368
rect 3142 12356 3148 12368
rect 3016 12328 3148 12356
rect 3016 12316 3022 12328
rect 3142 12316 3148 12328
rect 3200 12316 3206 12368
rect 5902 12316 5908 12368
rect 5960 12356 5966 12368
rect 6270 12356 6276 12368
rect 5960 12328 6276 12356
rect 5960 12316 5966 12328
rect 6270 12316 6276 12328
rect 6328 12316 6334 12368
rect 7006 12316 7012 12368
rect 7064 12365 7070 12368
rect 7064 12359 7128 12365
rect 7064 12325 7082 12359
rect 7116 12356 7128 12359
rect 8202 12356 8208 12368
rect 7116 12328 8208 12356
rect 7116 12325 7128 12328
rect 7064 12319 7128 12325
rect 7064 12316 7070 12319
rect 8202 12316 8208 12328
rect 8260 12316 8266 12368
rect 8570 12316 8576 12368
rect 8628 12356 8634 12368
rect 9309 12359 9367 12365
rect 9309 12356 9321 12359
rect 8628 12328 9321 12356
rect 8628 12316 8634 12328
rect 9309 12325 9321 12328
rect 9355 12325 9367 12359
rect 9309 12319 9367 12325
rect 10410 12316 10416 12368
rect 10468 12356 10474 12368
rect 10962 12356 10968 12368
rect 10468 12328 10968 12356
rect 10468 12316 10474 12328
rect 10962 12316 10968 12328
rect 11020 12316 11026 12368
rect 4525 12291 4583 12297
rect 4525 12257 4537 12291
rect 4571 12288 4583 12291
rect 4614 12288 4620 12300
rect 4571 12260 4620 12288
rect 4571 12257 4583 12260
rect 4525 12251 4583 12257
rect 4614 12248 4620 12260
rect 4672 12248 4678 12300
rect 5810 12288 5816 12300
rect 5771 12260 5816 12288
rect 5810 12248 5816 12260
rect 5868 12248 5874 12300
rect 8665 12291 8723 12297
rect 8665 12288 8677 12291
rect 8588 12260 8677 12288
rect 8588 12232 8616 12260
rect 8665 12257 8677 12260
rect 8711 12288 8723 12291
rect 10781 12291 10839 12297
rect 10781 12288 10793 12291
rect 8711 12260 10793 12288
rect 8711 12257 8723 12260
rect 8665 12251 8723 12257
rect 10781 12257 10793 12260
rect 10827 12288 10839 12291
rect 10870 12288 10876 12300
rect 10827 12260 10876 12288
rect 10827 12257 10839 12260
rect 10781 12251 10839 12257
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 11048 12291 11106 12297
rect 11048 12257 11060 12291
rect 11094 12288 11106 12291
rect 11330 12288 11336 12300
rect 11094 12260 11336 12288
rect 11094 12257 11106 12260
rect 11048 12251 11106 12257
rect 11330 12248 11336 12260
rect 11388 12248 11394 12300
rect 4706 12220 4712 12232
rect 4619 12192 4712 12220
rect 4706 12180 4712 12192
rect 4764 12220 4770 12232
rect 4890 12220 4896 12232
rect 4764 12192 4896 12220
rect 4764 12180 4770 12192
rect 4890 12180 4896 12192
rect 4948 12180 4954 12232
rect 5626 12180 5632 12232
rect 5684 12220 5690 12232
rect 5994 12220 6000 12232
rect 5684 12192 6000 12220
rect 5684 12180 5690 12192
rect 5994 12180 6000 12192
rect 6052 12180 6058 12232
rect 6822 12220 6828 12232
rect 6783 12192 6828 12220
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 8570 12180 8576 12232
rect 8628 12180 8634 12232
rect 9674 12180 9680 12232
rect 9732 12180 9738 12232
rect 9692 12152 9720 12180
rect 9953 12155 10011 12161
rect 9953 12152 9965 12155
rect 9692 12124 9965 12152
rect 9953 12121 9965 12124
rect 9999 12152 10011 12155
rect 10318 12152 10324 12164
rect 9999 12124 10324 12152
rect 9999 12121 10011 12124
rect 9953 12115 10011 12121
rect 10318 12112 10324 12124
rect 10376 12112 10382 12164
rect 2133 12087 2191 12093
rect 2133 12053 2145 12087
rect 2179 12084 2191 12087
rect 2498 12084 2504 12096
rect 2179 12056 2504 12084
rect 2179 12053 2191 12056
rect 2133 12047 2191 12053
rect 2498 12044 2504 12056
rect 2556 12084 2562 12096
rect 2958 12084 2964 12096
rect 2556 12056 2964 12084
rect 2556 12044 2562 12056
rect 2958 12044 2964 12056
rect 3016 12044 3022 12096
rect 3237 12087 3295 12093
rect 3237 12053 3249 12087
rect 3283 12084 3295 12087
rect 3510 12084 3516 12096
rect 3283 12056 3516 12084
rect 3283 12053 3295 12056
rect 3237 12047 3295 12053
rect 3510 12044 3516 12056
rect 3568 12084 3574 12096
rect 4065 12087 4123 12093
rect 4065 12084 4077 12087
rect 3568 12056 4077 12084
rect 3568 12044 3574 12056
rect 4065 12053 4077 12056
rect 4111 12053 4123 12087
rect 4065 12047 4123 12053
rect 5166 12044 5172 12096
rect 5224 12084 5230 12096
rect 5534 12084 5540 12096
rect 5224 12056 5540 12084
rect 5224 12044 5230 12056
rect 5534 12044 5540 12056
rect 5592 12084 5598 12096
rect 5629 12087 5687 12093
rect 5629 12084 5641 12087
rect 5592 12056 5641 12084
rect 5592 12044 5598 12056
rect 5629 12053 5641 12056
rect 5675 12053 5687 12087
rect 5629 12047 5687 12053
rect 7190 12044 7196 12096
rect 7248 12084 7254 12096
rect 8205 12087 8263 12093
rect 8205 12084 8217 12087
rect 7248 12056 8217 12084
rect 7248 12044 7254 12056
rect 8205 12053 8217 12056
rect 8251 12053 8263 12087
rect 8205 12047 8263 12053
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 10502 12084 10508 12096
rect 9732 12056 10508 12084
rect 9732 12044 9738 12056
rect 10502 12044 10508 12056
rect 10560 12044 10566 12096
rect 10962 12044 10968 12096
rect 11020 12084 11026 12096
rect 12161 12087 12219 12093
rect 12161 12084 12173 12087
rect 11020 12056 12173 12084
rect 11020 12044 11026 12056
rect 12161 12053 12173 12056
rect 12207 12053 12219 12087
rect 12161 12047 12219 12053
rect 1104 11994 14812 12016
rect 1104 11942 3648 11994
rect 3700 11942 3712 11994
rect 3764 11942 3776 11994
rect 3828 11942 3840 11994
rect 3892 11942 8982 11994
rect 9034 11942 9046 11994
rect 9098 11942 9110 11994
rect 9162 11942 9174 11994
rect 9226 11942 14315 11994
rect 14367 11942 14379 11994
rect 14431 11942 14443 11994
rect 14495 11942 14507 11994
rect 14559 11942 14812 11994
rect 1104 11920 14812 11942
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 3145 11883 3203 11889
rect 3145 11880 3157 11883
rect 3016 11852 3157 11880
rect 3016 11840 3022 11852
rect 3145 11849 3157 11852
rect 3191 11849 3203 11883
rect 3145 11843 3203 11849
rect 4338 11840 4344 11892
rect 4396 11880 4402 11892
rect 4614 11880 4620 11892
rect 4396 11852 4620 11880
rect 4396 11840 4402 11852
rect 4614 11840 4620 11852
rect 4672 11840 4678 11892
rect 5721 11883 5779 11889
rect 5721 11849 5733 11883
rect 5767 11880 5779 11883
rect 5810 11880 5816 11892
rect 5767 11852 5816 11880
rect 5767 11849 5779 11852
rect 5721 11843 5779 11849
rect 5810 11840 5816 11852
rect 5868 11840 5874 11892
rect 6914 11880 6920 11892
rect 6875 11852 6920 11880
rect 6914 11840 6920 11852
rect 6972 11840 6978 11892
rect 3053 11815 3111 11821
rect 3053 11781 3065 11815
rect 3099 11812 3111 11815
rect 3234 11812 3240 11824
rect 3099 11784 3240 11812
rect 3099 11781 3111 11784
rect 3053 11775 3111 11781
rect 3234 11772 3240 11784
rect 3292 11812 3298 11824
rect 3292 11784 3740 11812
rect 3292 11772 3298 11784
rect 3712 11753 3740 11784
rect 10502 11772 10508 11824
rect 10560 11812 10566 11824
rect 10781 11815 10839 11821
rect 10781 11812 10793 11815
rect 10560 11784 10793 11812
rect 10560 11772 10566 11784
rect 10781 11781 10793 11784
rect 10827 11781 10839 11815
rect 10781 11775 10839 11781
rect 10870 11772 10876 11824
rect 10928 11812 10934 11824
rect 12161 11815 12219 11821
rect 12161 11812 12173 11815
rect 10928 11784 12173 11812
rect 10928 11772 10934 11784
rect 12161 11781 12173 11784
rect 12207 11781 12219 11815
rect 12161 11775 12219 11781
rect 3697 11747 3755 11753
rect 3697 11713 3709 11747
rect 3743 11713 3755 11747
rect 3697 11707 3755 11713
rect 5626 11704 5632 11756
rect 5684 11744 5690 11756
rect 6178 11744 6184 11756
rect 5684 11716 6184 11744
rect 5684 11704 5690 11716
rect 6178 11704 6184 11716
rect 6236 11704 6242 11756
rect 7282 11704 7288 11756
rect 7340 11744 7346 11756
rect 7469 11747 7527 11753
rect 7469 11744 7481 11747
rect 7340 11716 7481 11744
rect 7340 11704 7346 11716
rect 7469 11713 7481 11716
rect 7515 11713 7527 11747
rect 7469 11707 7527 11713
rect 8481 11747 8539 11753
rect 8481 11713 8493 11747
rect 8527 11744 8539 11747
rect 8527 11716 8708 11744
rect 8527 11713 8539 11716
rect 8481 11707 8539 11713
rect 3510 11676 3516 11688
rect 3471 11648 3516 11676
rect 3510 11636 3516 11648
rect 3568 11636 3574 11688
rect 6273 11679 6331 11685
rect 6273 11645 6285 11679
rect 6319 11676 6331 11679
rect 7374 11676 7380 11688
rect 6319 11648 7380 11676
rect 6319 11645 6331 11648
rect 6273 11639 6331 11645
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 7558 11636 7564 11688
rect 7616 11676 7622 11688
rect 8294 11676 8300 11688
rect 7616 11648 8300 11676
rect 7616 11636 7622 11648
rect 8294 11636 8300 11648
rect 8352 11636 8358 11688
rect 8570 11676 8576 11688
rect 8531 11648 8576 11676
rect 8570 11636 8576 11648
rect 8628 11636 8634 11688
rect 8680 11676 8708 11716
rect 10042 11704 10048 11756
rect 10100 11744 10106 11756
rect 11241 11747 11299 11753
rect 11241 11744 11253 11747
rect 10100 11716 11253 11744
rect 10100 11704 10106 11716
rect 11241 11713 11253 11716
rect 11287 11713 11299 11747
rect 11241 11707 11299 11713
rect 11330 11704 11336 11756
rect 11388 11744 11394 11756
rect 11425 11747 11483 11753
rect 11425 11744 11437 11747
rect 11388 11716 11437 11744
rect 11388 11704 11394 11716
rect 11425 11713 11437 11716
rect 11471 11744 11483 11747
rect 11471 11716 11928 11744
rect 11471 11713 11483 11716
rect 11425 11707 11483 11713
rect 8840 11679 8898 11685
rect 8840 11676 8852 11679
rect 8680 11648 8852 11676
rect 8840 11645 8852 11648
rect 8886 11676 8898 11679
rect 10318 11676 10324 11688
rect 8886 11648 10324 11676
rect 8886 11645 8898 11648
rect 8840 11639 8898 11645
rect 10318 11636 10324 11648
rect 10376 11636 10382 11688
rect 7282 11608 7288 11620
rect 7195 11580 7288 11608
rect 7282 11568 7288 11580
rect 7340 11608 7346 11620
rect 7929 11611 7987 11617
rect 7929 11608 7941 11611
rect 7340 11580 7941 11608
rect 7340 11568 7346 11580
rect 7929 11577 7941 11580
rect 7975 11577 7987 11611
rect 7929 11571 7987 11577
rect 10689 11611 10747 11617
rect 10689 11577 10701 11611
rect 10735 11608 10747 11611
rect 11146 11608 11152 11620
rect 10735 11580 11152 11608
rect 10735 11577 10747 11580
rect 10689 11571 10747 11577
rect 11146 11568 11152 11580
rect 11204 11608 11210 11620
rect 11514 11608 11520 11620
rect 11204 11580 11520 11608
rect 11204 11568 11210 11580
rect 11514 11568 11520 11580
rect 11572 11568 11578 11620
rect 3602 11500 3608 11552
rect 3660 11540 3666 11552
rect 4249 11543 4307 11549
rect 3660 11512 3705 11540
rect 3660 11500 3666 11512
rect 4249 11509 4261 11543
rect 4295 11540 4307 11543
rect 4614 11540 4620 11552
rect 4295 11512 4620 11540
rect 4295 11509 4307 11512
rect 4249 11503 4307 11509
rect 4614 11500 4620 11512
rect 4672 11500 4678 11552
rect 4890 11540 4896 11552
rect 4851 11512 4896 11540
rect 4890 11500 4896 11512
rect 4948 11500 4954 11552
rect 6641 11543 6699 11549
rect 6641 11509 6653 11543
rect 6687 11540 6699 11543
rect 7006 11540 7012 11552
rect 6687 11512 7012 11540
rect 6687 11509 6699 11512
rect 6641 11503 6699 11509
rect 7006 11500 7012 11512
rect 7064 11540 7070 11552
rect 7834 11540 7840 11552
rect 7064 11512 7840 11540
rect 7064 11500 7070 11512
rect 7834 11500 7840 11512
rect 7892 11500 7898 11552
rect 9953 11543 10011 11549
rect 9953 11509 9965 11543
rect 9999 11540 10011 11543
rect 10134 11540 10140 11552
rect 9999 11512 10140 11540
rect 9999 11509 10011 11512
rect 9953 11503 10011 11509
rect 10134 11500 10140 11512
rect 10192 11500 10198 11552
rect 10318 11540 10324 11552
rect 10279 11512 10324 11540
rect 10318 11500 10324 11512
rect 10376 11500 10382 11552
rect 11900 11549 11928 11716
rect 11885 11543 11943 11549
rect 11885 11509 11897 11543
rect 11931 11540 11943 11543
rect 11974 11540 11980 11552
rect 11931 11512 11980 11540
rect 11931 11509 11943 11512
rect 11885 11503 11943 11509
rect 11974 11500 11980 11512
rect 12032 11500 12038 11552
rect 1104 11450 14812 11472
rect 1104 11398 6315 11450
rect 6367 11398 6379 11450
rect 6431 11398 6443 11450
rect 6495 11398 6507 11450
rect 6559 11398 11648 11450
rect 11700 11398 11712 11450
rect 11764 11398 11776 11450
rect 11828 11398 11840 11450
rect 11892 11398 14812 11450
rect 1104 11376 14812 11398
rect 2774 11296 2780 11348
rect 2832 11336 2838 11348
rect 3237 11339 3295 11345
rect 3237 11336 3249 11339
rect 2832 11308 3249 11336
rect 2832 11296 2838 11308
rect 3237 11305 3249 11308
rect 3283 11336 3295 11339
rect 3602 11336 3608 11348
rect 3283 11308 3608 11336
rect 3283 11305 3295 11308
rect 3237 11299 3295 11305
rect 3602 11296 3608 11308
rect 3660 11296 3666 11348
rect 6641 11339 6699 11345
rect 6641 11305 6653 11339
rect 6687 11336 6699 11339
rect 6822 11336 6828 11348
rect 6687 11308 6828 11336
rect 6687 11305 6699 11308
rect 6641 11299 6699 11305
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 7282 11336 7288 11348
rect 7243 11308 7288 11336
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 7466 11296 7472 11348
rect 7524 11336 7530 11348
rect 7745 11339 7803 11345
rect 7745 11336 7757 11339
rect 7524 11308 7757 11336
rect 7524 11296 7530 11308
rect 7745 11305 7757 11308
rect 7791 11305 7803 11339
rect 7745 11299 7803 11305
rect 8478 11296 8484 11348
rect 8536 11336 8542 11348
rect 9398 11336 9404 11348
rect 8536 11308 9404 11336
rect 8536 11296 8542 11308
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 9493 11339 9551 11345
rect 9493 11305 9505 11339
rect 9539 11336 9551 11339
rect 9582 11336 9588 11348
rect 9539 11308 9588 11336
rect 9539 11305 9551 11308
rect 9493 11299 9551 11305
rect 9582 11296 9588 11308
rect 9640 11296 9646 11348
rect 9766 11296 9772 11348
rect 9824 11336 9830 11348
rect 10042 11336 10048 11348
rect 9824 11308 10048 11336
rect 9824 11296 9830 11308
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 11054 11296 11060 11348
rect 11112 11336 11118 11348
rect 11241 11339 11299 11345
rect 11241 11336 11253 11339
rect 11112 11308 11253 11336
rect 11112 11296 11118 11308
rect 11241 11305 11253 11308
rect 11287 11305 11299 11339
rect 11241 11299 11299 11305
rect 7009 11271 7067 11277
rect 7009 11237 7021 11271
rect 7055 11268 7067 11271
rect 7190 11268 7196 11280
rect 7055 11240 7196 11268
rect 7055 11237 7067 11240
rect 7009 11231 7067 11237
rect 7190 11228 7196 11240
rect 7248 11228 7254 11280
rect 8386 11268 8392 11280
rect 8299 11240 8392 11268
rect 8386 11228 8392 11240
rect 8444 11268 8450 11280
rect 10134 11268 10140 11280
rect 8444 11240 10140 11268
rect 8444 11228 8450 11240
rect 10134 11228 10140 11240
rect 10192 11228 10198 11280
rect 10873 11271 10931 11277
rect 10873 11237 10885 11271
rect 10919 11268 10931 11271
rect 11146 11268 11152 11280
rect 10919 11240 11152 11268
rect 10919 11237 10931 11240
rect 10873 11231 10931 11237
rect 11146 11228 11152 11240
rect 11204 11228 11210 11280
rect 7558 11160 7564 11212
rect 7616 11200 7622 11212
rect 7653 11203 7711 11209
rect 7653 11200 7665 11203
rect 7616 11172 7665 11200
rect 7616 11160 7622 11172
rect 7653 11169 7665 11172
rect 7699 11200 7711 11203
rect 7742 11200 7748 11212
rect 7699 11172 7748 11200
rect 7699 11169 7711 11172
rect 7653 11163 7711 11169
rect 7742 11160 7748 11172
rect 7800 11160 7806 11212
rect 7834 11160 7840 11212
rect 7892 11200 7898 11212
rect 8294 11200 8300 11212
rect 7892 11172 8300 11200
rect 7892 11160 7898 11172
rect 8294 11160 8300 11172
rect 8352 11200 8358 11212
rect 8665 11203 8723 11209
rect 8665 11200 8677 11203
rect 8352 11172 8677 11200
rect 8352 11160 8358 11172
rect 8665 11169 8677 11172
rect 8711 11169 8723 11203
rect 8665 11163 8723 11169
rect 9398 11160 9404 11212
rect 9456 11200 9462 11212
rect 10045 11203 10103 11209
rect 10045 11200 10057 11203
rect 9456 11172 10057 11200
rect 9456 11160 9462 11172
rect 10045 11169 10057 11172
rect 10091 11169 10103 11203
rect 10152 11200 10180 11228
rect 11609 11203 11667 11209
rect 10152 11172 10272 11200
rect 10045 11163 10103 11169
rect 7926 11132 7932 11144
rect 7887 11104 7932 11132
rect 7926 11092 7932 11104
rect 7984 11092 7990 11144
rect 9306 11092 9312 11144
rect 9364 11132 9370 11144
rect 9766 11132 9772 11144
rect 9364 11104 9772 11132
rect 9364 11092 9370 11104
rect 9766 11092 9772 11104
rect 9824 11132 9830 11144
rect 10244 11141 10272 11172
rect 11609 11169 11621 11203
rect 11655 11200 11667 11203
rect 12342 11200 12348 11212
rect 11655 11172 12348 11200
rect 11655 11169 11667 11172
rect 11609 11163 11667 11169
rect 12342 11160 12348 11172
rect 12400 11200 12406 11212
rect 12434 11200 12440 11212
rect 12400 11172 12440 11200
rect 12400 11160 12406 11172
rect 12434 11160 12440 11172
rect 12492 11160 12498 11212
rect 10137 11135 10195 11141
rect 10137 11132 10149 11135
rect 9824 11104 10149 11132
rect 9824 11092 9830 11104
rect 10137 11101 10149 11104
rect 10183 11101 10195 11135
rect 10137 11095 10195 11101
rect 10229 11135 10287 11141
rect 10229 11101 10241 11135
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 11330 11092 11336 11144
rect 11388 11132 11394 11144
rect 11701 11135 11759 11141
rect 11701 11132 11713 11135
rect 11388 11104 11713 11132
rect 11388 11092 11394 11104
rect 11701 11101 11713 11104
rect 11747 11101 11759 11135
rect 11701 11095 11759 11101
rect 11885 11135 11943 11141
rect 11885 11101 11897 11135
rect 11931 11132 11943 11135
rect 11974 11132 11980 11144
rect 11931 11104 11980 11132
rect 11931 11101 11943 11104
rect 11885 11095 11943 11101
rect 11974 11092 11980 11104
rect 12032 11092 12038 11144
rect 3881 11067 3939 11073
rect 3881 11033 3893 11067
rect 3927 11064 3939 11067
rect 4062 11064 4068 11076
rect 3927 11036 4068 11064
rect 3927 11033 3939 11036
rect 3881 11027 3939 11033
rect 4062 11024 4068 11036
rect 4120 11024 4126 11076
rect 9677 11067 9735 11073
rect 9677 11064 9689 11067
rect 9600 11036 9689 11064
rect 9600 11008 9628 11036
rect 9677 11033 9689 11036
rect 9723 11033 9735 11067
rect 9677 11027 9735 11033
rect 9582 10956 9588 11008
rect 9640 10956 9646 11008
rect 1104 10906 14812 10928
rect 1104 10854 3648 10906
rect 3700 10854 3712 10906
rect 3764 10854 3776 10906
rect 3828 10854 3840 10906
rect 3892 10854 8982 10906
rect 9034 10854 9046 10906
rect 9098 10854 9110 10906
rect 9162 10854 9174 10906
rect 9226 10854 14315 10906
rect 14367 10854 14379 10906
rect 14431 10854 14443 10906
rect 14495 10854 14507 10906
rect 14559 10854 14812 10906
rect 1104 10832 14812 10854
rect 5810 10752 5816 10804
rect 5868 10792 5874 10804
rect 7466 10792 7472 10804
rect 5868 10764 7472 10792
rect 5868 10752 5874 10764
rect 7466 10752 7472 10764
rect 7524 10792 7530 10804
rect 7653 10795 7711 10801
rect 7653 10792 7665 10795
rect 7524 10764 7665 10792
rect 7524 10752 7530 10764
rect 7653 10761 7665 10764
rect 7699 10761 7711 10795
rect 7653 10755 7711 10761
rect 7926 10752 7932 10804
rect 7984 10792 7990 10804
rect 9309 10795 9367 10801
rect 9309 10792 9321 10795
rect 7984 10764 9321 10792
rect 7984 10752 7990 10764
rect 9309 10761 9321 10764
rect 9355 10761 9367 10795
rect 9309 10755 9367 10761
rect 10137 10795 10195 10801
rect 10137 10761 10149 10795
rect 10183 10792 10195 10795
rect 10594 10792 10600 10804
rect 10183 10764 10600 10792
rect 10183 10761 10195 10764
rect 10137 10755 10195 10761
rect 10594 10752 10600 10764
rect 10652 10752 10658 10804
rect 11333 10727 11391 10733
rect 11333 10693 11345 10727
rect 11379 10724 11391 10727
rect 12342 10724 12348 10736
rect 11379 10696 12348 10724
rect 11379 10693 11391 10696
rect 11333 10687 11391 10693
rect 12342 10684 12348 10696
rect 12400 10684 12406 10736
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4341 10659 4399 10665
rect 4341 10656 4353 10659
rect 4212 10628 4353 10656
rect 4212 10616 4218 10628
rect 4341 10625 4353 10628
rect 4387 10625 4399 10659
rect 4341 10619 4399 10625
rect 7834 10616 7840 10668
rect 7892 10656 7898 10668
rect 7929 10659 7987 10665
rect 7929 10656 7941 10659
rect 7892 10628 7941 10656
rect 7892 10616 7898 10628
rect 7929 10625 7941 10628
rect 7975 10625 7987 10659
rect 7929 10619 7987 10625
rect 10781 10659 10839 10665
rect 10781 10625 10793 10659
rect 10827 10656 10839 10659
rect 10962 10656 10968 10668
rect 10827 10628 10968 10656
rect 10827 10625 10839 10628
rect 10781 10619 10839 10625
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 1486 10588 1492 10600
rect 1443 10560 1492 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 1486 10548 1492 10560
rect 1544 10588 1550 10600
rect 2133 10591 2191 10597
rect 2133 10588 2145 10591
rect 1544 10560 2145 10588
rect 1544 10548 1550 10560
rect 2133 10557 2145 10560
rect 2179 10557 2191 10591
rect 2133 10551 2191 10557
rect 3697 10591 3755 10597
rect 3697 10557 3709 10591
rect 3743 10588 3755 10591
rect 4246 10588 4252 10600
rect 3743 10560 4252 10588
rect 3743 10557 3755 10560
rect 3697 10551 3755 10557
rect 4246 10548 4252 10560
rect 4304 10548 4310 10600
rect 3878 10480 3884 10532
rect 3936 10520 3942 10532
rect 4157 10523 4215 10529
rect 4157 10520 4169 10523
rect 3936 10492 4169 10520
rect 3936 10480 3942 10492
rect 4157 10489 4169 10492
rect 4203 10520 4215 10523
rect 4522 10520 4528 10532
rect 4203 10492 4528 10520
rect 4203 10489 4215 10492
rect 4157 10483 4215 10489
rect 4522 10480 4528 10492
rect 4580 10480 4586 10532
rect 2406 10412 2412 10464
rect 2464 10452 2470 10464
rect 3789 10455 3847 10461
rect 3789 10452 3801 10455
rect 2464 10424 3801 10452
rect 2464 10412 2470 10424
rect 3789 10421 3801 10424
rect 3835 10421 3847 10455
rect 3789 10415 3847 10421
rect 6825 10455 6883 10461
rect 6825 10421 6837 10455
rect 6871 10452 6883 10455
rect 6914 10452 6920 10464
rect 6871 10424 6920 10452
rect 6871 10421 6883 10424
rect 6825 10415 6883 10421
rect 6914 10412 6920 10424
rect 6972 10412 6978 10464
rect 7377 10455 7435 10461
rect 7377 10421 7389 10455
rect 7423 10452 7435 10455
rect 7558 10452 7564 10464
rect 7423 10424 7564 10452
rect 7423 10421 7435 10424
rect 7377 10415 7435 10421
rect 7558 10412 7564 10424
rect 7616 10412 7622 10464
rect 7944 10452 7972 10619
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 9674 10548 9680 10600
rect 9732 10548 9738 10600
rect 8196 10523 8254 10529
rect 8196 10489 8208 10523
rect 8242 10520 8254 10523
rect 8386 10520 8392 10532
rect 8242 10492 8392 10520
rect 8242 10489 8254 10492
rect 8196 10483 8254 10489
rect 8386 10480 8392 10492
rect 8444 10480 8450 10532
rect 9692 10520 9720 10548
rect 10962 10520 10968 10532
rect 9692 10492 10968 10520
rect 10962 10480 10968 10492
rect 11020 10480 11026 10532
rect 8110 10452 8116 10464
rect 7944 10424 8116 10452
rect 8110 10412 8116 10424
rect 8168 10412 8174 10464
rect 9674 10452 9680 10464
rect 9635 10424 9680 10452
rect 9674 10412 9680 10424
rect 9732 10412 9738 10464
rect 10502 10452 10508 10464
rect 10463 10424 10508 10452
rect 10502 10412 10508 10424
rect 10560 10412 10566 10464
rect 10594 10412 10600 10464
rect 10652 10452 10658 10464
rect 10652 10424 10697 10452
rect 10652 10412 10658 10424
rect 11330 10412 11336 10464
rect 11388 10452 11394 10464
rect 11609 10455 11667 10461
rect 11609 10452 11621 10455
rect 11388 10424 11621 10452
rect 11388 10412 11394 10424
rect 11609 10421 11621 10424
rect 11655 10421 11667 10455
rect 11974 10452 11980 10464
rect 11935 10424 11980 10452
rect 11609 10415 11667 10421
rect 11974 10412 11980 10424
rect 12032 10412 12038 10464
rect 1104 10362 14812 10384
rect 1104 10310 6315 10362
rect 6367 10310 6379 10362
rect 6431 10310 6443 10362
rect 6495 10310 6507 10362
rect 6559 10310 11648 10362
rect 11700 10310 11712 10362
rect 11764 10310 11776 10362
rect 11828 10310 11840 10362
rect 11892 10310 14812 10362
rect 1104 10288 14812 10310
rect 2406 10248 2412 10260
rect 2367 10220 2412 10248
rect 2406 10208 2412 10220
rect 2464 10208 2470 10260
rect 2498 10208 2504 10260
rect 2556 10248 2562 10260
rect 3878 10248 3884 10260
rect 2556 10220 3884 10248
rect 2556 10208 2562 10220
rect 3878 10208 3884 10220
rect 3936 10208 3942 10260
rect 5810 10248 5816 10260
rect 5771 10220 5816 10248
rect 5810 10208 5816 10220
rect 5868 10208 5874 10260
rect 7374 10208 7380 10260
rect 7432 10248 7438 10260
rect 7469 10251 7527 10257
rect 7469 10248 7481 10251
rect 7432 10220 7481 10248
rect 7432 10208 7438 10220
rect 7469 10217 7481 10220
rect 7515 10217 7527 10251
rect 7469 10211 7527 10217
rect 7929 10251 7987 10257
rect 7929 10217 7941 10251
rect 7975 10248 7987 10251
rect 8573 10251 8631 10257
rect 8573 10248 8585 10251
rect 7975 10220 8585 10248
rect 7975 10217 7987 10220
rect 7929 10211 7987 10217
rect 8573 10217 8585 10220
rect 8619 10248 8631 10251
rect 9582 10248 9588 10260
rect 8619 10220 9588 10248
rect 8619 10217 8631 10220
rect 8573 10211 8631 10217
rect 9582 10208 9588 10220
rect 9640 10208 9646 10260
rect 9769 10251 9827 10257
rect 9769 10217 9781 10251
rect 9815 10248 9827 10251
rect 10594 10248 10600 10260
rect 9815 10220 10600 10248
rect 9815 10217 9827 10220
rect 9769 10211 9827 10217
rect 10594 10208 10600 10220
rect 10652 10248 10658 10260
rect 11517 10251 11575 10257
rect 11517 10248 11529 10251
rect 10652 10220 11529 10248
rect 10652 10208 10658 10220
rect 11517 10217 11529 10220
rect 11563 10217 11575 10251
rect 11517 10211 11575 10217
rect 5721 10183 5779 10189
rect 5721 10149 5733 10183
rect 5767 10180 5779 10183
rect 5902 10180 5908 10192
rect 5767 10152 5908 10180
rect 5767 10149 5779 10152
rect 5721 10143 5779 10149
rect 5902 10140 5908 10152
rect 5960 10140 5966 10192
rect 6917 10183 6975 10189
rect 6917 10149 6929 10183
rect 6963 10180 6975 10183
rect 7190 10180 7196 10192
rect 6963 10152 7196 10180
rect 6963 10149 6975 10152
rect 6917 10143 6975 10149
rect 5258 10044 5264 10056
rect 5171 10016 5264 10044
rect 5258 10004 5264 10016
rect 5316 10044 5322 10056
rect 5997 10047 6055 10053
rect 5997 10044 6009 10047
rect 5316 10016 6009 10044
rect 5316 10004 5322 10016
rect 5997 10013 6009 10016
rect 6043 10044 6055 10047
rect 6932 10044 6960 10143
rect 7190 10140 7196 10152
rect 7248 10180 7254 10192
rect 7650 10180 7656 10192
rect 7248 10152 7656 10180
rect 7248 10140 7254 10152
rect 7650 10140 7656 10152
rect 7708 10140 7714 10192
rect 8386 10140 8392 10192
rect 8444 10180 8450 10192
rect 9033 10183 9091 10189
rect 9033 10180 9045 10183
rect 8444 10152 9045 10180
rect 8444 10140 8450 10152
rect 9033 10149 9045 10152
rect 9079 10149 9091 10183
rect 9033 10143 9091 10149
rect 9950 10140 9956 10192
rect 10008 10140 10014 10192
rect 10502 10140 10508 10192
rect 10560 10180 10566 10192
rect 11885 10183 11943 10189
rect 11885 10180 11897 10183
rect 10560 10152 11897 10180
rect 10560 10140 10566 10152
rect 11885 10149 11897 10152
rect 11931 10149 11943 10183
rect 11885 10143 11943 10149
rect 7098 10072 7104 10124
rect 7156 10112 7162 10124
rect 7742 10112 7748 10124
rect 7156 10084 7748 10112
rect 7156 10072 7162 10084
rect 7742 10072 7748 10084
rect 7800 10112 7806 10124
rect 7837 10115 7895 10121
rect 7837 10112 7849 10115
rect 7800 10084 7849 10112
rect 7800 10072 7806 10084
rect 7837 10081 7849 10084
rect 7883 10081 7895 10115
rect 9968 10112 9996 10140
rect 10134 10112 10140 10124
rect 9968 10084 10140 10112
rect 7837 10075 7895 10081
rect 10134 10072 10140 10084
rect 10192 10072 10198 10124
rect 10229 10115 10287 10121
rect 10229 10081 10241 10115
rect 10275 10112 10287 10115
rect 10275 10084 10732 10112
rect 10275 10081 10287 10084
rect 10229 10075 10287 10081
rect 10704 10056 10732 10084
rect 6043 10016 6960 10044
rect 7377 10047 7435 10053
rect 6043 10013 6055 10016
rect 5997 10007 6055 10013
rect 7377 10013 7389 10047
rect 7423 10044 7435 10047
rect 7926 10044 7932 10056
rect 7423 10016 7932 10044
rect 7423 10013 7435 10016
rect 7377 10007 7435 10013
rect 7926 10004 7932 10016
rect 7984 10044 7990 10056
rect 8113 10047 8171 10053
rect 8113 10044 8125 10047
rect 7984 10016 8125 10044
rect 7984 10004 7990 10016
rect 8113 10013 8125 10016
rect 8159 10044 8171 10047
rect 8294 10044 8300 10056
rect 8159 10016 8300 10044
rect 8159 10013 8171 10016
rect 8113 10007 8171 10013
rect 8294 10004 8300 10016
rect 8352 10004 8358 10056
rect 9950 10004 9956 10056
rect 10008 10044 10014 10056
rect 10318 10044 10324 10056
rect 10008 10016 10324 10044
rect 10008 10004 10014 10016
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 10686 10004 10692 10056
rect 10744 10004 10750 10056
rect 4614 9936 4620 9988
rect 4672 9976 4678 9988
rect 9306 9976 9312 9988
rect 4672 9948 9312 9976
rect 4672 9936 4678 9948
rect 9306 9936 9312 9948
rect 9364 9936 9370 9988
rect 10873 9979 10931 9985
rect 10873 9945 10885 9979
rect 10919 9976 10931 9979
rect 10962 9976 10968 9988
rect 10919 9948 10968 9976
rect 10919 9945 10931 9948
rect 10873 9939 10931 9945
rect 10962 9936 10968 9948
rect 11020 9976 11026 9988
rect 11422 9976 11428 9988
rect 11020 9948 11428 9976
rect 11020 9936 11026 9948
rect 11422 9936 11428 9948
rect 11480 9936 11486 9988
rect 5353 9911 5411 9917
rect 5353 9877 5365 9911
rect 5399 9908 5411 9911
rect 5534 9908 5540 9920
rect 5399 9880 5540 9908
rect 5399 9877 5411 9880
rect 5353 9871 5411 9877
rect 5534 9868 5540 9880
rect 5592 9868 5598 9920
rect 8478 9868 8484 9920
rect 8536 9908 8542 9920
rect 9398 9908 9404 9920
rect 8536 9880 9404 9908
rect 8536 9868 8542 9880
rect 9398 9868 9404 9880
rect 9456 9868 9462 9920
rect 11238 9908 11244 9920
rect 11199 9880 11244 9908
rect 11238 9868 11244 9880
rect 11296 9868 11302 9920
rect 1104 9818 14812 9840
rect 1104 9766 3648 9818
rect 3700 9766 3712 9818
rect 3764 9766 3776 9818
rect 3828 9766 3840 9818
rect 3892 9766 8982 9818
rect 9034 9766 9046 9818
rect 9098 9766 9110 9818
rect 9162 9766 9174 9818
rect 9226 9766 14315 9818
rect 14367 9766 14379 9818
rect 14431 9766 14443 9818
rect 14495 9766 14507 9818
rect 14559 9766 14812 9818
rect 1104 9744 14812 9766
rect 5810 9664 5816 9716
rect 5868 9704 5874 9716
rect 5905 9707 5963 9713
rect 5905 9704 5917 9707
rect 5868 9676 5917 9704
rect 5868 9664 5874 9676
rect 5905 9673 5917 9676
rect 5951 9673 5963 9707
rect 5905 9667 5963 9673
rect 7742 9664 7748 9716
rect 7800 9704 7806 9716
rect 7837 9707 7895 9713
rect 7837 9704 7849 9707
rect 7800 9676 7849 9704
rect 7800 9664 7806 9676
rect 7837 9673 7849 9676
rect 7883 9673 7895 9707
rect 7837 9667 7895 9673
rect 9398 9664 9404 9716
rect 9456 9704 9462 9716
rect 11146 9704 11152 9716
rect 9456 9676 11152 9704
rect 9456 9664 9462 9676
rect 11146 9664 11152 9676
rect 11204 9664 11210 9716
rect 2317 9639 2375 9645
rect 2317 9605 2329 9639
rect 2363 9636 2375 9639
rect 2682 9636 2688 9648
rect 2363 9608 2688 9636
rect 2363 9605 2375 9608
rect 2317 9599 2375 9605
rect 2682 9596 2688 9608
rect 2740 9596 2746 9648
rect 5994 9596 6000 9648
rect 6052 9636 6058 9648
rect 7098 9636 7104 9648
rect 6052 9608 7104 9636
rect 6052 9596 6058 9608
rect 7098 9596 7104 9608
rect 7156 9596 7162 9648
rect 7190 9596 7196 9648
rect 7248 9636 7254 9648
rect 9861 9639 9919 9645
rect 7248 9608 7512 9636
rect 7248 9596 7254 9608
rect 2406 9528 2412 9580
rect 2464 9568 2470 9580
rect 2777 9571 2835 9577
rect 2777 9568 2789 9571
rect 2464 9540 2789 9568
rect 2464 9528 2470 9540
rect 2777 9537 2789 9540
rect 2823 9537 2835 9571
rect 2777 9531 2835 9537
rect 2869 9571 2927 9577
rect 2869 9537 2881 9571
rect 2915 9537 2927 9571
rect 2869 9531 2927 9537
rect 2590 9460 2596 9512
rect 2648 9500 2654 9512
rect 2884 9500 2912 9531
rect 3418 9528 3424 9580
rect 3476 9568 3482 9580
rect 7484 9577 7512 9608
rect 9861 9605 9873 9639
rect 9907 9636 9919 9639
rect 9907 9608 11284 9636
rect 9907 9605 9919 9608
rect 9861 9599 9919 9605
rect 11256 9580 11284 9608
rect 12158 9596 12164 9648
rect 12216 9636 12222 9648
rect 12986 9636 12992 9648
rect 12216 9608 12992 9636
rect 12216 9596 12222 9608
rect 12986 9596 12992 9608
rect 13044 9596 13050 9648
rect 3881 9571 3939 9577
rect 3881 9568 3893 9571
rect 3476 9540 3893 9568
rect 3476 9528 3482 9540
rect 3881 9537 3893 9540
rect 3927 9537 3939 9571
rect 3881 9531 3939 9537
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9568 7527 9571
rect 7926 9568 7932 9580
rect 7515 9540 7932 9568
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 7926 9528 7932 9540
rect 7984 9528 7990 9580
rect 8110 9528 8116 9580
rect 8168 9568 8174 9580
rect 8386 9568 8392 9580
rect 8168 9540 8392 9568
rect 8168 9528 8174 9540
rect 8386 9528 8392 9540
rect 8444 9568 8450 9580
rect 8481 9571 8539 9577
rect 8481 9568 8493 9571
rect 8444 9540 8493 9568
rect 8444 9528 8450 9540
rect 8481 9537 8493 9540
rect 8527 9537 8539 9571
rect 8481 9531 8539 9537
rect 9674 9528 9680 9580
rect 9732 9568 9738 9580
rect 10134 9568 10140 9580
rect 9732 9540 10140 9568
rect 9732 9528 9738 9540
rect 10134 9528 10140 9540
rect 10192 9528 10198 9580
rect 10502 9568 10508 9580
rect 10463 9540 10508 9568
rect 10502 9528 10508 9540
rect 10560 9528 10566 9580
rect 11238 9568 11244 9580
rect 11199 9540 11244 9568
rect 11238 9528 11244 9540
rect 11296 9528 11302 9580
rect 2648 9472 3740 9500
rect 2648 9460 2654 9472
rect 2225 9367 2283 9373
rect 2225 9333 2237 9367
rect 2271 9364 2283 9367
rect 2682 9364 2688 9376
rect 2271 9336 2688 9364
rect 2271 9333 2283 9336
rect 2225 9327 2283 9333
rect 2682 9324 2688 9336
rect 2740 9324 2746 9376
rect 3418 9364 3424 9376
rect 3379 9336 3424 9364
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 3712 9364 3740 9472
rect 6638 9460 6644 9512
rect 6696 9460 6702 9512
rect 6914 9460 6920 9512
rect 6972 9500 6978 9512
rect 7193 9503 7251 9509
rect 7193 9500 7205 9503
rect 6972 9472 7205 9500
rect 6972 9460 6978 9472
rect 7193 9469 7205 9472
rect 7239 9469 7251 9503
rect 10520 9500 10548 9528
rect 11149 9503 11207 9509
rect 11149 9500 11161 9503
rect 10520 9472 11161 9500
rect 7193 9463 7251 9469
rect 11149 9469 11161 9472
rect 11195 9469 11207 9503
rect 11149 9463 11207 9469
rect 3789 9435 3847 9441
rect 3789 9401 3801 9435
rect 3835 9432 3847 9435
rect 4062 9432 4068 9444
rect 3835 9404 4068 9432
rect 3835 9401 3847 9404
rect 3789 9395 3847 9401
rect 4062 9392 4068 9404
rect 4120 9441 4126 9444
rect 4120 9435 4184 9441
rect 4120 9401 4138 9435
rect 4172 9432 4184 9435
rect 6656 9432 6684 9460
rect 7285 9435 7343 9441
rect 7285 9432 7297 9435
rect 4172 9404 4213 9432
rect 6564 9404 7297 9432
rect 4172 9401 4184 9404
rect 4120 9395 4184 9401
rect 4120 9392 4126 9395
rect 4890 9364 4896 9376
rect 3712 9336 4896 9364
rect 4890 9324 4896 9336
rect 4948 9364 4954 9376
rect 5261 9367 5319 9373
rect 5261 9364 5273 9367
rect 4948 9336 5273 9364
rect 4948 9324 4954 9336
rect 5261 9333 5273 9336
rect 5307 9333 5319 9367
rect 5261 9327 5319 9333
rect 5629 9367 5687 9373
rect 5629 9333 5641 9367
rect 5675 9364 5687 9367
rect 5902 9364 5908 9376
rect 5675 9336 5908 9364
rect 5675 9333 5687 9336
rect 5629 9327 5687 9333
rect 5902 9324 5908 9336
rect 5960 9324 5966 9376
rect 5994 9324 6000 9376
rect 6052 9364 6058 9376
rect 6564 9373 6592 9404
rect 7285 9401 7297 9404
rect 7331 9401 7343 9435
rect 7285 9395 7343 9401
rect 8389 9435 8447 9441
rect 8389 9401 8401 9435
rect 8435 9432 8447 9435
rect 8662 9432 8668 9444
rect 8435 9404 8668 9432
rect 8435 9401 8447 9404
rect 8389 9395 8447 9401
rect 8662 9392 8668 9404
rect 8720 9441 8726 9444
rect 8720 9435 8784 9441
rect 8720 9401 8738 9435
rect 8772 9401 8784 9435
rect 8720 9395 8784 9401
rect 11057 9435 11115 9441
rect 11057 9401 11069 9435
rect 11103 9432 11115 9435
rect 11422 9432 11428 9444
rect 11103 9404 11428 9432
rect 11103 9401 11115 9404
rect 11057 9395 11115 9401
rect 8720 9392 8726 9395
rect 11422 9392 11428 9404
rect 11480 9392 11486 9444
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 6052 9336 6561 9364
rect 6052 9324 6058 9336
rect 6549 9333 6561 9336
rect 6595 9333 6607 9367
rect 6549 9327 6607 9333
rect 6638 9324 6644 9376
rect 6696 9364 6702 9376
rect 6825 9367 6883 9373
rect 6825 9364 6837 9367
rect 6696 9336 6837 9364
rect 6696 9324 6702 9336
rect 6825 9333 6837 9336
rect 6871 9333 6883 9367
rect 10686 9364 10692 9376
rect 10647 9336 10692 9364
rect 6825 9327 6883 9333
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 1104 9274 14812 9296
rect 1104 9222 6315 9274
rect 6367 9222 6379 9274
rect 6431 9222 6443 9274
rect 6495 9222 6507 9274
rect 6559 9222 11648 9274
rect 11700 9222 11712 9274
rect 11764 9222 11776 9274
rect 11828 9222 11840 9274
rect 11892 9222 14812 9274
rect 1104 9200 14812 9222
rect 2409 9163 2467 9169
rect 2409 9129 2421 9163
rect 2455 9160 2467 9163
rect 2590 9160 2596 9172
rect 2455 9132 2596 9160
rect 2455 9129 2467 9132
rect 2409 9123 2467 9129
rect 2590 9120 2596 9132
rect 2648 9120 2654 9172
rect 6914 9160 6920 9172
rect 6875 9132 6920 9160
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 7742 9160 7748 9172
rect 7703 9132 7748 9160
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 8294 9160 8300 9172
rect 8255 9132 8300 9160
rect 8294 9120 8300 9132
rect 8352 9120 8358 9172
rect 9493 9163 9551 9169
rect 9493 9129 9505 9163
rect 9539 9160 9551 9163
rect 10686 9160 10692 9172
rect 9539 9132 10692 9160
rect 9539 9129 9551 9132
rect 9493 9123 9551 9129
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 11609 9163 11667 9169
rect 11609 9129 11621 9163
rect 11655 9160 11667 9163
rect 11974 9160 11980 9172
rect 11655 9132 11980 9160
rect 11655 9129 11667 9132
rect 11609 9123 11667 9129
rect 5258 9052 5264 9104
rect 5316 9101 5322 9104
rect 5316 9095 5380 9101
rect 5316 9061 5334 9095
rect 5368 9061 5380 9095
rect 5316 9055 5380 9061
rect 5316 9052 5322 9055
rect 5442 9052 5448 9104
rect 5500 9052 5506 9104
rect 9950 9092 9956 9104
rect 9911 9064 9956 9092
rect 9950 9052 9956 9064
rect 10008 9052 10014 9104
rect 10496 9095 10554 9101
rect 10496 9061 10508 9095
rect 10542 9092 10554 9095
rect 10962 9092 10968 9104
rect 10542 9064 10968 9092
rect 10542 9061 10554 9064
rect 10496 9055 10554 9061
rect 10962 9052 10968 9064
rect 11020 9092 11026 9104
rect 11146 9092 11152 9104
rect 11020 9064 11152 9092
rect 11020 9052 11026 9064
rect 11146 9052 11152 9064
rect 11204 9052 11210 9104
rect 5460 9024 5488 9052
rect 5092 8996 5488 9024
rect 5092 8965 5120 8996
rect 7098 8984 7104 9036
rect 7156 9024 7162 9036
rect 7653 9027 7711 9033
rect 7653 9024 7665 9027
rect 7156 8996 7665 9024
rect 7156 8984 7162 8996
rect 7653 8993 7665 8996
rect 7699 8993 7711 9027
rect 9968 9024 9996 9052
rect 11624 9024 11652 9123
rect 11974 9120 11980 9132
rect 12032 9120 12038 9172
rect 9968 8996 11652 9024
rect 7653 8987 7711 8993
rect 5077 8959 5135 8965
rect 5077 8956 5089 8959
rect 4908 8928 5089 8956
rect 2866 8780 2872 8832
rect 2924 8820 2930 8832
rect 3418 8820 3424 8832
rect 2924 8792 3424 8820
rect 2924 8780 2930 8792
rect 3418 8780 3424 8792
rect 3476 8820 3482 8832
rect 4908 8829 4936 8928
rect 5077 8925 5089 8928
rect 5123 8925 5135 8959
rect 7926 8956 7932 8968
rect 7887 8928 7932 8956
rect 5077 8919 5135 8925
rect 7926 8916 7932 8928
rect 7984 8916 7990 8968
rect 10229 8959 10287 8965
rect 10229 8925 10241 8959
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 4893 8823 4951 8829
rect 4893 8820 4905 8823
rect 3476 8792 4905 8820
rect 3476 8780 3482 8792
rect 4893 8789 4905 8792
rect 4939 8789 4951 8823
rect 6454 8820 6460 8832
rect 6415 8792 6460 8820
rect 4893 8783 4951 8789
rect 6454 8780 6460 8792
rect 6512 8780 6518 8832
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 7285 8823 7343 8829
rect 7285 8820 7297 8823
rect 6972 8792 7297 8820
rect 6972 8780 6978 8792
rect 7285 8789 7297 8792
rect 7331 8789 7343 8823
rect 7285 8783 7343 8789
rect 8386 8780 8392 8832
rect 8444 8820 8450 8832
rect 8665 8823 8723 8829
rect 8665 8820 8677 8823
rect 8444 8792 8677 8820
rect 8444 8780 8450 8792
rect 8665 8789 8677 8792
rect 8711 8789 8723 8823
rect 10244 8820 10272 8919
rect 10870 8820 10876 8832
rect 10244 8792 10876 8820
rect 8665 8783 8723 8789
rect 10870 8780 10876 8792
rect 10928 8820 10934 8832
rect 11146 8820 11152 8832
rect 10928 8792 11152 8820
rect 10928 8780 10934 8792
rect 11146 8780 11152 8792
rect 11204 8780 11210 8832
rect 1104 8730 14812 8752
rect 1104 8678 3648 8730
rect 3700 8678 3712 8730
rect 3764 8678 3776 8730
rect 3828 8678 3840 8730
rect 3892 8678 8982 8730
rect 9034 8678 9046 8730
rect 9098 8678 9110 8730
rect 9162 8678 9174 8730
rect 9226 8678 14315 8730
rect 14367 8678 14379 8730
rect 14431 8678 14443 8730
rect 14495 8678 14507 8730
rect 14559 8678 14812 8730
rect 1104 8656 14812 8678
rect 4062 8576 4068 8628
rect 4120 8616 4126 8628
rect 4157 8619 4215 8625
rect 4157 8616 4169 8619
rect 4120 8588 4169 8616
rect 4120 8576 4126 8588
rect 4157 8585 4169 8588
rect 4203 8585 4215 8619
rect 4157 8579 4215 8585
rect 5077 8619 5135 8625
rect 5077 8585 5089 8619
rect 5123 8616 5135 8619
rect 5258 8616 5264 8628
rect 5123 8588 5264 8616
rect 5123 8585 5135 8588
rect 5077 8579 5135 8585
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 6641 8619 6699 8625
rect 6641 8585 6653 8619
rect 6687 8616 6699 8619
rect 7098 8616 7104 8628
rect 6687 8588 7104 8616
rect 6687 8585 6699 8588
rect 6641 8579 6699 8585
rect 7098 8576 7104 8588
rect 7156 8576 7162 8628
rect 7926 8576 7932 8628
rect 7984 8616 7990 8628
rect 8481 8619 8539 8625
rect 8481 8616 8493 8619
rect 7984 8588 8493 8616
rect 7984 8576 7990 8588
rect 8481 8585 8493 8588
rect 8527 8585 8539 8619
rect 8481 8579 8539 8585
rect 10781 8619 10839 8625
rect 10781 8585 10793 8619
rect 10827 8616 10839 8619
rect 10962 8616 10968 8628
rect 10827 8588 10968 8616
rect 10827 8585 10839 8588
rect 10781 8579 10839 8585
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 6178 8508 6184 8560
rect 6236 8508 6242 8560
rect 8202 8548 8208 8560
rect 8163 8520 8208 8548
rect 8202 8508 8208 8520
rect 8260 8548 8266 8560
rect 8849 8551 8907 8557
rect 8849 8548 8861 8551
rect 8260 8520 8861 8548
rect 8260 8508 8266 8520
rect 8849 8517 8861 8520
rect 8895 8517 8907 8551
rect 8849 8511 8907 8517
rect 10413 8551 10471 8557
rect 10413 8517 10425 8551
rect 10459 8517 10471 8551
rect 10413 8511 10471 8517
rect 1578 8480 1584 8492
rect 1539 8452 1584 8480
rect 1578 8440 1584 8452
rect 1636 8440 1642 8492
rect 4709 8483 4767 8489
rect 4709 8449 4721 8483
rect 4755 8480 4767 8483
rect 5629 8483 5687 8489
rect 5629 8480 5641 8483
rect 4755 8452 5641 8480
rect 4755 8449 4767 8452
rect 4709 8443 4767 8449
rect 5629 8449 5641 8452
rect 5675 8480 5687 8483
rect 5718 8480 5724 8492
rect 5675 8452 5724 8480
rect 5675 8449 5687 8452
rect 5629 8443 5687 8449
rect 5718 8440 5724 8452
rect 5776 8440 5782 8492
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 6196 8480 6224 8508
rect 6454 8480 6460 8492
rect 5859 8452 6460 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 6454 8440 6460 8452
rect 6512 8480 6518 8492
rect 8864 8480 8892 8511
rect 10428 8480 10456 8511
rect 10962 8480 10968 8492
rect 6512 8452 6960 8480
rect 8864 8452 9168 8480
rect 10428 8452 10968 8480
rect 6512 8440 6518 8452
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 2777 8415 2835 8421
rect 1443 8384 2268 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 2240 8285 2268 8384
rect 2777 8381 2789 8415
rect 2823 8412 2835 8415
rect 2866 8412 2872 8424
rect 2823 8384 2872 8412
rect 2823 8381 2835 8384
rect 2777 8375 2835 8381
rect 2866 8372 2872 8384
rect 2924 8372 2930 8424
rect 5534 8412 5540 8424
rect 5495 8384 5540 8412
rect 5534 8372 5540 8384
rect 5592 8412 5598 8424
rect 6181 8415 6239 8421
rect 6181 8412 6193 8415
rect 5592 8384 6193 8412
rect 5592 8372 5598 8384
rect 6181 8381 6193 8384
rect 6227 8381 6239 8415
rect 6181 8375 6239 8381
rect 6825 8415 6883 8421
rect 6825 8381 6837 8415
rect 6871 8381 6883 8415
rect 6932 8412 6960 8452
rect 7081 8415 7139 8421
rect 7081 8412 7093 8415
rect 6932 8384 7093 8412
rect 6825 8375 6883 8381
rect 7081 8381 7093 8384
rect 7127 8381 7139 8415
rect 9030 8412 9036 8424
rect 8991 8384 9036 8412
rect 7081 8375 7139 8381
rect 2682 8344 2688 8356
rect 2643 8316 2688 8344
rect 2682 8304 2688 8316
rect 2740 8344 2746 8356
rect 3022 8347 3080 8353
rect 3022 8344 3034 8347
rect 2740 8316 3034 8344
rect 2740 8304 2746 8316
rect 3022 8313 3034 8316
rect 3068 8313 3080 8347
rect 6840 8344 6868 8375
rect 9030 8372 9036 8384
rect 9088 8372 9094 8424
rect 9140 8412 9168 8452
rect 10962 8440 10968 8452
rect 11020 8440 11026 8492
rect 9289 8415 9347 8421
rect 9289 8412 9301 8415
rect 9140 8384 9301 8412
rect 9289 8381 9301 8384
rect 9335 8381 9347 8415
rect 9289 8375 9347 8381
rect 8386 8344 8392 8356
rect 6840 8316 8392 8344
rect 3022 8307 3080 8313
rect 8386 8304 8392 8316
rect 8444 8304 8450 8356
rect 2225 8279 2283 8285
rect 2225 8245 2237 8279
rect 2271 8276 2283 8279
rect 2774 8276 2780 8288
rect 2271 8248 2780 8276
rect 2271 8245 2283 8248
rect 2225 8239 2283 8245
rect 2774 8236 2780 8248
rect 2832 8236 2838 8288
rect 5166 8276 5172 8288
rect 5127 8248 5172 8276
rect 5166 8236 5172 8248
rect 5224 8236 5230 8288
rect 11146 8276 11152 8288
rect 11107 8248 11152 8276
rect 11146 8236 11152 8248
rect 11204 8236 11210 8288
rect 1104 8186 14812 8208
rect 1104 8134 6315 8186
rect 6367 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 11648 8186
rect 11700 8134 11712 8186
rect 11764 8134 11776 8186
rect 11828 8134 11840 8186
rect 11892 8134 14812 8186
rect 1104 8112 14812 8134
rect 2225 8075 2283 8081
rect 2225 8041 2237 8075
rect 2271 8072 2283 8075
rect 2866 8072 2872 8084
rect 2271 8044 2872 8072
rect 2271 8041 2283 8044
rect 2225 8035 2283 8041
rect 2866 8032 2872 8044
rect 2924 8032 2930 8084
rect 5718 8032 5724 8084
rect 5776 8072 5782 8084
rect 6089 8075 6147 8081
rect 6089 8072 6101 8075
rect 5776 8044 6101 8072
rect 5776 8032 5782 8044
rect 6089 8041 6101 8044
rect 6135 8072 6147 8075
rect 6822 8072 6828 8084
rect 6135 8044 6828 8072
rect 6135 8041 6147 8044
rect 6089 8035 6147 8041
rect 6822 8032 6828 8044
rect 6880 8032 6886 8084
rect 7742 8072 7748 8084
rect 7703 8044 7748 8072
rect 7742 8032 7748 8044
rect 7800 8032 7806 8084
rect 10870 8032 10876 8084
rect 10928 8072 10934 8084
rect 11422 8072 11428 8084
rect 10928 8044 11428 8072
rect 10928 8032 10934 8044
rect 11422 8032 11428 8044
rect 11480 8032 11486 8084
rect 4522 7964 4528 8016
rect 4580 8004 4586 8016
rect 5997 8007 6055 8013
rect 5997 8004 6009 8007
rect 4580 7976 6009 8004
rect 4580 7964 4586 7976
rect 5997 7973 6009 7976
rect 6043 8004 6055 8007
rect 6638 8004 6644 8016
rect 6043 7976 6644 8004
rect 6043 7973 6055 7976
rect 5997 7967 6055 7973
rect 6638 7964 6644 7976
rect 6696 7964 6702 8016
rect 6730 7964 6736 8016
rect 6788 8004 6794 8016
rect 7760 8004 7788 8032
rect 6788 7976 7788 8004
rect 6788 7964 6794 7976
rect 7190 7936 7196 7948
rect 7151 7908 7196 7936
rect 7190 7896 7196 7908
rect 7248 7896 7254 7948
rect 11422 7945 11428 7948
rect 11416 7899 11428 7945
rect 11480 7936 11486 7948
rect 11480 7908 11516 7936
rect 11422 7896 11428 7899
rect 11480 7896 11486 7908
rect 4614 7868 4620 7880
rect 4575 7840 4620 7868
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 6178 7828 6184 7880
rect 6236 7868 6242 7880
rect 6825 7871 6883 7877
rect 6825 7868 6837 7871
rect 6236 7840 6837 7868
rect 6236 7828 6242 7840
rect 6825 7837 6837 7840
rect 6871 7837 6883 7871
rect 8386 7868 8392 7880
rect 6825 7831 6883 7837
rect 8128 7840 8392 7868
rect 5261 7803 5319 7809
rect 5261 7769 5273 7803
rect 5307 7800 5319 7803
rect 6196 7800 6224 7828
rect 5307 7772 6224 7800
rect 5307 7769 5319 7772
rect 5261 7763 5319 7769
rect 8128 7744 8156 7840
rect 8386 7828 8392 7840
rect 8444 7868 8450 7880
rect 9030 7868 9036 7880
rect 8444 7840 9036 7868
rect 8444 7828 8450 7840
rect 9030 7828 9036 7840
rect 9088 7828 9094 7880
rect 11146 7868 11152 7880
rect 11107 7840 11152 7868
rect 11146 7828 11152 7840
rect 11204 7828 11210 7880
rect 1670 7732 1676 7744
rect 1631 7704 1676 7732
rect 1670 7692 1676 7704
rect 1728 7692 1734 7744
rect 2866 7732 2872 7744
rect 2827 7704 2872 7732
rect 2866 7692 2872 7704
rect 2924 7692 2930 7744
rect 5626 7732 5632 7744
rect 5587 7704 5632 7732
rect 5626 7692 5632 7704
rect 5684 7692 5690 7744
rect 6914 7692 6920 7744
rect 6972 7732 6978 7744
rect 7377 7735 7435 7741
rect 7377 7732 7389 7735
rect 6972 7704 7389 7732
rect 6972 7692 6978 7704
rect 7377 7701 7389 7704
rect 7423 7701 7435 7735
rect 8110 7732 8116 7744
rect 8071 7704 8116 7732
rect 7377 7695 7435 7701
rect 8110 7692 8116 7704
rect 8168 7692 8174 7744
rect 12434 7692 12440 7744
rect 12492 7732 12498 7744
rect 12529 7735 12587 7741
rect 12529 7732 12541 7735
rect 12492 7704 12541 7732
rect 12492 7692 12498 7704
rect 12529 7701 12541 7704
rect 12575 7701 12587 7735
rect 12529 7695 12587 7701
rect 1104 7642 14812 7664
rect 1104 7590 3648 7642
rect 3700 7590 3712 7642
rect 3764 7590 3776 7642
rect 3828 7590 3840 7642
rect 3892 7590 8982 7642
rect 9034 7590 9046 7642
rect 9098 7590 9110 7642
rect 9162 7590 9174 7642
rect 9226 7590 14315 7642
rect 14367 7590 14379 7642
rect 14431 7590 14443 7642
rect 14495 7590 14507 7642
rect 14559 7590 14812 7642
rect 1104 7568 14812 7590
rect 2038 7488 2044 7540
rect 2096 7528 2102 7540
rect 2133 7531 2191 7537
rect 2133 7528 2145 7531
rect 2096 7500 2145 7528
rect 2096 7488 2102 7500
rect 2133 7497 2145 7500
rect 2179 7497 2191 7531
rect 2133 7491 2191 7497
rect 2593 7531 2651 7537
rect 2593 7497 2605 7531
rect 2639 7528 2651 7531
rect 2866 7528 2872 7540
rect 2639 7500 2872 7528
rect 2639 7497 2651 7500
rect 2593 7491 2651 7497
rect 2866 7488 2872 7500
rect 2924 7528 2930 7540
rect 3510 7528 3516 7540
rect 2924 7500 3516 7528
rect 2924 7488 2930 7500
rect 3510 7488 3516 7500
rect 3568 7488 3574 7540
rect 4522 7528 4528 7540
rect 4483 7500 4528 7528
rect 4522 7488 4528 7500
rect 4580 7488 4586 7540
rect 4893 7531 4951 7537
rect 4893 7497 4905 7531
rect 4939 7528 4951 7531
rect 5442 7528 5448 7540
rect 4939 7500 5448 7528
rect 4939 7497 4951 7500
rect 4893 7491 4951 7497
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 6089 7531 6147 7537
rect 6089 7497 6101 7531
rect 6135 7528 6147 7531
rect 6178 7528 6184 7540
rect 6135 7500 6184 7528
rect 6135 7497 6147 7500
rect 6089 7491 6147 7497
rect 6178 7488 6184 7500
rect 6236 7488 6242 7540
rect 7190 7528 7196 7540
rect 7151 7500 7196 7528
rect 7190 7488 7196 7500
rect 7248 7488 7254 7540
rect 8662 7528 8668 7540
rect 8623 7500 8668 7528
rect 8662 7488 8668 7500
rect 8720 7488 8726 7540
rect 11241 7531 11299 7537
rect 11241 7497 11253 7531
rect 11287 7528 11299 7531
rect 11422 7528 11428 7540
rect 11287 7500 11428 7528
rect 11287 7497 11299 7500
rect 11241 7491 11299 7497
rect 11422 7488 11428 7500
rect 11480 7488 11486 7540
rect 3329 7463 3387 7469
rect 3329 7429 3341 7463
rect 3375 7460 3387 7463
rect 4338 7460 4344 7472
rect 3375 7432 4344 7460
rect 3375 7429 3387 7432
rect 3329 7423 3387 7429
rect 1578 7392 1584 7404
rect 1539 7364 1584 7392
rect 1578 7352 1584 7364
rect 1636 7352 1642 7404
rect 3344 7392 3372 7423
rect 4338 7420 4344 7432
rect 4396 7420 4402 7472
rect 4982 7460 4988 7472
rect 4943 7432 4988 7460
rect 4982 7420 4988 7432
rect 5040 7420 5046 7472
rect 5460 7460 5488 7488
rect 5460 7432 5580 7460
rect 2700 7364 3372 7392
rect 4157 7395 4215 7401
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7324 1455 7327
rect 1670 7324 1676 7336
rect 1443 7296 1676 7324
rect 1443 7293 1455 7296
rect 1397 7287 1455 7293
rect 1670 7284 1676 7296
rect 1728 7284 1734 7336
rect 2700 7333 2728 7364
rect 4157 7361 4169 7395
rect 4203 7392 4215 7395
rect 5166 7392 5172 7404
rect 4203 7364 5172 7392
rect 4203 7361 4215 7364
rect 4157 7355 4215 7361
rect 5166 7352 5172 7364
rect 5224 7392 5230 7404
rect 5552 7401 5580 7432
rect 5445 7395 5503 7401
rect 5445 7392 5457 7395
rect 5224 7364 5457 7392
rect 5224 7352 5230 7364
rect 5445 7361 5457 7364
rect 5491 7361 5503 7395
rect 5445 7355 5503 7361
rect 5537 7395 5595 7401
rect 5537 7361 5549 7395
rect 5583 7361 5595 7395
rect 5537 7355 5595 7361
rect 2685 7327 2743 7333
rect 2685 7293 2697 7327
rect 2731 7293 2743 7327
rect 2685 7287 2743 7293
rect 5353 7327 5411 7333
rect 5353 7293 5365 7327
rect 5399 7324 5411 7327
rect 5626 7324 5632 7336
rect 5399 7296 5632 7324
rect 5399 7293 5411 7296
rect 5353 7287 5411 7293
rect 5626 7284 5632 7296
rect 5684 7284 5690 7336
rect 7285 7327 7343 7333
rect 7285 7293 7297 7327
rect 7331 7324 7343 7327
rect 8110 7324 8116 7336
rect 7331 7296 8116 7324
rect 7331 7293 7343 7296
rect 7285 7287 7343 7293
rect 8110 7284 8116 7296
rect 8168 7284 8174 7336
rect 6641 7259 6699 7265
rect 6641 7225 6653 7259
rect 6687 7256 6699 7259
rect 7552 7259 7610 7265
rect 7552 7256 7564 7259
rect 6687 7228 7564 7256
rect 6687 7225 6699 7228
rect 6641 7219 6699 7225
rect 7552 7225 7564 7228
rect 7598 7256 7610 7259
rect 7834 7256 7840 7268
rect 7598 7228 7840 7256
rect 7598 7225 7610 7228
rect 7552 7219 7610 7225
rect 7834 7216 7840 7228
rect 7892 7216 7898 7268
rect 2866 7188 2872 7200
rect 2827 7160 2872 7188
rect 2866 7148 2872 7160
rect 2924 7148 2930 7200
rect 8110 7148 8116 7200
rect 8168 7188 8174 7200
rect 8941 7191 8999 7197
rect 8941 7188 8953 7191
rect 8168 7160 8953 7188
rect 8168 7148 8174 7160
rect 8941 7157 8953 7160
rect 8987 7188 8999 7191
rect 9674 7188 9680 7200
rect 8987 7160 9680 7188
rect 8987 7157 8999 7160
rect 8941 7151 8999 7157
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 11609 7191 11667 7197
rect 11609 7157 11621 7191
rect 11655 7188 11667 7191
rect 12066 7188 12072 7200
rect 11655 7160 12072 7188
rect 11655 7157 11667 7160
rect 11609 7151 11667 7157
rect 12066 7148 12072 7160
rect 12124 7148 12130 7200
rect 1104 7098 14812 7120
rect 1104 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 11648 7098
rect 11700 7046 11712 7098
rect 11764 7046 11776 7098
rect 11828 7046 11840 7098
rect 11892 7046 14812 7098
rect 1104 7024 14812 7046
rect 4893 6987 4951 6993
rect 4893 6953 4905 6987
rect 4939 6984 4951 6987
rect 5626 6984 5632 6996
rect 4939 6956 5632 6984
rect 4939 6953 4951 6956
rect 4893 6947 4951 6953
rect 5626 6944 5632 6956
rect 5684 6944 5690 6996
rect 5718 6944 5724 6996
rect 5776 6984 5782 6996
rect 5776 6956 5821 6984
rect 5776 6944 5782 6956
rect 11146 6944 11152 6996
rect 11204 6944 11210 6996
rect 11422 6944 11428 6996
rect 11480 6984 11486 6996
rect 12345 6987 12403 6993
rect 12345 6984 12357 6987
rect 11480 6956 12357 6984
rect 11480 6944 11486 6956
rect 12345 6953 12357 6956
rect 12391 6953 12403 6987
rect 12345 6947 12403 6953
rect 8662 6916 8668 6928
rect 7576 6888 8668 6916
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 2130 6848 2136 6860
rect 1443 6820 2136 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 2130 6808 2136 6820
rect 2188 6808 2194 6860
rect 2498 6808 2504 6860
rect 2556 6848 2562 6860
rect 2685 6851 2743 6857
rect 2685 6848 2697 6851
rect 2556 6820 2697 6848
rect 2556 6808 2562 6820
rect 2685 6817 2697 6820
rect 2731 6817 2743 6851
rect 2685 6811 2743 6817
rect 4985 6851 5043 6857
rect 4985 6817 4997 6851
rect 5031 6848 5043 6851
rect 5350 6848 5356 6860
rect 5031 6820 5356 6848
rect 5031 6817 5043 6820
rect 4985 6811 5043 6817
rect 5350 6808 5356 6820
rect 5408 6848 5414 6860
rect 5626 6848 5632 6860
rect 5408 6820 5632 6848
rect 5408 6808 5414 6820
rect 5626 6808 5632 6820
rect 5684 6808 5690 6860
rect 5994 6808 6000 6860
rect 6052 6848 6058 6860
rect 6089 6851 6147 6857
rect 6089 6848 6101 6851
rect 6052 6820 6101 6848
rect 6052 6808 6058 6820
rect 6089 6817 6101 6820
rect 6135 6848 6147 6851
rect 6270 6848 6276 6860
rect 6135 6820 6276 6848
rect 6135 6817 6147 6820
rect 6089 6811 6147 6817
rect 6270 6808 6276 6820
rect 6328 6808 6334 6860
rect 6917 6851 6975 6857
rect 6917 6817 6929 6851
rect 6963 6848 6975 6851
rect 7466 6848 7472 6860
rect 6963 6820 7472 6848
rect 6963 6817 6975 6820
rect 6917 6811 6975 6817
rect 7466 6808 7472 6820
rect 7524 6848 7530 6860
rect 7576 6848 7604 6888
rect 8662 6876 8668 6888
rect 8720 6876 8726 6928
rect 11164 6916 11192 6944
rect 12066 6916 12072 6928
rect 10980 6888 12072 6916
rect 7524 6820 7604 6848
rect 7653 6851 7711 6857
rect 7524 6808 7530 6820
rect 7653 6817 7665 6851
rect 7699 6848 7711 6851
rect 7926 6848 7932 6860
rect 7699 6820 7932 6848
rect 7699 6817 7711 6820
rect 7653 6811 7711 6817
rect 7926 6808 7932 6820
rect 7984 6848 7990 6860
rect 9033 6851 9091 6857
rect 9033 6848 9045 6851
rect 7984 6820 9045 6848
rect 7984 6808 7990 6820
rect 9033 6817 9045 6820
rect 9079 6817 9091 6851
rect 9033 6811 9091 6817
rect 9677 6851 9735 6857
rect 9677 6817 9689 6851
rect 9723 6848 9735 6851
rect 9766 6848 9772 6860
rect 9723 6820 9772 6848
rect 9723 6817 9735 6820
rect 9677 6811 9735 6817
rect 9766 6808 9772 6820
rect 9824 6848 9830 6860
rect 10778 6848 10784 6860
rect 9824 6820 10784 6848
rect 9824 6808 9830 6820
rect 10778 6808 10784 6820
rect 10836 6808 10842 6860
rect 10980 6857 11008 6888
rect 12066 6876 12072 6888
rect 12124 6876 12130 6928
rect 10965 6851 11023 6857
rect 10965 6817 10977 6851
rect 11011 6817 11023 6851
rect 10965 6811 11023 6817
rect 11054 6808 11060 6860
rect 11112 6848 11118 6860
rect 11221 6851 11279 6857
rect 11221 6848 11233 6851
rect 11112 6820 11233 6848
rect 11112 6808 11118 6820
rect 11221 6817 11233 6820
rect 11267 6817 11279 6851
rect 11221 6811 11279 6817
rect 1578 6780 1584 6792
rect 1539 6752 1584 6780
rect 1578 6740 1584 6752
rect 1636 6740 1642 6792
rect 7742 6780 7748 6792
rect 7703 6752 7748 6780
rect 7742 6740 7748 6752
rect 7800 6740 7806 6792
rect 7834 6740 7840 6792
rect 7892 6780 7898 6792
rect 8113 6783 8171 6789
rect 7892 6752 7937 6780
rect 7892 6740 7898 6752
rect 8113 6749 8125 6783
rect 8159 6780 8171 6783
rect 8665 6783 8723 6789
rect 8665 6780 8677 6783
rect 8159 6752 8677 6780
rect 8159 6749 8171 6752
rect 8113 6743 8171 6749
rect 8665 6749 8677 6752
rect 8711 6749 8723 6783
rect 8665 6743 8723 6749
rect 7282 6712 7288 6724
rect 7195 6684 7288 6712
rect 7282 6672 7288 6684
rect 7340 6712 7346 6724
rect 9401 6715 9459 6721
rect 9401 6712 9413 6715
rect 7340 6684 9413 6712
rect 7340 6672 7346 6684
rect 9401 6681 9413 6684
rect 9447 6681 9459 6715
rect 9401 6675 9459 6681
rect 9674 6672 9680 6724
rect 9732 6712 9738 6724
rect 10229 6715 10287 6721
rect 10229 6712 10241 6715
rect 9732 6684 10241 6712
rect 9732 6672 9738 6684
rect 10229 6681 10241 6684
rect 10275 6681 10287 6715
rect 10229 6675 10287 6681
rect 2406 6644 2412 6656
rect 2367 6616 2412 6644
rect 2406 6604 2412 6616
rect 2464 6604 2470 6656
rect 2866 6644 2872 6656
rect 2827 6616 2872 6644
rect 2866 6604 2872 6616
rect 2924 6604 2930 6656
rect 3326 6644 3332 6656
rect 3287 6616 3332 6644
rect 3326 6604 3332 6616
rect 3384 6604 3390 6656
rect 3510 6604 3516 6656
rect 3568 6644 3574 6656
rect 3881 6647 3939 6653
rect 3881 6644 3893 6647
rect 3568 6616 3893 6644
rect 3568 6604 3574 6616
rect 3881 6613 3893 6616
rect 3927 6644 3939 6647
rect 4341 6647 4399 6653
rect 4341 6644 4353 6647
rect 3927 6616 4353 6644
rect 3927 6613 3939 6616
rect 3881 6607 3939 6613
rect 4341 6613 4353 6616
rect 4387 6644 4399 6647
rect 4798 6644 4804 6656
rect 4387 6616 4804 6644
rect 4387 6613 4399 6616
rect 4341 6607 4399 6613
rect 4798 6604 4804 6616
rect 4856 6604 4862 6656
rect 5169 6647 5227 6653
rect 5169 6613 5181 6647
rect 5215 6644 5227 6647
rect 5350 6644 5356 6656
rect 5215 6616 5356 6644
rect 5215 6613 5227 6616
rect 5169 6607 5227 6613
rect 5350 6604 5356 6616
rect 5408 6604 5414 6656
rect 5718 6604 5724 6656
rect 5776 6644 5782 6656
rect 6273 6647 6331 6653
rect 6273 6644 6285 6647
rect 5776 6616 6285 6644
rect 5776 6604 5782 6616
rect 6273 6613 6285 6616
rect 6319 6613 6331 6647
rect 6273 6607 6331 6613
rect 7742 6604 7748 6656
rect 7800 6644 7806 6656
rect 8113 6647 8171 6653
rect 8113 6644 8125 6647
rect 7800 6616 8125 6644
rect 7800 6604 7806 6616
rect 8113 6613 8125 6616
rect 8159 6613 8171 6647
rect 8294 6644 8300 6656
rect 8255 6616 8300 6644
rect 8113 6607 8171 6613
rect 8294 6604 8300 6616
rect 8352 6604 8358 6656
rect 9858 6644 9864 6656
rect 9819 6616 9864 6644
rect 9858 6604 9864 6616
rect 9916 6604 9922 6656
rect 1104 6554 14812 6576
rect 1104 6502 3648 6554
rect 3700 6502 3712 6554
rect 3764 6502 3776 6554
rect 3828 6502 3840 6554
rect 3892 6502 8982 6554
rect 9034 6502 9046 6554
rect 9098 6502 9110 6554
rect 9162 6502 9174 6554
rect 9226 6502 14315 6554
rect 14367 6502 14379 6554
rect 14431 6502 14443 6554
rect 14495 6502 14507 6554
rect 14559 6502 14812 6554
rect 1104 6480 14812 6502
rect 2041 6443 2099 6449
rect 2041 6409 2053 6443
rect 2087 6440 2099 6443
rect 2498 6440 2504 6452
rect 2087 6412 2504 6440
rect 2087 6409 2099 6412
rect 2041 6403 2099 6409
rect 2498 6400 2504 6412
rect 2556 6400 2562 6452
rect 5169 6443 5227 6449
rect 5169 6409 5181 6443
rect 5215 6440 5227 6443
rect 5442 6440 5448 6452
rect 5215 6412 5448 6440
rect 5215 6409 5227 6412
rect 5169 6403 5227 6409
rect 4154 6332 4160 6384
rect 4212 6372 4218 6384
rect 4709 6375 4767 6381
rect 4709 6372 4721 6375
rect 4212 6344 4721 6372
rect 4212 6332 4218 6344
rect 4709 6341 4721 6344
rect 4755 6341 4767 6375
rect 4709 6335 4767 6341
rect 2133 6239 2191 6245
rect 2133 6205 2145 6239
rect 2179 6236 2191 6239
rect 3510 6236 3516 6248
rect 2179 6208 3516 6236
rect 2179 6205 2191 6208
rect 2133 6199 2191 6205
rect 3510 6196 3516 6208
rect 3568 6196 3574 6248
rect 4525 6239 4583 6245
rect 4525 6205 4537 6239
rect 4571 6236 4583 6239
rect 5184 6236 5212 6403
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 5537 6443 5595 6449
rect 5537 6409 5549 6443
rect 5583 6440 5595 6443
rect 5626 6440 5632 6452
rect 5583 6412 5632 6440
rect 5583 6409 5595 6412
rect 5537 6403 5595 6409
rect 5626 6400 5632 6412
rect 5684 6400 5690 6452
rect 6822 6440 6828 6452
rect 6783 6412 6828 6440
rect 6822 6400 6828 6412
rect 6880 6400 6886 6452
rect 9033 6443 9091 6449
rect 9033 6409 9045 6443
rect 9079 6440 9091 6443
rect 9490 6440 9496 6452
rect 9079 6412 9496 6440
rect 9079 6409 9091 6412
rect 9033 6403 9091 6409
rect 6273 6375 6331 6381
rect 6273 6341 6285 6375
rect 6319 6372 6331 6375
rect 7006 6372 7012 6384
rect 6319 6344 7012 6372
rect 6319 6341 6331 6344
rect 6273 6335 6331 6341
rect 6288 6304 6316 6335
rect 7006 6332 7012 6344
rect 7064 6332 7070 6384
rect 7282 6304 7288 6316
rect 5644 6276 6316 6304
rect 7243 6276 7288 6304
rect 5644 6245 5672 6276
rect 7282 6264 7288 6276
rect 7340 6264 7346 6316
rect 7466 6304 7472 6316
rect 7427 6276 7472 6304
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 4571 6208 5212 6236
rect 5629 6239 5687 6245
rect 4571 6205 4583 6208
rect 4525 6199 4583 6205
rect 5629 6205 5641 6239
rect 5675 6205 5687 6239
rect 5629 6199 5687 6205
rect 5902 6196 5908 6248
rect 5960 6236 5966 6248
rect 6086 6236 6092 6248
rect 5960 6208 6092 6236
rect 5960 6196 5966 6208
rect 6086 6196 6092 6208
rect 6144 6196 6150 6248
rect 6178 6196 6184 6248
rect 6236 6236 6242 6248
rect 7193 6239 7251 6245
rect 7193 6236 7205 6239
rect 6236 6208 7205 6236
rect 6236 6196 6242 6208
rect 7193 6205 7205 6208
rect 7239 6205 7251 6239
rect 7193 6199 7251 6205
rect 8389 6239 8447 6245
rect 8389 6205 8401 6239
rect 8435 6236 8447 6239
rect 9048 6236 9076 6403
rect 9490 6400 9496 6412
rect 9548 6400 9554 6452
rect 9766 6440 9772 6452
rect 9727 6412 9772 6440
rect 9766 6400 9772 6412
rect 9824 6400 9830 6452
rect 11054 6400 11060 6452
rect 11112 6440 11118 6452
rect 11609 6443 11667 6449
rect 11609 6440 11621 6443
rect 11112 6412 11621 6440
rect 11112 6400 11118 6412
rect 11609 6409 11621 6412
rect 11655 6409 11667 6443
rect 11609 6403 11667 6409
rect 9674 6264 9680 6316
rect 9732 6304 9738 6316
rect 9953 6307 10011 6313
rect 9953 6304 9965 6307
rect 9732 6276 9965 6304
rect 9732 6264 9738 6276
rect 9953 6273 9965 6276
rect 9999 6273 10011 6307
rect 9953 6267 10011 6273
rect 8435 6208 9076 6236
rect 8435 6205 8447 6208
rect 8389 6199 8447 6205
rect 2222 6128 2228 6180
rect 2280 6168 2286 6180
rect 2378 6171 2436 6177
rect 2378 6168 2390 6171
rect 2280 6140 2390 6168
rect 2280 6128 2286 6140
rect 2378 6137 2390 6140
rect 2424 6137 2436 6171
rect 2378 6131 2436 6137
rect 4430 6128 4436 6180
rect 4488 6168 4494 6180
rect 5166 6168 5172 6180
rect 4488 6140 5172 6168
rect 4488 6128 4494 6140
rect 5166 6128 5172 6140
rect 5224 6128 5230 6180
rect 6270 6128 6276 6180
rect 6328 6168 6334 6180
rect 9398 6168 9404 6180
rect 6328 6140 6684 6168
rect 9311 6140 9404 6168
rect 6328 6128 6334 6140
rect 1670 6100 1676 6112
rect 1631 6072 1676 6100
rect 1670 6060 1676 6072
rect 1728 6060 1734 6112
rect 2682 6060 2688 6112
rect 2740 6100 2746 6112
rect 3050 6100 3056 6112
rect 2740 6072 3056 6100
rect 2740 6060 2746 6072
rect 3050 6060 3056 6072
rect 3108 6100 3114 6112
rect 3513 6103 3571 6109
rect 3513 6100 3525 6103
rect 3108 6072 3525 6100
rect 3108 6060 3114 6072
rect 3513 6069 3525 6072
rect 3559 6069 3571 6103
rect 4062 6100 4068 6112
rect 4023 6072 4068 6100
rect 3513 6063 3571 6069
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 4338 6100 4344 6112
rect 4299 6072 4344 6100
rect 4338 6060 4344 6072
rect 4396 6060 4402 6112
rect 5810 6100 5816 6112
rect 5771 6072 5816 6100
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 6656 6109 6684 6140
rect 9398 6128 9404 6140
rect 9456 6168 9462 6180
rect 10198 6171 10256 6177
rect 10198 6168 10210 6171
rect 9456 6140 10210 6168
rect 9456 6128 9462 6140
rect 10198 6137 10210 6140
rect 10244 6137 10256 6171
rect 10198 6131 10256 6137
rect 6641 6103 6699 6109
rect 6641 6069 6653 6103
rect 6687 6100 6699 6103
rect 6822 6100 6828 6112
rect 6687 6072 6828 6100
rect 6687 6069 6699 6072
rect 6641 6063 6699 6069
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 7558 6060 7564 6112
rect 7616 6100 7622 6112
rect 7834 6100 7840 6112
rect 7616 6072 7840 6100
rect 7616 6060 7622 6072
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 8297 6103 8355 6109
rect 8297 6069 8309 6103
rect 8343 6100 8355 6103
rect 8386 6100 8392 6112
rect 8343 6072 8392 6100
rect 8343 6069 8355 6072
rect 8297 6063 8355 6069
rect 8386 6060 8392 6072
rect 8444 6060 8450 6112
rect 8478 6060 8484 6112
rect 8536 6100 8542 6112
rect 8573 6103 8631 6109
rect 8573 6100 8585 6103
rect 8536 6072 8585 6100
rect 8536 6060 8542 6072
rect 8573 6069 8585 6072
rect 8619 6069 8631 6103
rect 11330 6100 11336 6112
rect 11291 6072 11336 6100
rect 8573 6063 8631 6069
rect 11330 6060 11336 6072
rect 11388 6060 11394 6112
rect 12066 6100 12072 6112
rect 12027 6072 12072 6100
rect 12066 6060 12072 6072
rect 12124 6060 12130 6112
rect 1104 6010 14812 6032
rect 1104 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 11648 6010
rect 11700 5958 11712 6010
rect 11764 5958 11776 6010
rect 11828 5958 11840 6010
rect 11892 5958 14812 6010
rect 1104 5936 14812 5958
rect 2409 5899 2467 5905
rect 2409 5865 2421 5899
rect 2455 5865 2467 5899
rect 2409 5859 2467 5865
rect 2777 5899 2835 5905
rect 2777 5865 2789 5899
rect 2823 5896 2835 5899
rect 3326 5896 3332 5908
rect 2823 5868 3332 5896
rect 2823 5865 2835 5868
rect 2777 5859 2835 5865
rect 1486 5788 1492 5840
rect 1544 5828 1550 5840
rect 2424 5828 2452 5859
rect 3326 5856 3332 5868
rect 3384 5896 3390 5908
rect 4246 5896 4252 5908
rect 3384 5868 4252 5896
rect 3384 5856 3390 5868
rect 4246 5856 4252 5868
rect 4304 5856 4310 5908
rect 4338 5856 4344 5908
rect 4396 5896 4402 5908
rect 6641 5899 6699 5905
rect 6641 5896 6653 5899
rect 4396 5868 6653 5896
rect 4396 5856 4402 5868
rect 6641 5865 6653 5868
rect 6687 5865 6699 5899
rect 6641 5859 6699 5865
rect 7837 5899 7895 5905
rect 7837 5865 7849 5899
rect 7883 5896 7895 5899
rect 7926 5896 7932 5908
rect 7883 5868 7932 5896
rect 7883 5865 7895 5868
rect 7837 5859 7895 5865
rect 7926 5856 7932 5868
rect 7984 5856 7990 5908
rect 8294 5896 8300 5908
rect 8255 5868 8300 5896
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 8570 5856 8576 5908
rect 8628 5896 8634 5908
rect 8941 5899 8999 5905
rect 8941 5896 8953 5899
rect 8628 5868 8953 5896
rect 8628 5856 8634 5868
rect 8941 5865 8953 5868
rect 8987 5896 8999 5899
rect 9030 5896 9036 5908
rect 8987 5868 9036 5896
rect 8987 5865 8999 5868
rect 8941 5859 8999 5865
rect 9030 5856 9036 5868
rect 9088 5856 9094 5908
rect 11054 5896 11060 5908
rect 11015 5868 11060 5896
rect 11054 5856 11060 5868
rect 11112 5856 11118 5908
rect 11146 5856 11152 5908
rect 11204 5896 11210 5908
rect 11425 5899 11483 5905
rect 11425 5896 11437 5899
rect 11204 5868 11437 5896
rect 11204 5856 11210 5868
rect 11425 5865 11437 5868
rect 11471 5865 11483 5899
rect 11425 5859 11483 5865
rect 5258 5828 5264 5840
rect 1544 5800 5264 5828
rect 1544 5788 1550 5800
rect 5258 5788 5264 5800
rect 5316 5788 5322 5840
rect 5994 5788 6000 5840
rect 6052 5828 6058 5840
rect 6822 5828 6828 5840
rect 6052 5800 6828 5828
rect 6052 5788 6058 5800
rect 6822 5788 6828 5800
rect 6880 5788 6886 5840
rect 8018 5788 8024 5840
rect 8076 5828 8082 5840
rect 8205 5831 8263 5837
rect 8205 5828 8217 5831
rect 8076 5800 8217 5828
rect 8076 5788 8082 5800
rect 8205 5797 8217 5800
rect 8251 5797 8263 5831
rect 8205 5791 8263 5797
rect 9766 5788 9772 5840
rect 9824 5828 9830 5840
rect 9944 5831 10002 5837
rect 9944 5828 9956 5831
rect 9824 5800 9956 5828
rect 9824 5788 9830 5800
rect 9944 5797 9956 5800
rect 9990 5828 10002 5831
rect 11330 5828 11336 5840
rect 9990 5800 11336 5828
rect 9990 5797 10002 5800
rect 9944 5791 10002 5797
rect 11330 5788 11336 5800
rect 11388 5788 11394 5840
rect 1946 5720 1952 5772
rect 2004 5760 2010 5772
rect 2406 5760 2412 5772
rect 2004 5732 2412 5760
rect 2004 5720 2010 5732
rect 2406 5720 2412 5732
rect 2464 5760 2470 5772
rect 4338 5769 4344 5772
rect 2869 5763 2927 5769
rect 2869 5760 2881 5763
rect 2464 5732 2881 5760
rect 2464 5720 2470 5732
rect 2869 5729 2881 5732
rect 2915 5729 2927 5763
rect 2869 5723 2927 5729
rect 3881 5763 3939 5769
rect 3881 5729 3893 5763
rect 3927 5760 3939 5763
rect 4332 5760 4344 5769
rect 3927 5732 4344 5760
rect 3927 5729 3939 5732
rect 3881 5723 3939 5729
rect 4332 5723 4344 5732
rect 4338 5720 4344 5723
rect 4396 5720 4402 5772
rect 6181 5763 6239 5769
rect 6181 5729 6193 5763
rect 6227 5760 6239 5763
rect 9677 5763 9735 5769
rect 6227 5732 6960 5760
rect 6227 5729 6239 5732
rect 6181 5723 6239 5729
rect 3050 5692 3056 5704
rect 3011 5664 3056 5692
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 5813 5695 5871 5701
rect 5813 5661 5825 5695
rect 5859 5692 5871 5695
rect 6730 5692 6736 5704
rect 5859 5664 6736 5692
rect 5859 5661 5871 5664
rect 5813 5655 5871 5661
rect 1854 5556 1860 5568
rect 1815 5528 1860 5556
rect 1854 5516 1860 5528
rect 1912 5516 1918 5568
rect 2222 5556 2228 5568
rect 2183 5528 2228 5556
rect 2222 5516 2228 5528
rect 2280 5516 2286 5568
rect 3510 5556 3516 5568
rect 3471 5528 3516 5556
rect 3510 5516 3516 5528
rect 3568 5516 3574 5568
rect 4080 5556 4108 5655
rect 6730 5652 6736 5664
rect 6788 5652 6794 5704
rect 6932 5701 6960 5732
rect 9677 5729 9689 5763
rect 9723 5760 9735 5763
rect 12066 5760 12072 5772
rect 9723 5732 12072 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 12066 5720 12072 5732
rect 12124 5720 12130 5772
rect 6917 5695 6975 5701
rect 6917 5661 6929 5695
rect 6963 5692 6975 5695
rect 7558 5692 7564 5704
rect 6963 5664 7564 5692
rect 6963 5661 6975 5664
rect 6917 5655 6975 5661
rect 7558 5652 7564 5664
rect 7616 5652 7622 5704
rect 7926 5652 7932 5704
rect 7984 5692 7990 5704
rect 8389 5695 8447 5701
rect 8389 5692 8401 5695
rect 7984 5664 8401 5692
rect 7984 5652 7990 5664
rect 8389 5661 8401 5664
rect 8435 5661 8447 5695
rect 8389 5655 8447 5661
rect 6270 5624 6276 5636
rect 6231 5596 6276 5624
rect 6270 5584 6276 5596
rect 6328 5584 6334 5636
rect 4798 5556 4804 5568
rect 4080 5528 4804 5556
rect 4798 5516 4804 5528
rect 4856 5516 4862 5568
rect 4982 5516 4988 5568
rect 5040 5556 5046 5568
rect 5445 5559 5503 5565
rect 5445 5556 5457 5559
rect 5040 5528 5457 5556
rect 5040 5516 5046 5528
rect 5445 5525 5457 5528
rect 5491 5525 5503 5559
rect 7282 5556 7288 5568
rect 7243 5528 7288 5556
rect 5445 5519 5503 5525
rect 7282 5516 7288 5528
rect 7340 5516 7346 5568
rect 7745 5559 7803 5565
rect 7745 5525 7757 5559
rect 7791 5556 7803 5559
rect 8202 5556 8208 5568
rect 7791 5528 8208 5556
rect 7791 5525 7803 5528
rect 7745 5519 7803 5525
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 9493 5559 9551 5565
rect 9493 5525 9505 5559
rect 9539 5556 9551 5559
rect 9582 5556 9588 5568
rect 9539 5528 9588 5556
rect 9539 5525 9551 5528
rect 9493 5519 9551 5525
rect 9582 5516 9588 5528
rect 9640 5516 9646 5568
rect 1104 5466 14812 5488
rect 1104 5414 3648 5466
rect 3700 5414 3712 5466
rect 3764 5414 3776 5466
rect 3828 5414 3840 5466
rect 3892 5414 8982 5466
rect 9034 5414 9046 5466
rect 9098 5414 9110 5466
rect 9162 5414 9174 5466
rect 9226 5414 14315 5466
rect 14367 5414 14379 5466
rect 14431 5414 14443 5466
rect 14495 5414 14507 5466
rect 14559 5414 14812 5466
rect 1104 5392 14812 5414
rect 1946 5352 1952 5364
rect 1907 5324 1952 5352
rect 1946 5312 1952 5324
rect 2004 5312 2010 5364
rect 3050 5352 3056 5364
rect 3011 5324 3056 5352
rect 3050 5312 3056 5324
rect 3108 5312 3114 5364
rect 4614 5352 4620 5364
rect 4575 5324 4620 5352
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 5534 5312 5540 5364
rect 5592 5352 5598 5364
rect 6181 5355 6239 5361
rect 6181 5352 6193 5355
rect 5592 5324 6193 5352
rect 5592 5312 5598 5324
rect 6181 5321 6193 5324
rect 6227 5352 6239 5355
rect 6457 5355 6515 5361
rect 6457 5352 6469 5355
rect 6227 5324 6469 5352
rect 6227 5321 6239 5324
rect 6181 5315 6239 5321
rect 6457 5321 6469 5324
rect 6503 5321 6515 5355
rect 6457 5315 6515 5321
rect 7929 5355 7987 5361
rect 7929 5321 7941 5355
rect 7975 5352 7987 5355
rect 8018 5352 8024 5364
rect 7975 5324 8024 5352
rect 7975 5321 7987 5324
rect 7929 5315 7987 5321
rect 8018 5312 8024 5324
rect 8076 5312 8082 5364
rect 8294 5312 8300 5364
rect 8352 5352 8358 5364
rect 8389 5355 8447 5361
rect 8389 5352 8401 5355
rect 8352 5324 8401 5352
rect 8352 5312 8358 5324
rect 8389 5321 8401 5324
rect 8435 5321 8447 5355
rect 9766 5352 9772 5364
rect 9727 5324 9772 5352
rect 8389 5315 8447 5321
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 9858 5312 9864 5364
rect 9916 5352 9922 5364
rect 10134 5352 10140 5364
rect 9916 5324 10140 5352
rect 9916 5312 9922 5324
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 10505 5355 10563 5361
rect 10505 5321 10517 5355
rect 10551 5352 10563 5355
rect 10594 5352 10600 5364
rect 10551 5324 10600 5352
rect 10551 5321 10563 5324
rect 10505 5315 10563 5321
rect 10594 5312 10600 5324
rect 10652 5312 10658 5364
rect 12066 5352 12072 5364
rect 12027 5324 12072 5352
rect 12066 5312 12072 5324
rect 12124 5312 12130 5364
rect 1765 5287 1823 5293
rect 1765 5253 1777 5287
rect 1811 5284 1823 5287
rect 2222 5284 2228 5296
rect 1811 5256 2228 5284
rect 1811 5253 1823 5256
rect 1765 5247 1823 5253
rect 2222 5244 2228 5256
rect 2280 5284 2286 5296
rect 4890 5284 4896 5296
rect 2280 5256 4896 5284
rect 2280 5244 2286 5256
rect 1854 5176 1860 5228
rect 1912 5216 1918 5228
rect 2406 5216 2412 5228
rect 1912 5188 2412 5216
rect 1912 5176 1918 5188
rect 2406 5176 2412 5188
rect 2464 5176 2470 5228
rect 2608 5225 2636 5256
rect 4890 5244 4896 5256
rect 4948 5244 4954 5296
rect 5166 5244 5172 5296
rect 5224 5284 5230 5296
rect 6365 5287 6423 5293
rect 6365 5284 6377 5287
rect 5224 5256 6377 5284
rect 5224 5244 5230 5256
rect 6365 5253 6377 5256
rect 6411 5284 6423 5287
rect 6549 5287 6607 5293
rect 6549 5284 6561 5287
rect 6411 5256 6561 5284
rect 6411 5253 6423 5256
rect 6365 5247 6423 5253
rect 6549 5253 6561 5256
rect 6595 5253 6607 5287
rect 6549 5247 6607 5253
rect 2593 5219 2651 5225
rect 2593 5185 2605 5219
rect 2639 5185 2651 5219
rect 2593 5179 2651 5185
rect 3510 5176 3516 5228
rect 3568 5216 3574 5228
rect 3973 5219 4031 5225
rect 3973 5216 3985 5219
rect 3568 5188 3985 5216
rect 3568 5176 3574 5188
rect 3973 5185 3985 5188
rect 4019 5185 4031 5219
rect 3973 5179 4031 5185
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5216 4215 5219
rect 4338 5216 4344 5228
rect 4203 5188 4344 5216
rect 4203 5185 4215 5188
rect 4157 5179 4215 5185
rect 4338 5176 4344 5188
rect 4396 5216 4402 5228
rect 5626 5216 5632 5228
rect 4396 5188 5632 5216
rect 4396 5176 4402 5188
rect 5626 5176 5632 5188
rect 5684 5216 5690 5228
rect 5721 5219 5779 5225
rect 5721 5216 5733 5219
rect 5684 5188 5733 5216
rect 5684 5176 5690 5188
rect 5721 5185 5733 5188
rect 5767 5216 5779 5219
rect 7282 5216 7288 5228
rect 5767 5188 7288 5216
rect 5767 5185 5779 5188
rect 5721 5179 5779 5185
rect 7282 5176 7288 5188
rect 7340 5216 7346 5228
rect 7377 5219 7435 5225
rect 7377 5216 7389 5219
rect 7340 5188 7389 5216
rect 7340 5176 7346 5188
rect 7377 5185 7389 5188
rect 7423 5185 7435 5219
rect 7377 5179 7435 5185
rect 9033 5219 9091 5225
rect 9033 5185 9045 5219
rect 9079 5216 9091 5219
rect 9306 5216 9312 5228
rect 9079 5188 9312 5216
rect 9079 5185 9091 5188
rect 9033 5179 9091 5185
rect 9306 5176 9312 5188
rect 9364 5176 9370 5228
rect 10137 5219 10195 5225
rect 10137 5185 10149 5219
rect 10183 5216 10195 5219
rect 11241 5219 11299 5225
rect 11241 5216 11253 5219
rect 10183 5188 11253 5216
rect 10183 5185 10195 5188
rect 10137 5179 10195 5185
rect 11241 5185 11253 5188
rect 11287 5216 11299 5219
rect 11422 5216 11428 5228
rect 11287 5188 11428 5216
rect 11287 5185 11299 5188
rect 11241 5179 11299 5185
rect 11422 5176 11428 5188
rect 11480 5176 11486 5228
rect 1670 5108 1676 5160
rect 1728 5148 1734 5160
rect 2317 5151 2375 5157
rect 2317 5148 2329 5151
rect 1728 5120 2329 5148
rect 1728 5108 1734 5120
rect 2317 5117 2329 5120
rect 2363 5117 2375 5151
rect 2317 5111 2375 5117
rect 3421 5151 3479 5157
rect 3421 5117 3433 5151
rect 3467 5148 3479 5151
rect 3467 5120 3924 5148
rect 3467 5117 3479 5120
rect 3421 5111 3479 5117
rect 2332 5080 2360 5111
rect 2332 5052 3556 5080
rect 3528 5021 3556 5052
rect 3896 5024 3924 5120
rect 4614 5108 4620 5160
rect 4672 5148 4678 5160
rect 5445 5151 5503 5157
rect 5445 5148 5457 5151
rect 4672 5120 5457 5148
rect 4672 5108 4678 5120
rect 5445 5117 5457 5120
rect 5491 5117 5503 5151
rect 5445 5111 5503 5117
rect 6365 5151 6423 5157
rect 6365 5117 6377 5151
rect 6411 5148 6423 5151
rect 7190 5148 7196 5160
rect 6411 5120 7196 5148
rect 6411 5117 6423 5120
rect 6365 5111 6423 5117
rect 7190 5108 7196 5120
rect 7248 5108 7254 5160
rect 8570 5108 8576 5160
rect 8628 5148 8634 5160
rect 8757 5151 8815 5157
rect 8757 5148 8769 5151
rect 8628 5120 8769 5148
rect 8628 5108 8634 5120
rect 8757 5117 8769 5120
rect 8803 5117 8815 5151
rect 8757 5111 8815 5117
rect 10594 5108 10600 5160
rect 10652 5148 10658 5160
rect 10965 5151 11023 5157
rect 10965 5148 10977 5151
rect 10652 5120 10977 5148
rect 10652 5108 10658 5120
rect 10965 5117 10977 5120
rect 11011 5117 11023 5151
rect 10965 5111 11023 5117
rect 4985 5083 5043 5089
rect 4985 5049 4997 5083
rect 5031 5080 5043 5083
rect 6457 5083 6515 5089
rect 5031 5052 5488 5080
rect 5031 5049 5043 5052
rect 4985 5043 5043 5049
rect 5460 5024 5488 5052
rect 6457 5049 6469 5083
rect 6503 5080 6515 5083
rect 7285 5083 7343 5089
rect 7285 5080 7297 5083
rect 6503 5052 7297 5080
rect 6503 5049 6515 5052
rect 6457 5043 6515 5049
rect 7285 5049 7297 5052
rect 7331 5049 7343 5083
rect 7285 5043 7343 5049
rect 10686 5040 10692 5092
rect 10744 5080 10750 5092
rect 11057 5083 11115 5089
rect 11057 5080 11069 5083
rect 10744 5052 11069 5080
rect 10744 5040 10750 5052
rect 11057 5049 11069 5052
rect 11103 5049 11115 5083
rect 11057 5043 11115 5049
rect 3513 5015 3571 5021
rect 3513 4981 3525 5015
rect 3559 4981 3571 5015
rect 3878 5012 3884 5024
rect 3839 4984 3884 5012
rect 3513 4975 3571 4981
rect 3878 4972 3884 4984
rect 3936 4972 3942 5024
rect 5074 5012 5080 5024
rect 5035 4984 5080 5012
rect 5074 4972 5080 4984
rect 5132 4972 5138 5024
rect 5442 4972 5448 5024
rect 5500 5012 5506 5024
rect 5537 5015 5595 5021
rect 5537 5012 5549 5015
rect 5500 4984 5549 5012
rect 5500 4972 5506 4984
rect 5537 4981 5549 4984
rect 5583 4981 5595 5015
rect 6822 5012 6828 5024
rect 6783 4984 6828 5012
rect 5537 4975 5595 4981
rect 6822 4972 6828 4984
rect 6880 4972 6886 5024
rect 8294 5012 8300 5024
rect 8255 4984 8300 5012
rect 8294 4972 8300 4984
rect 8352 5012 8358 5024
rect 8849 5015 8907 5021
rect 8849 5012 8861 5015
rect 8352 4984 8861 5012
rect 8352 4972 8358 4984
rect 8849 4981 8861 4984
rect 8895 4981 8907 5015
rect 10594 5012 10600 5024
rect 10555 4984 10600 5012
rect 8849 4975 8907 4981
rect 10594 4972 10600 4984
rect 10652 4972 10658 5024
rect 11514 4972 11520 5024
rect 11572 5012 11578 5024
rect 11609 5015 11667 5021
rect 11609 5012 11621 5015
rect 11572 4984 11621 5012
rect 11572 4972 11578 4984
rect 11609 4981 11621 4984
rect 11655 4981 11667 5015
rect 11609 4975 11667 4981
rect 12342 4972 12348 5024
rect 12400 5012 12406 5024
rect 12437 5015 12495 5021
rect 12437 5012 12449 5015
rect 12400 4984 12449 5012
rect 12400 4972 12406 4984
rect 12437 4981 12449 4984
rect 12483 4981 12495 5015
rect 12437 4975 12495 4981
rect 1104 4922 14812 4944
rect 1104 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 11648 4922
rect 11700 4870 11712 4922
rect 11764 4870 11776 4922
rect 11828 4870 11840 4922
rect 11892 4870 14812 4922
rect 1104 4848 14812 4870
rect 4246 4768 4252 4820
rect 4304 4808 4310 4820
rect 4341 4811 4399 4817
rect 4341 4808 4353 4811
rect 4304 4780 4353 4808
rect 4304 4768 4310 4780
rect 4341 4777 4353 4780
rect 4387 4777 4399 4811
rect 4341 4771 4399 4777
rect 4709 4811 4767 4817
rect 4709 4777 4721 4811
rect 4755 4808 4767 4811
rect 5074 4808 5080 4820
rect 4755 4780 5080 4808
rect 4755 4777 4767 4780
rect 4709 4771 4767 4777
rect 5074 4768 5080 4780
rect 5132 4808 5138 4820
rect 5721 4811 5779 4817
rect 5721 4808 5733 4811
rect 5132 4780 5733 4808
rect 5132 4768 5138 4780
rect 5721 4777 5733 4780
rect 5767 4777 5779 4811
rect 7558 4808 7564 4820
rect 7519 4780 7564 4808
rect 5721 4771 5779 4777
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 9033 4811 9091 4817
rect 9033 4777 9045 4811
rect 9079 4808 9091 4811
rect 9306 4808 9312 4820
rect 9079 4780 9312 4808
rect 9079 4777 9091 4780
rect 9033 4771 9091 4777
rect 9306 4768 9312 4780
rect 9364 4768 9370 4820
rect 9674 4768 9680 4820
rect 9732 4808 9738 4820
rect 10045 4811 10103 4817
rect 10045 4808 10057 4811
rect 9732 4780 10057 4808
rect 9732 4768 9738 4780
rect 10045 4777 10057 4780
rect 10091 4777 10103 4811
rect 10045 4771 10103 4777
rect 4801 4743 4859 4749
rect 4801 4709 4813 4743
rect 4847 4740 4859 4743
rect 5534 4740 5540 4752
rect 4847 4712 5540 4740
rect 4847 4709 4859 4712
rect 4801 4703 4859 4709
rect 5534 4700 5540 4712
rect 5592 4740 5598 4752
rect 6822 4740 6828 4752
rect 5592 4712 6828 4740
rect 5592 4700 5598 4712
rect 6822 4700 6828 4712
rect 6880 4700 6886 4752
rect 10060 4740 10088 4771
rect 10594 4768 10600 4820
rect 10652 4808 10658 4820
rect 11057 4811 11115 4817
rect 11057 4808 11069 4811
rect 10652 4780 11069 4808
rect 10652 4768 10658 4780
rect 11057 4777 11069 4780
rect 11103 4777 11115 4811
rect 11057 4771 11115 4777
rect 11241 4811 11299 4817
rect 11241 4777 11253 4811
rect 11287 4777 11299 4811
rect 11241 4771 11299 4777
rect 11256 4740 11284 4771
rect 11514 4768 11520 4820
rect 11572 4808 11578 4820
rect 11609 4811 11667 4817
rect 11609 4808 11621 4811
rect 11572 4780 11621 4808
rect 11572 4768 11578 4780
rect 11609 4777 11621 4780
rect 11655 4777 11667 4811
rect 11609 4771 11667 4777
rect 12158 4768 12164 4820
rect 12216 4808 12222 4820
rect 12437 4811 12495 4817
rect 12437 4808 12449 4811
rect 12216 4780 12449 4808
rect 12216 4768 12222 4780
rect 12437 4777 12449 4780
rect 12483 4808 12495 4811
rect 12618 4808 12624 4820
rect 12483 4780 12624 4808
rect 12483 4777 12495 4780
rect 12437 4771 12495 4777
rect 12618 4768 12624 4780
rect 12676 4768 12682 4820
rect 10060 4712 11284 4740
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4672 1455 4675
rect 1486 4672 1492 4684
rect 1443 4644 1492 4672
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 1486 4632 1492 4644
rect 1544 4632 1550 4684
rect 2314 4632 2320 4684
rect 2372 4672 2378 4684
rect 2685 4675 2743 4681
rect 2685 4672 2697 4675
rect 2372 4644 2697 4672
rect 2372 4632 2378 4644
rect 2685 4641 2697 4644
rect 2731 4641 2743 4675
rect 2685 4635 2743 4641
rect 3050 4632 3056 4684
rect 3108 4672 3114 4684
rect 3605 4675 3663 4681
rect 3605 4672 3617 4675
rect 3108 4644 3617 4672
rect 3108 4632 3114 4644
rect 3605 4641 3617 4644
rect 3651 4672 3663 4675
rect 4338 4672 4344 4684
rect 3651 4644 4344 4672
rect 3651 4641 3663 4644
rect 3605 4635 3663 4641
rect 4338 4632 4344 4644
rect 4396 4632 4402 4684
rect 5442 4672 5448 4684
rect 5355 4644 5448 4672
rect 5442 4632 5448 4644
rect 5500 4672 5506 4684
rect 5626 4672 5632 4684
rect 5500 4644 5632 4672
rect 5500 4632 5506 4644
rect 5626 4632 5632 4644
rect 5684 4632 5690 4684
rect 6178 4672 6184 4684
rect 6139 4644 6184 4672
rect 6178 4632 6184 4644
rect 6236 4632 6242 4684
rect 6454 4681 6460 4684
rect 6448 4672 6460 4681
rect 6415 4644 6460 4672
rect 6448 4635 6460 4644
rect 6454 4632 6460 4635
rect 6512 4632 6518 4684
rect 8389 4675 8447 4681
rect 8389 4641 8401 4675
rect 8435 4672 8447 4675
rect 8846 4672 8852 4684
rect 8435 4644 8852 4672
rect 8435 4641 8447 4644
rect 8389 4635 8447 4641
rect 8846 4632 8852 4644
rect 8904 4632 8910 4684
rect 9766 4632 9772 4684
rect 9824 4672 9830 4684
rect 9824 4644 10272 4672
rect 9824 4632 9830 4644
rect 1578 4604 1584 4616
rect 1539 4576 1584 4604
rect 1578 4564 1584 4576
rect 1636 4564 1642 4616
rect 4890 4604 4896 4616
rect 4851 4576 4896 4604
rect 4890 4564 4896 4576
rect 4948 4564 4954 4616
rect 8297 4607 8355 4613
rect 8297 4573 8309 4607
rect 8343 4604 8355 4607
rect 10134 4604 10140 4616
rect 8343 4576 10140 4604
rect 8343 4573 8355 4576
rect 8297 4567 8355 4573
rect 10134 4564 10140 4576
rect 10192 4564 10198 4616
rect 10244 4613 10272 4644
rect 11422 4632 11428 4684
rect 11480 4672 11486 4684
rect 11701 4675 11759 4681
rect 11701 4672 11713 4675
rect 11480 4644 11713 4672
rect 11480 4632 11486 4644
rect 11701 4641 11713 4644
rect 11747 4641 11759 4675
rect 12802 4672 12808 4684
rect 12763 4644 12808 4672
rect 11701 4635 11759 4641
rect 12802 4632 12808 4644
rect 12860 4632 12866 4684
rect 10229 4607 10287 4613
rect 10229 4573 10241 4607
rect 10275 4573 10287 4607
rect 11790 4604 11796 4616
rect 11751 4576 11796 4604
rect 10229 4567 10287 4573
rect 11790 4564 11796 4576
rect 11848 4604 11854 4616
rect 12250 4604 12256 4616
rect 11848 4576 12256 4604
rect 11848 4564 11854 4576
rect 12250 4564 12256 4576
rect 12308 4564 12314 4616
rect 2130 4496 2136 4548
rect 2188 4536 2194 4548
rect 2869 4539 2927 4545
rect 2869 4536 2881 4539
rect 2188 4508 2881 4536
rect 2188 4496 2194 4508
rect 2869 4505 2881 4508
rect 2915 4505 2927 4539
rect 2869 4499 2927 4505
rect 9677 4539 9735 4545
rect 9677 4505 9689 4539
rect 9723 4536 9735 4539
rect 9950 4536 9956 4548
rect 9723 4508 9956 4536
rect 9723 4505 9735 4508
rect 9677 4499 9735 4505
rect 9950 4496 9956 4508
rect 10008 4496 10014 4548
rect 12434 4496 12440 4548
rect 12492 4536 12498 4548
rect 12989 4539 13047 4545
rect 12989 4536 13001 4539
rect 12492 4508 13001 4536
rect 12492 4496 12498 4508
rect 12989 4505 13001 4508
rect 13035 4505 13047 4539
rect 12989 4499 13047 4505
rect 2501 4471 2559 4477
rect 2501 4437 2513 4471
rect 2547 4468 2559 4471
rect 2774 4468 2780 4480
rect 2547 4440 2780 4468
rect 2547 4437 2559 4440
rect 2501 4431 2559 4437
rect 2774 4428 2780 4440
rect 2832 4428 2838 4480
rect 7926 4468 7932 4480
rect 7887 4440 7932 4468
rect 7926 4428 7932 4440
rect 7984 4428 7990 4480
rect 8570 4468 8576 4480
rect 8531 4440 8576 4468
rect 8570 4428 8576 4440
rect 8628 4428 8634 4480
rect 9493 4471 9551 4477
rect 9493 4437 9505 4471
rect 9539 4468 9551 4471
rect 9582 4468 9588 4480
rect 9539 4440 9588 4468
rect 9539 4437 9551 4440
rect 9493 4431 9551 4437
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 10686 4468 10692 4480
rect 10647 4440 10692 4468
rect 10686 4428 10692 4440
rect 10744 4428 10750 4480
rect 1104 4378 14812 4400
rect 1104 4326 3648 4378
rect 3700 4326 3712 4378
rect 3764 4326 3776 4378
rect 3828 4326 3840 4378
rect 3892 4326 8982 4378
rect 9034 4326 9046 4378
rect 9098 4326 9110 4378
rect 9162 4326 9174 4378
rect 9226 4326 14315 4378
rect 14367 4326 14379 4378
rect 14431 4326 14443 4378
rect 14495 4326 14507 4378
rect 14559 4326 14812 4378
rect 1104 4304 14812 4326
rect 2041 4267 2099 4273
rect 2041 4233 2053 4267
rect 2087 4264 2099 4267
rect 2222 4264 2228 4276
rect 2087 4236 2228 4264
rect 2087 4233 2099 4236
rect 2041 4227 2099 4233
rect 2222 4224 2228 4236
rect 2280 4224 2286 4276
rect 3510 4224 3516 4276
rect 3568 4264 3574 4276
rect 3881 4267 3939 4273
rect 3881 4264 3893 4267
rect 3568 4236 3893 4264
rect 3568 4224 3574 4236
rect 3881 4233 3893 4236
rect 3927 4233 3939 4267
rect 3881 4227 3939 4233
rect 4890 4224 4896 4276
rect 4948 4264 4954 4276
rect 5261 4267 5319 4273
rect 5261 4264 5273 4267
rect 4948 4236 5273 4264
rect 4948 4224 4954 4236
rect 5261 4233 5273 4236
rect 5307 4233 5319 4267
rect 5261 4227 5319 4233
rect 7742 4224 7748 4276
rect 7800 4264 7806 4276
rect 7929 4267 7987 4273
rect 7929 4264 7941 4267
rect 7800 4236 7941 4264
rect 7800 4224 7806 4236
rect 7929 4233 7941 4236
rect 7975 4233 7987 4267
rect 7929 4227 7987 4233
rect 8846 4224 8852 4276
rect 8904 4264 8910 4276
rect 8941 4267 8999 4273
rect 8941 4264 8953 4267
rect 8904 4236 8953 4264
rect 8904 4224 8910 4236
rect 8941 4233 8953 4236
rect 8987 4233 8999 4267
rect 9766 4264 9772 4276
rect 9727 4236 9772 4264
rect 8941 4227 8999 4233
rect 9766 4224 9772 4236
rect 9824 4224 9830 4276
rect 10045 4267 10103 4273
rect 10045 4233 10057 4267
rect 10091 4264 10103 4267
rect 10134 4264 10140 4276
rect 10091 4236 10140 4264
rect 10091 4233 10103 4236
rect 10045 4227 10103 4233
rect 10134 4224 10140 4236
rect 10192 4224 10198 4276
rect 12802 4224 12808 4276
rect 12860 4264 12866 4276
rect 13449 4267 13507 4273
rect 13449 4264 13461 4267
rect 12860 4236 13461 4264
rect 12860 4224 12866 4236
rect 13449 4233 13461 4236
rect 13495 4233 13507 4267
rect 13449 4227 13507 4233
rect 2317 4199 2375 4205
rect 2317 4165 2329 4199
rect 2363 4165 2375 4199
rect 2317 4159 2375 4165
rect 198 4088 204 4140
rect 256 4128 262 4140
rect 2332 4128 2360 4159
rect 3142 4156 3148 4208
rect 3200 4196 3206 4208
rect 3697 4199 3755 4205
rect 3697 4196 3709 4199
rect 3200 4168 3709 4196
rect 3200 4156 3206 4168
rect 3697 4165 3709 4168
rect 3743 4196 3755 4199
rect 8294 4196 8300 4208
rect 3743 4168 8300 4196
rect 3743 4165 3755 4168
rect 3697 4159 3755 4165
rect 4356 4137 4384 4168
rect 8294 4156 8300 4168
rect 8352 4156 8358 4208
rect 11241 4199 11299 4205
rect 11241 4196 11253 4199
rect 9600 4168 11253 4196
rect 256 4100 2360 4128
rect 4341 4131 4399 4137
rect 256 4088 262 4100
rect 4341 4097 4353 4131
rect 4387 4097 4399 4131
rect 4341 4091 4399 4097
rect 4525 4131 4583 4137
rect 4525 4097 4537 4131
rect 4571 4128 4583 4131
rect 4982 4128 4988 4140
rect 4571 4100 4988 4128
rect 4571 4097 4583 4100
rect 4525 4091 4583 4097
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 5166 4088 5172 4140
rect 5224 4128 5230 4140
rect 6086 4128 6092 4140
rect 5224 4100 6092 4128
rect 5224 4088 5230 4100
rect 6086 4088 6092 4100
rect 6144 4128 6150 4140
rect 7377 4131 7435 4137
rect 7377 4128 7389 4131
rect 6144 4100 7389 4128
rect 6144 4088 6150 4100
rect 2133 4063 2191 4069
rect 2133 4029 2145 4063
rect 2179 4060 2191 4063
rect 2958 4060 2964 4072
rect 2179 4032 2964 4060
rect 2179 4029 2191 4032
rect 2133 4023 2191 4029
rect 1673 3995 1731 4001
rect 1673 3961 1685 3995
rect 1719 3992 1731 3995
rect 2774 3992 2780 4004
rect 1719 3964 2780 3992
rect 1719 3961 1731 3964
rect 1673 3955 1731 3961
rect 2774 3952 2780 3964
rect 2832 3952 2838 4004
rect 2685 3927 2743 3933
rect 2685 3893 2697 3927
rect 2731 3924 2743 3927
rect 2884 3924 2912 4032
rect 2958 4020 2964 4032
rect 3016 4020 3022 4072
rect 3421 4063 3479 4069
rect 3421 4029 3433 4063
rect 3467 4060 3479 4063
rect 4249 4063 4307 4069
rect 4249 4060 4261 4063
rect 3467 4032 4261 4060
rect 3467 4029 3479 4032
rect 3421 4023 3479 4029
rect 4249 4029 4261 4032
rect 4295 4060 4307 4063
rect 5445 4063 5503 4069
rect 5445 4060 5457 4063
rect 4295 4032 5457 4060
rect 4295 4029 4307 4032
rect 4249 4023 4307 4029
rect 5445 4029 5457 4032
rect 5491 4060 5503 4063
rect 5997 4063 6055 4069
rect 5997 4060 6009 4063
rect 5491 4032 6009 4060
rect 5491 4029 5503 4032
rect 5445 4023 5503 4029
rect 5997 4029 6009 4032
rect 6043 4060 6055 4063
rect 6270 4060 6276 4072
rect 6043 4032 6276 4060
rect 6043 4029 6055 4032
rect 5997 4023 6055 4029
rect 6270 4020 6276 4032
rect 6328 4020 6334 4072
rect 6840 4069 6868 4100
rect 7377 4097 7389 4100
rect 7423 4128 7435 4131
rect 7650 4128 7656 4140
rect 7423 4100 7656 4128
rect 7423 4097 7435 4100
rect 7377 4091 7435 4097
rect 7650 4088 7656 4100
rect 7708 4088 7714 4140
rect 7926 4088 7932 4140
rect 7984 4128 7990 4140
rect 8481 4131 8539 4137
rect 8481 4128 8493 4131
rect 7984 4100 8493 4128
rect 7984 4088 7990 4100
rect 8481 4097 8493 4100
rect 8527 4128 8539 4131
rect 8846 4128 8852 4140
rect 8527 4100 8852 4128
rect 8527 4097 8539 4100
rect 8481 4091 8539 4097
rect 8846 4088 8852 4100
rect 8904 4088 8910 4140
rect 9398 4128 9404 4140
rect 9359 4100 9404 4128
rect 9398 4088 9404 4100
rect 9456 4128 9462 4140
rect 9600 4128 9628 4168
rect 10612 4137 10640 4168
rect 11241 4165 11253 4168
rect 11287 4196 11299 4199
rect 11790 4196 11796 4208
rect 11287 4168 11796 4196
rect 11287 4165 11299 4168
rect 11241 4159 11299 4165
rect 11790 4156 11796 4168
rect 11848 4156 11854 4208
rect 11992 4168 12296 4196
rect 9456 4100 9628 4128
rect 10597 4131 10655 4137
rect 9456 4088 9462 4100
rect 10597 4097 10609 4131
rect 10643 4097 10655 4131
rect 11992 4128 12020 4168
rect 12268 4140 12296 4168
rect 12544 4168 13032 4196
rect 10597 4091 10655 4097
rect 11808 4100 12020 4128
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4060 6883 4063
rect 8297 4063 8355 4069
rect 6871 4032 6905 4060
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 8297 4029 8309 4063
rect 8343 4060 8355 4063
rect 8386 4060 8392 4072
rect 8343 4032 8392 4060
rect 8343 4029 8355 4032
rect 8297 4023 8355 4029
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 10134 4020 10140 4072
rect 10192 4060 10198 4072
rect 10502 4060 10508 4072
rect 10192 4032 10508 4060
rect 10192 4020 10198 4032
rect 10502 4020 10508 4032
rect 10560 4020 10566 4072
rect 11330 4020 11336 4072
rect 11388 4060 11394 4072
rect 11808 4069 11836 4100
rect 12250 4088 12256 4140
rect 12308 4128 12314 4140
rect 12544 4128 12572 4168
rect 12308 4100 12572 4128
rect 12308 4088 12314 4100
rect 12618 4088 12624 4140
rect 12676 4128 12682 4140
rect 13004 4137 13032 4168
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 12676 4100 12909 4128
rect 12676 4088 12682 4100
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 12897 4091 12955 4097
rect 12989 4131 13047 4137
rect 12989 4097 13001 4131
rect 13035 4097 13047 4131
rect 12989 4091 13047 4097
rect 11793 4063 11851 4069
rect 11793 4060 11805 4063
rect 11388 4032 11805 4060
rect 11388 4020 11394 4032
rect 11793 4029 11805 4032
rect 11839 4029 11851 4063
rect 11793 4023 11851 4029
rect 12161 4063 12219 4069
rect 12161 4029 12173 4063
rect 12207 4060 12219 4063
rect 12207 4032 12848 4060
rect 12207 4029 12219 4032
rect 12161 4023 12219 4029
rect 6454 3992 6460 4004
rect 6367 3964 6460 3992
rect 4982 3924 4988 3936
rect 2731 3896 2912 3924
rect 4943 3896 4988 3924
rect 2731 3893 2743 3896
rect 2685 3887 2743 3893
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 5626 3924 5632 3936
rect 5587 3896 5632 3924
rect 5626 3884 5632 3896
rect 5684 3884 5690 3936
rect 6086 3884 6092 3936
rect 6144 3924 6150 3936
rect 6380 3933 6408 3964
rect 6454 3952 6460 3964
rect 6512 3992 6518 4004
rect 7745 3995 7803 4001
rect 7745 3992 7757 3995
rect 6512 3964 7757 3992
rect 6512 3952 6518 3964
rect 7745 3961 7757 3964
rect 7791 3992 7803 3995
rect 7926 3992 7932 4004
rect 7791 3964 7932 3992
rect 7791 3961 7803 3964
rect 7745 3955 7803 3961
rect 7926 3952 7932 3964
rect 7984 3952 7990 4004
rect 9582 3952 9588 4004
rect 9640 3992 9646 4004
rect 10413 3995 10471 4001
rect 9640 3964 9812 3992
rect 9640 3952 9646 3964
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 6144 3896 6377 3924
rect 6144 3884 6150 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 7006 3924 7012 3936
rect 6967 3896 7012 3924
rect 6365 3887 6423 3893
rect 7006 3884 7012 3896
rect 7064 3884 7070 3936
rect 8202 3884 8208 3936
rect 8260 3924 8266 3936
rect 8389 3927 8447 3933
rect 8389 3924 8401 3927
rect 8260 3896 8401 3924
rect 8260 3884 8266 3896
rect 8389 3893 8401 3896
rect 8435 3893 8447 3927
rect 9784 3924 9812 3964
rect 10413 3961 10425 3995
rect 10459 3992 10471 3995
rect 10594 3992 10600 4004
rect 10459 3964 10600 3992
rect 10459 3961 10471 3964
rect 10413 3955 10471 3961
rect 10594 3952 10600 3964
rect 10652 3952 10658 4004
rect 11422 3952 11428 4004
rect 11480 3992 11486 4004
rect 11480 3964 12480 3992
rect 11480 3952 11486 3964
rect 10502 3924 10508 3936
rect 9784 3896 10508 3924
rect 8389 3887 8447 3893
rect 10502 3884 10508 3896
rect 10560 3884 10566 3936
rect 12452 3933 12480 3964
rect 12820 3933 12848 4032
rect 12437 3927 12495 3933
rect 12437 3893 12449 3927
rect 12483 3893 12495 3927
rect 12437 3887 12495 3893
rect 12805 3927 12863 3933
rect 12805 3893 12817 3927
rect 12851 3924 12863 3927
rect 12986 3924 12992 3936
rect 12851 3896 12992 3924
rect 12851 3893 12863 3896
rect 12805 3887 12863 3893
rect 12986 3884 12992 3896
rect 13044 3924 13050 3936
rect 15746 3924 15752 3936
rect 13044 3896 15752 3924
rect 13044 3884 13050 3896
rect 15746 3884 15752 3896
rect 15804 3884 15810 3936
rect 1104 3834 14812 3856
rect 1104 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 11648 3834
rect 11700 3782 11712 3834
rect 11764 3782 11776 3834
rect 11828 3782 11840 3834
rect 11892 3782 14812 3834
rect 1104 3760 14812 3782
rect 2406 3720 2412 3732
rect 2367 3692 2412 3720
rect 2406 3680 2412 3692
rect 2464 3680 2470 3732
rect 2774 3680 2780 3732
rect 2832 3720 2838 3732
rect 4065 3723 4123 3729
rect 4065 3720 4077 3723
rect 2832 3692 4077 3720
rect 2832 3680 2838 3692
rect 4065 3689 4077 3692
rect 4111 3689 4123 3723
rect 4065 3683 4123 3689
rect 4982 3680 4988 3732
rect 5040 3720 5046 3732
rect 5077 3723 5135 3729
rect 5077 3720 5089 3723
rect 5040 3692 5089 3720
rect 5040 3680 5046 3692
rect 5077 3689 5089 3692
rect 5123 3689 5135 3723
rect 5534 3720 5540 3732
rect 5495 3692 5540 3720
rect 5077 3683 5135 3689
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 6825 3723 6883 3729
rect 6825 3689 6837 3723
rect 6871 3720 6883 3723
rect 7098 3720 7104 3732
rect 6871 3692 7104 3720
rect 6871 3689 6883 3692
rect 6825 3683 6883 3689
rect 7098 3680 7104 3692
rect 7156 3680 7162 3732
rect 8021 3723 8079 3729
rect 8021 3689 8033 3723
rect 8067 3720 8079 3723
rect 8386 3720 8392 3732
rect 8067 3692 8392 3720
rect 8067 3689 8079 3692
rect 8021 3683 8079 3689
rect 8386 3680 8392 3692
rect 8444 3680 8450 3732
rect 9125 3723 9183 3729
rect 9125 3689 9137 3723
rect 9171 3720 9183 3723
rect 9306 3720 9312 3732
rect 9171 3692 9312 3720
rect 9171 3689 9183 3692
rect 9125 3683 9183 3689
rect 2317 3655 2375 3661
rect 2317 3621 2329 3655
rect 2363 3652 2375 3655
rect 3050 3652 3056 3664
rect 2363 3624 3056 3652
rect 2363 3621 2375 3624
rect 2317 3615 2375 3621
rect 3050 3612 3056 3624
rect 3108 3612 3114 3664
rect 3970 3612 3976 3664
rect 4028 3652 4034 3664
rect 4433 3655 4491 3661
rect 4433 3652 4445 3655
rect 4028 3624 4445 3652
rect 4028 3612 4034 3624
rect 4433 3621 4445 3624
rect 4479 3652 4491 3655
rect 5166 3652 5172 3664
rect 4479 3624 5172 3652
rect 4479 3621 4491 3624
rect 4433 3615 4491 3621
rect 5166 3612 5172 3624
rect 5224 3612 5230 3664
rect 5258 3612 5264 3664
rect 5316 3652 5322 3664
rect 5813 3655 5871 3661
rect 5813 3652 5825 3655
rect 5316 3624 5825 3652
rect 5316 3612 5322 3624
rect 5813 3621 5825 3624
rect 5859 3621 5871 3655
rect 5813 3615 5871 3621
rect 5902 3612 5908 3664
rect 5960 3652 5966 3664
rect 6917 3655 6975 3661
rect 6917 3652 6929 3655
rect 5960 3624 6929 3652
rect 5960 3612 5966 3624
rect 6917 3621 6929 3624
rect 6963 3621 6975 3655
rect 6917 3615 6975 3621
rect 7558 3612 7564 3664
rect 7616 3652 7622 3664
rect 7926 3652 7932 3664
rect 7616 3624 7932 3652
rect 7616 3612 7622 3624
rect 7926 3612 7932 3624
rect 7984 3652 7990 3664
rect 8481 3655 8539 3661
rect 8481 3652 8493 3655
rect 7984 3624 8493 3652
rect 7984 3612 7990 3624
rect 8481 3621 8493 3624
rect 8527 3621 8539 3655
rect 8481 3615 8539 3621
rect 4522 3584 4528 3596
rect 4435 3556 4528 3584
rect 4522 3544 4528 3556
rect 4580 3584 4586 3596
rect 7576 3584 7604 3612
rect 4580 3556 7604 3584
rect 4580 3544 4586 3556
rect 7650 3544 7656 3596
rect 7708 3584 7714 3596
rect 8389 3587 8447 3593
rect 8389 3584 8401 3587
rect 7708 3556 8401 3584
rect 7708 3544 7714 3556
rect 8389 3553 8401 3556
rect 8435 3553 8447 3587
rect 8389 3547 8447 3553
rect 2866 3516 2872 3528
rect 2827 3488 2872 3516
rect 2866 3476 2872 3488
rect 2924 3476 2930 3528
rect 3050 3516 3056 3528
rect 3011 3488 3056 3516
rect 3050 3476 3056 3488
rect 3108 3476 3114 3528
rect 4709 3519 4767 3525
rect 4709 3485 4721 3519
rect 4755 3516 4767 3519
rect 4982 3516 4988 3528
rect 4755 3488 4988 3516
rect 4755 3485 4767 3488
rect 4709 3479 4767 3485
rect 3326 3408 3332 3460
rect 3384 3448 3390 3460
rect 3513 3451 3571 3457
rect 3513 3448 3525 3451
rect 3384 3420 3525 3448
rect 3384 3408 3390 3420
rect 3513 3417 3525 3420
rect 3559 3448 3571 3451
rect 3881 3451 3939 3457
rect 3881 3448 3893 3451
rect 3559 3420 3893 3448
rect 3559 3417 3571 3420
rect 3513 3411 3571 3417
rect 3881 3417 3893 3420
rect 3927 3448 3939 3451
rect 4338 3448 4344 3460
rect 3927 3420 4344 3448
rect 3927 3417 3939 3420
rect 3881 3411 3939 3417
rect 4338 3408 4344 3420
rect 4396 3448 4402 3460
rect 4724 3448 4752 3479
rect 4982 3476 4988 3488
rect 5040 3476 5046 3528
rect 7009 3519 7067 3525
rect 7009 3516 7021 3519
rect 6288 3488 7021 3516
rect 4396 3420 4752 3448
rect 4396 3408 4402 3420
rect 1946 3380 1952 3392
rect 1907 3352 1952 3380
rect 1946 3340 1952 3352
rect 2004 3340 2010 3392
rect 3418 3340 3424 3392
rect 3476 3380 3482 3392
rect 6086 3380 6092 3392
rect 3476 3352 6092 3380
rect 3476 3340 3482 3352
rect 6086 3340 6092 3352
rect 6144 3380 6150 3392
rect 6288 3389 6316 3488
rect 7009 3485 7021 3488
rect 7055 3485 7067 3519
rect 7009 3479 7067 3485
rect 8665 3519 8723 3525
rect 8665 3485 8677 3519
rect 8711 3516 8723 3519
rect 9140 3516 9168 3683
rect 9306 3680 9312 3692
rect 9364 3680 9370 3732
rect 10137 3723 10195 3729
rect 10137 3689 10149 3723
rect 10183 3720 10195 3723
rect 10686 3720 10692 3732
rect 10183 3692 10692 3720
rect 10183 3689 10195 3692
rect 10137 3683 10195 3689
rect 10686 3680 10692 3692
rect 10744 3680 10750 3732
rect 10962 3680 10968 3732
rect 11020 3720 11026 3732
rect 11149 3723 11207 3729
rect 11149 3720 11161 3723
rect 11020 3692 11161 3720
rect 11020 3680 11026 3692
rect 11149 3689 11161 3692
rect 11195 3689 11207 3723
rect 11149 3683 11207 3689
rect 11514 3680 11520 3732
rect 11572 3720 11578 3732
rect 11701 3723 11759 3729
rect 11701 3720 11713 3723
rect 11572 3692 11713 3720
rect 11572 3680 11578 3692
rect 11701 3689 11713 3692
rect 11747 3689 11759 3723
rect 11701 3683 11759 3689
rect 12069 3723 12127 3729
rect 12069 3689 12081 3723
rect 12115 3720 12127 3723
rect 12342 3720 12348 3732
rect 12115 3692 12348 3720
rect 12115 3689 12127 3692
rect 12069 3683 12127 3689
rect 12342 3680 12348 3692
rect 12400 3680 12406 3732
rect 12710 3680 12716 3732
rect 12768 3720 12774 3732
rect 12768 3692 13308 3720
rect 12768 3680 12774 3692
rect 10042 3612 10048 3664
rect 10100 3652 10106 3664
rect 10597 3655 10655 3661
rect 10597 3652 10609 3655
rect 10100 3624 10609 3652
rect 10100 3612 10106 3624
rect 10597 3621 10609 3624
rect 10643 3621 10655 3655
rect 12802 3652 12808 3664
rect 10597 3615 10655 3621
rect 12176 3624 12808 3652
rect 10505 3587 10563 3593
rect 10505 3553 10517 3587
rect 10551 3553 10563 3587
rect 10505 3547 10563 3553
rect 8711 3488 9168 3516
rect 10045 3519 10103 3525
rect 8711 3485 8723 3488
rect 8665 3479 8723 3485
rect 10045 3485 10057 3519
rect 10091 3516 10103 3519
rect 10226 3516 10232 3528
rect 10091 3488 10232 3516
rect 10091 3485 10103 3488
rect 10045 3479 10103 3485
rect 6457 3451 6515 3457
rect 6457 3417 6469 3451
rect 6503 3448 6515 3451
rect 6730 3448 6736 3460
rect 6503 3420 6736 3448
rect 6503 3417 6515 3420
rect 6457 3411 6515 3417
rect 6730 3408 6736 3420
rect 6788 3408 6794 3460
rect 7561 3451 7619 3457
rect 7561 3417 7573 3451
rect 7607 3448 7619 3451
rect 7929 3451 7987 3457
rect 7929 3448 7941 3451
rect 7607 3420 7941 3448
rect 7607 3417 7619 3420
rect 7561 3411 7619 3417
rect 7929 3417 7941 3420
rect 7975 3448 7987 3451
rect 8386 3448 8392 3460
rect 7975 3420 8392 3448
rect 7975 3417 7987 3420
rect 7929 3411 7987 3417
rect 8386 3408 8392 3420
rect 8444 3448 8450 3460
rect 8680 3448 8708 3479
rect 10226 3476 10232 3488
rect 10284 3516 10290 3528
rect 10520 3516 10548 3547
rect 11422 3544 11428 3596
rect 11480 3584 11486 3596
rect 11517 3587 11575 3593
rect 11517 3584 11529 3587
rect 11480 3556 11529 3584
rect 11480 3544 11486 3556
rect 11517 3553 11529 3556
rect 11563 3553 11575 3587
rect 11517 3547 11575 3553
rect 12176 3528 12204 3624
rect 12802 3612 12808 3624
rect 12860 3612 12866 3664
rect 13280 3596 13308 3692
rect 13262 3584 13268 3596
rect 13175 3556 13268 3584
rect 13262 3544 13268 3556
rect 13320 3544 13326 3596
rect 10284 3488 10548 3516
rect 10781 3519 10839 3525
rect 10284 3476 10290 3488
rect 10781 3485 10793 3519
rect 10827 3516 10839 3519
rect 10962 3516 10968 3528
rect 10827 3488 10968 3516
rect 10827 3485 10839 3488
rect 10781 3479 10839 3485
rect 8444 3420 8708 3448
rect 9493 3451 9551 3457
rect 8444 3408 8450 3420
rect 9493 3417 9505 3451
rect 9539 3448 9551 3451
rect 10796 3448 10824 3479
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 12158 3516 12164 3528
rect 12119 3488 12164 3516
rect 12158 3476 12164 3488
rect 12216 3476 12222 3528
rect 12250 3476 12256 3528
rect 12308 3516 12314 3528
rect 12710 3516 12716 3528
rect 12308 3488 12716 3516
rect 12308 3476 12314 3488
rect 12710 3476 12716 3488
rect 12768 3476 12774 3528
rect 13446 3448 13452 3460
rect 9539 3420 10824 3448
rect 13407 3420 13452 3448
rect 9539 3417 9551 3420
rect 9493 3411 9551 3417
rect 13446 3408 13452 3420
rect 13504 3408 13510 3460
rect 6273 3383 6331 3389
rect 6273 3380 6285 3383
rect 6144 3352 6285 3380
rect 6144 3340 6150 3352
rect 6273 3349 6285 3352
rect 6319 3349 6331 3383
rect 13078 3380 13084 3392
rect 13039 3352 13084 3380
rect 6273 3343 6331 3349
rect 13078 3340 13084 3352
rect 13136 3340 13142 3392
rect 1104 3290 14812 3312
rect 1104 3238 3648 3290
rect 3700 3238 3712 3290
rect 3764 3238 3776 3290
rect 3828 3238 3840 3290
rect 3892 3238 8982 3290
rect 9034 3238 9046 3290
rect 9098 3238 9110 3290
rect 9162 3238 9174 3290
rect 9226 3238 14315 3290
rect 14367 3238 14379 3290
rect 14431 3238 14443 3290
rect 14495 3238 14507 3290
rect 14559 3238 14812 3290
rect 1104 3216 14812 3238
rect 3326 3176 3332 3188
rect 3287 3148 3332 3176
rect 3326 3136 3332 3148
rect 3384 3136 3390 3188
rect 3697 3179 3755 3185
rect 3697 3145 3709 3179
rect 3743 3176 3755 3179
rect 3970 3176 3976 3188
rect 3743 3148 3976 3176
rect 3743 3145 3755 3148
rect 3697 3139 3755 3145
rect 3970 3136 3976 3148
rect 4028 3136 4034 3188
rect 4065 3179 4123 3185
rect 4065 3145 4077 3179
rect 4111 3176 4123 3179
rect 4522 3176 4528 3188
rect 4111 3148 4528 3176
rect 4111 3145 4123 3148
rect 4065 3139 4123 3145
rect 4522 3136 4528 3148
rect 4580 3136 4586 3188
rect 5442 3136 5448 3188
rect 5500 3176 5506 3188
rect 5537 3179 5595 3185
rect 5537 3176 5549 3179
rect 5500 3148 5549 3176
rect 5500 3136 5506 3148
rect 5537 3145 5549 3148
rect 5583 3145 5595 3179
rect 5537 3139 5595 3145
rect 6181 3179 6239 3185
rect 6181 3145 6193 3179
rect 6227 3176 6239 3179
rect 6546 3176 6552 3188
rect 6227 3148 6552 3176
rect 6227 3145 6239 3148
rect 6181 3139 6239 3145
rect 6546 3136 6552 3148
rect 6604 3136 6610 3188
rect 7650 3176 7656 3188
rect 7611 3148 7656 3176
rect 7650 3136 7656 3148
rect 7708 3136 7714 3188
rect 7926 3136 7932 3188
rect 7984 3176 7990 3188
rect 8021 3179 8079 3185
rect 8021 3176 8033 3179
rect 7984 3148 8033 3176
rect 7984 3136 7990 3148
rect 8021 3145 8033 3148
rect 8067 3145 8079 3179
rect 8021 3139 8079 3145
rect 6457 3111 6515 3117
rect 6457 3077 6469 3111
rect 6503 3108 6515 3111
rect 6822 3108 6828 3120
rect 6503 3080 6828 3108
rect 6503 3077 6515 3080
rect 6457 3071 6515 3077
rect 6822 3068 6828 3080
rect 6880 3068 6886 3120
rect 8036 3040 8064 3139
rect 8846 3136 8852 3188
rect 8904 3176 8910 3188
rect 9585 3179 9643 3185
rect 9585 3176 9597 3179
rect 8904 3148 9597 3176
rect 8904 3136 8910 3148
rect 9585 3145 9597 3148
rect 9631 3145 9643 3179
rect 9585 3139 9643 3145
rect 9953 3179 10011 3185
rect 9953 3145 9965 3179
rect 9999 3176 10011 3179
rect 10042 3176 10048 3188
rect 9999 3148 10048 3176
rect 9999 3145 10011 3148
rect 9953 3139 10011 3145
rect 10042 3136 10048 3148
rect 10100 3136 10106 3188
rect 10134 3136 10140 3188
rect 10192 3176 10198 3188
rect 10229 3179 10287 3185
rect 10229 3176 10241 3179
rect 10192 3148 10241 3176
rect 10192 3136 10198 3148
rect 10229 3145 10241 3148
rect 10275 3145 10287 3179
rect 10229 3139 10287 3145
rect 11793 3179 11851 3185
rect 11793 3145 11805 3179
rect 11839 3176 11851 3179
rect 12158 3176 12164 3188
rect 11839 3148 12164 3176
rect 11839 3145 11851 3148
rect 11793 3139 11851 3145
rect 8036 3012 8340 3040
rect 1949 2975 2007 2981
rect 1949 2941 1961 2975
rect 1995 2972 2007 2975
rect 4157 2975 4215 2981
rect 4157 2972 4169 2975
rect 1995 2944 4169 2972
rect 1995 2941 2007 2944
rect 1949 2935 2007 2941
rect 4157 2941 4169 2944
rect 4203 2972 4215 2975
rect 4798 2972 4804 2984
rect 4203 2944 4804 2972
rect 4203 2941 4215 2944
rect 4157 2935 4215 2941
rect 4798 2932 4804 2944
rect 4856 2932 4862 2984
rect 6546 2932 6552 2984
rect 6604 2972 6610 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6604 2944 6837 2972
rect 6604 2932 6610 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 8110 2932 8116 2984
rect 8168 2972 8174 2984
rect 8205 2975 8263 2981
rect 8205 2972 8217 2975
rect 8168 2944 8217 2972
rect 8168 2932 8174 2944
rect 8205 2941 8217 2944
rect 8251 2941 8263 2975
rect 8312 2972 8340 3012
rect 8846 2972 8852 2984
rect 8312 2944 8852 2972
rect 8205 2935 8263 2941
rect 2216 2907 2274 2913
rect 2216 2873 2228 2907
rect 2262 2873 2274 2907
rect 2216 2867 2274 2873
rect 1857 2839 1915 2845
rect 1857 2805 1869 2839
rect 1903 2836 1915 2839
rect 2240 2836 2268 2867
rect 4338 2864 4344 2916
rect 4396 2913 4402 2916
rect 4396 2907 4460 2913
rect 4396 2873 4414 2907
rect 4448 2873 4460 2907
rect 8220 2904 8248 2935
rect 8846 2932 8852 2944
rect 8904 2932 8910 2984
rect 10244 2972 10272 3139
rect 12158 3136 12164 3148
rect 12216 3136 12222 3188
rect 12434 3136 12440 3188
rect 12492 3176 12498 3188
rect 12492 3148 12537 3176
rect 12492 3136 12498 3148
rect 13262 3136 13268 3188
rect 13320 3176 13326 3188
rect 13449 3179 13507 3185
rect 13449 3176 13461 3179
rect 13320 3148 13461 3176
rect 13320 3136 13326 3148
rect 13449 3145 13461 3148
rect 13495 3145 13507 3179
rect 13449 3139 13507 3145
rect 10413 3111 10471 3117
rect 10413 3077 10425 3111
rect 10459 3108 10471 3111
rect 13078 3108 13084 3120
rect 10459 3080 13084 3108
rect 10459 3077 10471 3080
rect 10413 3071 10471 3077
rect 10962 3040 10968 3052
rect 10923 3012 10968 3040
rect 10962 3000 10968 3012
rect 11020 3040 11026 3052
rect 11422 3040 11428 3052
rect 11020 3012 11428 3040
rect 11020 3000 11026 3012
rect 11422 3000 11428 3012
rect 11480 3000 11486 3052
rect 12161 3043 12219 3049
rect 12161 3009 12173 3043
rect 12207 3040 12219 3043
rect 12342 3040 12348 3052
rect 12207 3012 12348 3040
rect 12207 3009 12219 3012
rect 12161 3003 12219 3009
rect 12342 3000 12348 3012
rect 12400 3000 12406 3052
rect 12912 3049 12940 3080
rect 13078 3068 13084 3080
rect 13136 3068 13142 3120
rect 12897 3043 12955 3049
rect 12897 3009 12909 3043
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 12989 3043 13047 3049
rect 12989 3009 13001 3043
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 10873 2975 10931 2981
rect 10873 2972 10885 2975
rect 10244 2944 10885 2972
rect 8294 2904 8300 2916
rect 8220 2876 8300 2904
rect 4396 2867 4460 2873
rect 4396 2864 4402 2867
rect 8294 2864 8300 2876
rect 8352 2864 8358 2916
rect 8386 2864 8392 2916
rect 8444 2913 8450 2916
rect 8444 2907 8508 2913
rect 8444 2873 8462 2907
rect 8496 2873 8508 2907
rect 8444 2867 8508 2873
rect 8444 2864 8450 2867
rect 8570 2864 8576 2916
rect 8628 2904 8634 2916
rect 10244 2904 10272 2944
rect 10873 2941 10885 2944
rect 10919 2941 10931 2975
rect 10873 2935 10931 2941
rect 12710 2932 12716 2984
rect 12768 2972 12774 2984
rect 13004 2972 13032 3003
rect 12768 2944 13032 2972
rect 12768 2932 12774 2944
rect 10778 2904 10784 2916
rect 8628 2876 10272 2904
rect 10739 2876 10784 2904
rect 8628 2864 8634 2876
rect 10778 2864 10784 2876
rect 10836 2904 10842 2916
rect 11054 2904 11060 2916
rect 10836 2876 11060 2904
rect 10836 2864 10842 2876
rect 11054 2864 11060 2876
rect 11112 2864 11118 2916
rect 11146 2864 11152 2916
rect 11204 2904 11210 2916
rect 12158 2904 12164 2916
rect 11204 2876 12164 2904
rect 11204 2864 11210 2876
rect 12158 2864 12164 2876
rect 12216 2864 12222 2916
rect 12802 2904 12808 2916
rect 12763 2876 12808 2904
rect 12802 2864 12808 2876
rect 12860 2904 12866 2916
rect 13817 2907 13875 2913
rect 13817 2904 13829 2907
rect 12860 2876 13829 2904
rect 12860 2864 12866 2876
rect 13817 2873 13829 2876
rect 13863 2873 13875 2907
rect 13817 2867 13875 2873
rect 2682 2836 2688 2848
rect 1903 2808 2688 2836
rect 1903 2805 1915 2808
rect 1857 2799 1915 2805
rect 2682 2796 2688 2808
rect 2740 2796 2746 2848
rect 7006 2836 7012 2848
rect 6967 2808 7012 2836
rect 7006 2796 7012 2808
rect 7064 2796 7070 2848
rect 9490 2796 9496 2848
rect 9548 2836 9554 2848
rect 9674 2836 9680 2848
rect 9548 2808 9680 2836
rect 9548 2796 9554 2808
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 1104 2746 14812 2768
rect 1104 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 11648 2746
rect 11700 2694 11712 2746
rect 11764 2694 11776 2746
rect 11828 2694 11840 2746
rect 11892 2694 14812 2746
rect 1104 2672 14812 2694
rect 2409 2635 2467 2641
rect 2409 2601 2421 2635
rect 2455 2632 2467 2635
rect 2498 2632 2504 2644
rect 2455 2604 2504 2632
rect 2455 2601 2467 2604
rect 2409 2595 2467 2601
rect 2498 2592 2504 2604
rect 2556 2592 2562 2644
rect 2866 2592 2872 2644
rect 2924 2632 2930 2644
rect 4065 2635 4123 2641
rect 4065 2632 4077 2635
rect 2924 2604 4077 2632
rect 2924 2592 2930 2604
rect 4065 2601 4077 2604
rect 4111 2601 4123 2635
rect 4433 2635 4491 2641
rect 4433 2632 4445 2635
rect 4065 2595 4123 2601
rect 4172 2604 4445 2632
rect 2958 2524 2964 2576
rect 3016 2564 3022 2576
rect 3513 2567 3571 2573
rect 3513 2564 3525 2567
rect 3016 2536 3525 2564
rect 3016 2524 3022 2536
rect 3513 2533 3525 2536
rect 3559 2564 3571 2567
rect 4172 2564 4200 2604
rect 4433 2601 4445 2604
rect 4479 2632 4491 2635
rect 8113 2635 8171 2641
rect 4479 2604 4752 2632
rect 4479 2601 4491 2604
rect 4433 2595 4491 2601
rect 3559 2536 4200 2564
rect 3559 2533 3571 2536
rect 3513 2527 3571 2533
rect 4338 2524 4344 2576
rect 4396 2564 4402 2576
rect 4396 2536 4568 2564
rect 4396 2524 4402 2536
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2496 1455 2499
rect 1949 2499 2007 2505
rect 1949 2496 1961 2499
rect 1443 2468 1961 2496
rect 1443 2465 1455 2468
rect 1397 2459 1455 2465
rect 1949 2465 1961 2468
rect 1995 2496 2007 2499
rect 2777 2499 2835 2505
rect 2777 2496 2789 2499
rect 1995 2468 2789 2496
rect 1995 2465 2007 2468
rect 1949 2459 2007 2465
rect 2777 2465 2789 2468
rect 2823 2465 2835 2499
rect 4062 2496 4068 2508
rect 2777 2459 2835 2465
rect 2884 2468 4068 2496
rect 2884 2437 2912 2468
rect 4062 2456 4068 2468
rect 4120 2456 4126 2508
rect 4540 2496 4568 2536
rect 4540 2468 4660 2496
rect 2317 2431 2375 2437
rect 2317 2397 2329 2431
rect 2363 2428 2375 2431
rect 2869 2431 2927 2437
rect 2869 2428 2881 2431
rect 2363 2400 2881 2428
rect 2363 2397 2375 2400
rect 2317 2391 2375 2397
rect 2869 2397 2881 2400
rect 2915 2397 2927 2431
rect 2869 2391 2927 2397
rect 2961 2431 3019 2437
rect 2961 2397 2973 2431
rect 3007 2428 3019 2431
rect 3418 2428 3424 2440
rect 3007 2400 3424 2428
rect 3007 2397 3019 2400
rect 2961 2391 3019 2397
rect 1946 2320 1952 2372
rect 2004 2360 2010 2372
rect 2976 2360 3004 2391
rect 3418 2388 3424 2400
rect 3476 2388 3482 2440
rect 3881 2431 3939 2437
rect 3881 2397 3893 2431
rect 3927 2428 3939 2431
rect 4522 2428 4528 2440
rect 3927 2400 4528 2428
rect 3927 2397 3939 2400
rect 3881 2391 3939 2397
rect 4522 2388 4528 2400
rect 4580 2388 4586 2440
rect 4632 2437 4660 2468
rect 4617 2431 4675 2437
rect 4617 2397 4629 2431
rect 4663 2397 4675 2431
rect 4724 2428 4752 2604
rect 8113 2601 8125 2635
rect 8159 2632 8171 2635
rect 8202 2632 8208 2644
rect 8159 2604 8208 2632
rect 8159 2601 8171 2604
rect 8113 2595 8171 2601
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 8481 2635 8539 2641
rect 8481 2601 8493 2635
rect 8527 2632 8539 2635
rect 8662 2632 8668 2644
rect 8527 2604 8668 2632
rect 8527 2601 8539 2604
rect 8481 2595 8539 2601
rect 5537 2567 5595 2573
rect 5537 2533 5549 2567
rect 5583 2564 5595 2567
rect 7653 2567 7711 2573
rect 5583 2536 5948 2564
rect 5583 2533 5595 2536
rect 5537 2527 5595 2533
rect 5920 2508 5948 2536
rect 7653 2533 7665 2567
rect 7699 2564 7711 2567
rect 8496 2564 8524 2595
rect 8662 2592 8668 2604
rect 8720 2592 8726 2644
rect 10042 2632 10048 2644
rect 10003 2604 10048 2632
rect 10042 2592 10048 2604
rect 10100 2592 10106 2644
rect 11054 2632 11060 2644
rect 11015 2604 11060 2632
rect 11054 2592 11060 2604
rect 11112 2592 11118 2644
rect 11422 2632 11428 2644
rect 11383 2604 11428 2632
rect 11422 2592 11428 2604
rect 11480 2592 11486 2644
rect 11885 2635 11943 2641
rect 11885 2601 11897 2635
rect 11931 2632 11943 2635
rect 12066 2632 12072 2644
rect 11931 2604 12072 2632
rect 11931 2601 11943 2604
rect 11885 2595 11943 2601
rect 12066 2592 12072 2604
rect 12124 2592 12130 2644
rect 7699 2536 8524 2564
rect 8573 2567 8631 2573
rect 7699 2533 7711 2536
rect 7653 2527 7711 2533
rect 8573 2533 8585 2567
rect 8619 2564 8631 2567
rect 8754 2564 8760 2576
rect 8619 2536 8760 2564
rect 8619 2533 8631 2536
rect 8573 2527 8631 2533
rect 5169 2499 5227 2505
rect 5169 2465 5181 2499
rect 5215 2496 5227 2499
rect 5626 2496 5632 2508
rect 5215 2468 5632 2496
rect 5215 2465 5227 2468
rect 5169 2459 5227 2465
rect 5626 2456 5632 2468
rect 5684 2456 5690 2508
rect 5902 2456 5908 2508
rect 5960 2496 5966 2508
rect 6457 2499 6515 2505
rect 6457 2496 6469 2499
rect 5960 2468 6469 2496
rect 5960 2456 5966 2468
rect 6457 2465 6469 2468
rect 6503 2496 6515 2499
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 6503 2468 6929 2496
rect 6503 2465 6515 2468
rect 6457 2459 6515 2465
rect 6917 2465 6929 2468
rect 6963 2465 6975 2499
rect 6917 2459 6975 2465
rect 7668 2428 7696 2527
rect 8018 2496 8024 2508
rect 7931 2468 8024 2496
rect 8018 2456 8024 2468
rect 8076 2496 8082 2508
rect 8588 2496 8616 2527
rect 8754 2524 8760 2536
rect 8812 2524 8818 2576
rect 9217 2567 9275 2573
rect 9217 2533 9229 2567
rect 9263 2564 9275 2567
rect 9490 2564 9496 2576
rect 9263 2536 9496 2564
rect 9263 2533 9275 2536
rect 9217 2527 9275 2533
rect 9490 2524 9496 2536
rect 9548 2564 9554 2576
rect 10413 2567 10471 2573
rect 10413 2564 10425 2567
rect 9548 2536 10425 2564
rect 9548 2524 9554 2536
rect 10413 2533 10425 2536
rect 10459 2533 10471 2567
rect 10413 2527 10471 2533
rect 11146 2524 11152 2576
rect 11204 2564 11210 2576
rect 12161 2567 12219 2573
rect 12161 2564 12173 2567
rect 11204 2536 12173 2564
rect 11204 2524 11210 2536
rect 12161 2533 12173 2536
rect 12207 2533 12219 2567
rect 12161 2527 12219 2533
rect 8076 2468 8616 2496
rect 8076 2456 8082 2468
rect 9398 2456 9404 2508
rect 9456 2496 9462 2508
rect 9585 2499 9643 2505
rect 9585 2496 9597 2499
rect 9456 2468 9597 2496
rect 9456 2456 9462 2468
rect 9585 2465 9597 2468
rect 9631 2496 9643 2499
rect 9674 2496 9680 2508
rect 9631 2468 9680 2496
rect 9631 2465 9643 2468
rect 9585 2459 9643 2465
rect 9674 2456 9680 2468
rect 9732 2496 9738 2508
rect 10505 2499 10563 2505
rect 10505 2496 10517 2499
rect 9732 2468 10517 2496
rect 9732 2456 9738 2468
rect 10505 2465 10517 2468
rect 10551 2465 10563 2499
rect 12618 2496 12624 2508
rect 12579 2468 12624 2496
rect 10505 2459 10563 2465
rect 12618 2456 12624 2468
rect 12676 2496 12682 2508
rect 13173 2499 13231 2505
rect 13173 2496 13185 2499
rect 12676 2468 13185 2496
rect 12676 2456 12682 2468
rect 13173 2465 13185 2468
rect 13219 2465 13231 2499
rect 13173 2459 13231 2465
rect 4724 2400 7696 2428
rect 8665 2431 8723 2437
rect 4617 2391 4675 2397
rect 8665 2397 8677 2431
rect 8711 2397 8723 2431
rect 8665 2391 8723 2397
rect 10689 2431 10747 2437
rect 10689 2397 10701 2431
rect 10735 2428 10747 2431
rect 11422 2428 11428 2440
rect 10735 2400 11428 2428
rect 10735 2397 10747 2400
rect 10689 2391 10747 2397
rect 2004 2332 3004 2360
rect 2004 2320 2010 2332
rect 3970 2320 3976 2372
rect 4028 2360 4034 2372
rect 5813 2363 5871 2369
rect 5813 2360 5825 2363
rect 4028 2332 5825 2360
rect 4028 2320 4034 2332
rect 5813 2329 5825 2332
rect 5859 2329 5871 2363
rect 5813 2323 5871 2329
rect 8386 2320 8392 2372
rect 8444 2360 8450 2372
rect 8680 2360 8708 2391
rect 11422 2388 11428 2400
rect 11480 2388 11486 2440
rect 12802 2360 12808 2372
rect 8444 2332 8708 2360
rect 12763 2332 12808 2360
rect 8444 2320 8450 2332
rect 12802 2320 12808 2332
rect 12860 2320 12866 2372
rect 7098 2292 7104 2304
rect 7059 2264 7104 2292
rect 7098 2252 7104 2264
rect 7156 2252 7162 2304
rect 1104 2202 14812 2224
rect 1104 2150 3648 2202
rect 3700 2150 3712 2202
rect 3764 2150 3776 2202
rect 3828 2150 3840 2202
rect 3892 2150 8982 2202
rect 9034 2150 9046 2202
rect 9098 2150 9110 2202
rect 9162 2150 9174 2202
rect 9226 2150 14315 2202
rect 14367 2150 14379 2202
rect 14431 2150 14443 2202
rect 14495 2150 14507 2202
rect 14559 2150 14812 2202
rect 1104 2128 14812 2150
rect 9950 620 9956 672
rect 10008 660 10014 672
rect 10008 632 11008 660
rect 10008 620 10014 632
rect 10980 604 11008 632
rect 9858 552 9864 604
rect 9916 592 9922 604
rect 10594 592 10600 604
rect 9916 564 10600 592
rect 9916 552 9922 564
rect 10594 552 10600 564
rect 10652 552 10658 604
rect 10962 552 10968 604
rect 11020 552 11026 604
<< via1 >>
rect 11152 37680 11204 37732
rect 11796 37680 11848 37732
rect 6315 37510 6367 37562
rect 6379 37510 6431 37562
rect 6443 37510 6495 37562
rect 6507 37510 6559 37562
rect 11648 37510 11700 37562
rect 11712 37510 11764 37562
rect 11776 37510 11828 37562
rect 11840 37510 11892 37562
rect 3648 36966 3700 37018
rect 3712 36966 3764 37018
rect 3776 36966 3828 37018
rect 3840 36966 3892 37018
rect 8982 36966 9034 37018
rect 9046 36966 9098 37018
rect 9110 36966 9162 37018
rect 9174 36966 9226 37018
rect 14315 36966 14367 37018
rect 14379 36966 14431 37018
rect 14443 36966 14495 37018
rect 14507 36966 14559 37018
rect 4528 36864 4580 36916
rect 7932 36524 7984 36576
rect 6315 36422 6367 36474
rect 6379 36422 6431 36474
rect 6443 36422 6495 36474
rect 6507 36422 6559 36474
rect 11648 36422 11700 36474
rect 11712 36422 11764 36474
rect 11776 36422 11828 36474
rect 11840 36422 11892 36474
rect 4988 36363 5040 36372
rect 4988 36329 4997 36363
rect 4997 36329 5031 36363
rect 5031 36329 5040 36363
rect 4988 36320 5040 36329
rect 6184 36320 6236 36372
rect 5080 36184 5132 36236
rect 6736 36184 6788 36236
rect 3648 35878 3700 35930
rect 3712 35878 3764 35930
rect 3776 35878 3828 35930
rect 3840 35878 3892 35930
rect 8982 35878 9034 35930
rect 9046 35878 9098 35930
rect 9110 35878 9162 35930
rect 9174 35878 9226 35930
rect 14315 35878 14367 35930
rect 14379 35878 14431 35930
rect 14443 35878 14495 35930
rect 14507 35878 14559 35930
rect 5356 35776 5408 35828
rect 5724 35776 5776 35828
rect 6920 35776 6972 35828
rect 7748 35776 7800 35828
rect 9864 35751 9916 35760
rect 9864 35717 9873 35751
rect 9873 35717 9907 35751
rect 9907 35717 9916 35751
rect 9864 35708 9916 35717
rect 4988 35504 5040 35556
rect 5080 35479 5132 35488
rect 5080 35445 5089 35479
rect 5089 35445 5123 35479
rect 5123 35445 5132 35479
rect 5080 35436 5132 35445
rect 6184 35479 6236 35488
rect 6184 35445 6193 35479
rect 6193 35445 6227 35479
rect 6227 35445 6236 35479
rect 6184 35436 6236 35445
rect 6736 35436 6788 35488
rect 7656 35479 7708 35488
rect 7656 35445 7665 35479
rect 7665 35445 7699 35479
rect 7699 35445 7708 35479
rect 7656 35436 7708 35445
rect 7840 35436 7892 35488
rect 8852 35479 8904 35488
rect 8852 35445 8861 35479
rect 8861 35445 8895 35479
rect 8895 35445 8904 35479
rect 8852 35436 8904 35445
rect 10048 35436 10100 35488
rect 6315 35334 6367 35386
rect 6379 35334 6431 35386
rect 6443 35334 6495 35386
rect 6507 35334 6559 35386
rect 11648 35334 11700 35386
rect 11712 35334 11764 35386
rect 11776 35334 11828 35386
rect 11840 35334 11892 35386
rect 572 35232 624 35284
rect 4252 35275 4304 35284
rect 4252 35241 4261 35275
rect 4261 35241 4295 35275
rect 4295 35241 4304 35275
rect 4252 35232 4304 35241
rect 6644 35232 6696 35284
rect 7380 35232 7432 35284
rect 9772 35232 9824 35284
rect 10600 35232 10652 35284
rect 1952 35096 2004 35148
rect 2504 35139 2556 35148
rect 2504 35105 2513 35139
rect 2513 35105 2547 35139
rect 2547 35105 2556 35139
rect 2504 35096 2556 35105
rect 4068 35139 4120 35148
rect 4068 35105 4077 35139
rect 4077 35105 4111 35139
rect 4111 35105 4120 35139
rect 4068 35096 4120 35105
rect 5448 35139 5500 35148
rect 5448 35105 5457 35139
rect 5457 35105 5491 35139
rect 5491 35105 5500 35139
rect 5448 35096 5500 35105
rect 6920 35139 6972 35148
rect 6920 35105 6929 35139
rect 6929 35105 6963 35139
rect 6963 35105 6972 35139
rect 6920 35096 6972 35105
rect 7380 35096 7432 35148
rect 9312 35096 9364 35148
rect 7012 35071 7064 35080
rect 7012 35037 7021 35071
rect 7021 35037 7055 35071
rect 7055 35037 7064 35071
rect 7012 35028 7064 35037
rect 1400 34960 1452 35012
rect 9772 35028 9824 35080
rect 9864 34960 9916 35012
rect 2044 34935 2096 34944
rect 2044 34901 2053 34935
rect 2053 34901 2087 34935
rect 2087 34901 2096 34935
rect 2044 34892 2096 34901
rect 5724 34892 5776 34944
rect 7748 34935 7800 34944
rect 7748 34901 7757 34935
rect 7757 34901 7791 34935
rect 7791 34901 7800 34935
rect 7748 34892 7800 34901
rect 10140 34892 10192 34944
rect 10232 34892 10284 34944
rect 3648 34790 3700 34842
rect 3712 34790 3764 34842
rect 3776 34790 3828 34842
rect 3840 34790 3892 34842
rect 8982 34790 9034 34842
rect 9046 34790 9098 34842
rect 9110 34790 9162 34842
rect 9174 34790 9226 34842
rect 14315 34790 14367 34842
rect 14379 34790 14431 34842
rect 14443 34790 14495 34842
rect 14507 34790 14559 34842
rect 1952 34688 2004 34740
rect 2504 34731 2556 34740
rect 2504 34697 2513 34731
rect 2513 34697 2547 34731
rect 2547 34697 2556 34731
rect 2504 34688 2556 34697
rect 3240 34731 3292 34740
rect 3240 34697 3249 34731
rect 3249 34697 3283 34731
rect 3283 34697 3292 34731
rect 3240 34688 3292 34697
rect 4344 34731 4396 34740
rect 4344 34697 4353 34731
rect 4353 34697 4387 34731
rect 4387 34697 4396 34731
rect 4344 34688 4396 34697
rect 6920 34688 6972 34740
rect 8300 34688 8352 34740
rect 9772 34731 9824 34740
rect 9772 34697 9781 34731
rect 9781 34697 9815 34731
rect 9815 34697 9824 34731
rect 9772 34688 9824 34697
rect 3700 34663 3752 34672
rect 1584 34595 1636 34604
rect 1584 34561 1593 34595
rect 1593 34561 1627 34595
rect 1627 34561 1636 34595
rect 1584 34552 1636 34561
rect 2044 34552 2096 34604
rect 1768 34484 1820 34536
rect 3700 34629 3709 34663
rect 3709 34629 3743 34663
rect 3743 34629 3752 34663
rect 3700 34620 3752 34629
rect 3976 34620 4028 34672
rect 9864 34620 9916 34672
rect 3332 34552 3384 34604
rect 4344 34552 4396 34604
rect 4068 34527 4120 34536
rect 4068 34493 4077 34527
rect 4077 34493 4111 34527
rect 4111 34493 4120 34527
rect 4068 34484 4120 34493
rect 4252 34484 4304 34536
rect 2780 34416 2832 34468
rect 5448 34484 5500 34536
rect 7012 34527 7064 34536
rect 7012 34493 7021 34527
rect 7021 34493 7055 34527
rect 7055 34493 7064 34527
rect 7012 34484 7064 34493
rect 7380 34484 7432 34536
rect 7748 34484 7800 34536
rect 7840 34416 7892 34468
rect 8116 34416 8168 34468
rect 8760 34416 8812 34468
rect 10232 34416 10284 34468
rect 5264 34348 5316 34400
rect 7748 34348 7800 34400
rect 8208 34348 8260 34400
rect 9312 34391 9364 34400
rect 9312 34357 9321 34391
rect 9321 34357 9355 34391
rect 9355 34357 9364 34391
rect 9312 34348 9364 34357
rect 12164 34348 12216 34400
rect 6315 34246 6367 34298
rect 6379 34246 6431 34298
rect 6443 34246 6495 34298
rect 6507 34246 6559 34298
rect 11648 34246 11700 34298
rect 11712 34246 11764 34298
rect 11776 34246 11828 34298
rect 11840 34246 11892 34298
rect 2780 34144 2832 34196
rect 4344 34144 4396 34196
rect 6000 34187 6052 34196
rect 6000 34153 6009 34187
rect 6009 34153 6043 34187
rect 6043 34153 6052 34187
rect 6000 34144 6052 34153
rect 8760 34187 8812 34196
rect 8760 34153 8769 34187
rect 8769 34153 8803 34187
rect 8803 34153 8812 34187
rect 8760 34144 8812 34153
rect 9864 34187 9916 34196
rect 9864 34153 9873 34187
rect 9873 34153 9907 34187
rect 9907 34153 9916 34187
rect 9864 34144 9916 34153
rect 1492 34076 1544 34128
rect 5908 34119 5960 34128
rect 5908 34085 5917 34119
rect 5917 34085 5951 34119
rect 5951 34085 5960 34119
rect 5908 34076 5960 34085
rect 7564 34076 7616 34128
rect 12440 34076 12492 34128
rect 12716 34076 12768 34128
rect 2412 34008 2464 34060
rect 3056 34008 3108 34060
rect 3976 34008 4028 34060
rect 8116 34008 8168 34060
rect 10784 34051 10836 34060
rect 10784 34017 10793 34051
rect 10793 34017 10827 34051
rect 10827 34017 10836 34051
rect 10784 34008 10836 34017
rect 12348 34051 12400 34060
rect 12348 34017 12357 34051
rect 12357 34017 12391 34051
rect 12391 34017 12400 34051
rect 12348 34008 12400 34017
rect 6092 33983 6144 33992
rect 6092 33949 6101 33983
rect 6101 33949 6135 33983
rect 6135 33949 6144 33983
rect 6092 33940 6144 33949
rect 10876 33983 10928 33992
rect 10876 33949 10885 33983
rect 10885 33949 10919 33983
rect 10919 33949 10928 33983
rect 10876 33940 10928 33949
rect 7288 33872 7340 33924
rect 10692 33872 10744 33924
rect 11428 33940 11480 33992
rect 12256 33940 12308 33992
rect 5632 33804 5684 33856
rect 6092 33804 6144 33856
rect 7104 33804 7156 33856
rect 9404 33847 9456 33856
rect 9404 33813 9413 33847
rect 9413 33813 9447 33847
rect 9447 33813 9456 33847
rect 9404 33804 9456 33813
rect 9680 33804 9732 33856
rect 10784 33804 10836 33856
rect 12256 33804 12308 33856
rect 3648 33702 3700 33754
rect 3712 33702 3764 33754
rect 3776 33702 3828 33754
rect 3840 33702 3892 33754
rect 8982 33702 9034 33754
rect 9046 33702 9098 33754
rect 9110 33702 9162 33754
rect 9174 33702 9226 33754
rect 14315 33702 14367 33754
rect 14379 33702 14431 33754
rect 14443 33702 14495 33754
rect 14507 33702 14559 33754
rect 940 33600 992 33652
rect 6000 33600 6052 33652
rect 6552 33643 6604 33652
rect 6552 33609 6561 33643
rect 6561 33609 6595 33643
rect 6595 33609 6604 33643
rect 6552 33600 6604 33609
rect 2412 33575 2464 33584
rect 2412 33541 2421 33575
rect 2421 33541 2455 33575
rect 2455 33541 2464 33575
rect 2412 33532 2464 33541
rect 7104 33532 7156 33584
rect 9312 33575 9364 33584
rect 5908 33464 5960 33516
rect 7288 33507 7340 33516
rect 7288 33473 7297 33507
rect 7297 33473 7331 33507
rect 7331 33473 7340 33507
rect 7288 33464 7340 33473
rect 9312 33541 9321 33575
rect 9321 33541 9355 33575
rect 9355 33541 9364 33575
rect 9312 33532 9364 33541
rect 10876 33575 10928 33584
rect 10876 33541 10885 33575
rect 10885 33541 10919 33575
rect 10919 33541 10928 33575
rect 10876 33532 10928 33541
rect 9772 33464 9824 33516
rect 1952 33439 2004 33448
rect 1952 33405 1961 33439
rect 1961 33405 1995 33439
rect 1995 33405 2004 33439
rect 1952 33396 2004 33405
rect 5356 33396 5408 33448
rect 6552 33396 6604 33448
rect 7196 33439 7248 33448
rect 7196 33405 7205 33439
rect 7205 33405 7239 33439
rect 7239 33405 7248 33439
rect 7196 33396 7248 33405
rect 9680 33439 9732 33448
rect 9680 33405 9689 33439
rect 9689 33405 9723 33439
rect 9723 33405 9732 33439
rect 9680 33396 9732 33405
rect 11244 33396 11296 33448
rect 12900 33464 12952 33516
rect 4712 33328 4764 33380
rect 9404 33328 9456 33380
rect 12348 33328 12400 33380
rect 12716 33328 12768 33380
rect 13176 33328 13228 33380
rect 3056 33260 3108 33312
rect 3976 33303 4028 33312
rect 3976 33269 3985 33303
rect 3985 33269 4019 33303
rect 4019 33269 4028 33303
rect 3976 33260 4028 33269
rect 5632 33260 5684 33312
rect 6828 33303 6880 33312
rect 6828 33269 6837 33303
rect 6837 33269 6871 33303
rect 6871 33269 6880 33303
rect 6828 33260 6880 33269
rect 7288 33260 7340 33312
rect 7564 33260 7616 33312
rect 8116 33260 8168 33312
rect 9588 33260 9640 33312
rect 9864 33260 9916 33312
rect 10692 33260 10744 33312
rect 10876 33260 10928 33312
rect 11428 33260 11480 33312
rect 6315 33158 6367 33210
rect 6379 33158 6431 33210
rect 6443 33158 6495 33210
rect 6507 33158 6559 33210
rect 11648 33158 11700 33210
rect 11712 33158 11764 33210
rect 11776 33158 11828 33210
rect 11840 33158 11892 33210
rect 4160 33056 4212 33108
rect 5540 33056 5592 33108
rect 6828 33056 6880 33108
rect 7564 33056 7616 33108
rect 9312 33056 9364 33108
rect 10784 33056 10836 33108
rect 10876 33056 10928 33108
rect 12348 33056 12400 33108
rect 12716 33056 12768 33108
rect 12900 33099 12952 33108
rect 12900 33065 12909 33099
rect 12909 33065 12943 33099
rect 12943 33065 12952 33099
rect 12900 33056 12952 33065
rect 1676 33031 1728 33040
rect 1676 32997 1685 33031
rect 1685 32997 1719 33031
rect 1719 32997 1728 33031
rect 1676 32988 1728 32997
rect 1400 32963 1452 32972
rect 1400 32929 1409 32963
rect 1409 32929 1443 32963
rect 1443 32929 1452 32963
rect 1400 32920 1452 32929
rect 4160 32920 4212 32972
rect 5356 32963 5408 32972
rect 5356 32929 5365 32963
rect 5365 32929 5399 32963
rect 5399 32929 5408 32963
rect 5356 32920 5408 32929
rect 5632 32963 5684 32972
rect 5632 32929 5666 32963
rect 5666 32929 5684 32963
rect 5632 32920 5684 32929
rect 6184 32920 6236 32972
rect 7748 32920 7800 32972
rect 8116 32963 8168 32972
rect 8116 32929 8125 32963
rect 8125 32929 8159 32963
rect 8159 32929 8168 32963
rect 8116 32920 8168 32929
rect 8208 32963 8260 32972
rect 8208 32929 8217 32963
rect 8217 32929 8251 32963
rect 8251 32929 8260 32963
rect 8208 32920 8260 32929
rect 9680 32920 9732 32972
rect 10508 32963 10560 32972
rect 10508 32929 10542 32963
rect 10542 32929 10560 32963
rect 10508 32920 10560 32929
rect 12256 32920 12308 32972
rect 10232 32895 10284 32904
rect 10232 32861 10241 32895
rect 10241 32861 10275 32895
rect 10275 32861 10284 32895
rect 10232 32852 10284 32861
rect 12716 32852 12768 32904
rect 14648 32852 14700 32904
rect 6644 32784 6696 32836
rect 7104 32784 7156 32836
rect 8852 32784 8904 32836
rect 11520 32716 11572 32768
rect 3648 32614 3700 32666
rect 3712 32614 3764 32666
rect 3776 32614 3828 32666
rect 3840 32614 3892 32666
rect 8982 32614 9034 32666
rect 9046 32614 9098 32666
rect 9110 32614 9162 32666
rect 9174 32614 9226 32666
rect 14315 32614 14367 32666
rect 14379 32614 14431 32666
rect 14443 32614 14495 32666
rect 14507 32614 14559 32666
rect 1400 32512 1452 32564
rect 4160 32555 4212 32564
rect 4160 32521 4169 32555
rect 4169 32521 4203 32555
rect 4203 32521 4212 32555
rect 4160 32512 4212 32521
rect 5172 32555 5224 32564
rect 5172 32521 5181 32555
rect 5181 32521 5215 32555
rect 5215 32521 5224 32555
rect 5172 32512 5224 32521
rect 6184 32555 6236 32564
rect 6184 32521 6193 32555
rect 6193 32521 6227 32555
rect 6227 32521 6236 32555
rect 6184 32512 6236 32521
rect 6644 32555 6696 32564
rect 6644 32521 6653 32555
rect 6653 32521 6687 32555
rect 6687 32521 6696 32555
rect 6644 32512 6696 32521
rect 8116 32512 8168 32564
rect 8576 32555 8628 32564
rect 8576 32521 8585 32555
rect 8585 32521 8619 32555
rect 8619 32521 8628 32555
rect 8576 32512 8628 32521
rect 9680 32512 9732 32564
rect 8208 32487 8260 32496
rect 5540 32376 5592 32428
rect 7288 32376 7340 32428
rect 8208 32453 8217 32487
rect 8217 32453 8251 32487
rect 8251 32453 8260 32487
rect 8208 32444 8260 32453
rect 8300 32444 8352 32496
rect 9312 32419 9364 32428
rect 9312 32385 9321 32419
rect 9321 32385 9355 32419
rect 9355 32385 9364 32419
rect 9312 32376 9364 32385
rect 5264 32308 5316 32360
rect 8852 32308 8904 32360
rect 10508 32376 10560 32428
rect 12256 32512 12308 32564
rect 7748 32240 7800 32292
rect 9680 32240 9732 32292
rect 7472 32172 7524 32224
rect 8852 32172 8904 32224
rect 10324 32215 10376 32224
rect 10324 32181 10333 32215
rect 10333 32181 10367 32215
rect 10367 32181 10376 32215
rect 10324 32172 10376 32181
rect 6315 32070 6367 32122
rect 6379 32070 6431 32122
rect 6443 32070 6495 32122
rect 6507 32070 6559 32122
rect 11648 32070 11700 32122
rect 11712 32070 11764 32122
rect 11776 32070 11828 32122
rect 11840 32070 11892 32122
rect 5356 32011 5408 32020
rect 5356 31977 5365 32011
rect 5365 31977 5399 32011
rect 5399 31977 5408 32011
rect 5356 31968 5408 31977
rect 6184 31968 6236 32020
rect 7288 31968 7340 32020
rect 8576 32011 8628 32020
rect 8576 31977 8585 32011
rect 8585 31977 8619 32011
rect 8619 31977 8628 32011
rect 8576 31968 8628 31977
rect 9496 32011 9548 32020
rect 9496 31977 9505 32011
rect 9505 31977 9539 32011
rect 9539 31977 9548 32011
rect 9496 31968 9548 31977
rect 10324 31968 10376 32020
rect 10508 31968 10560 32020
rect 6644 31943 6696 31952
rect 6644 31909 6678 31943
rect 6678 31909 6696 31943
rect 6644 31900 6696 31909
rect 6920 31900 6972 31952
rect 10232 31900 10284 31952
rect 6184 31832 6236 31884
rect 10140 31875 10192 31884
rect 10140 31841 10149 31875
rect 10149 31841 10183 31875
rect 10183 31841 10192 31875
rect 10140 31832 10192 31841
rect 4896 31807 4948 31816
rect 4896 31773 4905 31807
rect 4905 31773 4939 31807
rect 4939 31773 4948 31807
rect 4896 31764 4948 31773
rect 10324 31807 10376 31816
rect 10324 31773 10333 31807
rect 10333 31773 10367 31807
rect 10367 31773 10376 31807
rect 10324 31764 10376 31773
rect 7012 31628 7064 31680
rect 8024 31671 8076 31680
rect 8024 31637 8033 31671
rect 8033 31637 8067 31671
rect 8067 31637 8076 31671
rect 8024 31628 8076 31637
rect 8852 31628 8904 31680
rect 9588 31628 9640 31680
rect 11520 31628 11572 31680
rect 3648 31526 3700 31578
rect 3712 31526 3764 31578
rect 3776 31526 3828 31578
rect 3840 31526 3892 31578
rect 8982 31526 9034 31578
rect 9046 31526 9098 31578
rect 9110 31526 9162 31578
rect 9174 31526 9226 31578
rect 14315 31526 14367 31578
rect 14379 31526 14431 31578
rect 14443 31526 14495 31578
rect 14507 31526 14559 31578
rect 8852 31424 8904 31476
rect 9404 31424 9456 31476
rect 6920 31356 6972 31408
rect 10324 31424 10376 31476
rect 9588 31356 9640 31408
rect 4160 31288 4212 31340
rect 5356 31331 5408 31340
rect 5356 31297 5365 31331
rect 5365 31297 5399 31331
rect 5399 31297 5408 31331
rect 5356 31288 5408 31297
rect 8024 31288 8076 31340
rect 9864 31331 9916 31340
rect 9864 31297 9873 31331
rect 9873 31297 9907 31331
rect 9907 31297 9916 31331
rect 9864 31288 9916 31297
rect 4896 31220 4948 31272
rect 8116 31263 8168 31272
rect 8116 31229 8125 31263
rect 8125 31229 8159 31263
rect 8159 31229 8168 31263
rect 8116 31220 8168 31229
rect 9496 31220 9548 31272
rect 5264 31195 5316 31204
rect 5264 31161 5273 31195
rect 5273 31161 5307 31195
rect 5307 31161 5316 31195
rect 5264 31152 5316 31161
rect 4804 31127 4856 31136
rect 4804 31093 4813 31127
rect 4813 31093 4847 31127
rect 4847 31093 4856 31127
rect 4804 31084 4856 31093
rect 6184 31084 6236 31136
rect 7104 31084 7156 31136
rect 7656 31152 7708 31204
rect 9680 31152 9732 31204
rect 9956 31152 10008 31204
rect 9588 31084 9640 31136
rect 10232 31127 10284 31136
rect 10232 31093 10241 31127
rect 10241 31093 10275 31127
rect 10275 31093 10284 31127
rect 10232 31084 10284 31093
rect 6315 30982 6367 31034
rect 6379 30982 6431 31034
rect 6443 30982 6495 31034
rect 6507 30982 6559 31034
rect 11648 30982 11700 31034
rect 11712 30982 11764 31034
rect 11776 30982 11828 31034
rect 11840 30982 11892 31034
rect 4896 30923 4948 30932
rect 4896 30889 4905 30923
rect 4905 30889 4939 30923
rect 4939 30889 4948 30923
rect 4896 30880 4948 30889
rect 8116 30880 8168 30932
rect 9312 30923 9364 30932
rect 9312 30889 9321 30923
rect 9321 30889 9355 30923
rect 9355 30889 9364 30923
rect 9312 30880 9364 30889
rect 10140 30880 10192 30932
rect 7472 30812 7524 30864
rect 8024 30812 8076 30864
rect 5080 30744 5132 30796
rect 5448 30787 5500 30796
rect 5448 30753 5457 30787
rect 5457 30753 5491 30787
rect 5491 30753 5500 30787
rect 5448 30744 5500 30753
rect 11980 30744 12032 30796
rect 5540 30719 5592 30728
rect 5540 30685 5549 30719
rect 5549 30685 5583 30719
rect 5583 30685 5592 30719
rect 5540 30676 5592 30685
rect 5356 30608 5408 30660
rect 2228 30540 2280 30592
rect 7288 30540 7340 30592
rect 10508 30540 10560 30592
rect 10784 30540 10836 30592
rect 11244 30540 11296 30592
rect 11520 30540 11572 30592
rect 12440 30540 12492 30592
rect 12900 30540 12952 30592
rect 3648 30438 3700 30490
rect 3712 30438 3764 30490
rect 3776 30438 3828 30490
rect 3840 30438 3892 30490
rect 8982 30438 9034 30490
rect 9046 30438 9098 30490
rect 9110 30438 9162 30490
rect 9174 30438 9226 30490
rect 14315 30438 14367 30490
rect 14379 30438 14431 30490
rect 14443 30438 14495 30490
rect 14507 30438 14559 30490
rect 10324 30336 10376 30388
rect 10692 30336 10744 30388
rect 4712 30311 4764 30320
rect 4712 30277 4721 30311
rect 4721 30277 4755 30311
rect 4755 30277 4764 30311
rect 4712 30268 4764 30277
rect 4804 30268 4856 30320
rect 10784 30311 10836 30320
rect 2412 30243 2464 30252
rect 2412 30209 2421 30243
rect 2421 30209 2455 30243
rect 2455 30209 2464 30243
rect 2412 30200 2464 30209
rect 5540 30200 5592 30252
rect 7288 30243 7340 30252
rect 7288 30209 7297 30243
rect 7297 30209 7331 30243
rect 7331 30209 7340 30243
rect 7288 30200 7340 30209
rect 10784 30277 10793 30311
rect 10793 30277 10827 30311
rect 10827 30277 10836 30311
rect 10784 30268 10836 30277
rect 10692 30243 10744 30252
rect 10692 30209 10701 30243
rect 10701 30209 10735 30243
rect 10735 30209 10744 30243
rect 12440 30268 12492 30320
rect 10692 30200 10744 30209
rect 13728 30200 13780 30252
rect 3332 30175 3384 30184
rect 3332 30141 3341 30175
rect 3341 30141 3375 30175
rect 3375 30141 3384 30175
rect 3332 30132 3384 30141
rect 7196 30175 7248 30184
rect 7196 30141 7205 30175
rect 7205 30141 7239 30175
rect 7239 30141 7248 30175
rect 7196 30132 7248 30141
rect 11244 30175 11296 30184
rect 11244 30141 11253 30175
rect 11253 30141 11287 30175
rect 11287 30141 11296 30175
rect 11244 30132 11296 30141
rect 12900 30132 12952 30184
rect 2136 30107 2188 30116
rect 2136 30073 2145 30107
rect 2145 30073 2179 30107
rect 2179 30073 2188 30107
rect 2136 30064 2188 30073
rect 4804 30064 4856 30116
rect 1768 30039 1820 30048
rect 1768 30005 1777 30039
rect 1777 30005 1811 30039
rect 1811 30005 1820 30039
rect 1768 29996 1820 30005
rect 2228 30039 2280 30048
rect 2228 30005 2237 30039
rect 2237 30005 2271 30039
rect 2271 30005 2280 30039
rect 2228 29996 2280 30005
rect 4528 29996 4580 30048
rect 5080 30039 5132 30048
rect 5080 30005 5089 30039
rect 5089 30005 5123 30039
rect 5123 30005 5132 30039
rect 5080 29996 5132 30005
rect 5632 29996 5684 30048
rect 6828 30039 6880 30048
rect 6828 30005 6837 30039
rect 6837 30005 6871 30039
rect 6871 30005 6880 30039
rect 6828 29996 6880 30005
rect 11152 30039 11204 30048
rect 11152 30005 11161 30039
rect 11161 30005 11195 30039
rect 11195 30005 11204 30039
rect 11152 29996 11204 30005
rect 11980 29996 12032 30048
rect 12532 29996 12584 30048
rect 12900 30039 12952 30048
rect 12900 30005 12909 30039
rect 12909 30005 12943 30039
rect 12943 30005 12952 30039
rect 12900 29996 12952 30005
rect 6315 29894 6367 29946
rect 6379 29894 6431 29946
rect 6443 29894 6495 29946
rect 6507 29894 6559 29946
rect 11648 29894 11700 29946
rect 11712 29894 11764 29946
rect 11776 29894 11828 29946
rect 11840 29894 11892 29946
rect 2136 29835 2188 29844
rect 2136 29801 2145 29835
rect 2145 29801 2179 29835
rect 2179 29801 2188 29835
rect 2136 29792 2188 29801
rect 4160 29835 4212 29844
rect 4160 29801 4169 29835
rect 4169 29801 4203 29835
rect 4203 29801 4212 29835
rect 4160 29792 4212 29801
rect 6644 29792 6696 29844
rect 7196 29792 7248 29844
rect 13728 29835 13780 29844
rect 13728 29801 13737 29835
rect 13737 29801 13771 29835
rect 13771 29801 13780 29835
rect 13728 29792 13780 29801
rect 1676 29767 1728 29776
rect 1676 29733 1685 29767
rect 1685 29733 1719 29767
rect 1719 29733 1728 29767
rect 1676 29724 1728 29733
rect 9312 29724 9364 29776
rect 1768 29656 1820 29708
rect 3332 29520 3384 29572
rect 4252 29520 4304 29572
rect 3516 29452 3568 29504
rect 4988 29656 5040 29708
rect 10232 29656 10284 29708
rect 4804 29631 4856 29640
rect 4804 29597 4813 29631
rect 4813 29597 4847 29631
rect 4847 29597 4856 29631
rect 4804 29588 4856 29597
rect 6000 29588 6052 29640
rect 6460 29631 6512 29640
rect 6460 29597 6469 29631
rect 6469 29597 6503 29631
rect 6503 29597 6512 29631
rect 12440 29656 12492 29708
rect 12992 29656 13044 29708
rect 6460 29588 6512 29597
rect 11520 29588 11572 29640
rect 12348 29631 12400 29640
rect 12348 29597 12357 29631
rect 12357 29597 12391 29631
rect 12391 29597 12400 29631
rect 12348 29588 12400 29597
rect 5908 29495 5960 29504
rect 5908 29461 5917 29495
rect 5917 29461 5951 29495
rect 5951 29461 5960 29495
rect 5908 29452 5960 29461
rect 8576 29452 8628 29504
rect 9956 29452 10008 29504
rect 3648 29350 3700 29402
rect 3712 29350 3764 29402
rect 3776 29350 3828 29402
rect 3840 29350 3892 29402
rect 8982 29350 9034 29402
rect 9046 29350 9098 29402
rect 9110 29350 9162 29402
rect 9174 29350 9226 29402
rect 14315 29350 14367 29402
rect 14379 29350 14431 29402
rect 14443 29350 14495 29402
rect 14507 29350 14559 29402
rect 1768 29248 1820 29300
rect 4804 29248 4856 29300
rect 6644 29248 6696 29300
rect 9312 29248 9364 29300
rect 9956 29291 10008 29300
rect 9956 29257 9965 29291
rect 9965 29257 9999 29291
rect 9999 29257 10008 29291
rect 9956 29248 10008 29257
rect 10968 29248 11020 29300
rect 8576 29155 8628 29164
rect 8576 29121 8585 29155
rect 8585 29121 8619 29155
rect 8619 29121 8628 29155
rect 8576 29112 8628 29121
rect 3424 29044 3476 29096
rect 6000 29087 6052 29096
rect 6000 29053 6009 29087
rect 6009 29053 6043 29087
rect 6043 29053 6052 29087
rect 6000 29044 6052 29053
rect 8300 29044 8352 29096
rect 9588 29112 9640 29164
rect 4068 28976 4120 29028
rect 5172 28976 5224 29028
rect 4620 28908 4672 28960
rect 5264 28908 5316 28960
rect 6460 28976 6512 29028
rect 11244 29248 11296 29300
rect 11244 29112 11296 29164
rect 11888 29180 11940 29232
rect 12348 29180 12400 29232
rect 11980 29112 12032 29164
rect 11520 28976 11572 29028
rect 7656 28951 7708 28960
rect 7656 28917 7665 28951
rect 7665 28917 7699 28951
rect 7699 28917 7708 28951
rect 7656 28908 7708 28917
rect 8116 28951 8168 28960
rect 8116 28917 8125 28951
rect 8125 28917 8159 28951
rect 8159 28917 8168 28951
rect 8116 28908 8168 28917
rect 9680 28908 9732 28960
rect 10968 28908 11020 28960
rect 12164 28976 12216 29028
rect 14188 29044 14240 29096
rect 6315 28806 6367 28858
rect 6379 28806 6431 28858
rect 6443 28806 6495 28858
rect 6507 28806 6559 28858
rect 11648 28806 11700 28858
rect 11712 28806 11764 28858
rect 11776 28806 11828 28858
rect 11840 28806 11892 28858
rect 3700 28747 3752 28756
rect 3700 28713 3709 28747
rect 3709 28713 3743 28747
rect 3743 28713 3752 28747
rect 3700 28704 3752 28713
rect 4068 28704 4120 28756
rect 4804 28704 4856 28756
rect 5540 28704 5592 28756
rect 7656 28704 7708 28756
rect 9588 28704 9640 28756
rect 11152 28704 11204 28756
rect 12072 28704 12124 28756
rect 12992 28747 13044 28756
rect 12992 28713 13001 28747
rect 13001 28713 13035 28747
rect 13035 28713 13044 28747
rect 12992 28704 13044 28713
rect 9680 28636 9732 28688
rect 10232 28636 10284 28688
rect 5264 28568 5316 28620
rect 8392 28611 8444 28620
rect 8392 28577 8401 28611
rect 8401 28577 8435 28611
rect 8435 28577 8444 28611
rect 8392 28568 8444 28577
rect 12348 28611 12400 28620
rect 12348 28577 12357 28611
rect 12357 28577 12391 28611
rect 12391 28577 12400 28611
rect 12348 28568 12400 28577
rect 8484 28543 8536 28552
rect 8484 28509 8493 28543
rect 8493 28509 8527 28543
rect 8527 28509 8536 28543
rect 8484 28500 8536 28509
rect 9404 28500 9456 28552
rect 9680 28543 9732 28552
rect 9680 28509 9689 28543
rect 9689 28509 9723 28543
rect 9723 28509 9732 28543
rect 9680 28500 9732 28509
rect 11980 28500 12032 28552
rect 12440 28500 12492 28552
rect 4988 28364 5040 28416
rect 5264 28407 5316 28416
rect 5264 28373 5273 28407
rect 5273 28373 5307 28407
rect 5307 28373 5316 28407
rect 5264 28364 5316 28373
rect 5448 28364 5500 28416
rect 6184 28364 6236 28416
rect 6828 28364 6880 28416
rect 3648 28262 3700 28314
rect 3712 28262 3764 28314
rect 3776 28262 3828 28314
rect 3840 28262 3892 28314
rect 8982 28262 9034 28314
rect 9046 28262 9098 28314
rect 9110 28262 9162 28314
rect 9174 28262 9226 28314
rect 14315 28262 14367 28314
rect 14379 28262 14431 28314
rect 14443 28262 14495 28314
rect 14507 28262 14559 28314
rect 3516 28160 3568 28212
rect 4252 28160 4304 28212
rect 5448 28160 5500 28212
rect 6000 28160 6052 28212
rect 6184 28160 6236 28212
rect 8576 28160 8628 28212
rect 10784 28203 10836 28212
rect 10784 28169 10793 28203
rect 10793 28169 10827 28203
rect 10827 28169 10836 28203
rect 10784 28160 10836 28169
rect 12072 28203 12124 28212
rect 12072 28169 12081 28203
rect 12081 28169 12115 28203
rect 12115 28169 12124 28203
rect 12072 28160 12124 28169
rect 8852 28135 8904 28144
rect 8852 28101 8861 28135
rect 8861 28101 8895 28135
rect 8895 28101 8904 28135
rect 8852 28092 8904 28101
rect 10692 28135 10744 28144
rect 10692 28101 10701 28135
rect 10701 28101 10735 28135
rect 10735 28101 10744 28135
rect 10692 28092 10744 28101
rect 1584 28067 1636 28076
rect 1584 28033 1593 28067
rect 1593 28033 1627 28067
rect 1627 28033 1636 28067
rect 1584 28024 1636 28033
rect 4068 28067 4120 28076
rect 4068 28033 4077 28067
rect 4077 28033 4111 28067
rect 4111 28033 4120 28067
rect 4068 28024 4120 28033
rect 4160 28067 4212 28076
rect 4160 28033 4169 28067
rect 4169 28033 4203 28067
rect 4203 28033 4212 28067
rect 4160 28024 4212 28033
rect 5264 28024 5316 28076
rect 6000 28024 6052 28076
rect 4620 27956 4672 28008
rect 5724 27956 5776 28008
rect 6828 27999 6880 28008
rect 6828 27965 6837 27999
rect 6837 27965 6871 27999
rect 6871 27965 6880 27999
rect 6828 27956 6880 27965
rect 9404 27956 9456 28008
rect 12072 28024 12124 28076
rect 12348 28024 12400 28076
rect 5080 27931 5132 27940
rect 5080 27897 5089 27931
rect 5089 27897 5123 27931
rect 5123 27897 5132 27931
rect 5080 27888 5132 27897
rect 5540 27931 5592 27940
rect 5540 27897 5549 27931
rect 5549 27897 5583 27931
rect 5583 27897 5592 27931
rect 5540 27888 5592 27897
rect 7012 27888 7064 27940
rect 8484 27888 8536 27940
rect 9588 27888 9640 27940
rect 11428 27888 11480 27940
rect 2228 27863 2280 27872
rect 2228 27829 2237 27863
rect 2237 27829 2271 27863
rect 2271 27829 2280 27863
rect 2228 27820 2280 27829
rect 5172 27863 5224 27872
rect 5172 27829 5181 27863
rect 5181 27829 5215 27863
rect 5215 27829 5224 27863
rect 5172 27820 5224 27829
rect 6000 27820 6052 27872
rect 8852 27820 8904 27872
rect 9312 27820 9364 27872
rect 9496 27863 9548 27872
rect 9496 27829 9505 27863
rect 9505 27829 9539 27863
rect 9539 27829 9548 27863
rect 11244 27863 11296 27872
rect 9496 27820 9548 27829
rect 11244 27829 11253 27863
rect 11253 27829 11287 27863
rect 11287 27829 11296 27863
rect 11244 27820 11296 27829
rect 6315 27718 6367 27770
rect 6379 27718 6431 27770
rect 6443 27718 6495 27770
rect 6507 27718 6559 27770
rect 11648 27718 11700 27770
rect 11712 27718 11764 27770
rect 11776 27718 11828 27770
rect 11840 27718 11892 27770
rect 4068 27616 4120 27668
rect 4712 27616 4764 27668
rect 5540 27616 5592 27668
rect 8392 27616 8444 27668
rect 3056 27548 3108 27600
rect 3332 27548 3384 27600
rect 11244 27616 11296 27668
rect 12072 27659 12124 27668
rect 12072 27625 12081 27659
rect 12081 27625 12115 27659
rect 12115 27625 12124 27659
rect 12072 27616 12124 27625
rect 12440 27659 12492 27668
rect 12440 27625 12449 27659
rect 12449 27625 12483 27659
rect 12483 27625 12492 27659
rect 12440 27616 12492 27625
rect 5816 27523 5868 27532
rect 5816 27489 5825 27523
rect 5825 27489 5859 27523
rect 5859 27489 5868 27523
rect 5816 27480 5868 27489
rect 6644 27480 6696 27532
rect 8208 27480 8260 27532
rect 5540 27412 5592 27464
rect 6000 27455 6052 27464
rect 6000 27421 6009 27455
rect 6009 27421 6043 27455
rect 6043 27421 6052 27455
rect 6000 27412 6052 27421
rect 6828 27412 6880 27464
rect 5356 27276 5408 27328
rect 8208 27276 8260 27328
rect 8392 27319 8444 27328
rect 8392 27285 8401 27319
rect 8401 27285 8435 27319
rect 8435 27285 8444 27319
rect 8392 27276 8444 27285
rect 8668 27276 8720 27328
rect 9496 27276 9548 27328
rect 10232 27319 10284 27328
rect 10232 27285 10241 27319
rect 10241 27285 10275 27319
rect 10275 27285 10284 27319
rect 10232 27276 10284 27285
rect 10692 27319 10744 27328
rect 10692 27285 10701 27319
rect 10701 27285 10735 27319
rect 10735 27285 10744 27319
rect 10692 27276 10744 27285
rect 11428 27319 11480 27328
rect 11428 27285 11437 27319
rect 11437 27285 11471 27319
rect 11471 27285 11480 27319
rect 11428 27276 11480 27285
rect 3648 27174 3700 27226
rect 3712 27174 3764 27226
rect 3776 27174 3828 27226
rect 3840 27174 3892 27226
rect 8982 27174 9034 27226
rect 9046 27174 9098 27226
rect 9110 27174 9162 27226
rect 9174 27174 9226 27226
rect 14315 27174 14367 27226
rect 14379 27174 14431 27226
rect 14443 27174 14495 27226
rect 14507 27174 14559 27226
rect 4988 27115 5040 27124
rect 4988 27081 4997 27115
rect 4997 27081 5031 27115
rect 5031 27081 5040 27115
rect 4988 27072 5040 27081
rect 6644 27115 6696 27124
rect 6644 27081 6653 27115
rect 6653 27081 6687 27115
rect 6687 27081 6696 27115
rect 6644 27072 6696 27081
rect 7012 27115 7064 27124
rect 7012 27081 7021 27115
rect 7021 27081 7055 27115
rect 7055 27081 7064 27115
rect 7012 27072 7064 27081
rect 7196 27115 7248 27124
rect 7196 27081 7205 27115
rect 7205 27081 7239 27115
rect 7239 27081 7248 27115
rect 7196 27072 7248 27081
rect 8208 27115 8260 27124
rect 8208 27081 8217 27115
rect 8217 27081 8251 27115
rect 8251 27081 8260 27115
rect 8208 27072 8260 27081
rect 11244 27072 11296 27124
rect 12808 27072 12860 27124
rect 6000 27004 6052 27056
rect 5172 26936 5224 26988
rect 5356 26911 5408 26920
rect 5356 26877 5365 26911
rect 5365 26877 5399 26911
rect 5399 26877 5408 26911
rect 5356 26868 5408 26877
rect 8392 26936 8444 26988
rect 12440 26936 12492 26988
rect 7564 26911 7616 26920
rect 4988 26800 5040 26852
rect 7564 26877 7573 26911
rect 7573 26877 7607 26911
rect 7607 26877 7616 26911
rect 7564 26868 7616 26877
rect 8116 26868 8168 26920
rect 12900 26868 12952 26920
rect 7288 26800 7340 26852
rect 5540 26732 5592 26784
rect 10140 26775 10192 26784
rect 10140 26741 10149 26775
rect 10149 26741 10183 26775
rect 10183 26741 10192 26775
rect 10140 26732 10192 26741
rect 10692 26732 10744 26784
rect 6315 26630 6367 26682
rect 6379 26630 6431 26682
rect 6443 26630 6495 26682
rect 6507 26630 6559 26682
rect 11648 26630 11700 26682
rect 11712 26630 11764 26682
rect 11776 26630 11828 26682
rect 11840 26630 11892 26682
rect 4068 26528 4120 26580
rect 4988 26571 5040 26580
rect 4988 26537 4997 26571
rect 4997 26537 5031 26571
rect 5031 26537 5040 26571
rect 4988 26528 5040 26537
rect 7564 26571 7616 26580
rect 7564 26537 7573 26571
rect 7573 26537 7607 26571
rect 7607 26537 7616 26571
rect 7564 26528 7616 26537
rect 10140 26528 10192 26580
rect 11428 26528 11480 26580
rect 12992 26528 13044 26580
rect 10324 26460 10376 26512
rect 10784 26503 10836 26512
rect 10784 26469 10793 26503
rect 10793 26469 10827 26503
rect 10827 26469 10836 26503
rect 10784 26460 10836 26469
rect 10416 26392 10468 26444
rect 11152 26392 11204 26444
rect 11980 26392 12032 26444
rect 11060 26324 11112 26376
rect 12440 26324 12492 26376
rect 9404 26256 9456 26308
rect 5816 26188 5868 26240
rect 7012 26188 7064 26240
rect 7288 26231 7340 26240
rect 7288 26197 7297 26231
rect 7297 26197 7331 26231
rect 7331 26197 7340 26231
rect 7288 26188 7340 26197
rect 8576 26231 8628 26240
rect 8576 26197 8585 26231
rect 8585 26197 8619 26231
rect 8619 26197 8628 26231
rect 8576 26188 8628 26197
rect 9588 26188 9640 26240
rect 3648 26086 3700 26138
rect 3712 26086 3764 26138
rect 3776 26086 3828 26138
rect 3840 26086 3892 26138
rect 8982 26086 9034 26138
rect 9046 26086 9098 26138
rect 9110 26086 9162 26138
rect 9174 26086 9226 26138
rect 14315 26086 14367 26138
rect 14379 26086 14431 26138
rect 14443 26086 14495 26138
rect 14507 26086 14559 26138
rect 6828 25984 6880 26036
rect 10232 25984 10284 26036
rect 10692 25984 10744 26036
rect 10784 25984 10836 26036
rect 11980 26027 12032 26036
rect 11980 25993 11989 26027
rect 11989 25993 12023 26027
rect 12023 25993 12032 26027
rect 11980 25984 12032 25993
rect 12440 25984 12492 26036
rect 10968 25916 11020 25968
rect 11152 25916 11204 25968
rect 9312 25891 9364 25900
rect 9312 25857 9321 25891
rect 9321 25857 9355 25891
rect 9355 25857 9364 25891
rect 9312 25848 9364 25857
rect 9404 25848 9456 25900
rect 9772 25848 9824 25900
rect 11060 25891 11112 25900
rect 11060 25857 11069 25891
rect 11069 25857 11103 25891
rect 11103 25857 11112 25891
rect 11060 25848 11112 25857
rect 5632 25780 5684 25832
rect 8576 25780 8628 25832
rect 10416 25780 10468 25832
rect 10508 25780 10560 25832
rect 9588 25712 9640 25764
rect 10600 25712 10652 25764
rect 10968 25712 11020 25764
rect 6000 25644 6052 25696
rect 6184 25644 6236 25696
rect 8852 25687 8904 25696
rect 8852 25653 8861 25687
rect 8861 25653 8895 25687
rect 8895 25653 8904 25687
rect 8852 25644 8904 25653
rect 9956 25644 10008 25696
rect 11244 25644 11296 25696
rect 12992 25687 13044 25696
rect 12992 25653 13001 25687
rect 13001 25653 13035 25687
rect 13035 25653 13044 25687
rect 12992 25644 13044 25653
rect 6315 25542 6367 25594
rect 6379 25542 6431 25594
rect 6443 25542 6495 25594
rect 6507 25542 6559 25594
rect 11648 25542 11700 25594
rect 11712 25542 11764 25594
rect 11776 25542 11828 25594
rect 11840 25542 11892 25594
rect 7288 25440 7340 25492
rect 8852 25440 8904 25492
rect 9312 25440 9364 25492
rect 10508 25440 10560 25492
rect 11060 25483 11112 25492
rect 11060 25449 11069 25483
rect 11069 25449 11103 25483
rect 11103 25449 11112 25483
rect 11060 25440 11112 25449
rect 12440 25440 12492 25492
rect 4344 25415 4396 25424
rect 4344 25381 4353 25415
rect 4353 25381 4387 25415
rect 4387 25381 4396 25415
rect 4344 25372 4396 25381
rect 6184 25415 6236 25424
rect 6184 25381 6193 25415
rect 6193 25381 6227 25415
rect 6227 25381 6236 25415
rect 6184 25372 6236 25381
rect 9956 25372 10008 25424
rect 11428 25372 11480 25424
rect 4068 25347 4120 25356
rect 4068 25313 4077 25347
rect 4077 25313 4111 25347
rect 4111 25313 4120 25347
rect 4068 25304 4120 25313
rect 6828 25304 6880 25356
rect 7564 25304 7616 25356
rect 10232 25304 10284 25356
rect 11888 25304 11940 25356
rect 6276 25279 6328 25288
rect 6276 25245 6285 25279
rect 6285 25245 6319 25279
rect 6319 25245 6328 25279
rect 6276 25236 6328 25245
rect 8300 25236 8352 25288
rect 10324 25279 10376 25288
rect 10324 25245 10333 25279
rect 10333 25245 10367 25279
rect 10367 25245 10376 25279
rect 10324 25236 10376 25245
rect 5264 25100 5316 25152
rect 5540 25100 5592 25152
rect 7656 25143 7708 25152
rect 7656 25109 7665 25143
rect 7665 25109 7699 25143
rect 7699 25109 7708 25143
rect 7656 25100 7708 25109
rect 3648 24998 3700 25050
rect 3712 24998 3764 25050
rect 3776 24998 3828 25050
rect 3840 24998 3892 25050
rect 8982 24998 9034 25050
rect 9046 24998 9098 25050
rect 9110 24998 9162 25050
rect 9174 24998 9226 25050
rect 14315 24998 14367 25050
rect 14379 24998 14431 25050
rect 14443 24998 14495 25050
rect 14507 24998 14559 25050
rect 6184 24939 6236 24948
rect 6184 24905 6193 24939
rect 6193 24905 6227 24939
rect 6227 24905 6236 24939
rect 6184 24896 6236 24905
rect 7564 24939 7616 24948
rect 7564 24905 7573 24939
rect 7573 24905 7607 24939
rect 7607 24905 7616 24939
rect 7564 24896 7616 24905
rect 6276 24828 6328 24880
rect 6736 24828 6788 24880
rect 7656 24828 7708 24880
rect 9772 24896 9824 24948
rect 10508 24896 10560 24948
rect 10692 24896 10744 24948
rect 11428 24896 11480 24948
rect 11888 24939 11940 24948
rect 11888 24905 11897 24939
rect 11897 24905 11931 24939
rect 11931 24905 11940 24939
rect 11888 24896 11940 24905
rect 5356 24803 5408 24812
rect 5356 24769 5365 24803
rect 5365 24769 5399 24803
rect 5399 24769 5408 24803
rect 5356 24760 5408 24769
rect 8300 24760 8352 24812
rect 8760 24760 8812 24812
rect 5448 24692 5500 24744
rect 7932 24735 7984 24744
rect 7932 24701 7941 24735
rect 7941 24701 7975 24735
rect 7975 24701 7984 24735
rect 7932 24692 7984 24701
rect 4068 24624 4120 24676
rect 10324 24760 10376 24812
rect 9128 24735 9180 24744
rect 9128 24701 9137 24735
rect 9137 24701 9171 24735
rect 9171 24701 9180 24735
rect 9128 24692 9180 24701
rect 9220 24692 9272 24744
rect 9312 24624 9364 24676
rect 5264 24599 5316 24608
rect 5264 24565 5273 24599
rect 5273 24565 5307 24599
rect 5307 24565 5316 24599
rect 5264 24556 5316 24565
rect 6828 24556 6880 24608
rect 8024 24599 8076 24608
rect 8024 24565 8033 24599
rect 8033 24565 8067 24599
rect 8067 24565 8076 24599
rect 8024 24556 8076 24565
rect 9772 24556 9824 24608
rect 6315 24454 6367 24506
rect 6379 24454 6431 24506
rect 6443 24454 6495 24506
rect 6507 24454 6559 24506
rect 11648 24454 11700 24506
rect 11712 24454 11764 24506
rect 11776 24454 11828 24506
rect 11840 24454 11892 24506
rect 6184 24352 6236 24404
rect 6736 24352 6788 24404
rect 7564 24352 7616 24404
rect 9220 24352 9272 24404
rect 9680 24395 9732 24404
rect 9680 24361 9689 24395
rect 9689 24361 9723 24395
rect 9723 24361 9732 24395
rect 9680 24352 9732 24361
rect 11244 24395 11296 24404
rect 11244 24361 11253 24395
rect 11253 24361 11287 24395
rect 11287 24361 11296 24395
rect 11244 24352 11296 24361
rect 12256 24352 12308 24404
rect 6276 24327 6328 24336
rect 6276 24293 6285 24327
rect 6285 24293 6319 24327
rect 6319 24293 6328 24327
rect 6276 24284 6328 24293
rect 6920 24284 6972 24336
rect 7472 24284 7524 24336
rect 10784 24284 10836 24336
rect 11428 24284 11480 24336
rect 6092 24216 6144 24268
rect 4804 24191 4856 24200
rect 4804 24157 4813 24191
rect 4813 24157 4847 24191
rect 4847 24157 4856 24191
rect 4804 24148 4856 24157
rect 5540 24148 5592 24200
rect 4436 24055 4488 24064
rect 4436 24021 4445 24055
rect 4445 24021 4479 24055
rect 4479 24021 4488 24055
rect 4436 24012 4488 24021
rect 7196 24012 7248 24064
rect 9956 24148 10008 24200
rect 10416 24216 10468 24268
rect 10324 24191 10376 24200
rect 10324 24157 10333 24191
rect 10333 24157 10367 24191
rect 10367 24157 10376 24191
rect 10324 24148 10376 24157
rect 11520 24148 11572 24200
rect 9128 24080 9180 24132
rect 8392 24012 8444 24064
rect 3648 23910 3700 23962
rect 3712 23910 3764 23962
rect 3776 23910 3828 23962
rect 3840 23910 3892 23962
rect 8982 23910 9034 23962
rect 9046 23910 9098 23962
rect 9110 23910 9162 23962
rect 9174 23910 9226 23962
rect 14315 23910 14367 23962
rect 14379 23910 14431 23962
rect 14443 23910 14495 23962
rect 14507 23910 14559 23962
rect 5816 23808 5868 23860
rect 6092 23808 6144 23860
rect 6276 23851 6328 23860
rect 6276 23817 6285 23851
rect 6285 23817 6319 23851
rect 6319 23817 6328 23851
rect 6276 23808 6328 23817
rect 7472 23808 7524 23860
rect 5632 23740 5684 23792
rect 6736 23740 6788 23792
rect 8024 23808 8076 23860
rect 10508 23851 10560 23860
rect 10508 23817 10517 23851
rect 10517 23817 10551 23851
rect 10551 23817 10560 23851
rect 10508 23808 10560 23817
rect 10784 23808 10836 23860
rect 11152 23808 11204 23860
rect 11428 23808 11480 23860
rect 11520 23808 11572 23860
rect 8852 23783 8904 23792
rect 8852 23749 8861 23783
rect 8861 23749 8895 23783
rect 8895 23749 8904 23783
rect 8852 23740 8904 23749
rect 4436 23672 4488 23724
rect 5724 23672 5776 23724
rect 6092 23672 6144 23724
rect 12256 23740 12308 23792
rect 4712 23579 4764 23588
rect 4712 23545 4721 23579
rect 4721 23545 4755 23579
rect 4755 23545 4764 23579
rect 4712 23536 4764 23545
rect 9864 23672 9916 23724
rect 10324 23672 10376 23724
rect 10784 23672 10836 23724
rect 11060 23672 11112 23724
rect 11428 23672 11480 23724
rect 9404 23647 9456 23656
rect 5080 23536 5132 23588
rect 5448 23536 5500 23588
rect 5724 23536 5776 23588
rect 6552 23536 6604 23588
rect 4344 23511 4396 23520
rect 4344 23477 4353 23511
rect 4353 23477 4387 23511
rect 4387 23477 4396 23511
rect 4344 23468 4396 23477
rect 5540 23511 5592 23520
rect 5540 23477 5549 23511
rect 5549 23477 5583 23511
rect 5583 23477 5592 23511
rect 5540 23468 5592 23477
rect 9404 23613 9413 23647
rect 9413 23613 9447 23647
rect 9447 23613 9456 23647
rect 9404 23604 9456 23613
rect 7196 23536 7248 23588
rect 7564 23468 7616 23520
rect 9956 23468 10008 23520
rect 6315 23366 6367 23418
rect 6379 23366 6431 23418
rect 6443 23366 6495 23418
rect 6507 23366 6559 23418
rect 11648 23366 11700 23418
rect 11712 23366 11764 23418
rect 11776 23366 11828 23418
rect 11840 23366 11892 23418
rect 4712 23264 4764 23316
rect 6644 23307 6696 23316
rect 6644 23273 6653 23307
rect 6653 23273 6687 23307
rect 6687 23273 6696 23307
rect 6644 23264 6696 23273
rect 6920 23307 6972 23316
rect 6920 23273 6929 23307
rect 6929 23273 6963 23307
rect 6963 23273 6972 23307
rect 6920 23264 6972 23273
rect 7472 23307 7524 23316
rect 7472 23273 7481 23307
rect 7481 23273 7515 23307
rect 7515 23273 7524 23307
rect 7472 23264 7524 23273
rect 9404 23264 9456 23316
rect 9864 23307 9916 23316
rect 9864 23273 9873 23307
rect 9873 23273 9907 23307
rect 9907 23273 9916 23307
rect 9864 23264 9916 23273
rect 5540 23239 5592 23248
rect 5540 23205 5574 23239
rect 5574 23205 5592 23239
rect 5540 23196 5592 23205
rect 5632 23196 5684 23248
rect 4068 23128 4120 23180
rect 7840 23171 7892 23180
rect 7840 23137 7849 23171
rect 7849 23137 7883 23171
rect 7883 23137 7892 23171
rect 7840 23128 7892 23137
rect 8208 23128 8260 23180
rect 4252 22924 4304 22976
rect 6644 23060 6696 23112
rect 8024 23103 8076 23112
rect 8024 23069 8033 23103
rect 8033 23069 8067 23103
rect 8067 23069 8076 23103
rect 8024 23060 8076 23069
rect 7472 22924 7524 22976
rect 8392 22924 8444 22976
rect 3648 22822 3700 22874
rect 3712 22822 3764 22874
rect 3776 22822 3828 22874
rect 3840 22822 3892 22874
rect 8982 22822 9034 22874
rect 9046 22822 9098 22874
rect 9110 22822 9162 22874
rect 9174 22822 9226 22874
rect 14315 22822 14367 22874
rect 14379 22822 14431 22874
rect 14443 22822 14495 22874
rect 14507 22822 14559 22874
rect 3424 22763 3476 22772
rect 3424 22729 3433 22763
rect 3433 22729 3467 22763
rect 3467 22729 3476 22763
rect 3424 22720 3476 22729
rect 4068 22720 4120 22772
rect 4436 22720 4488 22772
rect 6828 22763 6880 22772
rect 6828 22729 6837 22763
rect 6837 22729 6871 22763
rect 6871 22729 6880 22763
rect 6828 22720 6880 22729
rect 8024 22720 8076 22772
rect 8484 22720 8536 22772
rect 4068 22584 4120 22636
rect 4252 22627 4304 22636
rect 4252 22593 4261 22627
rect 4261 22593 4295 22627
rect 4295 22593 4304 22627
rect 4252 22584 4304 22593
rect 6920 22516 6972 22568
rect 7288 22559 7340 22568
rect 7288 22525 7297 22559
rect 7297 22525 7331 22559
rect 7331 22525 7340 22559
rect 7288 22516 7340 22525
rect 4436 22448 4488 22500
rect 6644 22491 6696 22500
rect 6644 22457 6653 22491
rect 6653 22457 6687 22491
rect 6687 22457 6696 22491
rect 6644 22448 6696 22457
rect 5540 22380 5592 22432
rect 5724 22380 5776 22432
rect 6920 22380 6972 22432
rect 7564 22516 7616 22568
rect 8208 22423 8260 22432
rect 8208 22389 8217 22423
rect 8217 22389 8251 22423
rect 8251 22389 8260 22423
rect 8208 22380 8260 22389
rect 10232 22380 10284 22432
rect 6315 22278 6367 22330
rect 6379 22278 6431 22330
rect 6443 22278 6495 22330
rect 6507 22278 6559 22330
rect 11648 22278 11700 22330
rect 11712 22278 11764 22330
rect 11776 22278 11828 22330
rect 11840 22278 11892 22330
rect 4436 22176 4488 22228
rect 6000 22176 6052 22228
rect 7564 22219 7616 22228
rect 7564 22185 7573 22219
rect 7573 22185 7607 22219
rect 7607 22185 7616 22219
rect 7564 22176 7616 22185
rect 7840 22176 7892 22228
rect 4068 22108 4120 22160
rect 6276 22108 6328 22160
rect 7104 22108 7156 22160
rect 4160 22040 4212 22092
rect 5908 22040 5960 22092
rect 10324 22040 10376 22092
rect 4068 22015 4120 22024
rect 4068 21981 4077 22015
rect 4077 21981 4111 22015
rect 4111 21981 4120 22015
rect 4068 21972 4120 21981
rect 6920 22015 6972 22024
rect 6920 21981 6929 22015
rect 6929 21981 6963 22015
rect 6963 21981 6972 22015
rect 6920 21972 6972 21981
rect 10232 22015 10284 22024
rect 10232 21981 10241 22015
rect 10241 21981 10275 22015
rect 10275 21981 10284 22015
rect 10232 21972 10284 21981
rect 7564 21904 7616 21956
rect 5724 21879 5776 21888
rect 5724 21845 5733 21879
rect 5733 21845 5767 21879
rect 5767 21845 5776 21879
rect 5724 21836 5776 21845
rect 8484 21836 8536 21888
rect 9956 21836 10008 21888
rect 3648 21734 3700 21786
rect 3712 21734 3764 21786
rect 3776 21734 3828 21786
rect 3840 21734 3892 21786
rect 8982 21734 9034 21786
rect 9046 21734 9098 21786
rect 9110 21734 9162 21786
rect 9174 21734 9226 21786
rect 14315 21734 14367 21786
rect 14379 21734 14431 21786
rect 14443 21734 14495 21786
rect 14507 21734 14559 21786
rect 4068 21632 4120 21684
rect 4804 21675 4856 21684
rect 4804 21641 4813 21675
rect 4813 21641 4847 21675
rect 4847 21641 4856 21675
rect 4804 21632 4856 21641
rect 4988 21632 5040 21684
rect 5172 21632 5224 21684
rect 5540 21632 5592 21684
rect 6276 21675 6328 21684
rect 6276 21641 6285 21675
rect 6285 21641 6319 21675
rect 6319 21641 6328 21675
rect 6276 21632 6328 21641
rect 7472 21632 7524 21684
rect 10324 21675 10376 21684
rect 10324 21641 10333 21675
rect 10333 21641 10367 21675
rect 10367 21641 10376 21675
rect 10324 21632 10376 21641
rect 1584 21539 1636 21548
rect 1584 21505 1593 21539
rect 1593 21505 1627 21539
rect 1627 21505 1636 21539
rect 1584 21496 1636 21505
rect 5172 21496 5224 21548
rect 5356 21539 5408 21548
rect 5356 21505 5365 21539
rect 5365 21505 5399 21539
rect 5399 21505 5408 21539
rect 5356 21496 5408 21505
rect 5724 21496 5776 21548
rect 4344 21428 4396 21480
rect 6736 21428 6788 21480
rect 8484 21471 8536 21480
rect 8484 21437 8493 21471
rect 8493 21437 8527 21471
rect 8527 21437 8536 21471
rect 8484 21428 8536 21437
rect 4988 21360 5040 21412
rect 5724 21360 5776 21412
rect 7104 21403 7156 21412
rect 7104 21369 7113 21403
rect 7113 21369 7147 21403
rect 7147 21369 7156 21403
rect 7104 21360 7156 21369
rect 7564 21360 7616 21412
rect 8852 21360 8904 21412
rect 2412 21292 2464 21344
rect 4160 21335 4212 21344
rect 4160 21301 4169 21335
rect 4169 21301 4203 21335
rect 4203 21301 4212 21335
rect 4160 21292 4212 21301
rect 7472 21335 7524 21344
rect 7472 21301 7481 21335
rect 7481 21301 7515 21335
rect 7515 21301 7524 21335
rect 7472 21292 7524 21301
rect 9404 21292 9456 21344
rect 10232 21292 10284 21344
rect 11980 21292 12032 21344
rect 6315 21190 6367 21242
rect 6379 21190 6431 21242
rect 6443 21190 6495 21242
rect 6507 21190 6559 21242
rect 11648 21190 11700 21242
rect 11712 21190 11764 21242
rect 11776 21190 11828 21242
rect 11840 21190 11892 21242
rect 2596 21088 2648 21140
rect 4068 21088 4120 21140
rect 5172 21131 5224 21140
rect 5172 21097 5181 21131
rect 5181 21097 5215 21131
rect 5215 21097 5224 21131
rect 5172 21088 5224 21097
rect 6736 21088 6788 21140
rect 8852 21088 8904 21140
rect 11244 21088 11296 21140
rect 1676 21063 1728 21072
rect 1676 21029 1685 21063
rect 1685 21029 1719 21063
rect 1719 21029 1728 21063
rect 1676 21020 1728 21029
rect 5356 21020 5408 21072
rect 5448 21020 5500 21072
rect 8760 21020 8812 21072
rect 9956 21063 10008 21072
rect 9956 21029 9990 21063
rect 9990 21029 10008 21063
rect 9956 21020 10008 21029
rect 12072 21020 12124 21072
rect 3976 20952 4028 21004
rect 7104 20952 7156 21004
rect 7472 20952 7524 21004
rect 8208 20952 8260 21004
rect 8484 20952 8536 21004
rect 10232 20952 10284 21004
rect 11980 20952 12032 21004
rect 1676 20884 1728 20936
rect 6920 20884 6972 20936
rect 7656 20884 7708 20936
rect 8024 20927 8076 20936
rect 8024 20893 8033 20927
rect 8033 20893 8067 20927
rect 8067 20893 8076 20927
rect 8024 20884 8076 20893
rect 7380 20791 7432 20800
rect 7380 20757 7389 20791
rect 7389 20757 7423 20791
rect 7423 20757 7432 20791
rect 7380 20748 7432 20757
rect 9588 20748 9640 20800
rect 12532 20748 12584 20800
rect 3648 20646 3700 20698
rect 3712 20646 3764 20698
rect 3776 20646 3828 20698
rect 3840 20646 3892 20698
rect 8982 20646 9034 20698
rect 9046 20646 9098 20698
rect 9110 20646 9162 20698
rect 9174 20646 9226 20698
rect 14315 20646 14367 20698
rect 14379 20646 14431 20698
rect 14443 20646 14495 20698
rect 14507 20646 14559 20698
rect 5908 20587 5960 20596
rect 5908 20553 5917 20587
rect 5917 20553 5951 20587
rect 5951 20553 5960 20587
rect 5908 20544 5960 20553
rect 6828 20544 6880 20596
rect 8300 20544 8352 20596
rect 2596 20451 2648 20460
rect 2596 20417 2605 20451
rect 2605 20417 2639 20451
rect 2639 20417 2648 20451
rect 2596 20408 2648 20417
rect 8024 20476 8076 20528
rect 9404 20544 9456 20596
rect 9772 20544 9824 20596
rect 10232 20544 10284 20596
rect 12440 20519 12492 20528
rect 12440 20485 12449 20519
rect 12449 20485 12483 20519
rect 12483 20485 12492 20519
rect 12440 20476 12492 20485
rect 5540 20340 5592 20392
rect 5908 20340 5960 20392
rect 6092 20340 6144 20392
rect 6828 20340 6880 20392
rect 9956 20408 10008 20460
rect 10876 20408 10928 20460
rect 12256 20451 12308 20460
rect 12256 20417 12265 20451
rect 12265 20417 12299 20451
rect 12299 20417 12308 20451
rect 12900 20451 12952 20460
rect 12256 20408 12308 20417
rect 12900 20417 12909 20451
rect 12909 20417 12943 20451
rect 12943 20417 12952 20451
rect 12900 20408 12952 20417
rect 9864 20340 9916 20392
rect 10232 20383 10284 20392
rect 10232 20349 10241 20383
rect 10241 20349 10275 20383
rect 10275 20349 10284 20383
rect 10232 20340 10284 20349
rect 3516 20272 3568 20324
rect 1676 20247 1728 20256
rect 1676 20213 1685 20247
rect 1685 20213 1719 20247
rect 1719 20213 1728 20247
rect 1676 20204 1728 20213
rect 2964 20204 3016 20256
rect 4160 20204 4212 20256
rect 9772 20272 9824 20324
rect 7288 20204 7340 20256
rect 8300 20247 8352 20256
rect 8300 20213 8309 20247
rect 8309 20213 8343 20247
rect 8343 20213 8352 20247
rect 8300 20204 8352 20213
rect 9680 20204 9732 20256
rect 10324 20247 10376 20256
rect 10324 20213 10333 20247
rect 10333 20213 10367 20247
rect 10367 20213 10376 20247
rect 10324 20204 10376 20213
rect 11336 20204 11388 20256
rect 12072 20340 12124 20392
rect 13176 20340 13228 20392
rect 6315 20102 6367 20154
rect 6379 20102 6431 20154
rect 6443 20102 6495 20154
rect 6507 20102 6559 20154
rect 11648 20102 11700 20154
rect 11712 20102 11764 20154
rect 11776 20102 11828 20154
rect 11840 20102 11892 20154
rect 2412 20043 2464 20052
rect 2412 20009 2421 20043
rect 2421 20009 2455 20043
rect 2455 20009 2464 20043
rect 2412 20000 2464 20009
rect 6092 20043 6144 20052
rect 6092 20009 6101 20043
rect 6101 20009 6135 20043
rect 6135 20009 6144 20043
rect 6092 20000 6144 20009
rect 2872 19975 2924 19984
rect 2872 19941 2881 19975
rect 2881 19941 2915 19975
rect 2915 19941 2924 19975
rect 2872 19932 2924 19941
rect 2780 19907 2832 19916
rect 2780 19873 2789 19907
rect 2789 19873 2823 19907
rect 2823 19873 2832 19907
rect 2780 19864 2832 19873
rect 4804 19864 4856 19916
rect 5264 19864 5316 19916
rect 5540 19864 5592 19916
rect 6460 19907 6512 19916
rect 6460 19873 6469 19907
rect 6469 19873 6503 19907
rect 6503 19873 6512 19907
rect 6460 19864 6512 19873
rect 2964 19839 3016 19848
rect 2964 19805 2973 19839
rect 2973 19805 3007 19839
rect 3007 19805 3016 19839
rect 2964 19796 3016 19805
rect 5172 19839 5224 19848
rect 5172 19805 5181 19839
rect 5181 19805 5215 19839
rect 5215 19805 5224 19839
rect 5172 19796 5224 19805
rect 7380 20000 7432 20052
rect 7840 20000 7892 20052
rect 8852 20000 8904 20052
rect 10324 20000 10376 20052
rect 12440 20000 12492 20052
rect 10876 19932 10928 19984
rect 11888 19932 11940 19984
rect 12164 19932 12216 19984
rect 7288 19907 7340 19916
rect 7288 19873 7297 19907
rect 7297 19873 7331 19907
rect 7331 19873 7340 19907
rect 7288 19864 7340 19873
rect 6092 19728 6144 19780
rect 7472 19796 7524 19848
rect 8208 19839 8260 19848
rect 8208 19805 8217 19839
rect 8217 19805 8251 19839
rect 8251 19805 8260 19839
rect 8208 19796 8260 19805
rect 8300 19839 8352 19848
rect 8300 19805 8309 19839
rect 8309 19805 8343 19839
rect 8343 19805 8352 19839
rect 8300 19796 8352 19805
rect 9956 19796 10008 19848
rect 10508 19796 10560 19848
rect 7012 19728 7064 19780
rect 10232 19728 10284 19780
rect 11796 19864 11848 19916
rect 11612 19839 11664 19848
rect 11612 19805 11621 19839
rect 11621 19805 11655 19839
rect 11655 19805 11664 19839
rect 11612 19796 11664 19805
rect 12348 19796 12400 19848
rect 12624 19864 12676 19916
rect 12992 19907 13044 19916
rect 12992 19873 13001 19907
rect 13001 19873 13035 19907
rect 13035 19873 13044 19907
rect 12992 19864 13044 19873
rect 12532 19796 12584 19848
rect 13084 19839 13136 19848
rect 13084 19805 13093 19839
rect 13093 19805 13127 19839
rect 13127 19805 13136 19839
rect 13084 19796 13136 19805
rect 13176 19839 13228 19848
rect 13176 19805 13185 19839
rect 13185 19805 13219 19839
rect 13219 19805 13228 19839
rect 13176 19796 13228 19805
rect 11520 19728 11572 19780
rect 4252 19660 4304 19712
rect 7472 19660 7524 19712
rect 8760 19703 8812 19712
rect 8760 19669 8769 19703
rect 8769 19669 8803 19703
rect 8803 19669 8812 19703
rect 8760 19660 8812 19669
rect 10508 19703 10560 19712
rect 10508 19669 10517 19703
rect 10517 19669 10551 19703
rect 10551 19669 10560 19703
rect 10508 19660 10560 19669
rect 10876 19703 10928 19712
rect 10876 19669 10885 19703
rect 10885 19669 10919 19703
rect 10919 19669 10928 19703
rect 10876 19660 10928 19669
rect 12164 19660 12216 19712
rect 3648 19558 3700 19610
rect 3712 19558 3764 19610
rect 3776 19558 3828 19610
rect 3840 19558 3892 19610
rect 8982 19558 9034 19610
rect 9046 19558 9098 19610
rect 9110 19558 9162 19610
rect 9174 19558 9226 19610
rect 14315 19558 14367 19610
rect 14379 19558 14431 19610
rect 14443 19558 14495 19610
rect 14507 19558 14559 19610
rect 10324 19456 10376 19508
rect 11520 19499 11572 19508
rect 11520 19465 11529 19499
rect 11529 19465 11563 19499
rect 11563 19465 11572 19499
rect 11520 19456 11572 19465
rect 2780 19388 2832 19440
rect 8208 19388 8260 19440
rect 10416 19388 10468 19440
rect 1400 19295 1452 19304
rect 1400 19261 1409 19295
rect 1409 19261 1443 19295
rect 1443 19261 1452 19295
rect 1400 19252 1452 19261
rect 1676 19295 1728 19304
rect 1676 19261 1685 19295
rect 1685 19261 1719 19295
rect 1719 19261 1728 19295
rect 1676 19252 1728 19261
rect 2964 19320 3016 19372
rect 4252 19363 4304 19372
rect 4252 19329 4261 19363
rect 4261 19329 4295 19363
rect 4295 19329 4304 19363
rect 4252 19320 4304 19329
rect 8024 19363 8076 19372
rect 3516 19252 3568 19304
rect 8024 19329 8033 19363
rect 8033 19329 8067 19363
rect 8067 19329 8076 19363
rect 8024 19320 8076 19329
rect 8852 19320 8904 19372
rect 11612 19388 11664 19440
rect 12532 19320 12584 19372
rect 12992 19363 13044 19372
rect 7196 19295 7248 19304
rect 7196 19261 7205 19295
rect 7205 19261 7239 19295
rect 7239 19261 7248 19295
rect 7196 19252 7248 19261
rect 7932 19252 7984 19304
rect 8760 19252 8812 19304
rect 10416 19295 10468 19304
rect 10416 19261 10425 19295
rect 10425 19261 10459 19295
rect 10459 19261 10468 19295
rect 10416 19252 10468 19261
rect 10876 19252 10928 19304
rect 12992 19329 13001 19363
rect 13001 19329 13035 19363
rect 13035 19329 13044 19363
rect 12992 19320 13044 19329
rect 5264 19227 5316 19236
rect 5264 19193 5273 19227
rect 5273 19193 5307 19227
rect 5307 19193 5316 19227
rect 5264 19184 5316 19193
rect 8852 19227 8904 19236
rect 8852 19193 8861 19227
rect 8861 19193 8895 19227
rect 8895 19193 8904 19227
rect 8852 19184 8904 19193
rect 2872 19159 2924 19168
rect 2872 19125 2881 19159
rect 2881 19125 2915 19159
rect 2915 19125 2924 19159
rect 2872 19116 2924 19125
rect 3976 19116 4028 19168
rect 4160 19159 4212 19168
rect 4160 19125 4169 19159
rect 4169 19125 4203 19159
rect 4203 19125 4212 19159
rect 4160 19116 4212 19125
rect 4804 19159 4856 19168
rect 4804 19125 4813 19159
rect 4813 19125 4847 19159
rect 4847 19125 4856 19159
rect 4804 19116 4856 19125
rect 5356 19159 5408 19168
rect 5356 19125 5365 19159
rect 5365 19125 5399 19159
rect 5399 19125 5408 19159
rect 5356 19116 5408 19125
rect 6092 19159 6144 19168
rect 6092 19125 6101 19159
rect 6101 19125 6135 19159
rect 6135 19125 6144 19159
rect 6092 19116 6144 19125
rect 6828 19116 6880 19168
rect 8116 19116 8168 19168
rect 8484 19159 8536 19168
rect 8484 19125 8493 19159
rect 8493 19125 8527 19159
rect 8527 19125 8536 19159
rect 8484 19116 8536 19125
rect 10508 19159 10560 19168
rect 10508 19125 10517 19159
rect 10517 19125 10551 19159
rect 10551 19125 10560 19159
rect 10508 19116 10560 19125
rect 11336 19116 11388 19168
rect 11520 19116 11572 19168
rect 11980 19116 12032 19168
rect 12440 19159 12492 19168
rect 12440 19125 12449 19159
rect 12449 19125 12483 19159
rect 12483 19125 12492 19159
rect 12440 19116 12492 19125
rect 12624 19116 12676 19168
rect 6315 19014 6367 19066
rect 6379 19014 6431 19066
rect 6443 19014 6495 19066
rect 6507 19014 6559 19066
rect 11648 19014 11700 19066
rect 11712 19014 11764 19066
rect 11776 19014 11828 19066
rect 11840 19014 11892 19066
rect 1400 18912 1452 18964
rect 2780 18912 2832 18964
rect 2872 18912 2924 18964
rect 5356 18912 5408 18964
rect 6000 18955 6052 18964
rect 6000 18921 6009 18955
rect 6009 18921 6043 18955
rect 6043 18921 6052 18955
rect 6000 18912 6052 18921
rect 8024 18912 8076 18964
rect 8208 18912 8260 18964
rect 9680 18955 9732 18964
rect 9680 18921 9689 18955
rect 9689 18921 9723 18955
rect 9723 18921 9732 18955
rect 9680 18912 9732 18921
rect 10140 18955 10192 18964
rect 10140 18921 10149 18955
rect 10149 18921 10183 18955
rect 10183 18921 10192 18955
rect 10140 18912 10192 18921
rect 12992 18955 13044 18964
rect 12992 18921 13001 18955
rect 13001 18921 13035 18955
rect 13035 18921 13044 18955
rect 12992 18912 13044 18921
rect 3516 18844 3568 18896
rect 4620 18844 4672 18896
rect 5540 18887 5592 18896
rect 5540 18853 5549 18887
rect 5549 18853 5583 18887
rect 5583 18853 5592 18887
rect 5540 18844 5592 18853
rect 5632 18844 5684 18896
rect 10232 18844 10284 18896
rect 10692 18844 10744 18896
rect 4344 18708 4396 18760
rect 7380 18776 7432 18828
rect 9864 18776 9916 18828
rect 10048 18819 10100 18828
rect 10048 18785 10057 18819
rect 10057 18785 10091 18819
rect 10091 18785 10100 18819
rect 10048 18776 10100 18785
rect 10600 18776 10652 18828
rect 10876 18776 10928 18828
rect 11336 18776 11388 18828
rect 12072 18844 12124 18896
rect 13084 18844 13136 18896
rect 4712 18708 4764 18760
rect 6828 18708 6880 18760
rect 9312 18708 9364 18760
rect 11704 18751 11756 18760
rect 11704 18717 11713 18751
rect 11713 18717 11747 18751
rect 11747 18717 11756 18751
rect 11704 18708 11756 18717
rect 4160 18640 4212 18692
rect 8392 18640 8444 18692
rect 10600 18640 10652 18692
rect 11244 18640 11296 18692
rect 12072 18708 12124 18760
rect 12992 18708 13044 18760
rect 3240 18615 3292 18624
rect 3240 18581 3249 18615
rect 3249 18581 3283 18615
rect 3283 18581 3292 18615
rect 3240 18572 3292 18581
rect 6736 18615 6788 18624
rect 6736 18581 6745 18615
rect 6745 18581 6779 18615
rect 6779 18581 6788 18615
rect 6736 18572 6788 18581
rect 10692 18615 10744 18624
rect 10692 18581 10701 18615
rect 10701 18581 10735 18615
rect 10735 18581 10744 18615
rect 10692 18572 10744 18581
rect 3648 18470 3700 18522
rect 3712 18470 3764 18522
rect 3776 18470 3828 18522
rect 3840 18470 3892 18522
rect 8982 18470 9034 18522
rect 9046 18470 9098 18522
rect 9110 18470 9162 18522
rect 9174 18470 9226 18522
rect 14315 18470 14367 18522
rect 14379 18470 14431 18522
rect 14443 18470 14495 18522
rect 14507 18470 14559 18522
rect 4712 18368 4764 18420
rect 5632 18411 5684 18420
rect 5632 18377 5641 18411
rect 5641 18377 5675 18411
rect 5675 18377 5684 18411
rect 5632 18368 5684 18377
rect 6000 18411 6052 18420
rect 6000 18377 6009 18411
rect 6009 18377 6043 18411
rect 6043 18377 6052 18411
rect 6000 18368 6052 18377
rect 6736 18368 6788 18420
rect 8300 18368 8352 18420
rect 10140 18368 10192 18420
rect 11704 18368 11756 18420
rect 12072 18411 12124 18420
rect 12072 18377 12081 18411
rect 12081 18377 12115 18411
rect 12115 18377 12124 18411
rect 12072 18368 12124 18377
rect 8024 18300 8076 18352
rect 8576 18300 8628 18352
rect 9312 18343 9364 18352
rect 9312 18309 9321 18343
rect 9321 18309 9355 18343
rect 9355 18309 9364 18343
rect 9312 18300 9364 18309
rect 3240 18164 3292 18216
rect 6736 18164 6788 18216
rect 10600 18232 10652 18284
rect 9772 18164 9824 18216
rect 10324 18164 10376 18216
rect 4068 18096 4120 18148
rect 10232 18096 10284 18148
rect 10692 18139 10744 18148
rect 10692 18105 10701 18139
rect 10701 18105 10735 18139
rect 10735 18105 10744 18139
rect 10692 18096 10744 18105
rect 3792 18028 3844 18080
rect 3976 18028 4028 18080
rect 5172 18028 5224 18080
rect 5540 18028 5592 18080
rect 6092 18028 6144 18080
rect 9864 18028 9916 18080
rect 10324 18071 10376 18080
rect 10324 18037 10333 18071
rect 10333 18037 10367 18071
rect 10367 18037 10376 18071
rect 10324 18028 10376 18037
rect 11336 18028 11388 18080
rect 6315 17926 6367 17978
rect 6379 17926 6431 17978
rect 6443 17926 6495 17978
rect 6507 17926 6559 17978
rect 11648 17926 11700 17978
rect 11712 17926 11764 17978
rect 11776 17926 11828 17978
rect 11840 17926 11892 17978
rect 4344 17867 4396 17876
rect 4344 17833 4353 17867
rect 4353 17833 4387 17867
rect 4387 17833 4396 17867
rect 4344 17824 4396 17833
rect 4620 17867 4672 17876
rect 4620 17833 4629 17867
rect 4629 17833 4663 17867
rect 4663 17833 4672 17867
rect 4620 17824 4672 17833
rect 5540 17824 5592 17876
rect 6828 17824 6880 17876
rect 7840 17867 7892 17876
rect 7840 17833 7849 17867
rect 7849 17833 7883 17867
rect 7883 17833 7892 17867
rect 7840 17824 7892 17833
rect 8484 17867 8536 17876
rect 8484 17833 8493 17867
rect 8493 17833 8527 17867
rect 8527 17833 8536 17867
rect 8484 17824 8536 17833
rect 10324 17824 10376 17876
rect 10784 17824 10836 17876
rect 3792 17799 3844 17808
rect 3792 17765 3801 17799
rect 3801 17765 3835 17799
rect 3835 17765 3844 17799
rect 3792 17756 3844 17765
rect 8392 17799 8444 17808
rect 8392 17765 8401 17799
rect 8401 17765 8435 17799
rect 8435 17765 8444 17799
rect 8392 17756 8444 17765
rect 2780 17731 2832 17740
rect 2780 17697 2789 17731
rect 2789 17697 2823 17731
rect 2823 17697 2832 17731
rect 2780 17688 2832 17697
rect 2872 17663 2924 17672
rect 2872 17629 2881 17663
rect 2881 17629 2915 17663
rect 2915 17629 2924 17663
rect 2872 17620 2924 17629
rect 5080 17688 5132 17740
rect 10876 17688 10928 17740
rect 4068 17620 4120 17672
rect 4988 17663 5040 17672
rect 4988 17629 4997 17663
rect 4997 17629 5031 17663
rect 5031 17629 5040 17663
rect 4988 17620 5040 17629
rect 8576 17663 8628 17672
rect 8576 17629 8585 17663
rect 8585 17629 8619 17663
rect 8619 17629 8628 17663
rect 8576 17620 8628 17629
rect 10324 17620 10376 17672
rect 11520 17620 11572 17672
rect 7472 17552 7524 17604
rect 10416 17595 10468 17604
rect 10416 17561 10425 17595
rect 10425 17561 10459 17595
rect 10459 17561 10468 17595
rect 10416 17552 10468 17561
rect 4988 17484 5040 17536
rect 6736 17484 6788 17536
rect 7380 17484 7432 17536
rect 10600 17484 10652 17536
rect 3648 17382 3700 17434
rect 3712 17382 3764 17434
rect 3776 17382 3828 17434
rect 3840 17382 3892 17434
rect 8982 17382 9034 17434
rect 9046 17382 9098 17434
rect 9110 17382 9162 17434
rect 9174 17382 9226 17434
rect 14315 17382 14367 17434
rect 14379 17382 14431 17434
rect 14443 17382 14495 17434
rect 14507 17382 14559 17434
rect 2780 17280 2832 17332
rect 4620 17280 4672 17332
rect 7288 17280 7340 17332
rect 8484 17323 8536 17332
rect 5632 17212 5684 17264
rect 5816 17212 5868 17264
rect 3976 17144 4028 17196
rect 2872 17076 2924 17128
rect 4160 17076 4212 17128
rect 8484 17289 8493 17323
rect 8493 17289 8527 17323
rect 8527 17289 8536 17323
rect 8484 17280 8536 17289
rect 10876 17280 10928 17332
rect 12348 17280 12400 17332
rect 8392 17212 8444 17264
rect 8576 17144 8628 17196
rect 10600 17187 10652 17196
rect 10600 17153 10609 17187
rect 10609 17153 10643 17187
rect 10643 17153 10652 17187
rect 10600 17144 10652 17153
rect 4252 17008 4304 17060
rect 4988 17008 5040 17060
rect 3976 16940 4028 16992
rect 5080 16983 5132 16992
rect 5080 16949 5089 16983
rect 5089 16949 5123 16983
rect 5123 16949 5132 16983
rect 5080 16940 5132 16949
rect 5724 16940 5776 16992
rect 7564 16983 7616 16992
rect 7564 16949 7573 16983
rect 7573 16949 7607 16983
rect 7607 16949 7616 16983
rect 7564 16940 7616 16949
rect 9680 16940 9732 16992
rect 9956 16983 10008 16992
rect 9956 16949 9965 16983
rect 9965 16949 9999 16983
rect 9999 16949 10008 16983
rect 9956 16940 10008 16949
rect 10048 16940 10100 16992
rect 6315 16838 6367 16890
rect 6379 16838 6431 16890
rect 6443 16838 6495 16890
rect 6507 16838 6559 16890
rect 11648 16838 11700 16890
rect 11712 16838 11764 16890
rect 11776 16838 11828 16890
rect 11840 16838 11892 16890
rect 3976 16736 4028 16788
rect 5080 16779 5132 16788
rect 5080 16745 5089 16779
rect 5089 16745 5123 16779
rect 5123 16745 5132 16779
rect 5080 16736 5132 16745
rect 10048 16779 10100 16788
rect 10048 16745 10057 16779
rect 10057 16745 10091 16779
rect 10091 16745 10100 16779
rect 10048 16736 10100 16745
rect 10784 16779 10836 16788
rect 10784 16745 10793 16779
rect 10793 16745 10827 16779
rect 10827 16745 10836 16779
rect 10784 16736 10836 16745
rect 6092 16668 6144 16720
rect 10324 16668 10376 16720
rect 12440 16736 12492 16788
rect 12624 16736 12676 16788
rect 5448 16643 5500 16652
rect 5448 16609 5457 16643
rect 5457 16609 5491 16643
rect 5491 16609 5500 16643
rect 5448 16600 5500 16609
rect 5724 16600 5776 16652
rect 5908 16643 5960 16652
rect 5908 16609 5942 16643
rect 5942 16609 5960 16643
rect 5908 16600 5960 16609
rect 7656 16600 7708 16652
rect 8208 16643 8260 16652
rect 8208 16609 8217 16643
rect 8217 16609 8251 16643
rect 8251 16609 8260 16643
rect 8208 16600 8260 16609
rect 10600 16600 10652 16652
rect 8300 16575 8352 16584
rect 8300 16541 8309 16575
rect 8309 16541 8343 16575
rect 8343 16541 8352 16575
rect 8300 16532 8352 16541
rect 8392 16575 8444 16584
rect 8392 16541 8401 16575
rect 8401 16541 8435 16575
rect 8435 16541 8444 16575
rect 8392 16532 8444 16541
rect 7012 16464 7064 16516
rect 9312 16464 9364 16516
rect 7840 16439 7892 16448
rect 7840 16405 7849 16439
rect 7849 16405 7883 16439
rect 7883 16405 7892 16439
rect 7840 16396 7892 16405
rect 10324 16396 10376 16448
rect 11336 16396 11388 16448
rect 3648 16294 3700 16346
rect 3712 16294 3764 16346
rect 3776 16294 3828 16346
rect 3840 16294 3892 16346
rect 8982 16294 9034 16346
rect 9046 16294 9098 16346
rect 9110 16294 9162 16346
rect 9174 16294 9226 16346
rect 14315 16294 14367 16346
rect 14379 16294 14431 16346
rect 14443 16294 14495 16346
rect 14507 16294 14559 16346
rect 4160 16192 4212 16244
rect 5908 16192 5960 16244
rect 11336 16235 11388 16244
rect 11336 16201 11345 16235
rect 11345 16201 11379 16235
rect 11379 16201 11388 16235
rect 11336 16192 11388 16201
rect 1584 16099 1636 16108
rect 1584 16065 1593 16099
rect 1593 16065 1627 16099
rect 1627 16065 1636 16099
rect 1584 16056 1636 16065
rect 5080 16056 5132 16108
rect 7012 16099 7064 16108
rect 7012 16065 7021 16099
rect 7021 16065 7055 16099
rect 7055 16065 7064 16099
rect 7012 16056 7064 16065
rect 9220 16099 9272 16108
rect 9220 16065 9229 16099
rect 9229 16065 9263 16099
rect 9263 16065 9272 16099
rect 9220 16056 9272 16065
rect 9312 15988 9364 16040
rect 7656 15920 7708 15972
rect 2228 15895 2280 15904
rect 2228 15861 2237 15895
rect 2237 15861 2271 15895
rect 2271 15861 2280 15895
rect 2228 15852 2280 15861
rect 5080 15852 5132 15904
rect 7104 15852 7156 15904
rect 8852 15852 8904 15904
rect 10600 15895 10652 15904
rect 10600 15861 10609 15895
rect 10609 15861 10643 15895
rect 10643 15861 10652 15895
rect 10600 15852 10652 15861
rect 6315 15750 6367 15802
rect 6379 15750 6431 15802
rect 6443 15750 6495 15802
rect 6507 15750 6559 15802
rect 11648 15750 11700 15802
rect 11712 15750 11764 15802
rect 11776 15750 11828 15802
rect 11840 15750 11892 15802
rect 5540 15648 5592 15700
rect 8208 15648 8260 15700
rect 9220 15691 9272 15700
rect 9220 15657 9229 15691
rect 9229 15657 9263 15691
rect 9263 15657 9272 15691
rect 9220 15648 9272 15657
rect 9956 15648 10008 15700
rect 11060 15648 11112 15700
rect 6920 15555 6972 15564
rect 6920 15521 6929 15555
rect 6929 15521 6963 15555
rect 6963 15521 6972 15555
rect 6920 15512 6972 15521
rect 7012 15487 7064 15496
rect 7012 15453 7021 15487
rect 7021 15453 7055 15487
rect 7055 15453 7064 15487
rect 7012 15444 7064 15453
rect 7104 15487 7156 15496
rect 7104 15453 7113 15487
rect 7113 15453 7147 15487
rect 7147 15453 7156 15487
rect 7104 15444 7156 15453
rect 9956 15444 10008 15496
rect 5448 15419 5500 15428
rect 5448 15385 5457 15419
rect 5457 15385 5491 15419
rect 5491 15385 5500 15419
rect 5448 15376 5500 15385
rect 5816 15376 5868 15428
rect 6828 15376 6880 15428
rect 10324 15376 10376 15428
rect 5080 15351 5132 15360
rect 5080 15317 5089 15351
rect 5089 15317 5123 15351
rect 5123 15317 5132 15351
rect 5080 15308 5132 15317
rect 5540 15308 5592 15360
rect 5724 15351 5776 15360
rect 5724 15317 5733 15351
rect 5733 15317 5767 15351
rect 5767 15317 5776 15351
rect 5724 15308 5776 15317
rect 8208 15308 8260 15360
rect 8392 15308 8444 15360
rect 10508 15308 10560 15360
rect 3648 15206 3700 15258
rect 3712 15206 3764 15258
rect 3776 15206 3828 15258
rect 3840 15206 3892 15258
rect 8982 15206 9034 15258
rect 9046 15206 9098 15258
rect 9110 15206 9162 15258
rect 9174 15206 9226 15258
rect 14315 15206 14367 15258
rect 14379 15206 14431 15258
rect 14443 15206 14495 15258
rect 14507 15206 14559 15258
rect 6828 15104 6880 15156
rect 7840 15104 7892 15156
rect 9956 15147 10008 15156
rect 9956 15113 9965 15147
rect 9965 15113 9999 15147
rect 9999 15113 10008 15147
rect 9956 15104 10008 15113
rect 11060 15147 11112 15156
rect 11060 15113 11069 15147
rect 11069 15113 11103 15147
rect 11103 15113 11112 15147
rect 11060 15104 11112 15113
rect 6920 15036 6972 15088
rect 9404 15036 9456 15088
rect 7196 14968 7248 15020
rect 7656 15011 7708 15020
rect 7656 14977 7665 15011
rect 7665 14977 7699 15011
rect 7699 14977 7708 15011
rect 7656 14968 7708 14977
rect 10600 14968 10652 15020
rect 3148 14943 3200 14952
rect 3148 14909 3157 14943
rect 3157 14909 3191 14943
rect 3191 14909 3200 14943
rect 3148 14900 3200 14909
rect 5540 14900 5592 14952
rect 7840 14900 7892 14952
rect 10140 14900 10192 14952
rect 3976 14832 4028 14884
rect 7656 14832 7708 14884
rect 4620 14764 4672 14816
rect 6315 14662 6367 14714
rect 6379 14662 6431 14714
rect 6443 14662 6495 14714
rect 6507 14662 6559 14714
rect 11648 14662 11700 14714
rect 11712 14662 11764 14714
rect 11776 14662 11828 14714
rect 11840 14662 11892 14714
rect 3148 14603 3200 14612
rect 3148 14569 3157 14603
rect 3157 14569 3191 14603
rect 3191 14569 3200 14603
rect 3148 14560 3200 14569
rect 4528 14560 4580 14612
rect 5356 14560 5408 14612
rect 7196 14603 7248 14612
rect 7196 14569 7205 14603
rect 7205 14569 7239 14603
rect 7239 14569 7248 14603
rect 7196 14560 7248 14569
rect 7656 14603 7708 14612
rect 7656 14569 7665 14603
rect 7665 14569 7699 14603
rect 7699 14569 7708 14603
rect 7656 14560 7708 14569
rect 7932 14560 7984 14612
rect 9680 14560 9732 14612
rect 9956 14560 10008 14612
rect 10140 14560 10192 14612
rect 10508 14560 10560 14612
rect 10324 14535 10376 14544
rect 10324 14501 10333 14535
rect 10333 14501 10367 14535
rect 10367 14501 10376 14535
rect 10324 14492 10376 14501
rect 4896 14467 4948 14476
rect 4896 14433 4905 14467
rect 4905 14433 4939 14467
rect 4939 14433 4948 14467
rect 4896 14424 4948 14433
rect 7564 14467 7616 14476
rect 7564 14433 7573 14467
rect 7573 14433 7607 14467
rect 7607 14433 7616 14467
rect 7564 14424 7616 14433
rect 8116 14467 8168 14476
rect 8116 14433 8125 14467
rect 8125 14433 8159 14467
rect 8159 14433 8168 14467
rect 8116 14424 8168 14433
rect 4068 14288 4120 14340
rect 5540 14399 5592 14408
rect 5540 14365 5549 14399
rect 5549 14365 5583 14399
rect 5583 14365 5592 14399
rect 5540 14356 5592 14365
rect 8208 14399 8260 14408
rect 8208 14365 8217 14399
rect 8217 14365 8251 14399
rect 8251 14365 8260 14399
rect 8208 14356 8260 14365
rect 3332 14220 3384 14272
rect 4712 14220 4764 14272
rect 5816 14220 5868 14272
rect 6828 14220 6880 14272
rect 8300 14220 8352 14272
rect 3648 14118 3700 14170
rect 3712 14118 3764 14170
rect 3776 14118 3828 14170
rect 3840 14118 3892 14170
rect 8982 14118 9034 14170
rect 9046 14118 9098 14170
rect 9110 14118 9162 14170
rect 9174 14118 9226 14170
rect 14315 14118 14367 14170
rect 14379 14118 14431 14170
rect 14443 14118 14495 14170
rect 14507 14118 14559 14170
rect 3424 14016 3476 14068
rect 4528 14059 4580 14068
rect 4528 14025 4537 14059
rect 4537 14025 4571 14059
rect 4571 14025 4580 14059
rect 4528 14016 4580 14025
rect 7564 14016 7616 14068
rect 7932 14016 7984 14068
rect 8760 14016 8812 14068
rect 4160 13948 4212 14000
rect 8116 13991 8168 14000
rect 8116 13957 8125 13991
rect 8125 13957 8159 13991
rect 8159 13957 8168 13991
rect 8116 13948 8168 13957
rect 5540 13923 5592 13932
rect 5540 13889 5549 13923
rect 5549 13889 5583 13923
rect 5583 13889 5592 13923
rect 5540 13880 5592 13889
rect 9680 13880 9732 13932
rect 2780 13855 2832 13864
rect 2780 13821 2789 13855
rect 2789 13821 2823 13855
rect 2823 13821 2832 13855
rect 2780 13812 2832 13821
rect 3332 13812 3384 13864
rect 5264 13812 5316 13864
rect 5448 13855 5500 13864
rect 5448 13821 5457 13855
rect 5457 13821 5491 13855
rect 5491 13821 5500 13855
rect 5448 13812 5500 13821
rect 8208 13812 8260 13864
rect 5172 13744 5224 13796
rect 5540 13744 5592 13796
rect 11060 13812 11112 13864
rect 11244 13744 11296 13796
rect 3976 13676 4028 13728
rect 4804 13676 4856 13728
rect 5448 13676 5500 13728
rect 10140 13676 10192 13728
rect 6315 13574 6367 13626
rect 6379 13574 6431 13626
rect 6443 13574 6495 13626
rect 6507 13574 6559 13626
rect 11648 13574 11700 13626
rect 11712 13574 11764 13626
rect 11776 13574 11828 13626
rect 11840 13574 11892 13626
rect 4068 13472 4120 13524
rect 1676 13447 1728 13456
rect 1676 13413 1685 13447
rect 1685 13413 1719 13447
rect 1719 13413 1728 13447
rect 1676 13404 1728 13413
rect 4896 13472 4948 13524
rect 8300 13472 8352 13524
rect 1400 13379 1452 13388
rect 1400 13345 1409 13379
rect 1409 13345 1443 13379
rect 1443 13345 1452 13379
rect 1400 13336 1452 13345
rect 4620 13336 4672 13388
rect 2228 13175 2280 13184
rect 2228 13141 2237 13175
rect 2237 13141 2271 13175
rect 2271 13141 2280 13175
rect 2228 13132 2280 13141
rect 2780 13132 2832 13184
rect 3148 13132 3200 13184
rect 6736 13404 6788 13456
rect 7840 13336 7892 13388
rect 8852 13472 8904 13524
rect 9312 13472 9364 13524
rect 9680 13515 9732 13524
rect 9680 13481 9689 13515
rect 9689 13481 9723 13515
rect 9723 13481 9732 13515
rect 9680 13472 9732 13481
rect 11244 13515 11296 13524
rect 11244 13481 11253 13515
rect 11253 13481 11287 13515
rect 11287 13481 11296 13515
rect 11244 13472 11296 13481
rect 8576 13336 8628 13388
rect 10048 13379 10100 13388
rect 10048 13345 10057 13379
rect 10057 13345 10091 13379
rect 10091 13345 10100 13379
rect 10048 13336 10100 13345
rect 11612 13379 11664 13388
rect 11612 13345 11621 13379
rect 11621 13345 11655 13379
rect 11655 13345 11664 13379
rect 11612 13336 11664 13345
rect 11704 13379 11756 13388
rect 11704 13345 11713 13379
rect 11713 13345 11747 13379
rect 11747 13345 11756 13379
rect 11704 13336 11756 13345
rect 12256 13336 12308 13388
rect 10140 13311 10192 13320
rect 5172 13132 5224 13184
rect 5908 13175 5960 13184
rect 5908 13141 5917 13175
rect 5917 13141 5951 13175
rect 5951 13141 5960 13175
rect 5908 13132 5960 13141
rect 6092 13132 6144 13184
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 10324 13311 10376 13320
rect 10324 13277 10333 13311
rect 10333 13277 10367 13311
rect 10367 13277 10376 13311
rect 10324 13268 10376 13277
rect 11796 13311 11848 13320
rect 11796 13277 11805 13311
rect 11805 13277 11839 13311
rect 11839 13277 11848 13311
rect 11796 13268 11848 13277
rect 7656 13132 7708 13184
rect 8392 13200 8444 13252
rect 8116 13175 8168 13184
rect 8116 13141 8125 13175
rect 8125 13141 8159 13175
rect 8159 13141 8168 13175
rect 8116 13132 8168 13141
rect 3648 13030 3700 13082
rect 3712 13030 3764 13082
rect 3776 13030 3828 13082
rect 3840 13030 3892 13082
rect 8982 13030 9034 13082
rect 9046 13030 9098 13082
rect 9110 13030 9162 13082
rect 9174 13030 9226 13082
rect 14315 13030 14367 13082
rect 14379 13030 14431 13082
rect 14443 13030 14495 13082
rect 14507 13030 14559 13082
rect 3148 12971 3200 12980
rect 3148 12937 3157 12971
rect 3157 12937 3191 12971
rect 3191 12937 3200 12971
rect 3148 12928 3200 12937
rect 3240 12928 3292 12980
rect 3976 12928 4028 12980
rect 5264 12928 5316 12980
rect 7840 12971 7892 12980
rect 2688 12835 2740 12844
rect 2688 12801 2697 12835
rect 2697 12801 2731 12835
rect 2731 12801 2740 12835
rect 2688 12792 2740 12801
rect 2228 12724 2280 12776
rect 4620 12903 4672 12912
rect 4620 12869 4629 12903
rect 4629 12869 4663 12903
rect 4663 12869 4672 12903
rect 4620 12860 4672 12869
rect 5908 12792 5960 12844
rect 7840 12937 7849 12971
rect 7849 12937 7883 12971
rect 7883 12937 7892 12971
rect 7840 12928 7892 12937
rect 8116 12928 8168 12980
rect 8392 12971 8444 12980
rect 8392 12937 8401 12971
rect 8401 12937 8435 12971
rect 8435 12937 8444 12971
rect 8392 12928 8444 12937
rect 10140 12928 10192 12980
rect 10600 12971 10652 12980
rect 10600 12937 10609 12971
rect 10609 12937 10643 12971
rect 10643 12937 10652 12971
rect 10600 12928 10652 12937
rect 11336 12928 11388 12980
rect 11796 12928 11848 12980
rect 7104 12860 7156 12912
rect 7656 12792 7708 12844
rect 11704 12903 11756 12912
rect 11704 12869 11713 12903
rect 11713 12869 11747 12903
rect 11747 12869 11756 12903
rect 11704 12860 11756 12869
rect 8484 12792 8536 12844
rect 8852 12792 8904 12844
rect 11612 12792 11664 12844
rect 4068 12724 4120 12776
rect 4804 12724 4856 12776
rect 5540 12767 5592 12776
rect 5540 12733 5549 12767
rect 5549 12733 5583 12767
rect 5583 12733 5592 12767
rect 5540 12724 5592 12733
rect 6736 12724 6788 12776
rect 6828 12724 6880 12776
rect 8576 12767 8628 12776
rect 8576 12733 8585 12767
rect 8585 12733 8619 12767
rect 8619 12733 8628 12767
rect 8576 12724 8628 12733
rect 9036 12724 9088 12776
rect 9588 12724 9640 12776
rect 7104 12656 7156 12708
rect 8668 12656 8720 12708
rect 8852 12656 8904 12708
rect 2044 12631 2096 12640
rect 2044 12597 2053 12631
rect 2053 12597 2087 12631
rect 2087 12597 2096 12631
rect 2044 12588 2096 12597
rect 2504 12631 2556 12640
rect 2504 12597 2513 12631
rect 2513 12597 2547 12631
rect 2547 12597 2556 12631
rect 4068 12631 4120 12640
rect 2504 12588 2556 12597
rect 4068 12597 4077 12631
rect 4077 12597 4111 12631
rect 4111 12597 4120 12631
rect 4068 12588 4120 12597
rect 5540 12588 5592 12640
rect 5724 12588 5776 12640
rect 9680 12588 9732 12640
rect 10324 12631 10376 12640
rect 10324 12597 10333 12631
rect 10333 12597 10367 12631
rect 10367 12597 10376 12631
rect 10324 12588 10376 12597
rect 6315 12486 6367 12538
rect 6379 12486 6431 12538
rect 6443 12486 6495 12538
rect 6507 12486 6559 12538
rect 11648 12486 11700 12538
rect 11712 12486 11764 12538
rect 11776 12486 11828 12538
rect 11840 12486 11892 12538
rect 1400 12384 1452 12436
rect 4068 12384 4120 12436
rect 4252 12384 4304 12436
rect 4528 12384 4580 12436
rect 4804 12384 4856 12436
rect 5540 12384 5592 12436
rect 6828 12384 6880 12436
rect 9036 12427 9088 12436
rect 9036 12393 9045 12427
rect 9045 12393 9079 12427
rect 9079 12393 9088 12427
rect 9036 12384 9088 12393
rect 10048 12384 10100 12436
rect 2964 12316 3016 12368
rect 3148 12316 3200 12368
rect 5908 12316 5960 12368
rect 6276 12316 6328 12368
rect 7012 12316 7064 12368
rect 8208 12316 8260 12368
rect 8576 12316 8628 12368
rect 10416 12316 10468 12368
rect 10968 12316 11020 12368
rect 4620 12248 4672 12300
rect 5816 12291 5868 12300
rect 5816 12257 5825 12291
rect 5825 12257 5859 12291
rect 5859 12257 5868 12291
rect 5816 12248 5868 12257
rect 10876 12248 10928 12300
rect 11336 12248 11388 12300
rect 4712 12223 4764 12232
rect 4712 12189 4721 12223
rect 4721 12189 4755 12223
rect 4755 12189 4764 12223
rect 4712 12180 4764 12189
rect 4896 12180 4948 12232
rect 5632 12180 5684 12232
rect 6000 12180 6052 12232
rect 6828 12223 6880 12232
rect 6828 12189 6837 12223
rect 6837 12189 6871 12223
rect 6871 12189 6880 12223
rect 6828 12180 6880 12189
rect 8576 12180 8628 12232
rect 9680 12180 9732 12232
rect 10324 12112 10376 12164
rect 2504 12044 2556 12096
rect 2964 12044 3016 12096
rect 3516 12044 3568 12096
rect 5172 12044 5224 12096
rect 5540 12044 5592 12096
rect 7196 12044 7248 12096
rect 9680 12044 9732 12096
rect 10508 12044 10560 12096
rect 10968 12044 11020 12096
rect 3648 11942 3700 11994
rect 3712 11942 3764 11994
rect 3776 11942 3828 11994
rect 3840 11942 3892 11994
rect 8982 11942 9034 11994
rect 9046 11942 9098 11994
rect 9110 11942 9162 11994
rect 9174 11942 9226 11994
rect 14315 11942 14367 11994
rect 14379 11942 14431 11994
rect 14443 11942 14495 11994
rect 14507 11942 14559 11994
rect 2964 11840 3016 11892
rect 4344 11840 4396 11892
rect 4620 11883 4672 11892
rect 4620 11849 4629 11883
rect 4629 11849 4663 11883
rect 4663 11849 4672 11883
rect 4620 11840 4672 11849
rect 5816 11840 5868 11892
rect 6920 11883 6972 11892
rect 6920 11849 6929 11883
rect 6929 11849 6963 11883
rect 6963 11849 6972 11883
rect 6920 11840 6972 11849
rect 3240 11772 3292 11824
rect 10508 11772 10560 11824
rect 10876 11772 10928 11824
rect 5632 11704 5684 11756
rect 6184 11704 6236 11756
rect 7288 11704 7340 11756
rect 3516 11679 3568 11688
rect 3516 11645 3525 11679
rect 3525 11645 3559 11679
rect 3559 11645 3568 11679
rect 3516 11636 3568 11645
rect 7380 11679 7432 11688
rect 7380 11645 7389 11679
rect 7389 11645 7423 11679
rect 7423 11645 7432 11679
rect 7380 11636 7432 11645
rect 7564 11636 7616 11688
rect 8300 11636 8352 11688
rect 8576 11679 8628 11688
rect 8576 11645 8585 11679
rect 8585 11645 8619 11679
rect 8619 11645 8628 11679
rect 8576 11636 8628 11645
rect 10048 11704 10100 11756
rect 11336 11704 11388 11756
rect 10324 11636 10376 11688
rect 7288 11611 7340 11620
rect 7288 11577 7297 11611
rect 7297 11577 7331 11611
rect 7331 11577 7340 11611
rect 7288 11568 7340 11577
rect 11152 11611 11204 11620
rect 11152 11577 11161 11611
rect 11161 11577 11195 11611
rect 11195 11577 11204 11611
rect 11152 11568 11204 11577
rect 11520 11568 11572 11620
rect 3608 11543 3660 11552
rect 3608 11509 3617 11543
rect 3617 11509 3651 11543
rect 3651 11509 3660 11543
rect 3608 11500 3660 11509
rect 4620 11500 4672 11552
rect 4896 11543 4948 11552
rect 4896 11509 4905 11543
rect 4905 11509 4939 11543
rect 4939 11509 4948 11543
rect 4896 11500 4948 11509
rect 7012 11500 7064 11552
rect 7840 11500 7892 11552
rect 10140 11500 10192 11552
rect 10324 11543 10376 11552
rect 10324 11509 10333 11543
rect 10333 11509 10367 11543
rect 10367 11509 10376 11543
rect 10324 11500 10376 11509
rect 11980 11500 12032 11552
rect 6315 11398 6367 11450
rect 6379 11398 6431 11450
rect 6443 11398 6495 11450
rect 6507 11398 6559 11450
rect 11648 11398 11700 11450
rect 11712 11398 11764 11450
rect 11776 11398 11828 11450
rect 11840 11398 11892 11450
rect 2780 11296 2832 11348
rect 3608 11296 3660 11348
rect 6828 11296 6880 11348
rect 7288 11339 7340 11348
rect 7288 11305 7297 11339
rect 7297 11305 7331 11339
rect 7331 11305 7340 11339
rect 7288 11296 7340 11305
rect 7472 11296 7524 11348
rect 8484 11296 8536 11348
rect 9404 11296 9456 11348
rect 9588 11296 9640 11348
rect 9772 11296 9824 11348
rect 10048 11296 10100 11348
rect 11060 11296 11112 11348
rect 7196 11228 7248 11280
rect 8392 11271 8444 11280
rect 8392 11237 8401 11271
rect 8401 11237 8435 11271
rect 8435 11237 8444 11271
rect 8392 11228 8444 11237
rect 10140 11228 10192 11280
rect 11152 11228 11204 11280
rect 7564 11160 7616 11212
rect 7748 11160 7800 11212
rect 7840 11160 7892 11212
rect 8300 11160 8352 11212
rect 9404 11160 9456 11212
rect 7932 11135 7984 11144
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 9312 11092 9364 11144
rect 9772 11092 9824 11144
rect 12348 11160 12400 11212
rect 12440 11160 12492 11212
rect 11336 11092 11388 11144
rect 11980 11092 12032 11144
rect 4068 11024 4120 11076
rect 9588 10956 9640 11008
rect 3648 10854 3700 10906
rect 3712 10854 3764 10906
rect 3776 10854 3828 10906
rect 3840 10854 3892 10906
rect 8982 10854 9034 10906
rect 9046 10854 9098 10906
rect 9110 10854 9162 10906
rect 9174 10854 9226 10906
rect 14315 10854 14367 10906
rect 14379 10854 14431 10906
rect 14443 10854 14495 10906
rect 14507 10854 14559 10906
rect 5816 10752 5868 10804
rect 7472 10752 7524 10804
rect 7932 10752 7984 10804
rect 10600 10752 10652 10804
rect 12348 10684 12400 10736
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 4160 10616 4212 10668
rect 7840 10616 7892 10668
rect 1492 10548 1544 10600
rect 4252 10591 4304 10600
rect 4252 10557 4261 10591
rect 4261 10557 4295 10591
rect 4295 10557 4304 10591
rect 4252 10548 4304 10557
rect 3884 10480 3936 10532
rect 4528 10480 4580 10532
rect 2412 10412 2464 10464
rect 6920 10412 6972 10464
rect 7564 10412 7616 10464
rect 10968 10616 11020 10668
rect 9680 10548 9732 10600
rect 8392 10480 8444 10532
rect 10968 10480 11020 10532
rect 8116 10412 8168 10464
rect 9680 10455 9732 10464
rect 9680 10421 9689 10455
rect 9689 10421 9723 10455
rect 9723 10421 9732 10455
rect 9680 10412 9732 10421
rect 10508 10455 10560 10464
rect 10508 10421 10517 10455
rect 10517 10421 10551 10455
rect 10551 10421 10560 10455
rect 10508 10412 10560 10421
rect 10600 10455 10652 10464
rect 10600 10421 10609 10455
rect 10609 10421 10643 10455
rect 10643 10421 10652 10455
rect 10600 10412 10652 10421
rect 11336 10412 11388 10464
rect 11980 10455 12032 10464
rect 11980 10421 11989 10455
rect 11989 10421 12023 10455
rect 12023 10421 12032 10455
rect 11980 10412 12032 10421
rect 6315 10310 6367 10362
rect 6379 10310 6431 10362
rect 6443 10310 6495 10362
rect 6507 10310 6559 10362
rect 11648 10310 11700 10362
rect 11712 10310 11764 10362
rect 11776 10310 11828 10362
rect 11840 10310 11892 10362
rect 2412 10251 2464 10260
rect 2412 10217 2421 10251
rect 2421 10217 2455 10251
rect 2455 10217 2464 10251
rect 2412 10208 2464 10217
rect 2504 10208 2556 10260
rect 3884 10251 3936 10260
rect 3884 10217 3893 10251
rect 3893 10217 3927 10251
rect 3927 10217 3936 10251
rect 3884 10208 3936 10217
rect 5816 10251 5868 10260
rect 5816 10217 5825 10251
rect 5825 10217 5859 10251
rect 5859 10217 5868 10251
rect 5816 10208 5868 10217
rect 7380 10208 7432 10260
rect 9588 10208 9640 10260
rect 10600 10208 10652 10260
rect 5908 10140 5960 10192
rect 5264 10047 5316 10056
rect 5264 10013 5273 10047
rect 5273 10013 5307 10047
rect 5307 10013 5316 10047
rect 5264 10004 5316 10013
rect 7196 10140 7248 10192
rect 7656 10140 7708 10192
rect 8392 10140 8444 10192
rect 9956 10140 10008 10192
rect 10508 10140 10560 10192
rect 7104 10072 7156 10124
rect 7748 10072 7800 10124
rect 10140 10115 10192 10124
rect 10140 10081 10149 10115
rect 10149 10081 10183 10115
rect 10183 10081 10192 10115
rect 10140 10072 10192 10081
rect 7932 10004 7984 10056
rect 8300 10004 8352 10056
rect 9956 10004 10008 10056
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 10692 10004 10744 10056
rect 4620 9936 4672 9988
rect 9312 9936 9364 9988
rect 10968 9936 11020 9988
rect 11428 9936 11480 9988
rect 5540 9868 5592 9920
rect 8484 9868 8536 9920
rect 9404 9911 9456 9920
rect 9404 9877 9413 9911
rect 9413 9877 9447 9911
rect 9447 9877 9456 9911
rect 9404 9868 9456 9877
rect 11244 9911 11296 9920
rect 11244 9877 11253 9911
rect 11253 9877 11287 9911
rect 11287 9877 11296 9911
rect 11244 9868 11296 9877
rect 3648 9766 3700 9818
rect 3712 9766 3764 9818
rect 3776 9766 3828 9818
rect 3840 9766 3892 9818
rect 8982 9766 9034 9818
rect 9046 9766 9098 9818
rect 9110 9766 9162 9818
rect 9174 9766 9226 9818
rect 14315 9766 14367 9818
rect 14379 9766 14431 9818
rect 14443 9766 14495 9818
rect 14507 9766 14559 9818
rect 5816 9664 5868 9716
rect 7748 9664 7800 9716
rect 9404 9664 9456 9716
rect 11152 9664 11204 9716
rect 2688 9596 2740 9648
rect 6000 9596 6052 9648
rect 7104 9596 7156 9648
rect 7196 9596 7248 9648
rect 2412 9528 2464 9580
rect 2596 9460 2648 9512
rect 3424 9528 3476 9580
rect 12164 9596 12216 9648
rect 12992 9596 13044 9648
rect 7932 9528 7984 9580
rect 8116 9528 8168 9580
rect 8392 9528 8444 9580
rect 9680 9528 9732 9580
rect 10140 9571 10192 9580
rect 10140 9537 10149 9571
rect 10149 9537 10183 9571
rect 10183 9537 10192 9571
rect 10140 9528 10192 9537
rect 10508 9571 10560 9580
rect 10508 9537 10517 9571
rect 10517 9537 10551 9571
rect 10551 9537 10560 9571
rect 10508 9528 10560 9537
rect 11244 9571 11296 9580
rect 11244 9537 11253 9571
rect 11253 9537 11287 9571
rect 11287 9537 11296 9571
rect 11244 9528 11296 9537
rect 2688 9367 2740 9376
rect 2688 9333 2697 9367
rect 2697 9333 2731 9367
rect 2731 9333 2740 9367
rect 2688 9324 2740 9333
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 6644 9460 6696 9512
rect 6920 9460 6972 9512
rect 4068 9392 4120 9444
rect 4896 9324 4948 9376
rect 5908 9324 5960 9376
rect 6000 9324 6052 9376
rect 8668 9392 8720 9444
rect 11428 9392 11480 9444
rect 6644 9324 6696 9376
rect 10692 9367 10744 9376
rect 10692 9333 10701 9367
rect 10701 9333 10735 9367
rect 10735 9333 10744 9367
rect 10692 9324 10744 9333
rect 6315 9222 6367 9274
rect 6379 9222 6431 9274
rect 6443 9222 6495 9274
rect 6507 9222 6559 9274
rect 11648 9222 11700 9274
rect 11712 9222 11764 9274
rect 11776 9222 11828 9274
rect 11840 9222 11892 9274
rect 2596 9120 2648 9172
rect 6920 9163 6972 9172
rect 6920 9129 6929 9163
rect 6929 9129 6963 9163
rect 6963 9129 6972 9163
rect 6920 9120 6972 9129
rect 7748 9163 7800 9172
rect 7748 9129 7757 9163
rect 7757 9129 7791 9163
rect 7791 9129 7800 9163
rect 7748 9120 7800 9129
rect 8300 9163 8352 9172
rect 8300 9129 8309 9163
rect 8309 9129 8343 9163
rect 8343 9129 8352 9163
rect 8300 9120 8352 9129
rect 10692 9120 10744 9172
rect 5264 9052 5316 9104
rect 5448 9052 5500 9104
rect 9956 9095 10008 9104
rect 9956 9061 9965 9095
rect 9965 9061 9999 9095
rect 9999 9061 10008 9095
rect 9956 9052 10008 9061
rect 10968 9052 11020 9104
rect 11152 9052 11204 9104
rect 7104 8984 7156 9036
rect 11980 9120 12032 9172
rect 2872 8780 2924 8832
rect 3424 8780 3476 8832
rect 7932 8959 7984 8968
rect 7932 8925 7941 8959
rect 7941 8925 7975 8959
rect 7975 8925 7984 8959
rect 7932 8916 7984 8925
rect 6460 8823 6512 8832
rect 6460 8789 6469 8823
rect 6469 8789 6503 8823
rect 6503 8789 6512 8823
rect 6460 8780 6512 8789
rect 6920 8780 6972 8832
rect 8392 8780 8444 8832
rect 10876 8780 10928 8832
rect 11152 8780 11204 8832
rect 3648 8678 3700 8730
rect 3712 8678 3764 8730
rect 3776 8678 3828 8730
rect 3840 8678 3892 8730
rect 8982 8678 9034 8730
rect 9046 8678 9098 8730
rect 9110 8678 9162 8730
rect 9174 8678 9226 8730
rect 14315 8678 14367 8730
rect 14379 8678 14431 8730
rect 14443 8678 14495 8730
rect 14507 8678 14559 8730
rect 4068 8576 4120 8628
rect 5264 8576 5316 8628
rect 7104 8576 7156 8628
rect 7932 8576 7984 8628
rect 10968 8576 11020 8628
rect 6184 8508 6236 8560
rect 8208 8551 8260 8560
rect 8208 8517 8217 8551
rect 8217 8517 8251 8551
rect 8251 8517 8260 8551
rect 8208 8508 8260 8517
rect 1584 8483 1636 8492
rect 1584 8449 1593 8483
rect 1593 8449 1627 8483
rect 1627 8449 1636 8483
rect 1584 8440 1636 8449
rect 5724 8440 5776 8492
rect 6460 8440 6512 8492
rect 2872 8372 2924 8424
rect 5540 8415 5592 8424
rect 5540 8381 5549 8415
rect 5549 8381 5583 8415
rect 5583 8381 5592 8415
rect 5540 8372 5592 8381
rect 9036 8415 9088 8424
rect 2688 8347 2740 8356
rect 2688 8313 2697 8347
rect 2697 8313 2731 8347
rect 2731 8313 2740 8347
rect 2688 8304 2740 8313
rect 9036 8381 9045 8415
rect 9045 8381 9079 8415
rect 9079 8381 9088 8415
rect 9036 8372 9088 8381
rect 10968 8440 11020 8492
rect 8392 8304 8444 8356
rect 2780 8236 2832 8288
rect 5172 8279 5224 8288
rect 5172 8245 5181 8279
rect 5181 8245 5215 8279
rect 5215 8245 5224 8279
rect 5172 8236 5224 8245
rect 11152 8279 11204 8288
rect 11152 8245 11161 8279
rect 11161 8245 11195 8279
rect 11195 8245 11204 8279
rect 11152 8236 11204 8245
rect 6315 8134 6367 8186
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 11648 8134 11700 8186
rect 11712 8134 11764 8186
rect 11776 8134 11828 8186
rect 11840 8134 11892 8186
rect 2872 8032 2924 8084
rect 5724 8032 5776 8084
rect 6828 8032 6880 8084
rect 7748 8075 7800 8084
rect 7748 8041 7757 8075
rect 7757 8041 7791 8075
rect 7791 8041 7800 8075
rect 7748 8032 7800 8041
rect 10876 8032 10928 8084
rect 11428 8032 11480 8084
rect 4528 7964 4580 8016
rect 6644 7964 6696 8016
rect 6736 7964 6788 8016
rect 7196 7939 7248 7948
rect 7196 7905 7205 7939
rect 7205 7905 7239 7939
rect 7239 7905 7248 7939
rect 7196 7896 7248 7905
rect 11428 7939 11480 7948
rect 11428 7905 11462 7939
rect 11462 7905 11480 7939
rect 11428 7896 11480 7905
rect 4620 7871 4672 7880
rect 4620 7837 4629 7871
rect 4629 7837 4663 7871
rect 4663 7837 4672 7871
rect 4620 7828 4672 7837
rect 6184 7871 6236 7880
rect 6184 7837 6193 7871
rect 6193 7837 6227 7871
rect 6227 7837 6236 7871
rect 6184 7828 6236 7837
rect 8392 7828 8444 7880
rect 9036 7871 9088 7880
rect 9036 7837 9045 7871
rect 9045 7837 9079 7871
rect 9079 7837 9088 7871
rect 9036 7828 9088 7837
rect 11152 7871 11204 7880
rect 11152 7837 11161 7871
rect 11161 7837 11195 7871
rect 11195 7837 11204 7871
rect 11152 7828 11204 7837
rect 1676 7735 1728 7744
rect 1676 7701 1685 7735
rect 1685 7701 1719 7735
rect 1719 7701 1728 7735
rect 1676 7692 1728 7701
rect 2872 7735 2924 7744
rect 2872 7701 2881 7735
rect 2881 7701 2915 7735
rect 2915 7701 2924 7735
rect 2872 7692 2924 7701
rect 5632 7735 5684 7744
rect 5632 7701 5641 7735
rect 5641 7701 5675 7735
rect 5675 7701 5684 7735
rect 5632 7692 5684 7701
rect 6920 7692 6972 7744
rect 8116 7735 8168 7744
rect 8116 7701 8125 7735
rect 8125 7701 8159 7735
rect 8159 7701 8168 7735
rect 8116 7692 8168 7701
rect 12440 7692 12492 7744
rect 3648 7590 3700 7642
rect 3712 7590 3764 7642
rect 3776 7590 3828 7642
rect 3840 7590 3892 7642
rect 8982 7590 9034 7642
rect 9046 7590 9098 7642
rect 9110 7590 9162 7642
rect 9174 7590 9226 7642
rect 14315 7590 14367 7642
rect 14379 7590 14431 7642
rect 14443 7590 14495 7642
rect 14507 7590 14559 7642
rect 2044 7488 2096 7540
rect 2872 7488 2924 7540
rect 3516 7488 3568 7540
rect 4528 7531 4580 7540
rect 4528 7497 4537 7531
rect 4537 7497 4571 7531
rect 4571 7497 4580 7531
rect 4528 7488 4580 7497
rect 5448 7488 5500 7540
rect 6184 7488 6236 7540
rect 7196 7531 7248 7540
rect 7196 7497 7205 7531
rect 7205 7497 7239 7531
rect 7239 7497 7248 7531
rect 7196 7488 7248 7497
rect 8668 7531 8720 7540
rect 8668 7497 8677 7531
rect 8677 7497 8711 7531
rect 8711 7497 8720 7531
rect 8668 7488 8720 7497
rect 11428 7488 11480 7540
rect 1584 7395 1636 7404
rect 1584 7361 1593 7395
rect 1593 7361 1627 7395
rect 1627 7361 1636 7395
rect 1584 7352 1636 7361
rect 4344 7420 4396 7472
rect 4988 7463 5040 7472
rect 4988 7429 4997 7463
rect 4997 7429 5031 7463
rect 5031 7429 5040 7463
rect 4988 7420 5040 7429
rect 1676 7284 1728 7336
rect 5172 7352 5224 7404
rect 5632 7284 5684 7336
rect 8116 7284 8168 7336
rect 7840 7216 7892 7268
rect 2872 7191 2924 7200
rect 2872 7157 2881 7191
rect 2881 7157 2915 7191
rect 2915 7157 2924 7191
rect 2872 7148 2924 7157
rect 8116 7148 8168 7200
rect 9680 7148 9732 7200
rect 12072 7148 12124 7200
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 11648 7046 11700 7098
rect 11712 7046 11764 7098
rect 11776 7046 11828 7098
rect 11840 7046 11892 7098
rect 5632 6944 5684 6996
rect 5724 6987 5776 6996
rect 5724 6953 5733 6987
rect 5733 6953 5767 6987
rect 5767 6953 5776 6987
rect 5724 6944 5776 6953
rect 11152 6944 11204 6996
rect 11428 6944 11480 6996
rect 2136 6808 2188 6860
rect 2504 6808 2556 6860
rect 5356 6808 5408 6860
rect 5632 6808 5684 6860
rect 6000 6808 6052 6860
rect 6276 6808 6328 6860
rect 7472 6808 7524 6860
rect 8668 6876 8720 6928
rect 7932 6808 7984 6860
rect 9772 6808 9824 6860
rect 10784 6808 10836 6860
rect 12072 6876 12124 6928
rect 11060 6808 11112 6860
rect 1584 6783 1636 6792
rect 1584 6749 1593 6783
rect 1593 6749 1627 6783
rect 1627 6749 1636 6783
rect 1584 6740 1636 6749
rect 7748 6783 7800 6792
rect 7748 6749 7757 6783
rect 7757 6749 7791 6783
rect 7791 6749 7800 6783
rect 7748 6740 7800 6749
rect 7840 6783 7892 6792
rect 7840 6749 7849 6783
rect 7849 6749 7883 6783
rect 7883 6749 7892 6783
rect 7840 6740 7892 6749
rect 7288 6715 7340 6724
rect 7288 6681 7297 6715
rect 7297 6681 7331 6715
rect 7331 6681 7340 6715
rect 7288 6672 7340 6681
rect 9680 6672 9732 6724
rect 2412 6647 2464 6656
rect 2412 6613 2421 6647
rect 2421 6613 2455 6647
rect 2455 6613 2464 6647
rect 2412 6604 2464 6613
rect 2872 6647 2924 6656
rect 2872 6613 2881 6647
rect 2881 6613 2915 6647
rect 2915 6613 2924 6647
rect 2872 6604 2924 6613
rect 3332 6647 3384 6656
rect 3332 6613 3341 6647
rect 3341 6613 3375 6647
rect 3375 6613 3384 6647
rect 3332 6604 3384 6613
rect 3516 6604 3568 6656
rect 4804 6604 4856 6656
rect 5356 6604 5408 6656
rect 5724 6604 5776 6656
rect 7748 6604 7800 6656
rect 8300 6647 8352 6656
rect 8300 6613 8309 6647
rect 8309 6613 8343 6647
rect 8343 6613 8352 6647
rect 8300 6604 8352 6613
rect 9864 6647 9916 6656
rect 9864 6613 9873 6647
rect 9873 6613 9907 6647
rect 9907 6613 9916 6647
rect 9864 6604 9916 6613
rect 3648 6502 3700 6554
rect 3712 6502 3764 6554
rect 3776 6502 3828 6554
rect 3840 6502 3892 6554
rect 8982 6502 9034 6554
rect 9046 6502 9098 6554
rect 9110 6502 9162 6554
rect 9174 6502 9226 6554
rect 14315 6502 14367 6554
rect 14379 6502 14431 6554
rect 14443 6502 14495 6554
rect 14507 6502 14559 6554
rect 2504 6400 2556 6452
rect 4160 6332 4212 6384
rect 3516 6196 3568 6248
rect 5448 6400 5500 6452
rect 5632 6400 5684 6452
rect 6828 6443 6880 6452
rect 6828 6409 6837 6443
rect 6837 6409 6871 6443
rect 6871 6409 6880 6443
rect 6828 6400 6880 6409
rect 7012 6332 7064 6384
rect 7288 6307 7340 6316
rect 7288 6273 7297 6307
rect 7297 6273 7331 6307
rect 7331 6273 7340 6307
rect 7288 6264 7340 6273
rect 7472 6307 7524 6316
rect 7472 6273 7481 6307
rect 7481 6273 7515 6307
rect 7515 6273 7524 6307
rect 7472 6264 7524 6273
rect 5908 6196 5960 6248
rect 6092 6196 6144 6248
rect 6184 6196 6236 6248
rect 9496 6400 9548 6452
rect 9772 6443 9824 6452
rect 9772 6409 9781 6443
rect 9781 6409 9815 6443
rect 9815 6409 9824 6443
rect 9772 6400 9824 6409
rect 11060 6400 11112 6452
rect 9680 6264 9732 6316
rect 2228 6128 2280 6180
rect 4436 6128 4488 6180
rect 5172 6128 5224 6180
rect 6276 6128 6328 6180
rect 9404 6171 9456 6180
rect 1676 6103 1728 6112
rect 1676 6069 1685 6103
rect 1685 6069 1719 6103
rect 1719 6069 1728 6103
rect 1676 6060 1728 6069
rect 2688 6060 2740 6112
rect 3056 6060 3108 6112
rect 4068 6103 4120 6112
rect 4068 6069 4077 6103
rect 4077 6069 4111 6103
rect 4111 6069 4120 6103
rect 4068 6060 4120 6069
rect 4344 6103 4396 6112
rect 4344 6069 4353 6103
rect 4353 6069 4387 6103
rect 4387 6069 4396 6103
rect 4344 6060 4396 6069
rect 5816 6103 5868 6112
rect 5816 6069 5825 6103
rect 5825 6069 5859 6103
rect 5859 6069 5868 6103
rect 5816 6060 5868 6069
rect 9404 6137 9413 6171
rect 9413 6137 9447 6171
rect 9447 6137 9456 6171
rect 9404 6128 9456 6137
rect 6828 6060 6880 6112
rect 7564 6060 7616 6112
rect 7840 6103 7892 6112
rect 7840 6069 7849 6103
rect 7849 6069 7883 6103
rect 7883 6069 7892 6103
rect 7840 6060 7892 6069
rect 8392 6060 8444 6112
rect 8484 6060 8536 6112
rect 11336 6103 11388 6112
rect 11336 6069 11345 6103
rect 11345 6069 11379 6103
rect 11379 6069 11388 6103
rect 11336 6060 11388 6069
rect 12072 6103 12124 6112
rect 12072 6069 12081 6103
rect 12081 6069 12115 6103
rect 12115 6069 12124 6103
rect 12072 6060 12124 6069
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 11648 5958 11700 6010
rect 11712 5958 11764 6010
rect 11776 5958 11828 6010
rect 11840 5958 11892 6010
rect 1492 5788 1544 5840
rect 3332 5856 3384 5908
rect 4252 5856 4304 5908
rect 4344 5856 4396 5908
rect 7932 5856 7984 5908
rect 8300 5899 8352 5908
rect 8300 5865 8309 5899
rect 8309 5865 8343 5899
rect 8343 5865 8352 5899
rect 8300 5856 8352 5865
rect 8576 5856 8628 5908
rect 9036 5856 9088 5908
rect 11060 5899 11112 5908
rect 11060 5865 11069 5899
rect 11069 5865 11103 5899
rect 11103 5865 11112 5899
rect 11060 5856 11112 5865
rect 11152 5856 11204 5908
rect 5264 5788 5316 5840
rect 6000 5788 6052 5840
rect 6828 5788 6880 5840
rect 8024 5788 8076 5840
rect 9772 5788 9824 5840
rect 11336 5788 11388 5840
rect 1952 5720 2004 5772
rect 2412 5720 2464 5772
rect 4344 5763 4396 5772
rect 4344 5729 4378 5763
rect 4378 5729 4396 5763
rect 4344 5720 4396 5729
rect 3056 5695 3108 5704
rect 3056 5661 3065 5695
rect 3065 5661 3099 5695
rect 3099 5661 3108 5695
rect 3056 5652 3108 5661
rect 6736 5695 6788 5704
rect 1860 5559 1912 5568
rect 1860 5525 1869 5559
rect 1869 5525 1903 5559
rect 1903 5525 1912 5559
rect 1860 5516 1912 5525
rect 2228 5559 2280 5568
rect 2228 5525 2237 5559
rect 2237 5525 2271 5559
rect 2271 5525 2280 5559
rect 2228 5516 2280 5525
rect 3516 5559 3568 5568
rect 3516 5525 3525 5559
rect 3525 5525 3559 5559
rect 3559 5525 3568 5559
rect 3516 5516 3568 5525
rect 6736 5661 6745 5695
rect 6745 5661 6779 5695
rect 6779 5661 6788 5695
rect 6736 5652 6788 5661
rect 12072 5720 12124 5772
rect 7564 5652 7616 5704
rect 7932 5652 7984 5704
rect 6276 5627 6328 5636
rect 6276 5593 6285 5627
rect 6285 5593 6319 5627
rect 6319 5593 6328 5627
rect 6276 5584 6328 5593
rect 4804 5516 4856 5568
rect 4988 5516 5040 5568
rect 7288 5559 7340 5568
rect 7288 5525 7297 5559
rect 7297 5525 7331 5559
rect 7331 5525 7340 5559
rect 7288 5516 7340 5525
rect 8208 5516 8260 5568
rect 9588 5516 9640 5568
rect 3648 5414 3700 5466
rect 3712 5414 3764 5466
rect 3776 5414 3828 5466
rect 3840 5414 3892 5466
rect 8982 5414 9034 5466
rect 9046 5414 9098 5466
rect 9110 5414 9162 5466
rect 9174 5414 9226 5466
rect 14315 5414 14367 5466
rect 14379 5414 14431 5466
rect 14443 5414 14495 5466
rect 14507 5414 14559 5466
rect 1952 5355 2004 5364
rect 1952 5321 1961 5355
rect 1961 5321 1995 5355
rect 1995 5321 2004 5355
rect 1952 5312 2004 5321
rect 3056 5355 3108 5364
rect 3056 5321 3065 5355
rect 3065 5321 3099 5355
rect 3099 5321 3108 5355
rect 3056 5312 3108 5321
rect 4620 5355 4672 5364
rect 4620 5321 4629 5355
rect 4629 5321 4663 5355
rect 4663 5321 4672 5355
rect 4620 5312 4672 5321
rect 5540 5312 5592 5364
rect 8024 5312 8076 5364
rect 8300 5312 8352 5364
rect 9772 5355 9824 5364
rect 9772 5321 9781 5355
rect 9781 5321 9815 5355
rect 9815 5321 9824 5355
rect 9772 5312 9824 5321
rect 9864 5312 9916 5364
rect 10140 5312 10192 5364
rect 10600 5312 10652 5364
rect 12072 5355 12124 5364
rect 12072 5321 12081 5355
rect 12081 5321 12115 5355
rect 12115 5321 12124 5355
rect 12072 5312 12124 5321
rect 2228 5244 2280 5296
rect 1860 5176 1912 5228
rect 2412 5219 2464 5228
rect 2412 5185 2421 5219
rect 2421 5185 2455 5219
rect 2455 5185 2464 5219
rect 2412 5176 2464 5185
rect 4896 5244 4948 5296
rect 5172 5244 5224 5296
rect 3516 5176 3568 5228
rect 4344 5176 4396 5228
rect 5632 5176 5684 5228
rect 7288 5176 7340 5228
rect 9312 5176 9364 5228
rect 11428 5176 11480 5228
rect 1676 5108 1728 5160
rect 4620 5108 4672 5160
rect 7196 5151 7248 5160
rect 7196 5117 7205 5151
rect 7205 5117 7239 5151
rect 7239 5117 7248 5151
rect 7196 5108 7248 5117
rect 8576 5108 8628 5160
rect 10600 5108 10652 5160
rect 10692 5040 10744 5092
rect 3884 5015 3936 5024
rect 3884 4981 3893 5015
rect 3893 4981 3927 5015
rect 3927 4981 3936 5015
rect 3884 4972 3936 4981
rect 5080 5015 5132 5024
rect 5080 4981 5089 5015
rect 5089 4981 5123 5015
rect 5123 4981 5132 5015
rect 5080 4972 5132 4981
rect 5448 4972 5500 5024
rect 6828 5015 6880 5024
rect 6828 4981 6837 5015
rect 6837 4981 6871 5015
rect 6871 4981 6880 5015
rect 6828 4972 6880 4981
rect 8300 5015 8352 5024
rect 8300 4981 8309 5015
rect 8309 4981 8343 5015
rect 8343 4981 8352 5015
rect 8300 4972 8352 4981
rect 10600 5015 10652 5024
rect 10600 4981 10609 5015
rect 10609 4981 10643 5015
rect 10643 4981 10652 5015
rect 10600 4972 10652 4981
rect 11520 4972 11572 5024
rect 12348 4972 12400 5024
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 11648 4870 11700 4922
rect 11712 4870 11764 4922
rect 11776 4870 11828 4922
rect 11840 4870 11892 4922
rect 4252 4768 4304 4820
rect 5080 4768 5132 4820
rect 7564 4811 7616 4820
rect 7564 4777 7573 4811
rect 7573 4777 7607 4811
rect 7607 4777 7616 4811
rect 7564 4768 7616 4777
rect 9312 4768 9364 4820
rect 9680 4768 9732 4820
rect 5540 4700 5592 4752
rect 6828 4700 6880 4752
rect 10600 4768 10652 4820
rect 11520 4768 11572 4820
rect 12164 4768 12216 4820
rect 12624 4768 12676 4820
rect 1492 4632 1544 4684
rect 2320 4632 2372 4684
rect 3056 4632 3108 4684
rect 4344 4632 4396 4684
rect 5448 4675 5500 4684
rect 5448 4641 5457 4675
rect 5457 4641 5491 4675
rect 5491 4641 5500 4675
rect 5448 4632 5500 4641
rect 5632 4632 5684 4684
rect 6184 4675 6236 4684
rect 6184 4641 6193 4675
rect 6193 4641 6227 4675
rect 6227 4641 6236 4675
rect 6184 4632 6236 4641
rect 6460 4675 6512 4684
rect 6460 4641 6494 4675
rect 6494 4641 6512 4675
rect 6460 4632 6512 4641
rect 8852 4632 8904 4684
rect 9772 4632 9824 4684
rect 1584 4607 1636 4616
rect 1584 4573 1593 4607
rect 1593 4573 1627 4607
rect 1627 4573 1636 4607
rect 1584 4564 1636 4573
rect 4896 4607 4948 4616
rect 4896 4573 4905 4607
rect 4905 4573 4939 4607
rect 4939 4573 4948 4607
rect 4896 4564 4948 4573
rect 10140 4607 10192 4616
rect 10140 4573 10149 4607
rect 10149 4573 10183 4607
rect 10183 4573 10192 4607
rect 10140 4564 10192 4573
rect 11428 4632 11480 4684
rect 12808 4675 12860 4684
rect 12808 4641 12817 4675
rect 12817 4641 12851 4675
rect 12851 4641 12860 4675
rect 12808 4632 12860 4641
rect 11796 4607 11848 4616
rect 11796 4573 11805 4607
rect 11805 4573 11839 4607
rect 11839 4573 11848 4607
rect 11796 4564 11848 4573
rect 12256 4564 12308 4616
rect 2136 4496 2188 4548
rect 9956 4496 10008 4548
rect 12440 4496 12492 4548
rect 2780 4428 2832 4480
rect 7932 4471 7984 4480
rect 7932 4437 7941 4471
rect 7941 4437 7975 4471
rect 7975 4437 7984 4471
rect 7932 4428 7984 4437
rect 8576 4471 8628 4480
rect 8576 4437 8585 4471
rect 8585 4437 8619 4471
rect 8619 4437 8628 4471
rect 8576 4428 8628 4437
rect 9588 4428 9640 4480
rect 10692 4471 10744 4480
rect 10692 4437 10701 4471
rect 10701 4437 10735 4471
rect 10735 4437 10744 4471
rect 10692 4428 10744 4437
rect 3648 4326 3700 4378
rect 3712 4326 3764 4378
rect 3776 4326 3828 4378
rect 3840 4326 3892 4378
rect 8982 4326 9034 4378
rect 9046 4326 9098 4378
rect 9110 4326 9162 4378
rect 9174 4326 9226 4378
rect 14315 4326 14367 4378
rect 14379 4326 14431 4378
rect 14443 4326 14495 4378
rect 14507 4326 14559 4378
rect 2228 4224 2280 4276
rect 3516 4224 3568 4276
rect 4896 4224 4948 4276
rect 7748 4224 7800 4276
rect 8852 4224 8904 4276
rect 9772 4267 9824 4276
rect 9772 4233 9781 4267
rect 9781 4233 9815 4267
rect 9815 4233 9824 4267
rect 9772 4224 9824 4233
rect 10140 4224 10192 4276
rect 12808 4224 12860 4276
rect 204 4088 256 4140
rect 3148 4156 3200 4208
rect 8300 4156 8352 4208
rect 4988 4088 5040 4140
rect 5172 4088 5224 4140
rect 6092 4088 6144 4140
rect 2780 3952 2832 4004
rect 2964 4020 3016 4072
rect 6276 4020 6328 4072
rect 7656 4088 7708 4140
rect 7932 4088 7984 4140
rect 8852 4088 8904 4140
rect 9404 4131 9456 4140
rect 9404 4097 9413 4131
rect 9413 4097 9447 4131
rect 9447 4097 9456 4131
rect 11796 4156 11848 4208
rect 9404 4088 9456 4097
rect 8392 4020 8444 4072
rect 10140 4020 10192 4072
rect 10508 4020 10560 4072
rect 11336 4020 11388 4072
rect 12256 4088 12308 4140
rect 12624 4088 12676 4140
rect 4988 3927 5040 3936
rect 4988 3893 4997 3927
rect 4997 3893 5031 3927
rect 5031 3893 5040 3927
rect 4988 3884 5040 3893
rect 5632 3927 5684 3936
rect 5632 3893 5641 3927
rect 5641 3893 5675 3927
rect 5675 3893 5684 3927
rect 5632 3884 5684 3893
rect 6092 3884 6144 3936
rect 6460 3952 6512 4004
rect 7932 3952 7984 4004
rect 9588 3952 9640 4004
rect 7012 3927 7064 3936
rect 7012 3893 7021 3927
rect 7021 3893 7055 3927
rect 7055 3893 7064 3927
rect 7012 3884 7064 3893
rect 8208 3884 8260 3936
rect 10600 3952 10652 4004
rect 11428 3952 11480 4004
rect 10508 3927 10560 3936
rect 10508 3893 10517 3927
rect 10517 3893 10551 3927
rect 10551 3893 10560 3927
rect 10508 3884 10560 3893
rect 12992 3884 13044 3936
rect 15752 3884 15804 3936
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 11648 3782 11700 3834
rect 11712 3782 11764 3834
rect 11776 3782 11828 3834
rect 11840 3782 11892 3834
rect 2412 3723 2464 3732
rect 2412 3689 2421 3723
rect 2421 3689 2455 3723
rect 2455 3689 2464 3723
rect 2412 3680 2464 3689
rect 2780 3723 2832 3732
rect 2780 3689 2789 3723
rect 2789 3689 2823 3723
rect 2823 3689 2832 3723
rect 2780 3680 2832 3689
rect 4988 3680 5040 3732
rect 5540 3723 5592 3732
rect 5540 3689 5549 3723
rect 5549 3689 5583 3723
rect 5583 3689 5592 3723
rect 5540 3680 5592 3689
rect 7104 3680 7156 3732
rect 8392 3680 8444 3732
rect 3056 3612 3108 3664
rect 3976 3612 4028 3664
rect 5172 3612 5224 3664
rect 5264 3612 5316 3664
rect 5908 3612 5960 3664
rect 7564 3612 7616 3664
rect 7932 3612 7984 3664
rect 4528 3587 4580 3596
rect 4528 3553 4537 3587
rect 4537 3553 4571 3587
rect 4571 3553 4580 3587
rect 4528 3544 4580 3553
rect 7656 3544 7708 3596
rect 2872 3519 2924 3528
rect 2872 3485 2881 3519
rect 2881 3485 2915 3519
rect 2915 3485 2924 3519
rect 2872 3476 2924 3485
rect 3056 3519 3108 3528
rect 3056 3485 3065 3519
rect 3065 3485 3099 3519
rect 3099 3485 3108 3519
rect 3056 3476 3108 3485
rect 3332 3408 3384 3460
rect 4344 3408 4396 3460
rect 4988 3476 5040 3528
rect 1952 3383 2004 3392
rect 1952 3349 1961 3383
rect 1961 3349 1995 3383
rect 1995 3349 2004 3383
rect 1952 3340 2004 3349
rect 3424 3340 3476 3392
rect 6092 3340 6144 3392
rect 9312 3680 9364 3732
rect 10692 3680 10744 3732
rect 10968 3680 11020 3732
rect 11520 3680 11572 3732
rect 12348 3680 12400 3732
rect 12716 3680 12768 3732
rect 10048 3612 10100 3664
rect 6736 3408 6788 3460
rect 8392 3408 8444 3460
rect 10232 3476 10284 3528
rect 11428 3544 11480 3596
rect 12808 3612 12860 3664
rect 13268 3587 13320 3596
rect 13268 3553 13277 3587
rect 13277 3553 13311 3587
rect 13311 3553 13320 3587
rect 13268 3544 13320 3553
rect 10968 3476 11020 3528
rect 12164 3519 12216 3528
rect 12164 3485 12173 3519
rect 12173 3485 12207 3519
rect 12207 3485 12216 3519
rect 12164 3476 12216 3485
rect 12256 3519 12308 3528
rect 12256 3485 12265 3519
rect 12265 3485 12299 3519
rect 12299 3485 12308 3519
rect 12716 3519 12768 3528
rect 12256 3476 12308 3485
rect 12716 3485 12725 3519
rect 12725 3485 12759 3519
rect 12759 3485 12768 3519
rect 12716 3476 12768 3485
rect 13452 3451 13504 3460
rect 13452 3417 13461 3451
rect 13461 3417 13495 3451
rect 13495 3417 13504 3451
rect 13452 3408 13504 3417
rect 13084 3383 13136 3392
rect 13084 3349 13093 3383
rect 13093 3349 13127 3383
rect 13127 3349 13136 3383
rect 13084 3340 13136 3349
rect 3648 3238 3700 3290
rect 3712 3238 3764 3290
rect 3776 3238 3828 3290
rect 3840 3238 3892 3290
rect 8982 3238 9034 3290
rect 9046 3238 9098 3290
rect 9110 3238 9162 3290
rect 9174 3238 9226 3290
rect 14315 3238 14367 3290
rect 14379 3238 14431 3290
rect 14443 3238 14495 3290
rect 14507 3238 14559 3290
rect 3332 3179 3384 3188
rect 3332 3145 3341 3179
rect 3341 3145 3375 3179
rect 3375 3145 3384 3179
rect 3332 3136 3384 3145
rect 3976 3136 4028 3188
rect 4528 3136 4580 3188
rect 5448 3136 5500 3188
rect 6552 3136 6604 3188
rect 7656 3179 7708 3188
rect 7656 3145 7665 3179
rect 7665 3145 7699 3179
rect 7699 3145 7708 3179
rect 7656 3136 7708 3145
rect 7932 3136 7984 3188
rect 6828 3068 6880 3120
rect 8852 3136 8904 3188
rect 10048 3136 10100 3188
rect 10140 3136 10192 3188
rect 4804 2932 4856 2984
rect 6552 2932 6604 2984
rect 8116 2932 8168 2984
rect 4344 2864 4396 2916
rect 8852 2932 8904 2984
rect 12164 3136 12216 3188
rect 12440 3179 12492 3188
rect 12440 3145 12449 3179
rect 12449 3145 12483 3179
rect 12483 3145 12492 3179
rect 12440 3136 12492 3145
rect 13268 3136 13320 3188
rect 10968 3043 11020 3052
rect 10968 3009 10977 3043
rect 10977 3009 11011 3043
rect 11011 3009 11020 3043
rect 10968 3000 11020 3009
rect 11428 3000 11480 3052
rect 12348 3000 12400 3052
rect 13084 3068 13136 3120
rect 8300 2864 8352 2916
rect 8392 2864 8444 2916
rect 8576 2864 8628 2916
rect 12716 2932 12768 2984
rect 10784 2907 10836 2916
rect 10784 2873 10793 2907
rect 10793 2873 10827 2907
rect 10827 2873 10836 2907
rect 10784 2864 10836 2873
rect 11060 2864 11112 2916
rect 11152 2864 11204 2916
rect 12164 2864 12216 2916
rect 12808 2907 12860 2916
rect 12808 2873 12817 2907
rect 12817 2873 12851 2907
rect 12851 2873 12860 2907
rect 12808 2864 12860 2873
rect 2688 2796 2740 2848
rect 7012 2839 7064 2848
rect 7012 2805 7021 2839
rect 7021 2805 7055 2839
rect 7055 2805 7064 2839
rect 7012 2796 7064 2805
rect 9496 2796 9548 2848
rect 9680 2796 9732 2848
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 11648 2694 11700 2746
rect 11712 2694 11764 2746
rect 11776 2694 11828 2746
rect 11840 2694 11892 2746
rect 2504 2592 2556 2644
rect 2872 2592 2924 2644
rect 2964 2524 3016 2576
rect 4344 2524 4396 2576
rect 4068 2456 4120 2508
rect 1952 2320 2004 2372
rect 3424 2388 3476 2440
rect 4528 2431 4580 2440
rect 4528 2397 4537 2431
rect 4537 2397 4571 2431
rect 4571 2397 4580 2431
rect 4528 2388 4580 2397
rect 8208 2592 8260 2644
rect 8668 2592 8720 2644
rect 10048 2635 10100 2644
rect 10048 2601 10057 2635
rect 10057 2601 10091 2635
rect 10091 2601 10100 2635
rect 10048 2592 10100 2601
rect 11060 2635 11112 2644
rect 11060 2601 11069 2635
rect 11069 2601 11103 2635
rect 11103 2601 11112 2635
rect 11060 2592 11112 2601
rect 11428 2635 11480 2644
rect 11428 2601 11437 2635
rect 11437 2601 11471 2635
rect 11471 2601 11480 2635
rect 11428 2592 11480 2601
rect 12072 2592 12124 2644
rect 5632 2499 5684 2508
rect 5632 2465 5641 2499
rect 5641 2465 5675 2499
rect 5675 2465 5684 2499
rect 5632 2456 5684 2465
rect 5908 2456 5960 2508
rect 8024 2499 8076 2508
rect 8024 2465 8033 2499
rect 8033 2465 8067 2499
rect 8067 2465 8076 2499
rect 8760 2524 8812 2576
rect 9496 2524 9548 2576
rect 11152 2524 11204 2576
rect 8024 2456 8076 2465
rect 9404 2456 9456 2508
rect 9680 2456 9732 2508
rect 12624 2499 12676 2508
rect 12624 2465 12633 2499
rect 12633 2465 12667 2499
rect 12667 2465 12676 2499
rect 12624 2456 12676 2465
rect 3976 2320 4028 2372
rect 8392 2320 8444 2372
rect 11428 2388 11480 2440
rect 12808 2363 12860 2372
rect 12808 2329 12817 2363
rect 12817 2329 12851 2363
rect 12851 2329 12860 2363
rect 12808 2320 12860 2329
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 7104 2252 7156 2261
rect 3648 2150 3700 2202
rect 3712 2150 3764 2202
rect 3776 2150 3828 2202
rect 3840 2150 3892 2202
rect 8982 2150 9034 2202
rect 9046 2150 9098 2202
rect 9110 2150 9162 2202
rect 9174 2150 9226 2202
rect 14315 2150 14367 2202
rect 14379 2150 14431 2202
rect 14443 2150 14495 2202
rect 14507 2150 14559 2202
rect 9956 620 10008 672
rect 9864 552 9916 604
rect 10600 552 10652 604
rect 10968 552 11020 604
<< metal2 >>
rect 202 39520 258 40000
rect 570 39520 626 40000
rect 938 39520 994 40000
rect 1398 39520 1454 40000
rect 1766 39520 1822 40000
rect 2134 39520 2190 40000
rect 2594 39520 2650 40000
rect 2962 39520 3018 40000
rect 3330 39520 3386 40000
rect 3790 39520 3846 40000
rect 4158 39520 4214 40000
rect 4526 39520 4582 40000
rect 4986 39520 5042 40000
rect 5354 39520 5410 40000
rect 5722 39520 5778 40000
rect 6182 39520 6238 40000
rect 6550 39520 6606 40000
rect 6918 39520 6974 40000
rect 7378 39520 7434 40000
rect 7746 39520 7802 40000
rect 8206 39520 8262 40000
rect 8574 39520 8630 40000
rect 8942 39520 8998 40000
rect 9402 39520 9458 40000
rect 9770 39520 9826 40000
rect 10138 39520 10194 40000
rect 10598 39520 10654 40000
rect 10966 39522 11022 40000
rect 10966 39520 11100 39522
rect 11334 39520 11390 40000
rect 11794 39520 11850 40000
rect 12162 39520 12218 40000
rect 12530 39520 12586 40000
rect 12990 39520 13046 40000
rect 13358 39520 13414 40000
rect 13726 39522 13782 40000
rect 13648 39520 13782 39522
rect 14186 39520 14242 40000
rect 14554 39520 14610 40000
rect 14922 39520 14978 40000
rect 15382 39520 15438 40000
rect 15750 39520 15806 40000
rect 216 34785 244 39520
rect 584 35290 612 39520
rect 572 35284 624 35290
rect 572 35226 624 35232
rect 202 34776 258 34785
rect 202 34711 258 34720
rect 952 33658 980 39520
rect 1412 35018 1440 39520
rect 1582 38720 1638 38729
rect 1582 38655 1638 38664
rect 1490 36408 1546 36417
rect 1490 36343 1546 36352
rect 1400 35012 1452 35018
rect 1400 34954 1452 34960
rect 1504 34134 1532 36343
rect 1596 34610 1624 38655
rect 1584 34604 1636 34610
rect 1584 34546 1636 34552
rect 1780 34542 1808 39520
rect 1952 35148 2004 35154
rect 1952 35090 2004 35096
rect 1964 34746 1992 35090
rect 2148 35057 2176 39520
rect 2608 35329 2636 39520
rect 2976 35737 3004 39520
rect 2962 35728 3018 35737
rect 2962 35663 3018 35672
rect 2594 35320 2650 35329
rect 2594 35255 2650 35264
rect 2504 35148 2556 35154
rect 2504 35090 2556 35096
rect 2134 35048 2190 35057
rect 2134 34983 2190 34992
rect 2044 34944 2096 34950
rect 2044 34886 2096 34892
rect 1952 34740 2004 34746
rect 1952 34682 2004 34688
rect 1768 34536 1820 34542
rect 1768 34478 1820 34484
rect 1964 34241 1992 34682
rect 2056 34610 2084 34886
rect 2516 34746 2544 35090
rect 3238 34776 3294 34785
rect 2504 34740 2556 34746
rect 3238 34711 3240 34720
rect 2504 34682 2556 34688
rect 3292 34711 3294 34720
rect 3240 34682 3292 34688
rect 2044 34604 2096 34610
rect 2044 34546 2096 34552
rect 1950 34232 2006 34241
rect 1950 34167 2006 34176
rect 1492 34128 1544 34134
rect 1492 34070 1544 34076
rect 1674 34096 1730 34105
rect 1674 34031 1730 34040
rect 940 33652 992 33658
rect 940 33594 992 33600
rect 1688 33046 1716 34031
rect 2056 33969 2084 34546
rect 2516 34105 2544 34682
rect 3344 34610 3372 39520
rect 3804 37210 3832 39520
rect 3804 37182 4016 37210
rect 3622 37020 3918 37040
rect 3678 37018 3702 37020
rect 3758 37018 3782 37020
rect 3838 37018 3862 37020
rect 3700 36966 3702 37018
rect 3764 36966 3776 37018
rect 3838 36966 3840 37018
rect 3678 36964 3702 36966
rect 3758 36964 3782 36966
rect 3838 36964 3862 36966
rect 3622 36944 3918 36964
rect 3622 35932 3918 35952
rect 3678 35930 3702 35932
rect 3758 35930 3782 35932
rect 3838 35930 3862 35932
rect 3700 35878 3702 35930
rect 3764 35878 3776 35930
rect 3838 35878 3840 35930
rect 3678 35876 3702 35878
rect 3758 35876 3782 35878
rect 3838 35876 3862 35878
rect 3622 35856 3918 35876
rect 3622 34844 3918 34864
rect 3678 34842 3702 34844
rect 3758 34842 3782 34844
rect 3838 34842 3862 34844
rect 3700 34790 3702 34842
rect 3764 34790 3776 34842
rect 3838 34790 3840 34842
rect 3678 34788 3702 34790
rect 3758 34788 3782 34790
rect 3838 34788 3862 34790
rect 3622 34768 3918 34788
rect 3988 34678 4016 37182
rect 4068 35148 4120 35154
rect 4068 35090 4120 35096
rect 3700 34672 3752 34678
rect 3698 34640 3700 34649
rect 3976 34672 4028 34678
rect 3752 34640 3754 34649
rect 3332 34604 3384 34610
rect 3976 34614 4028 34620
rect 3698 34575 3754 34584
rect 3332 34546 3384 34552
rect 4080 34542 4108 35090
rect 4068 34536 4120 34542
rect 4068 34478 4120 34484
rect 2780 34468 2832 34474
rect 2780 34410 2832 34416
rect 2792 34202 2820 34410
rect 2780 34196 2832 34202
rect 2780 34138 2832 34144
rect 2502 34096 2558 34105
rect 2412 34060 2464 34066
rect 2502 34031 2558 34040
rect 3056 34060 3108 34066
rect 2412 34002 2464 34008
rect 3056 34002 3108 34008
rect 3976 34060 4028 34066
rect 3976 34002 4028 34008
rect 2042 33960 2098 33969
rect 2042 33895 2098 33904
rect 2424 33590 2452 34002
rect 2412 33584 2464 33590
rect 2410 33552 2412 33561
rect 2464 33552 2466 33561
rect 2410 33487 2466 33496
rect 1952 33448 2004 33454
rect 1952 33390 2004 33396
rect 1676 33040 1728 33046
rect 1398 33008 1454 33017
rect 1676 32982 1728 32988
rect 1398 32943 1400 32952
rect 1452 32943 1454 32952
rect 1400 32914 1452 32920
rect 1412 32570 1440 32914
rect 1400 32564 1452 32570
rect 1400 32506 1452 32512
rect 1674 31648 1730 31657
rect 1674 31583 1730 31592
rect 1688 29782 1716 31583
rect 1964 30841 1992 33390
rect 3068 33318 3096 34002
rect 3622 33756 3918 33776
rect 3678 33754 3702 33756
rect 3758 33754 3782 33756
rect 3838 33754 3862 33756
rect 3700 33702 3702 33754
rect 3764 33702 3776 33754
rect 3838 33702 3840 33754
rect 3678 33700 3702 33702
rect 3758 33700 3782 33702
rect 3838 33700 3862 33702
rect 3622 33680 3918 33700
rect 3988 33318 4016 34002
rect 3056 33312 3108 33318
rect 3056 33254 3108 33260
rect 3976 33312 4028 33318
rect 3976 33254 4028 33260
rect 1950 30832 2006 30841
rect 1950 30767 2006 30776
rect 2228 30592 2280 30598
rect 2228 30534 2280 30540
rect 2134 30152 2190 30161
rect 2134 30087 2136 30096
rect 2188 30087 2190 30096
rect 2136 30058 2188 30064
rect 1768 30048 1820 30054
rect 1768 29990 1820 29996
rect 1676 29776 1728 29782
rect 1676 29718 1728 29724
rect 1780 29714 1808 29990
rect 2148 29850 2176 30058
rect 2240 30054 2268 30534
rect 2410 30288 2466 30297
rect 2410 30223 2412 30232
rect 2464 30223 2466 30232
rect 2412 30194 2464 30200
rect 2228 30048 2280 30054
rect 2226 30016 2228 30025
rect 2280 30016 2282 30025
rect 2226 29951 2282 29960
rect 2136 29844 2188 29850
rect 2136 29786 2188 29792
rect 1768 29708 1820 29714
rect 1768 29650 1820 29656
rect 1780 29306 1808 29650
rect 1768 29300 1820 29306
rect 1768 29242 1820 29248
rect 1582 28928 1638 28937
rect 1582 28863 1638 28872
rect 1596 28082 1624 28863
rect 1584 28076 1636 28082
rect 1584 28018 1636 28024
rect 2228 27872 2280 27878
rect 2228 27814 2280 27820
rect 2240 27577 2268 27814
rect 3068 27606 3096 33254
rect 3622 32668 3918 32688
rect 3678 32666 3702 32668
rect 3758 32666 3782 32668
rect 3838 32666 3862 32668
rect 3700 32614 3702 32666
rect 3764 32614 3776 32666
rect 3838 32614 3840 32666
rect 3678 32612 3702 32614
rect 3758 32612 3782 32614
rect 3838 32612 3862 32614
rect 3622 32592 3918 32612
rect 3622 31580 3918 31600
rect 3678 31578 3702 31580
rect 3758 31578 3782 31580
rect 3838 31578 3862 31580
rect 3700 31526 3702 31578
rect 3764 31526 3776 31578
rect 3838 31526 3840 31578
rect 3678 31524 3702 31526
rect 3758 31524 3782 31526
rect 3838 31524 3862 31526
rect 3622 31504 3918 31524
rect 3622 30492 3918 30512
rect 3678 30490 3702 30492
rect 3758 30490 3782 30492
rect 3838 30490 3862 30492
rect 3700 30438 3702 30490
rect 3764 30438 3776 30490
rect 3838 30438 3840 30490
rect 3678 30436 3702 30438
rect 3758 30436 3782 30438
rect 3838 30436 3862 30438
rect 3622 30416 3918 30436
rect 3332 30184 3384 30190
rect 3332 30126 3384 30132
rect 3344 29578 3372 30126
rect 3332 29572 3384 29578
rect 3332 29514 3384 29520
rect 3516 29504 3568 29510
rect 3516 29446 3568 29452
rect 3424 29096 3476 29102
rect 3424 29038 3476 29044
rect 3056 27600 3108 27606
rect 2226 27568 2282 27577
rect 3056 27542 3108 27548
rect 3332 27600 3384 27606
rect 3332 27542 3384 27548
rect 2226 27503 2282 27512
rect 1582 24576 1638 24585
rect 1582 24511 1638 24520
rect 1596 21554 1624 24511
rect 1674 22264 1730 22273
rect 1674 22199 1730 22208
rect 1584 21548 1636 21554
rect 1584 21490 1636 21496
rect 1688 21078 1716 22199
rect 2412 21344 2464 21350
rect 2412 21286 2464 21292
rect 1676 21072 1728 21078
rect 1676 21014 1728 21020
rect 1676 20936 1728 20942
rect 1676 20878 1728 20884
rect 1398 20360 1454 20369
rect 1398 20295 1454 20304
rect 1412 19310 1440 20295
rect 1688 20262 1716 20878
rect 1676 20256 1728 20262
rect 1674 20224 1676 20233
rect 1728 20224 1730 20233
rect 1674 20159 1730 20168
rect 2424 20058 2452 21286
rect 2596 21140 2648 21146
rect 2596 21082 2648 21088
rect 2608 20466 2636 21082
rect 2596 20460 2648 20466
rect 2596 20402 2648 20408
rect 2964 20256 3016 20262
rect 2964 20198 3016 20204
rect 2412 20052 2464 20058
rect 2412 19994 2464 20000
rect 2872 19984 2924 19990
rect 1674 19952 1730 19961
rect 2872 19926 2924 19932
rect 1674 19887 1730 19896
rect 2780 19916 2832 19922
rect 1688 19310 1716 19887
rect 2780 19858 2832 19864
rect 2792 19446 2820 19858
rect 2780 19440 2832 19446
rect 2780 19382 2832 19388
rect 1400 19304 1452 19310
rect 1400 19246 1452 19252
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 1412 18970 1440 19246
rect 2792 18970 2820 19382
rect 2884 19174 2912 19926
rect 2976 19854 3004 20198
rect 2964 19848 3016 19854
rect 2964 19790 3016 19796
rect 2976 19378 3004 19790
rect 2964 19372 3016 19378
rect 2964 19314 3016 19320
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 2884 18970 2912 19110
rect 1400 18964 1452 18970
rect 1400 18906 1452 18912
rect 2780 18964 2832 18970
rect 2780 18906 2832 18912
rect 2872 18964 2924 18970
rect 2872 18906 2924 18912
rect 3240 18624 3292 18630
rect 3240 18566 3292 18572
rect 3252 18222 3280 18566
rect 3240 18216 3292 18222
rect 3240 18158 3292 18164
rect 3344 18057 3372 27542
rect 3436 22778 3464 29038
rect 3528 28218 3556 29446
rect 3622 29404 3918 29424
rect 3678 29402 3702 29404
rect 3758 29402 3782 29404
rect 3838 29402 3862 29404
rect 3700 29350 3702 29402
rect 3764 29350 3776 29402
rect 3838 29350 3840 29402
rect 3678 29348 3702 29350
rect 3758 29348 3782 29350
rect 3838 29348 3862 29350
rect 3622 29328 3918 29348
rect 3698 29064 3754 29073
rect 3698 28999 3754 29008
rect 3712 28762 3740 28999
rect 3700 28756 3752 28762
rect 3700 28698 3752 28704
rect 3622 28316 3918 28336
rect 3678 28314 3702 28316
rect 3758 28314 3782 28316
rect 3838 28314 3862 28316
rect 3700 28262 3702 28314
rect 3764 28262 3776 28314
rect 3838 28262 3840 28314
rect 3678 28260 3702 28262
rect 3758 28260 3782 28262
rect 3838 28260 3862 28262
rect 3622 28240 3918 28260
rect 3516 28212 3568 28218
rect 3516 28154 3568 28160
rect 3622 27228 3918 27248
rect 3678 27226 3702 27228
rect 3758 27226 3782 27228
rect 3838 27226 3862 27228
rect 3700 27174 3702 27226
rect 3764 27174 3776 27226
rect 3838 27174 3840 27226
rect 3678 27172 3702 27174
rect 3758 27172 3782 27174
rect 3838 27172 3862 27174
rect 3622 27152 3918 27172
rect 3622 26140 3918 26160
rect 3678 26138 3702 26140
rect 3758 26138 3782 26140
rect 3838 26138 3862 26140
rect 3700 26086 3702 26138
rect 3764 26086 3776 26138
rect 3838 26086 3840 26138
rect 3678 26084 3702 26086
rect 3758 26084 3782 26086
rect 3838 26084 3862 26086
rect 3622 26064 3918 26084
rect 3622 25052 3918 25072
rect 3678 25050 3702 25052
rect 3758 25050 3782 25052
rect 3838 25050 3862 25052
rect 3700 24998 3702 25050
rect 3764 24998 3776 25050
rect 3838 24998 3840 25050
rect 3678 24996 3702 24998
rect 3758 24996 3782 24998
rect 3838 24996 3862 24998
rect 3622 24976 3918 24996
rect 3622 23964 3918 23984
rect 3678 23962 3702 23964
rect 3758 23962 3782 23964
rect 3838 23962 3862 23964
rect 3700 23910 3702 23962
rect 3764 23910 3776 23962
rect 3838 23910 3840 23962
rect 3678 23908 3702 23910
rect 3758 23908 3782 23910
rect 3838 23908 3862 23910
rect 3622 23888 3918 23908
rect 3622 22876 3918 22896
rect 3678 22874 3702 22876
rect 3758 22874 3782 22876
rect 3838 22874 3862 22876
rect 3700 22822 3702 22874
rect 3764 22822 3776 22874
rect 3838 22822 3840 22874
rect 3678 22820 3702 22822
rect 3758 22820 3782 22822
rect 3838 22820 3862 22822
rect 3622 22800 3918 22820
rect 3424 22772 3476 22778
rect 3424 22714 3476 22720
rect 3622 21788 3918 21808
rect 3678 21786 3702 21788
rect 3758 21786 3782 21788
rect 3838 21786 3862 21788
rect 3700 21734 3702 21786
rect 3764 21734 3776 21786
rect 3838 21734 3840 21786
rect 3678 21732 3702 21734
rect 3758 21732 3782 21734
rect 3838 21732 3862 21734
rect 3622 21712 3918 21732
rect 3988 21010 4016 33254
rect 4080 30569 4108 34478
rect 4172 33114 4200 39520
rect 4540 36922 4568 39520
rect 4528 36916 4580 36922
rect 4528 36858 4580 36864
rect 5000 36378 5028 39520
rect 4988 36372 5040 36378
rect 4988 36314 5040 36320
rect 5080 36236 5132 36242
rect 5080 36178 5132 36184
rect 4988 35556 5040 35562
rect 4988 35498 5040 35504
rect 4250 35320 4306 35329
rect 4250 35255 4252 35264
rect 4304 35255 4306 35264
rect 4252 35226 4304 35232
rect 4342 35048 4398 35057
rect 4342 34983 4398 34992
rect 4356 34746 4384 34983
rect 4344 34740 4396 34746
rect 4344 34682 4396 34688
rect 4344 34604 4396 34610
rect 4344 34546 4396 34552
rect 4252 34536 4304 34542
rect 4252 34478 4304 34484
rect 4160 33108 4212 33114
rect 4160 33050 4212 33056
rect 4160 32972 4212 32978
rect 4160 32914 4212 32920
rect 4172 32570 4200 32914
rect 4160 32564 4212 32570
rect 4160 32506 4212 32512
rect 4172 32337 4200 32506
rect 4158 32328 4214 32337
rect 4158 32263 4214 32272
rect 4264 32212 4292 34478
rect 4356 34202 4384 34546
rect 4344 34196 4396 34202
rect 4344 34138 4396 34144
rect 4894 34096 4950 34105
rect 4894 34031 4950 34040
rect 4908 33833 4936 34031
rect 4894 33824 4950 33833
rect 4894 33759 4950 33768
rect 4712 33380 4764 33386
rect 4712 33322 4764 33328
rect 4172 32184 4292 32212
rect 4172 31668 4200 32184
rect 4172 31640 4384 31668
rect 4160 31340 4212 31346
rect 4160 31282 4212 31288
rect 4066 30560 4122 30569
rect 4066 30495 4122 30504
rect 4172 30138 4200 31282
rect 4080 30110 4200 30138
rect 4080 29034 4108 30110
rect 4158 30016 4214 30025
rect 4158 29951 4214 29960
rect 4172 29850 4200 29951
rect 4160 29844 4212 29850
rect 4160 29786 4212 29792
rect 4252 29572 4304 29578
rect 4252 29514 4304 29520
rect 4068 29028 4120 29034
rect 4068 28970 4120 28976
rect 4080 28914 4108 28970
rect 4080 28886 4200 28914
rect 4068 28756 4120 28762
rect 4068 28698 4120 28704
rect 4080 28082 4108 28698
rect 4172 28082 4200 28886
rect 4264 28218 4292 29514
rect 4252 28212 4304 28218
rect 4252 28154 4304 28160
rect 4068 28076 4120 28082
rect 4068 28018 4120 28024
rect 4160 28076 4212 28082
rect 4160 28018 4212 28024
rect 4172 27962 4200 28018
rect 4080 27934 4200 27962
rect 4080 27674 4108 27934
rect 4068 27668 4120 27674
rect 4068 27610 4120 27616
rect 4080 26586 4108 27610
rect 4356 27112 4384 31640
rect 4724 30326 4752 33322
rect 4896 31816 4948 31822
rect 4896 31758 4948 31764
rect 4908 31278 4936 31758
rect 4896 31272 4948 31278
rect 4896 31214 4948 31220
rect 4804 31136 4856 31142
rect 4804 31078 4856 31084
rect 4816 30433 4844 31078
rect 4908 30938 4936 31214
rect 4896 30932 4948 30938
rect 4896 30874 4948 30880
rect 4802 30424 4858 30433
rect 4802 30359 4858 30368
rect 4712 30320 4764 30326
rect 4710 30288 4712 30297
rect 4804 30320 4856 30326
rect 4764 30288 4766 30297
rect 4804 30262 4856 30268
rect 4710 30223 4766 30232
rect 4816 30122 4844 30262
rect 4804 30116 4856 30122
rect 4804 30058 4856 30064
rect 4528 30048 4580 30054
rect 4528 29990 4580 29996
rect 4540 27282 4568 29990
rect 4816 29646 4844 30058
rect 5000 29866 5028 35498
rect 5092 35494 5120 36178
rect 5368 35834 5396 39520
rect 5736 35834 5764 39520
rect 6196 36378 6224 39520
rect 6564 37754 6592 39520
rect 6564 37726 6684 37754
rect 6289 37564 6585 37584
rect 6345 37562 6369 37564
rect 6425 37562 6449 37564
rect 6505 37562 6529 37564
rect 6367 37510 6369 37562
rect 6431 37510 6443 37562
rect 6505 37510 6507 37562
rect 6345 37508 6369 37510
rect 6425 37508 6449 37510
rect 6505 37508 6529 37510
rect 6289 37488 6585 37508
rect 6289 36476 6585 36496
rect 6345 36474 6369 36476
rect 6425 36474 6449 36476
rect 6505 36474 6529 36476
rect 6367 36422 6369 36474
rect 6431 36422 6443 36474
rect 6505 36422 6507 36474
rect 6345 36420 6369 36422
rect 6425 36420 6449 36422
rect 6505 36420 6529 36422
rect 6289 36400 6585 36420
rect 6184 36372 6236 36378
rect 6184 36314 6236 36320
rect 5356 35828 5408 35834
rect 5356 35770 5408 35776
rect 5724 35828 5776 35834
rect 5724 35770 5776 35776
rect 5080 35488 5132 35494
rect 5080 35430 5132 35436
rect 6184 35488 6236 35494
rect 6184 35430 6236 35436
rect 5092 32212 5120 35430
rect 5448 35148 5500 35154
rect 5448 35090 5500 35096
rect 5460 34542 5488 35090
rect 5724 34944 5776 34950
rect 5724 34886 5776 34892
rect 5448 34536 5500 34542
rect 5448 34478 5500 34484
rect 5264 34400 5316 34406
rect 5264 34342 5316 34348
rect 5170 34096 5226 34105
rect 5170 34031 5226 34040
rect 5184 32570 5212 34031
rect 5172 32564 5224 32570
rect 5172 32506 5224 32512
rect 5276 32366 5304 34342
rect 5356 33448 5408 33454
rect 5356 33390 5408 33396
rect 5368 32978 5396 33390
rect 5356 32972 5408 32978
rect 5356 32914 5408 32920
rect 5264 32360 5316 32366
rect 5264 32302 5316 32308
rect 5092 32184 5304 32212
rect 5276 31668 5304 32184
rect 5368 32026 5396 32914
rect 5356 32020 5408 32026
rect 5356 31962 5408 31968
rect 5184 31640 5304 31668
rect 5080 30796 5132 30802
rect 5080 30738 5132 30744
rect 5092 30054 5120 30738
rect 5080 30048 5132 30054
rect 5080 29990 5132 29996
rect 4908 29838 5028 29866
rect 4804 29640 4856 29646
rect 4804 29582 4856 29588
rect 4816 29306 4844 29582
rect 4804 29300 4856 29306
rect 4804 29242 4856 29248
rect 4620 28960 4672 28966
rect 4620 28902 4672 28908
rect 4632 28014 4660 28902
rect 4816 28762 4844 29242
rect 4804 28756 4856 28762
rect 4804 28698 4856 28704
rect 4620 28008 4672 28014
rect 4620 27950 4672 27956
rect 4632 27441 4660 27950
rect 4712 27668 4764 27674
rect 4712 27610 4764 27616
rect 4618 27432 4674 27441
rect 4618 27367 4674 27376
rect 4540 27254 4660 27282
rect 4172 27084 4384 27112
rect 4068 26580 4120 26586
rect 4068 26522 4120 26528
rect 4068 25356 4120 25362
rect 4068 25298 4120 25304
rect 4080 24682 4108 25298
rect 4068 24676 4120 24682
rect 4068 24618 4120 24624
rect 4172 23769 4200 27084
rect 4342 27024 4398 27033
rect 4342 26959 4398 26968
rect 4356 25430 4384 26959
rect 4344 25424 4396 25430
rect 4344 25366 4396 25372
rect 4436 24064 4488 24070
rect 4436 24006 4488 24012
rect 4158 23760 4214 23769
rect 4448 23730 4476 24006
rect 4158 23695 4214 23704
rect 4436 23724 4488 23730
rect 4068 23180 4120 23186
rect 4068 23122 4120 23128
rect 4080 22778 4108 23122
rect 4068 22772 4120 22778
rect 4068 22714 4120 22720
rect 4068 22636 4120 22642
rect 4068 22578 4120 22584
rect 4080 22166 4108 22578
rect 4172 22216 4200 23695
rect 4436 23666 4488 23672
rect 4344 23520 4396 23526
rect 4344 23462 4396 23468
rect 4252 22976 4304 22982
rect 4252 22918 4304 22924
rect 4264 22642 4292 22918
rect 4252 22636 4304 22642
rect 4252 22578 4304 22584
rect 4172 22188 4292 22216
rect 4068 22160 4120 22166
rect 4068 22102 4120 22108
rect 4080 22030 4108 22102
rect 4160 22092 4212 22098
rect 4160 22034 4212 22040
rect 4068 22024 4120 22030
rect 4068 21966 4120 21972
rect 4080 21690 4108 21966
rect 4068 21684 4120 21690
rect 4068 21626 4120 21632
rect 4080 21146 4108 21626
rect 4172 21350 4200 22034
rect 4160 21344 4212 21350
rect 4264 21332 4292 22188
rect 4356 21486 4384 23462
rect 4448 22778 4476 23666
rect 4436 22772 4488 22778
rect 4436 22714 4488 22720
rect 4448 22506 4476 22714
rect 4436 22500 4488 22506
rect 4436 22442 4488 22448
rect 4448 22234 4476 22442
rect 4436 22228 4488 22234
rect 4436 22170 4488 22176
rect 4344 21480 4396 21486
rect 4344 21422 4396 21428
rect 4264 21304 4384 21332
rect 4160 21286 4212 21292
rect 4068 21140 4120 21146
rect 4068 21082 4120 21088
rect 3976 21004 4028 21010
rect 3976 20946 4028 20952
rect 3622 20700 3918 20720
rect 3678 20698 3702 20700
rect 3758 20698 3782 20700
rect 3838 20698 3862 20700
rect 3700 20646 3702 20698
rect 3764 20646 3776 20698
rect 3838 20646 3840 20698
rect 3678 20644 3702 20646
rect 3758 20644 3782 20646
rect 3838 20644 3862 20646
rect 3622 20624 3918 20644
rect 3516 20324 3568 20330
rect 3516 20266 3568 20272
rect 3528 19310 3556 20266
rect 4172 20262 4200 21286
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 4252 19712 4304 19718
rect 4252 19654 4304 19660
rect 3622 19612 3918 19632
rect 3678 19610 3702 19612
rect 3758 19610 3782 19612
rect 3838 19610 3862 19612
rect 3700 19558 3702 19610
rect 3764 19558 3776 19610
rect 3838 19558 3840 19610
rect 3678 19556 3702 19558
rect 3758 19556 3782 19558
rect 3838 19556 3862 19558
rect 3622 19536 3918 19556
rect 4264 19378 4292 19654
rect 4252 19372 4304 19378
rect 4252 19314 4304 19320
rect 3516 19304 3568 19310
rect 3516 19246 3568 19252
rect 3528 18902 3556 19246
rect 3976 19168 4028 19174
rect 3976 19110 4028 19116
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 3516 18896 3568 18902
rect 3516 18838 3568 18844
rect 3622 18524 3918 18544
rect 3678 18522 3702 18524
rect 3758 18522 3782 18524
rect 3838 18522 3862 18524
rect 3700 18470 3702 18522
rect 3764 18470 3776 18522
rect 3838 18470 3840 18522
rect 3678 18468 3702 18470
rect 3758 18468 3782 18470
rect 3838 18468 3862 18470
rect 3622 18448 3918 18468
rect 3988 18086 4016 19110
rect 4172 18698 4200 19110
rect 4356 18850 4384 21304
rect 4632 21162 4660 27254
rect 4724 23594 4752 27610
rect 4804 24200 4856 24206
rect 4804 24142 4856 24148
rect 4816 23633 4844 24142
rect 4802 23624 4858 23633
rect 4712 23588 4764 23594
rect 4802 23559 4858 23568
rect 4712 23530 4764 23536
rect 4724 23322 4752 23530
rect 4712 23316 4764 23322
rect 4712 23258 4764 23264
rect 4264 18822 4384 18850
rect 4448 21134 4660 21162
rect 4160 18692 4212 18698
rect 4160 18634 4212 18640
rect 4068 18148 4120 18154
rect 4068 18090 4120 18096
rect 3792 18080 3844 18086
rect 3054 18048 3110 18057
rect 3054 17983 3110 17992
rect 3330 18048 3386 18057
rect 3792 18022 3844 18028
rect 3976 18080 4028 18086
rect 3976 18022 4028 18028
rect 3330 17983 3386 17992
rect 2778 17776 2834 17785
rect 2778 17711 2780 17720
rect 2832 17711 2834 17720
rect 2780 17682 2832 17688
rect 1582 17640 1638 17649
rect 1582 17575 1638 17584
rect 1596 16114 1624 17575
rect 2792 17338 2820 17682
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2884 17134 2912 17614
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 1584 16108 1636 16114
rect 1584 16050 1636 16056
rect 2228 15904 2280 15910
rect 2226 15872 2228 15881
rect 2280 15872 2282 15881
rect 2226 15807 2282 15816
rect 1674 15192 1730 15201
rect 1674 15127 1730 15136
rect 1688 13462 1716 15127
rect 3068 14498 3096 17983
rect 3804 17814 3832 18022
rect 3792 17808 3844 17814
rect 3792 17750 3844 17756
rect 3622 17436 3918 17456
rect 3678 17434 3702 17436
rect 3758 17434 3782 17436
rect 3838 17434 3862 17436
rect 3700 17382 3702 17434
rect 3764 17382 3776 17434
rect 3838 17382 3840 17434
rect 3678 17380 3702 17382
rect 3758 17380 3782 17382
rect 3838 17380 3862 17382
rect 3622 17360 3918 17380
rect 3988 17202 4016 18022
rect 4080 17678 4108 18090
rect 4068 17672 4120 17678
rect 4068 17614 4120 17620
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 4160 17128 4212 17134
rect 3974 17096 4030 17105
rect 4160 17070 4212 17076
rect 3974 17031 4030 17040
rect 3988 16998 4016 17031
rect 3976 16992 4028 16998
rect 3976 16934 4028 16940
rect 3988 16794 4016 16934
rect 3976 16788 4028 16794
rect 3976 16730 4028 16736
rect 3622 16348 3918 16368
rect 3678 16346 3702 16348
rect 3758 16346 3782 16348
rect 3838 16346 3862 16348
rect 3700 16294 3702 16346
rect 3764 16294 3776 16346
rect 3838 16294 3840 16346
rect 3678 16292 3702 16294
rect 3758 16292 3782 16294
rect 3838 16292 3862 16294
rect 3622 16272 3918 16292
rect 4172 16250 4200 17070
rect 4264 17066 4292 18822
rect 4344 18760 4396 18766
rect 4344 18702 4396 18708
rect 4356 17882 4384 18702
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4252 17060 4304 17066
rect 4252 17002 4304 17008
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 3622 15260 3918 15280
rect 3678 15258 3702 15260
rect 3758 15258 3782 15260
rect 3838 15258 3862 15260
rect 3700 15206 3702 15258
rect 3764 15206 3776 15258
rect 3838 15206 3840 15258
rect 3678 15204 3702 15206
rect 3758 15204 3782 15206
rect 3838 15204 3862 15206
rect 3622 15184 3918 15204
rect 3148 14952 3200 14958
rect 3148 14894 3200 14900
rect 3160 14618 3188 14894
rect 3976 14884 4028 14890
rect 3976 14826 4028 14832
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 2976 14470 3096 14498
rect 2780 13864 2832 13870
rect 2318 13832 2374 13841
rect 2780 13806 2832 13812
rect 2318 13767 2374 13776
rect 1676 13456 1728 13462
rect 1398 13424 1454 13433
rect 1676 13398 1728 13404
rect 1398 13359 1400 13368
rect 1452 13359 1454 13368
rect 1400 13330 1452 13336
rect 1412 12442 1440 13330
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 1582 12880 1638 12889
rect 1582 12815 1638 12824
rect 1400 12436 1452 12442
rect 1400 12378 1452 12384
rect 1596 10674 1624 12815
rect 2240 12782 2268 13126
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1492 10600 1544 10606
rect 1492 10542 1544 10548
rect 1582 10568 1638 10577
rect 1504 6905 1532 10542
rect 1582 10503 1638 10512
rect 1596 8498 1624 10503
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1582 8120 1638 8129
rect 1582 8055 1638 8064
rect 1596 7410 1624 8055
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1688 7449 1716 7686
rect 2056 7546 2084 12582
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 1674 7440 1730 7449
rect 1584 7404 1636 7410
rect 2056 7426 2084 7482
rect 2056 7398 2176 7426
rect 1674 7375 1730 7384
rect 1584 7346 1636 7352
rect 1688 7342 1716 7375
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 1490 6896 1546 6905
rect 2148 6866 2176 7398
rect 1490 6831 1546 6840
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 1584 6792 1636 6798
rect 1398 6760 1454 6769
rect 1584 6734 1636 6740
rect 1398 6695 1454 6704
rect 570 4312 626 4321
rect 570 4247 626 4256
rect 204 4140 256 4146
rect 204 4082 256 4088
rect 216 480 244 4082
rect 584 480 612 4247
rect 938 3632 994 3641
rect 938 3567 994 3576
rect 952 480 980 3567
rect 1412 480 1440 6695
rect 1492 5840 1544 5846
rect 1596 5817 1624 6734
rect 2228 6180 2280 6186
rect 2228 6122 2280 6128
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1492 5782 1544 5788
rect 1582 5808 1638 5817
rect 1504 4690 1532 5782
rect 1582 5743 1638 5752
rect 1688 5166 1716 6054
rect 1952 5772 2004 5778
rect 1952 5714 2004 5720
rect 1860 5568 1912 5574
rect 1860 5510 1912 5516
rect 1872 5234 1900 5510
rect 1964 5370 1992 5714
rect 2240 5574 2268 6122
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 2240 5302 2268 5510
rect 2228 5296 2280 5302
rect 2228 5238 2280 5244
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 1676 5160 1728 5166
rect 1676 5102 1728 5108
rect 2332 4690 2360 13767
rect 2792 13190 2820 13806
rect 2780 13184 2832 13190
rect 2780 13126 2832 13132
rect 2686 12880 2742 12889
rect 2686 12815 2688 12824
rect 2740 12815 2742 12824
rect 2688 12786 2740 12792
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 2516 12102 2544 12582
rect 2976 12374 3004 14470
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 3344 14090 3372 14214
rect 3622 14172 3918 14192
rect 3678 14170 3702 14172
rect 3758 14170 3782 14172
rect 3838 14170 3862 14172
rect 3700 14118 3702 14170
rect 3764 14118 3776 14170
rect 3838 14118 3840 14170
rect 3678 14116 3702 14118
rect 3758 14116 3782 14118
rect 3838 14116 3862 14118
rect 3622 14096 3918 14116
rect 3344 14074 3464 14090
rect 3344 14068 3476 14074
rect 3344 14062 3424 14068
rect 3344 13870 3372 14062
rect 3424 14010 3476 14016
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 3988 13734 4016 14826
rect 4068 14340 4120 14346
rect 4068 14282 4120 14288
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3160 12986 3188 13126
rect 3622 13084 3918 13104
rect 3678 13082 3702 13084
rect 3758 13082 3782 13084
rect 3838 13082 3862 13084
rect 3700 13030 3702 13082
rect 3764 13030 3776 13082
rect 3838 13030 3840 13082
rect 3678 13028 3702 13030
rect 3758 13028 3782 13030
rect 3838 13028 3862 13030
rect 3622 13008 3918 13028
rect 3988 12986 4016 13670
rect 4080 13530 4108 14282
rect 4160 14000 4212 14006
rect 4160 13942 4212 13948
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 2964 12368 3016 12374
rect 2964 12310 3016 12316
rect 3148 12368 3200 12374
rect 3148 12310 3200 12316
rect 2504 12096 2556 12102
rect 2504 12038 2556 12044
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 2976 11898 3004 12038
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2792 11098 2820 11290
rect 2700 11070 2820 11098
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2424 10266 2452 10406
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2424 9586 2452 10202
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 2516 6866 2544 10202
rect 2700 9654 2728 11070
rect 2688 9648 2740 9654
rect 2688 9590 2740 9596
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2608 9178 2636 9454
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 2700 8945 2728 9318
rect 2686 8936 2742 8945
rect 2686 8871 2742 8880
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2884 8430 2912 8774
rect 2872 8424 2924 8430
rect 2778 8392 2834 8401
rect 2688 8356 2740 8362
rect 2872 8366 2924 8372
rect 2778 8327 2834 8336
rect 2688 8298 2740 8304
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2424 5778 2452 6598
rect 2516 6458 2544 6802
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2700 6118 2728 8298
rect 2792 8294 2820 8327
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 2884 8090 2912 8366
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 2884 7750 2912 8026
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2884 7546 2912 7686
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2884 6769 2912 7142
rect 2870 6760 2926 6769
rect 2870 6695 2926 6704
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2688 6112 2740 6118
rect 2594 6080 2650 6089
rect 2688 6054 2740 6060
rect 2594 6015 2650 6024
rect 2412 5772 2464 5778
rect 2412 5714 2464 5720
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 1492 4684 1544 4690
rect 1492 4626 1544 4632
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1596 3505 1624 4558
rect 2136 4548 2188 4554
rect 2136 4490 2188 4496
rect 1582 3496 1638 3505
rect 1582 3431 1638 3440
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 1766 2816 1822 2825
rect 1766 2751 1822 2760
rect 1780 480 1808 2751
rect 1964 2378 1992 3334
rect 1952 2372 2004 2378
rect 1952 2314 2004 2320
rect 2148 480 2176 4490
rect 2332 4298 2360 4626
rect 2240 4282 2360 4298
rect 2228 4276 2360 4282
rect 2280 4270 2360 4276
rect 2228 4218 2280 4224
rect 2424 3738 2452 5170
rect 2608 4570 2636 6015
rect 2516 4542 2636 4570
rect 2412 3732 2464 3738
rect 2412 3674 2464 3680
rect 2516 2650 2544 4542
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2792 4162 2820 4422
rect 2884 4321 2912 6598
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 3068 5710 3096 6054
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 3068 5370 3096 5646
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 2870 4312 2926 4321
rect 2870 4247 2926 4256
rect 2792 4134 2912 4162
rect 2780 4004 2832 4010
rect 2780 3946 2832 3952
rect 2792 3738 2820 3946
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 2884 3534 2912 4134
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2594 2952 2650 2961
rect 2594 2887 2650 2896
rect 2504 2644 2556 2650
rect 2504 2586 2556 2592
rect 2608 480 2636 2887
rect 2688 2848 2740 2854
rect 2740 2808 2820 2836
rect 2688 2790 2740 2796
rect 2792 1193 2820 2808
rect 2884 2650 2912 3470
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 2976 2582 3004 4014
rect 3068 3670 3096 4626
rect 3160 4214 3188 12310
rect 3252 11830 3280 12922
rect 4080 12782 4108 13466
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 4068 12640 4120 12646
rect 4172 12628 4200 13942
rect 4120 12600 4200 12628
rect 4068 12582 4120 12588
rect 4080 12442 4108 12582
rect 4264 12442 4292 17002
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 3240 11824 3292 11830
rect 3240 11766 3292 11772
rect 3528 11694 3556 12038
rect 3622 11996 3918 12016
rect 3678 11994 3702 11996
rect 3758 11994 3782 11996
rect 3838 11994 3862 11996
rect 3700 11942 3702 11994
rect 3764 11942 3776 11994
rect 3838 11942 3840 11994
rect 3678 11940 3702 11942
rect 3758 11940 3782 11942
rect 3838 11940 3862 11942
rect 3622 11920 3918 11940
rect 4344 11892 4396 11898
rect 4344 11834 4396 11840
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3620 11354 3648 11494
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 3622 10908 3918 10928
rect 3678 10906 3702 10908
rect 3758 10906 3782 10908
rect 3838 10906 3862 10908
rect 3700 10854 3702 10906
rect 3764 10854 3776 10906
rect 3838 10854 3840 10906
rect 3678 10852 3702 10854
rect 3758 10852 3782 10854
rect 3838 10852 3862 10854
rect 3622 10832 3918 10852
rect 4080 10690 4108 11018
rect 4080 10674 4200 10690
rect 4080 10668 4212 10674
rect 4080 10662 4160 10668
rect 3884 10532 3936 10538
rect 3884 10474 3936 10480
rect 3896 10266 3924 10474
rect 3884 10260 3936 10266
rect 3884 10202 3936 10208
rect 3622 9820 3918 9840
rect 3678 9818 3702 9820
rect 3758 9818 3782 9820
rect 3838 9818 3862 9820
rect 3700 9766 3702 9818
rect 3764 9766 3776 9818
rect 3838 9766 3840 9818
rect 3678 9764 3702 9766
rect 3758 9764 3782 9766
rect 3838 9764 3862 9766
rect 3622 9744 3918 9764
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3436 9382 3464 9522
rect 4080 9450 4108 10662
rect 4160 10610 4212 10616
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4264 10033 4292 10542
rect 4250 10024 4306 10033
rect 4250 9959 4306 9968
rect 4068 9444 4120 9450
rect 4068 9386 4120 9392
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3436 8838 3464 9318
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3622 8732 3918 8752
rect 3678 8730 3702 8732
rect 3758 8730 3782 8732
rect 3838 8730 3862 8732
rect 3700 8678 3702 8730
rect 3764 8678 3776 8730
rect 3838 8678 3840 8730
rect 3678 8676 3702 8678
rect 3758 8676 3782 8678
rect 3838 8676 3862 8678
rect 3622 8656 3918 8676
rect 4080 8634 4108 9386
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 3622 7644 3918 7664
rect 3678 7642 3702 7644
rect 3758 7642 3782 7644
rect 3838 7642 3862 7644
rect 3700 7590 3702 7642
rect 3764 7590 3776 7642
rect 3838 7590 3840 7642
rect 3678 7588 3702 7590
rect 3758 7588 3782 7590
rect 3838 7588 3862 7590
rect 3622 7568 3918 7588
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3528 6662 3556 7482
rect 4356 7478 4384 11834
rect 4344 7472 4396 7478
rect 4344 7414 4396 7420
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3344 5914 3372 6598
rect 3528 6254 3556 6598
rect 3622 6556 3918 6576
rect 3678 6554 3702 6556
rect 3758 6554 3782 6556
rect 3838 6554 3862 6556
rect 3700 6502 3702 6554
rect 3764 6502 3776 6554
rect 3838 6502 3840 6554
rect 3678 6500 3702 6502
rect 3758 6500 3782 6502
rect 3838 6500 3862 6502
rect 3622 6480 3918 6500
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 4080 5817 4108 6054
rect 4066 5808 4122 5817
rect 4066 5743 4122 5752
rect 3516 5568 3568 5574
rect 3516 5510 3568 5516
rect 3528 5234 3556 5510
rect 3622 5468 3918 5488
rect 3678 5466 3702 5468
rect 3758 5466 3782 5468
rect 3838 5466 3862 5468
rect 3700 5414 3702 5466
rect 3764 5414 3776 5466
rect 3838 5414 3840 5466
rect 3678 5412 3702 5414
rect 3758 5412 3782 5414
rect 3838 5412 3862 5414
rect 3622 5392 3918 5412
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 3528 4282 3556 5170
rect 3884 5024 3936 5030
rect 3882 4992 3884 5001
rect 3936 4992 3938 5001
rect 3882 4927 3938 4936
rect 3622 4380 3918 4400
rect 3678 4378 3702 4380
rect 3758 4378 3782 4380
rect 3838 4378 3862 4380
rect 3700 4326 3702 4378
rect 3764 4326 3776 4378
rect 3838 4326 3840 4378
rect 3678 4324 3702 4326
rect 3758 4324 3782 4326
rect 3838 4324 3862 4326
rect 3622 4304 3918 4324
rect 3516 4276 3568 4282
rect 3516 4218 3568 4224
rect 3148 4208 3200 4214
rect 3148 4150 3200 4156
rect 3056 3664 3108 3670
rect 3056 3606 3108 3612
rect 3976 3664 4028 3670
rect 3976 3606 4028 3612
rect 3068 3534 3096 3606
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 3332 3460 3384 3466
rect 3332 3402 3384 3408
rect 3344 3194 3372 3402
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 2964 2576 3016 2582
rect 2964 2518 3016 2524
rect 3436 2446 3464 3334
rect 3622 3292 3918 3312
rect 3678 3290 3702 3292
rect 3758 3290 3782 3292
rect 3838 3290 3862 3292
rect 3700 3238 3702 3290
rect 3764 3238 3776 3290
rect 3838 3238 3840 3290
rect 3678 3236 3702 3238
rect 3758 3236 3782 3238
rect 3838 3236 3862 3238
rect 3622 3216 3918 3236
rect 3988 3194 4016 3606
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 4066 2680 4122 2689
rect 4066 2615 4122 2624
rect 4080 2514 4108 2615
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 3424 2440 3476 2446
rect 2962 2408 3018 2417
rect 3424 2382 3476 2388
rect 2962 2343 3018 2352
rect 3976 2372 4028 2378
rect 2778 1184 2834 1193
rect 2778 1119 2834 1128
rect 2976 480 3004 2343
rect 3976 2314 4028 2320
rect 3622 2204 3918 2224
rect 3678 2202 3702 2204
rect 3758 2202 3782 2204
rect 3838 2202 3862 2204
rect 3700 2150 3702 2202
rect 3764 2150 3776 2202
rect 3838 2150 3840 2202
rect 3678 2148 3702 2150
rect 3758 2148 3782 2150
rect 3838 2148 3862 2150
rect 3622 2128 3918 2148
rect 3330 1456 3386 1465
rect 3330 1391 3386 1400
rect 3344 480 3372 1391
rect 3988 1170 4016 2314
rect 3804 1142 4016 1170
rect 3804 480 3832 1142
rect 4172 480 4200 6326
rect 4448 6186 4476 21134
rect 4724 19281 4752 23258
rect 4802 22128 4858 22137
rect 4802 22063 4858 22072
rect 4816 21690 4844 22063
rect 4804 21684 4856 21690
rect 4804 21626 4856 21632
rect 4804 19916 4856 19922
rect 4908 19904 4936 29838
rect 4988 29708 5040 29714
rect 4988 29650 5040 29656
rect 5000 28422 5028 29650
rect 5184 29034 5212 31640
rect 5356 31340 5408 31346
rect 5356 31282 5408 31288
rect 5262 31240 5318 31249
rect 5262 31175 5264 31184
rect 5316 31175 5318 31184
rect 5264 31146 5316 31152
rect 5262 30832 5318 30841
rect 5262 30767 5318 30776
rect 5276 30138 5304 30767
rect 5368 30666 5396 31282
rect 5460 30802 5488 34478
rect 5632 33856 5684 33862
rect 5632 33798 5684 33804
rect 5644 33318 5672 33798
rect 5632 33312 5684 33318
rect 5632 33254 5684 33260
rect 5540 33108 5592 33114
rect 5540 33050 5592 33056
rect 5552 32434 5580 33050
rect 5644 32978 5672 33254
rect 5736 33017 5764 34886
rect 5814 34640 5870 34649
rect 5814 34575 5870 34584
rect 5722 33008 5778 33017
rect 5632 32972 5684 32978
rect 5722 32943 5778 32952
rect 5632 32914 5684 32920
rect 5828 32858 5856 34575
rect 5906 34504 5962 34513
rect 5906 34439 5962 34448
rect 5920 34134 5948 34439
rect 5998 34232 6054 34241
rect 5998 34167 6000 34176
rect 6052 34167 6054 34176
rect 6000 34138 6052 34144
rect 5908 34128 5960 34134
rect 5908 34070 5960 34076
rect 5920 33522 5948 34070
rect 6012 33658 6040 34138
rect 6092 33992 6144 33998
rect 6092 33934 6144 33940
rect 6104 33862 6132 33934
rect 6092 33856 6144 33862
rect 6092 33798 6144 33804
rect 6196 33674 6224 35430
rect 6289 35388 6585 35408
rect 6345 35386 6369 35388
rect 6425 35386 6449 35388
rect 6505 35386 6529 35388
rect 6367 35334 6369 35386
rect 6431 35334 6443 35386
rect 6505 35334 6507 35386
rect 6345 35332 6369 35334
rect 6425 35332 6449 35334
rect 6505 35332 6529 35334
rect 6289 35312 6585 35332
rect 6656 35290 6684 37726
rect 6736 36236 6788 36242
rect 6736 36178 6788 36184
rect 6748 35494 6776 36178
rect 6932 35834 6960 39520
rect 6920 35828 6972 35834
rect 6920 35770 6972 35776
rect 6736 35488 6788 35494
rect 6736 35430 6788 35436
rect 6644 35284 6696 35290
rect 6644 35226 6696 35232
rect 6289 34300 6585 34320
rect 6345 34298 6369 34300
rect 6425 34298 6449 34300
rect 6505 34298 6529 34300
rect 6367 34246 6369 34298
rect 6431 34246 6443 34298
rect 6505 34246 6507 34298
rect 6345 34244 6369 34246
rect 6425 34244 6449 34246
rect 6505 34244 6529 34246
rect 6289 34224 6585 34244
rect 6550 33824 6606 33833
rect 6550 33759 6606 33768
rect 6000 33652 6052 33658
rect 6000 33594 6052 33600
rect 6104 33646 6224 33674
rect 6564 33658 6592 33759
rect 6552 33652 6604 33658
rect 5908 33516 5960 33522
rect 5908 33458 5960 33464
rect 6012 33425 6040 33594
rect 5998 33416 6054 33425
rect 5998 33351 6054 33360
rect 5736 32830 5856 32858
rect 5906 32872 5962 32881
rect 5540 32428 5592 32434
rect 5540 32370 5592 32376
rect 5736 31770 5764 32830
rect 5906 32807 5962 32816
rect 5716 31742 5764 31770
rect 5716 31668 5744 31742
rect 5716 31640 5764 31668
rect 5538 30832 5594 30841
rect 5448 30796 5500 30802
rect 5538 30767 5594 30776
rect 5448 30738 5500 30744
rect 5552 30734 5580 30767
rect 5540 30728 5592 30734
rect 5540 30670 5592 30676
rect 5356 30660 5408 30666
rect 5356 30602 5408 30608
rect 5368 30240 5396 30602
rect 5552 30410 5580 30670
rect 5552 30382 5672 30410
rect 5540 30252 5592 30258
rect 5368 30212 5540 30240
rect 5540 30194 5592 30200
rect 5276 30110 5396 30138
rect 5172 29028 5224 29034
rect 5172 28970 5224 28976
rect 5264 28960 5316 28966
rect 5264 28902 5316 28908
rect 5276 28626 5304 28902
rect 5264 28620 5316 28626
rect 5264 28562 5316 28568
rect 5276 28422 5304 28562
rect 4988 28416 5040 28422
rect 4988 28358 5040 28364
rect 5264 28416 5316 28422
rect 5264 28358 5316 28364
rect 5000 27130 5028 28358
rect 5276 28082 5304 28358
rect 5264 28076 5316 28082
rect 5264 28018 5316 28024
rect 5080 27940 5132 27946
rect 5080 27882 5132 27888
rect 4988 27124 5040 27130
rect 4988 27066 5040 27072
rect 4988 26852 5040 26858
rect 4988 26794 5040 26800
rect 5000 26586 5028 26794
rect 4988 26580 5040 26586
rect 4988 26522 5040 26528
rect 5092 23594 5120 27882
rect 5172 27872 5224 27878
rect 5172 27814 5224 27820
rect 5184 26994 5212 27814
rect 5368 27418 5396 30110
rect 5552 28762 5580 30194
rect 5644 30054 5672 30382
rect 5632 30048 5684 30054
rect 5632 29990 5684 29996
rect 5540 28756 5592 28762
rect 5540 28698 5592 28704
rect 5538 28656 5594 28665
rect 5538 28591 5594 28600
rect 5448 28416 5500 28422
rect 5448 28358 5500 28364
rect 5460 28218 5488 28358
rect 5448 28212 5500 28218
rect 5448 28154 5500 28160
rect 5552 27946 5580 28591
rect 5540 27940 5592 27946
rect 5540 27882 5592 27888
rect 5552 27674 5580 27882
rect 5540 27668 5592 27674
rect 5540 27610 5592 27616
rect 5540 27464 5592 27470
rect 5368 27412 5540 27418
rect 5368 27406 5592 27412
rect 5368 27390 5580 27406
rect 5356 27328 5408 27334
rect 5356 27270 5408 27276
rect 5172 26988 5224 26994
rect 5172 26930 5224 26936
rect 5368 26926 5396 27270
rect 5356 26920 5408 26926
rect 5356 26862 5408 26868
rect 5552 26790 5580 27390
rect 5540 26784 5592 26790
rect 5540 26726 5592 26732
rect 5552 25242 5580 26726
rect 5644 25922 5672 29990
rect 5736 28014 5764 31640
rect 5920 29594 5948 32807
rect 5998 30560 6054 30569
rect 5998 30495 6054 30504
rect 6012 29646 6040 30495
rect 5828 29566 5948 29594
rect 6000 29640 6052 29646
rect 6000 29582 6052 29588
rect 5724 28008 5776 28014
rect 5724 27950 5776 27956
rect 5828 27538 5856 29566
rect 5908 29504 5960 29510
rect 5908 29446 5960 29452
rect 5920 29073 5948 29446
rect 6012 29102 6040 29582
rect 6000 29096 6052 29102
rect 5906 29064 5962 29073
rect 6000 29038 6052 29044
rect 5906 28999 5962 29008
rect 6012 28218 6040 29038
rect 6000 28212 6052 28218
rect 6000 28154 6052 28160
rect 6000 28076 6052 28082
rect 6000 28018 6052 28024
rect 6012 27878 6040 28018
rect 6000 27872 6052 27878
rect 6000 27814 6052 27820
rect 5816 27532 5868 27538
rect 5816 27474 5868 27480
rect 5828 26246 5856 27474
rect 6012 27470 6040 27814
rect 6000 27464 6052 27470
rect 6000 27406 6052 27412
rect 6012 27062 6040 27406
rect 6000 27056 6052 27062
rect 6000 26998 6052 27004
rect 5816 26240 5868 26246
rect 5816 26182 5868 26188
rect 5644 25894 5764 25922
rect 5632 25832 5684 25838
rect 5632 25774 5684 25780
rect 5184 25214 5580 25242
rect 5080 23588 5132 23594
rect 5080 23530 5132 23536
rect 5184 21690 5212 25214
rect 5264 25152 5316 25158
rect 5264 25094 5316 25100
rect 5540 25152 5592 25158
rect 5540 25094 5592 25100
rect 5276 24614 5304 25094
rect 5552 24834 5580 25094
rect 5356 24812 5408 24818
rect 5356 24754 5408 24760
rect 5460 24806 5580 24834
rect 5368 24721 5396 24754
rect 5460 24750 5488 24806
rect 5448 24744 5500 24750
rect 5354 24712 5410 24721
rect 5448 24686 5500 24692
rect 5354 24647 5410 24656
rect 5264 24608 5316 24614
rect 5264 24550 5316 24556
rect 5276 23225 5304 24550
rect 5540 24200 5592 24206
rect 5540 24142 5592 24148
rect 5448 23588 5500 23594
rect 5448 23530 5500 23536
rect 5262 23216 5318 23225
rect 5262 23151 5318 23160
rect 5262 23080 5318 23089
rect 5262 23015 5318 23024
rect 4988 21684 5040 21690
rect 4988 21626 5040 21632
rect 5172 21684 5224 21690
rect 5172 21626 5224 21632
rect 5000 21418 5028 21626
rect 5172 21548 5224 21554
rect 5172 21490 5224 21496
rect 4988 21412 5040 21418
rect 4988 21354 5040 21360
rect 5184 21146 5212 21490
rect 5172 21140 5224 21146
rect 5172 21082 5224 21088
rect 5276 19922 5304 23015
rect 5356 21548 5408 21554
rect 5356 21490 5408 21496
rect 5368 21078 5396 21490
rect 5460 21078 5488 23530
rect 5552 23526 5580 24142
rect 5644 23798 5672 25774
rect 5632 23792 5684 23798
rect 5632 23734 5684 23740
rect 5540 23520 5592 23526
rect 5540 23462 5592 23468
rect 5552 23254 5580 23462
rect 5644 23254 5672 23734
rect 5736 23730 5764 25894
rect 6000 25696 6052 25702
rect 6000 25638 6052 25644
rect 5816 23860 5868 23866
rect 5816 23802 5868 23808
rect 5724 23724 5776 23730
rect 5724 23666 5776 23672
rect 5724 23588 5776 23594
rect 5724 23530 5776 23536
rect 5540 23248 5592 23254
rect 5540 23190 5592 23196
rect 5632 23248 5684 23254
rect 5632 23190 5684 23196
rect 5552 22438 5580 23190
rect 5736 23066 5764 23530
rect 5644 23038 5764 23066
rect 5540 22432 5592 22438
rect 5540 22374 5592 22380
rect 5540 21684 5592 21690
rect 5540 21626 5592 21632
rect 5356 21072 5408 21078
rect 5356 21014 5408 21020
rect 5448 21072 5500 21078
rect 5448 21014 5500 21020
rect 5552 20398 5580 21626
rect 5540 20392 5592 20398
rect 5540 20334 5592 20340
rect 4856 19876 4936 19904
rect 5264 19916 5316 19922
rect 4804 19858 4856 19864
rect 5264 19858 5316 19864
rect 5540 19916 5592 19922
rect 5540 19858 5592 19864
rect 4710 19272 4766 19281
rect 4710 19207 4766 19216
rect 4816 19174 4844 19858
rect 5172 19848 5224 19854
rect 5172 19790 5224 19796
rect 5078 19272 5134 19281
rect 5078 19207 5134 19216
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4620 18896 4672 18902
rect 4620 18838 4672 18844
rect 4632 17882 4660 18838
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4724 18426 4752 18702
rect 4712 18420 4764 18426
rect 4712 18362 4764 18368
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 4632 17338 4660 17818
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4528 14612 4580 14618
rect 4528 14554 4580 14560
rect 4540 14074 4568 14554
rect 4528 14068 4580 14074
rect 4528 14010 4580 14016
rect 4632 13394 4660 14758
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4632 12918 4660 13330
rect 4620 12912 4672 12918
rect 4618 12880 4620 12889
rect 4672 12880 4674 12889
rect 4618 12815 4674 12824
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4540 11540 4568 12378
rect 4618 12336 4674 12345
rect 4618 12271 4620 12280
rect 4672 12271 4674 12280
rect 4620 12242 4672 12248
rect 4632 11898 4660 12242
rect 4724 12238 4752 14214
rect 4816 13734 4844 19110
rect 5092 17898 5120 19207
rect 5184 18086 5212 19790
rect 5276 19242 5304 19858
rect 5264 19236 5316 19242
rect 5264 19178 5316 19184
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 5092 17870 5212 17898
rect 5080 17740 5132 17746
rect 5080 17682 5132 17688
rect 4988 17672 5040 17678
rect 4988 17614 5040 17620
rect 5000 17542 5028 17614
rect 4988 17536 5040 17542
rect 4988 17478 5040 17484
rect 5000 17066 5028 17478
rect 4988 17060 5040 17066
rect 4988 17002 5040 17008
rect 5092 16998 5120 17682
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 5092 16794 5120 16934
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 5092 16114 5120 16730
rect 5080 16108 5132 16114
rect 5080 16050 5132 16056
rect 5080 15904 5132 15910
rect 5080 15846 5132 15852
rect 5092 15366 5120 15846
rect 5080 15360 5132 15366
rect 5080 15302 5132 15308
rect 4896 14476 4948 14482
rect 4896 14418 4948 14424
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4908 13530 4936 14418
rect 4896 13524 4948 13530
rect 4896 13466 4948 13472
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4816 12442 4844 12718
rect 4804 12436 4856 12442
rect 4804 12378 4856 12384
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4908 11558 4936 12174
rect 4620 11552 4672 11558
rect 4540 11512 4620 11540
rect 4620 11494 4672 11500
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4526 10704 4582 10713
rect 4526 10639 4582 10648
rect 4540 10538 4568 10639
rect 4528 10532 4580 10538
rect 4528 10474 4580 10480
rect 4632 9994 4660 11494
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 4908 9382 4936 11494
rect 5092 10713 5120 15302
rect 5184 13802 5212 17870
rect 5276 13870 5304 19178
rect 5356 19168 5408 19174
rect 5356 19110 5408 19116
rect 5368 18970 5396 19110
rect 5356 18964 5408 18970
rect 5356 18906 5408 18912
rect 5552 18902 5580 19858
rect 5644 18902 5672 23038
rect 5724 22432 5776 22438
rect 5724 22374 5776 22380
rect 5736 21894 5764 22374
rect 5724 21888 5776 21894
rect 5724 21830 5776 21836
rect 5736 21554 5764 21830
rect 5724 21548 5776 21554
rect 5724 21490 5776 21496
rect 5724 21412 5776 21418
rect 5724 21354 5776 21360
rect 5540 18896 5592 18902
rect 5540 18838 5592 18844
rect 5632 18896 5684 18902
rect 5736 18873 5764 21354
rect 5632 18838 5684 18844
rect 5722 18864 5778 18873
rect 5644 18426 5672 18838
rect 5722 18799 5778 18808
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5552 17882 5580 18022
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5644 17354 5672 18362
rect 5552 17326 5672 17354
rect 5552 16776 5580 17326
rect 5828 17270 5856 23802
rect 6012 22234 6040 25638
rect 6104 24274 6132 33646
rect 6552 33594 6604 33600
rect 6564 33454 6592 33594
rect 6552 33448 6604 33454
rect 6552 33390 6604 33396
rect 6289 33212 6585 33232
rect 6345 33210 6369 33212
rect 6425 33210 6449 33212
rect 6505 33210 6529 33212
rect 6367 33158 6369 33210
rect 6431 33158 6443 33210
rect 6505 33158 6507 33210
rect 6345 33156 6369 33158
rect 6425 33156 6449 33158
rect 6505 33156 6529 33158
rect 6289 33136 6585 33156
rect 6184 32972 6236 32978
rect 6184 32914 6236 32920
rect 6196 32570 6224 32914
rect 6644 32836 6696 32842
rect 6644 32778 6696 32784
rect 6656 32570 6684 32778
rect 6184 32564 6236 32570
rect 6184 32506 6236 32512
rect 6644 32564 6696 32570
rect 6644 32506 6696 32512
rect 6289 32124 6585 32144
rect 6345 32122 6369 32124
rect 6425 32122 6449 32124
rect 6505 32122 6529 32124
rect 6367 32070 6369 32122
rect 6431 32070 6443 32122
rect 6505 32070 6507 32122
rect 6345 32068 6369 32070
rect 6425 32068 6449 32070
rect 6505 32068 6529 32070
rect 6289 32048 6585 32068
rect 6184 32020 6236 32026
rect 6184 31962 6236 31968
rect 6196 31890 6224 31962
rect 6656 31958 6684 32506
rect 6644 31952 6696 31958
rect 6644 31894 6696 31900
rect 6184 31884 6236 31890
rect 6184 31826 6236 31832
rect 6196 31142 6224 31826
rect 6184 31136 6236 31142
rect 6184 31078 6236 31084
rect 6196 28422 6224 31078
rect 6289 31036 6585 31056
rect 6345 31034 6369 31036
rect 6425 31034 6449 31036
rect 6505 31034 6529 31036
rect 6367 30982 6369 31034
rect 6431 30982 6443 31034
rect 6505 30982 6507 31034
rect 6345 30980 6369 30982
rect 6425 30980 6449 30982
rect 6505 30980 6529 30982
rect 6289 30960 6585 30980
rect 6642 30288 6698 30297
rect 6642 30223 6698 30232
rect 6289 29948 6585 29968
rect 6345 29946 6369 29948
rect 6425 29946 6449 29948
rect 6505 29946 6529 29948
rect 6367 29894 6369 29946
rect 6431 29894 6443 29946
rect 6505 29894 6507 29946
rect 6345 29892 6369 29894
rect 6425 29892 6449 29894
rect 6505 29892 6529 29894
rect 6289 29872 6585 29892
rect 6656 29850 6684 30223
rect 6644 29844 6696 29850
rect 6644 29786 6696 29792
rect 6460 29640 6512 29646
rect 6460 29582 6512 29588
rect 6472 29034 6500 29582
rect 6656 29306 6684 29786
rect 6644 29300 6696 29306
rect 6644 29242 6696 29248
rect 6460 29028 6512 29034
rect 6460 28970 6512 28976
rect 6289 28860 6585 28880
rect 6345 28858 6369 28860
rect 6425 28858 6449 28860
rect 6505 28858 6529 28860
rect 6367 28806 6369 28858
rect 6431 28806 6443 28858
rect 6505 28806 6507 28858
rect 6345 28804 6369 28806
rect 6425 28804 6449 28806
rect 6505 28804 6529 28806
rect 6289 28784 6585 28804
rect 6184 28416 6236 28422
rect 6184 28358 6236 28364
rect 6184 28212 6236 28218
rect 6184 28154 6236 28160
rect 6196 25702 6224 28154
rect 6289 27772 6585 27792
rect 6345 27770 6369 27772
rect 6425 27770 6449 27772
rect 6505 27770 6529 27772
rect 6367 27718 6369 27770
rect 6431 27718 6443 27770
rect 6505 27718 6507 27770
rect 6345 27716 6369 27718
rect 6425 27716 6449 27718
rect 6505 27716 6529 27718
rect 6289 27696 6585 27716
rect 6656 27656 6684 29242
rect 6748 28529 6776 35430
rect 7392 35290 7420 39520
rect 7760 35834 7788 39520
rect 7932 36576 7984 36582
rect 7932 36518 7984 36524
rect 7748 35828 7800 35834
rect 7748 35770 7800 35776
rect 7656 35488 7708 35494
rect 7656 35430 7708 35436
rect 7840 35488 7892 35494
rect 7840 35430 7892 35436
rect 7380 35284 7432 35290
rect 7380 35226 7432 35232
rect 6920 35148 6972 35154
rect 6920 35090 6972 35096
rect 7380 35148 7432 35154
rect 7380 35090 7432 35096
rect 6932 34746 6960 35090
rect 7012 35080 7064 35086
rect 7012 35022 7064 35028
rect 6920 34740 6972 34746
rect 6920 34682 6972 34688
rect 7024 34542 7052 35022
rect 7392 34542 7420 35090
rect 7012 34536 7064 34542
rect 7012 34478 7064 34484
rect 7380 34536 7432 34542
rect 7380 34478 7432 34484
rect 7024 34105 7052 34478
rect 7010 34096 7066 34105
rect 7010 34031 7066 34040
rect 7194 34096 7250 34105
rect 7194 34031 7250 34040
rect 7104 33856 7156 33862
rect 7104 33798 7156 33804
rect 7116 33590 7144 33798
rect 7104 33584 7156 33590
rect 7104 33526 7156 33532
rect 6828 33312 6880 33318
rect 6828 33254 6880 33260
rect 6840 33114 6868 33254
rect 6828 33108 6880 33114
rect 6828 33050 6880 33056
rect 7116 32842 7144 33526
rect 7208 33454 7236 34031
rect 7288 33924 7340 33930
rect 7288 33866 7340 33872
rect 7300 33522 7328 33866
rect 7288 33516 7340 33522
rect 7288 33458 7340 33464
rect 7196 33448 7248 33454
rect 7196 33390 7248 33396
rect 7288 33312 7340 33318
rect 7392 33289 7420 34478
rect 7564 34128 7616 34134
rect 7564 34070 7616 34076
rect 7576 33318 7604 34070
rect 7564 33312 7616 33318
rect 7288 33254 7340 33260
rect 7378 33280 7434 33289
rect 7104 32836 7156 32842
rect 7104 32778 7156 32784
rect 7300 32434 7328 33254
rect 7564 33254 7616 33260
rect 7378 33215 7434 33224
rect 7288 32428 7340 32434
rect 7288 32370 7340 32376
rect 7300 32026 7328 32370
rect 7288 32020 7340 32026
rect 7288 31962 7340 31968
rect 6920 31952 6972 31958
rect 6920 31894 6972 31900
rect 6932 31634 6960 31894
rect 7012 31680 7064 31686
rect 6932 31628 7012 31634
rect 6932 31622 7064 31628
rect 6932 31606 7052 31622
rect 6932 31414 6960 31606
rect 6920 31408 6972 31414
rect 6920 31350 6972 31356
rect 7104 31136 7156 31142
rect 7104 31078 7156 31084
rect 6826 30152 6882 30161
rect 6826 30087 6882 30096
rect 6840 30054 6868 30087
rect 6828 30048 6880 30054
rect 6828 29990 6880 29996
rect 6734 28520 6790 28529
rect 6734 28455 6790 28464
rect 6828 28416 6880 28422
rect 6828 28358 6880 28364
rect 6840 28014 6868 28358
rect 6828 28008 6880 28014
rect 6828 27950 6880 27956
rect 6656 27628 6776 27656
rect 6644 27532 6696 27538
rect 6644 27474 6696 27480
rect 6656 27130 6684 27474
rect 6644 27124 6696 27130
rect 6644 27066 6696 27072
rect 6642 27024 6698 27033
rect 6642 26959 6698 26968
rect 6289 26684 6585 26704
rect 6345 26682 6369 26684
rect 6425 26682 6449 26684
rect 6505 26682 6529 26684
rect 6367 26630 6369 26682
rect 6431 26630 6443 26682
rect 6505 26630 6507 26682
rect 6345 26628 6369 26630
rect 6425 26628 6449 26630
rect 6505 26628 6529 26630
rect 6289 26608 6585 26628
rect 6184 25696 6236 25702
rect 6184 25638 6236 25644
rect 6289 25596 6585 25616
rect 6345 25594 6369 25596
rect 6425 25594 6449 25596
rect 6505 25594 6529 25596
rect 6367 25542 6369 25594
rect 6431 25542 6443 25594
rect 6505 25542 6507 25594
rect 6345 25540 6369 25542
rect 6425 25540 6449 25542
rect 6505 25540 6529 25542
rect 6289 25520 6585 25540
rect 6184 25424 6236 25430
rect 6184 25366 6236 25372
rect 6196 24954 6224 25366
rect 6276 25288 6328 25294
rect 6276 25230 6328 25236
rect 6184 24948 6236 24954
rect 6184 24890 6236 24896
rect 6196 24410 6224 24890
rect 6288 24886 6316 25230
rect 6276 24880 6328 24886
rect 6276 24822 6328 24828
rect 6289 24508 6585 24528
rect 6345 24506 6369 24508
rect 6425 24506 6449 24508
rect 6505 24506 6529 24508
rect 6367 24454 6369 24506
rect 6431 24454 6443 24506
rect 6505 24454 6507 24506
rect 6345 24452 6369 24454
rect 6425 24452 6449 24454
rect 6505 24452 6529 24454
rect 6289 24432 6585 24452
rect 6184 24404 6236 24410
rect 6184 24346 6236 24352
rect 6276 24336 6328 24342
rect 6276 24278 6328 24284
rect 6092 24268 6144 24274
rect 6092 24210 6144 24216
rect 6104 23866 6132 24210
rect 6288 23866 6316 24278
rect 6656 23882 6684 26959
rect 6748 25480 6776 27628
rect 6840 27470 6868 27950
rect 7012 27940 7064 27946
rect 7012 27882 7064 27888
rect 6828 27464 6880 27470
rect 6828 27406 6880 27412
rect 6840 26042 6868 27406
rect 7024 27130 7052 27882
rect 7012 27124 7064 27130
rect 7012 27066 7064 27072
rect 7012 26240 7064 26246
rect 7012 26182 7064 26188
rect 6828 26036 6880 26042
rect 6828 25978 6880 25984
rect 6748 25452 6960 25480
rect 6828 25356 6880 25362
rect 6828 25298 6880 25304
rect 6736 24880 6788 24886
rect 6736 24822 6788 24828
rect 6748 24410 6776 24822
rect 6840 24614 6868 25298
rect 6828 24608 6880 24614
rect 6828 24550 6880 24556
rect 6736 24404 6788 24410
rect 6736 24346 6788 24352
rect 6092 23860 6144 23866
rect 6276 23860 6328 23866
rect 6092 23802 6144 23808
rect 6196 23820 6276 23848
rect 6092 23724 6144 23730
rect 6092 23666 6144 23672
rect 6000 22228 6052 22234
rect 6000 22170 6052 22176
rect 5908 22092 5960 22098
rect 5908 22034 5960 22040
rect 5920 20602 5948 22034
rect 5908 20596 5960 20602
rect 5908 20538 5960 20544
rect 6104 20398 6132 23666
rect 5908 20392 5960 20398
rect 5908 20334 5960 20340
rect 6092 20392 6144 20398
rect 6092 20334 6144 20340
rect 5632 17264 5684 17270
rect 5632 17206 5684 17212
rect 5816 17264 5868 17270
rect 5816 17206 5868 17212
rect 5368 16748 5580 16776
rect 5368 14618 5396 16748
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5460 15434 5488 16594
rect 5538 15872 5594 15881
rect 5538 15807 5594 15816
rect 5552 15706 5580 15807
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5448 15428 5500 15434
rect 5448 15370 5500 15376
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5552 14958 5580 15302
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5356 14612 5408 14618
rect 5356 14554 5408 14560
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5172 13796 5224 13802
rect 5172 13738 5224 13744
rect 5262 13288 5318 13297
rect 5262 13223 5318 13232
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 5184 12102 5212 13126
rect 5276 12986 5304 13223
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 5078 10704 5134 10713
rect 5078 10639 5134 10648
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 5276 9110 5304 9998
rect 5264 9104 5316 9110
rect 5264 9046 5316 9052
rect 5276 8634 5304 9046
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 4528 8016 4580 8022
rect 4528 7958 4580 7964
rect 4540 7546 4568 7958
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4436 6180 4488 6186
rect 4436 6122 4488 6128
rect 4344 6112 4396 6118
rect 4342 6080 4344 6089
rect 4396 6080 4398 6089
rect 4342 6015 4398 6024
rect 4356 5914 4384 6015
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4264 4826 4292 5850
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4356 5234 4384 5714
rect 4434 5672 4490 5681
rect 4434 5607 4490 5616
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 4356 4690 4384 5170
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4344 3460 4396 3466
rect 4344 3402 4396 3408
rect 4356 2922 4384 3402
rect 4344 2916 4396 2922
rect 4344 2858 4396 2864
rect 4356 2582 4384 2858
rect 4344 2576 4396 2582
rect 4344 2518 4396 2524
rect 4448 2122 4476 5607
rect 4632 5370 4660 7822
rect 4988 7472 5040 7478
rect 4986 7440 4988 7449
rect 5040 7440 5042 7449
rect 5184 7410 5212 8230
rect 4986 7375 5042 7384
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5368 6866 5396 14554
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5552 13938 5580 14350
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5448 13864 5500 13870
rect 5446 13832 5448 13841
rect 5500 13832 5502 13841
rect 5446 13767 5502 13776
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5448 13728 5500 13734
rect 5448 13670 5500 13676
rect 5460 12889 5488 13670
rect 5446 12880 5502 12889
rect 5446 12815 5502 12824
rect 5552 12782 5580 13738
rect 5540 12776 5592 12782
rect 5540 12718 5592 12724
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5552 12442 5580 12582
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5644 12238 5672 17206
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 5736 16658 5764 16934
rect 5920 16833 5948 20334
rect 6090 20224 6146 20233
rect 6090 20159 6146 20168
rect 6104 20058 6132 20159
rect 6092 20052 6144 20058
rect 6092 19994 6144 20000
rect 6092 19780 6144 19786
rect 6092 19722 6144 19728
rect 6104 19174 6132 19722
rect 6092 19168 6144 19174
rect 6092 19110 6144 19116
rect 6000 18964 6052 18970
rect 6000 18906 6052 18912
rect 6012 18426 6040 18906
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 6104 18086 6132 19110
rect 6092 18080 6144 18086
rect 6092 18022 6144 18028
rect 5906 16824 5962 16833
rect 5906 16759 5962 16768
rect 6104 16726 6132 18022
rect 6092 16720 6144 16726
rect 6092 16662 6144 16668
rect 5724 16652 5776 16658
rect 5724 16594 5776 16600
rect 5908 16652 5960 16658
rect 5908 16594 5960 16600
rect 5736 15366 5764 16594
rect 5920 16250 5948 16594
rect 5908 16244 5960 16250
rect 5908 16186 5960 16192
rect 5816 15428 5868 15434
rect 5816 15370 5868 15376
rect 5724 15360 5776 15366
rect 5724 15302 5776 15308
rect 5828 14278 5856 15370
rect 6196 14600 6224 23820
rect 6276 23802 6328 23808
rect 6564 23854 6684 23882
rect 6564 23594 6592 23854
rect 6748 23798 6776 24346
rect 6736 23792 6788 23798
rect 6656 23740 6736 23746
rect 6656 23734 6788 23740
rect 6656 23718 6776 23734
rect 6552 23588 6604 23594
rect 6552 23530 6604 23536
rect 6289 23420 6585 23440
rect 6345 23418 6369 23420
rect 6425 23418 6449 23420
rect 6505 23418 6529 23420
rect 6367 23366 6369 23418
rect 6431 23366 6443 23418
rect 6505 23366 6507 23418
rect 6345 23364 6369 23366
rect 6425 23364 6449 23366
rect 6505 23364 6529 23366
rect 6289 23344 6585 23364
rect 6656 23322 6684 23718
rect 6644 23316 6696 23322
rect 6644 23258 6696 23264
rect 6656 23118 6684 23258
rect 6644 23112 6696 23118
rect 6644 23054 6696 23060
rect 6840 22778 6868 24550
rect 6932 24342 6960 25452
rect 6920 24336 6972 24342
rect 6920 24278 6972 24284
rect 6918 23624 6974 23633
rect 6918 23559 6974 23568
rect 6932 23322 6960 23559
rect 6920 23316 6972 23322
rect 6920 23258 6972 23264
rect 6828 22772 6880 22778
rect 6828 22714 6880 22720
rect 6932 22574 6960 23258
rect 7024 23236 7052 26182
rect 7116 23361 7144 31078
rect 7288 30592 7340 30598
rect 7288 30534 7340 30540
rect 7194 30424 7250 30433
rect 7194 30359 7250 30368
rect 7208 30190 7236 30359
rect 7300 30258 7328 30534
rect 7288 30252 7340 30258
rect 7288 30194 7340 30200
rect 7196 30184 7248 30190
rect 7196 30126 7248 30132
rect 7208 29850 7236 30126
rect 7196 29844 7248 29850
rect 7196 29786 7248 29792
rect 7194 27568 7250 27577
rect 7194 27503 7250 27512
rect 7208 27130 7236 27503
rect 7196 27124 7248 27130
rect 7196 27066 7248 27072
rect 7288 26852 7340 26858
rect 7288 26794 7340 26800
rect 7300 26246 7328 26794
rect 7288 26240 7340 26246
rect 7288 26182 7340 26188
rect 7300 25498 7328 26182
rect 7288 25492 7340 25498
rect 7288 25434 7340 25440
rect 7196 24064 7248 24070
rect 7196 24006 7248 24012
rect 7208 23594 7236 24006
rect 7196 23588 7248 23594
rect 7196 23530 7248 23536
rect 7102 23352 7158 23361
rect 7102 23287 7158 23296
rect 7024 23208 7144 23236
rect 6920 22568 6972 22574
rect 6920 22510 6972 22516
rect 6644 22500 6696 22506
rect 6644 22442 6696 22448
rect 6289 22332 6585 22352
rect 6345 22330 6369 22332
rect 6425 22330 6449 22332
rect 6505 22330 6529 22332
rect 6367 22278 6369 22330
rect 6431 22278 6443 22330
rect 6505 22278 6507 22330
rect 6345 22276 6369 22278
rect 6425 22276 6449 22278
rect 6505 22276 6529 22278
rect 6289 22256 6585 22276
rect 6276 22160 6328 22166
rect 6276 22102 6328 22108
rect 6288 21690 6316 22102
rect 6276 21684 6328 21690
rect 6276 21626 6328 21632
rect 6289 21244 6585 21264
rect 6345 21242 6369 21244
rect 6425 21242 6449 21244
rect 6505 21242 6529 21244
rect 6367 21190 6369 21242
rect 6431 21190 6443 21242
rect 6505 21190 6507 21242
rect 6345 21188 6369 21190
rect 6425 21188 6449 21190
rect 6505 21188 6529 21190
rect 6289 21168 6585 21188
rect 6289 20156 6585 20176
rect 6345 20154 6369 20156
rect 6425 20154 6449 20156
rect 6505 20154 6529 20156
rect 6367 20102 6369 20154
rect 6431 20102 6443 20154
rect 6505 20102 6507 20154
rect 6345 20100 6369 20102
rect 6425 20100 6449 20102
rect 6505 20100 6529 20102
rect 6289 20080 6585 20100
rect 6460 19916 6512 19922
rect 6460 19858 6512 19864
rect 6472 19825 6500 19858
rect 6458 19816 6514 19825
rect 6458 19751 6514 19760
rect 6289 19068 6585 19088
rect 6345 19066 6369 19068
rect 6425 19066 6449 19068
rect 6505 19066 6529 19068
rect 6367 19014 6369 19066
rect 6431 19014 6443 19066
rect 6505 19014 6507 19066
rect 6345 19012 6369 19014
rect 6425 19012 6449 19014
rect 6505 19012 6529 19014
rect 6289 18992 6585 19012
rect 6289 17980 6585 18000
rect 6345 17978 6369 17980
rect 6425 17978 6449 17980
rect 6505 17978 6529 17980
rect 6367 17926 6369 17978
rect 6431 17926 6443 17978
rect 6505 17926 6507 17978
rect 6345 17924 6369 17926
rect 6425 17924 6449 17926
rect 6505 17924 6529 17926
rect 6289 17904 6585 17924
rect 6289 16892 6585 16912
rect 6345 16890 6369 16892
rect 6425 16890 6449 16892
rect 6505 16890 6529 16892
rect 6367 16838 6369 16890
rect 6431 16838 6443 16890
rect 6505 16838 6507 16890
rect 6345 16836 6369 16838
rect 6425 16836 6449 16838
rect 6505 16836 6529 16838
rect 6289 16816 6585 16836
rect 6289 15804 6585 15824
rect 6345 15802 6369 15804
rect 6425 15802 6449 15804
rect 6505 15802 6529 15804
rect 6367 15750 6369 15802
rect 6431 15750 6443 15802
rect 6505 15750 6507 15802
rect 6345 15748 6369 15750
rect 6425 15748 6449 15750
rect 6505 15748 6529 15750
rect 6289 15728 6585 15748
rect 6289 14716 6585 14736
rect 6345 14714 6369 14716
rect 6425 14714 6449 14716
rect 6505 14714 6529 14716
rect 6367 14662 6369 14714
rect 6431 14662 6443 14714
rect 6505 14662 6507 14714
rect 6345 14660 6369 14662
rect 6425 14660 6449 14662
rect 6505 14660 6529 14662
rect 6289 14640 6585 14660
rect 6012 14572 6224 14600
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5540 12096 5592 12102
rect 5460 12056 5540 12084
rect 5460 9110 5488 12056
rect 5540 12038 5592 12044
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 5446 8528 5502 8537
rect 5446 8463 5502 8472
rect 5460 7546 5488 8463
rect 5552 8430 5580 9862
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5644 7834 5672 11698
rect 5736 8498 5764 12582
rect 5828 12306 5856 14214
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 5920 12850 5948 13126
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 6012 12458 6040 14572
rect 6090 13832 6146 13841
rect 6090 13767 6146 13776
rect 6104 13274 6132 13767
rect 6289 13628 6585 13648
rect 6345 13626 6369 13628
rect 6425 13626 6449 13628
rect 6505 13626 6529 13628
rect 6367 13574 6369 13626
rect 6431 13574 6443 13626
rect 6505 13574 6507 13626
rect 6345 13572 6369 13574
rect 6425 13572 6449 13574
rect 6505 13572 6529 13574
rect 6289 13552 6585 13572
rect 6104 13246 6224 13274
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 5920 12430 6040 12458
rect 5920 12374 5948 12430
rect 5908 12368 5960 12374
rect 5908 12310 5960 12316
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 5828 11898 5856 12242
rect 6000 12232 6052 12238
rect 5906 12200 5962 12209
rect 6000 12174 6052 12180
rect 5906 12135 5962 12144
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5828 10266 5856 10746
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5828 9722 5856 10202
rect 5920 10198 5948 12135
rect 5908 10192 5960 10198
rect 5908 10134 5960 10140
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5552 7806 5672 7834
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 4816 5574 4844 6598
rect 5172 6180 5224 6186
rect 5172 6122 5224 6128
rect 4804 5568 4856 5574
rect 4802 5536 4804 5545
rect 4988 5568 5040 5574
rect 4856 5536 4858 5545
rect 4802 5471 4858 5480
rect 4908 5528 4988 5556
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4632 5166 4660 5306
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4540 3194 4568 3538
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4816 2990 4844 5471
rect 4908 5302 4936 5528
rect 4988 5510 5040 5516
rect 5184 5302 5212 6122
rect 5264 5840 5316 5846
rect 5264 5782 5316 5788
rect 4896 5296 4948 5302
rect 4896 5238 4948 5244
rect 5172 5296 5224 5302
rect 5172 5238 5224 5244
rect 4908 4622 4936 5238
rect 5080 5024 5132 5030
rect 5080 4966 5132 4972
rect 5092 4826 5120 4966
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4908 4282 4936 4558
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 5078 4176 5134 4185
rect 4988 4140 5040 4146
rect 5078 4111 5134 4120
rect 5172 4140 5224 4146
rect 4988 4082 5040 4088
rect 5000 3942 5028 4082
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 5000 3738 5028 3878
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 5000 3534 5028 3674
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 4540 2281 4568 2382
rect 4526 2272 4582 2281
rect 4526 2207 4582 2216
rect 5092 2122 5120 4111
rect 5172 4082 5224 4088
rect 5184 3670 5212 4082
rect 5276 3670 5304 5782
rect 5172 3664 5224 3670
rect 5172 3606 5224 3612
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 4448 2094 4568 2122
rect 4540 480 4568 2094
rect 5000 2094 5120 2122
rect 5000 480 5028 2094
rect 5368 480 5396 6598
rect 5448 6452 5500 6458
rect 5552 6440 5580 7806
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5644 7342 5672 7686
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5644 7002 5672 7278
rect 5736 7002 5764 8026
rect 5632 6996 5684 7002
rect 5632 6938 5684 6944
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5644 6769 5672 6802
rect 5630 6760 5686 6769
rect 5630 6695 5686 6704
rect 5644 6458 5672 6695
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5500 6412 5580 6440
rect 5448 6394 5500 6400
rect 5552 5370 5580 6412
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5446 5264 5502 5273
rect 5446 5199 5502 5208
rect 5632 5228 5684 5234
rect 5460 5030 5488 5199
rect 5632 5170 5684 5176
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5540 4752 5592 4758
rect 5540 4694 5592 4700
rect 5448 4684 5500 4690
rect 5448 4626 5500 4632
rect 5460 3194 5488 4626
rect 5552 3738 5580 4694
rect 5644 4690 5672 5170
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5644 2825 5672 3878
rect 5630 2816 5686 2825
rect 5630 2751 5686 2760
rect 5630 2544 5686 2553
rect 5630 2479 5632 2488
rect 5684 2479 5686 2488
rect 5632 2450 5684 2456
rect 5736 480 5764 6598
rect 5828 6338 5856 9658
rect 5920 9382 5948 10134
rect 6012 9654 6040 12174
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 5920 7449 5948 9318
rect 5906 7440 5962 7449
rect 5906 7375 5962 7384
rect 6012 6866 6040 9318
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 5828 6310 6040 6338
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5828 5681 5856 6054
rect 5814 5672 5870 5681
rect 5814 5607 5870 5616
rect 5920 3670 5948 6190
rect 6012 6100 6040 6310
rect 6104 6254 6132 13126
rect 6196 11762 6224 13246
rect 6289 12540 6585 12560
rect 6345 12538 6369 12540
rect 6425 12538 6449 12540
rect 6505 12538 6529 12540
rect 6367 12486 6369 12538
rect 6431 12486 6443 12538
rect 6505 12486 6507 12538
rect 6345 12484 6369 12486
rect 6425 12484 6449 12486
rect 6505 12484 6529 12486
rect 6289 12464 6585 12484
rect 6276 12368 6328 12374
rect 6276 12310 6328 12316
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 6288 11642 6316 12310
rect 6196 11614 6316 11642
rect 6196 9489 6224 11614
rect 6289 11452 6585 11472
rect 6345 11450 6369 11452
rect 6425 11450 6449 11452
rect 6505 11450 6529 11452
rect 6367 11398 6369 11450
rect 6431 11398 6443 11450
rect 6505 11398 6507 11450
rect 6345 11396 6369 11398
rect 6425 11396 6449 11398
rect 6505 11396 6529 11398
rect 6289 11376 6585 11396
rect 6289 10364 6585 10384
rect 6345 10362 6369 10364
rect 6425 10362 6449 10364
rect 6505 10362 6529 10364
rect 6367 10310 6369 10362
rect 6431 10310 6443 10362
rect 6505 10310 6507 10362
rect 6345 10308 6369 10310
rect 6425 10308 6449 10310
rect 6505 10308 6529 10310
rect 6289 10288 6585 10308
rect 6656 9518 6684 22442
rect 6920 22432 6972 22438
rect 6920 22374 6972 22380
rect 6932 22030 6960 22374
rect 7116 22166 7144 23208
rect 7286 22672 7342 22681
rect 7286 22607 7342 22616
rect 7300 22574 7328 22607
rect 7288 22568 7340 22574
rect 7288 22510 7340 22516
rect 7104 22160 7156 22166
rect 7392 22114 7420 33215
rect 7576 33114 7604 33254
rect 7564 33108 7616 33114
rect 7564 33050 7616 33056
rect 7562 32328 7618 32337
rect 7562 32263 7618 32272
rect 7472 32224 7524 32230
rect 7472 32166 7524 32172
rect 7484 30870 7512 32166
rect 7472 30864 7524 30870
rect 7472 30806 7524 30812
rect 7576 28642 7604 32263
rect 7668 31210 7696 35430
rect 7748 34944 7800 34950
rect 7748 34886 7800 34892
rect 7760 34542 7788 34886
rect 7748 34536 7800 34542
rect 7748 34478 7800 34484
rect 7852 34474 7880 35430
rect 7840 34468 7892 34474
rect 7840 34410 7892 34416
rect 7748 34400 7800 34406
rect 7800 34348 7880 34354
rect 7748 34342 7880 34348
rect 7760 34326 7880 34342
rect 7748 32972 7800 32978
rect 7748 32914 7800 32920
rect 7760 32473 7788 32914
rect 7746 32464 7802 32473
rect 7746 32399 7802 32408
rect 7760 32298 7788 32399
rect 7748 32292 7800 32298
rect 7748 32234 7800 32240
rect 7852 32178 7880 34326
rect 7760 32150 7880 32178
rect 7656 31204 7708 31210
rect 7656 31146 7708 31152
rect 7656 28960 7708 28966
rect 7656 28902 7708 28908
rect 7668 28762 7696 28902
rect 7760 28801 7788 32150
rect 7944 31804 7972 36518
rect 8116 34468 8168 34474
rect 8116 34410 8168 34416
rect 8128 34066 8156 34410
rect 8220 34406 8248 39520
rect 8482 35048 8538 35057
rect 8482 34983 8538 34992
rect 8300 34740 8352 34746
rect 8300 34682 8352 34688
rect 8208 34400 8260 34406
rect 8208 34342 8260 34348
rect 8116 34060 8168 34066
rect 8116 34002 8168 34008
rect 8128 33318 8156 34002
rect 8116 33312 8168 33318
rect 8116 33254 8168 33260
rect 8206 33008 8262 33017
rect 8116 32972 8168 32978
rect 8206 32943 8208 32952
rect 8116 32914 8168 32920
rect 8260 32943 8262 32952
rect 8208 32914 8260 32920
rect 8128 32570 8156 32914
rect 8116 32564 8168 32570
rect 8116 32506 8168 32512
rect 8220 32502 8248 32914
rect 8312 32502 8340 34682
rect 8208 32496 8260 32502
rect 8208 32438 8260 32444
rect 8300 32496 8352 32502
rect 8300 32438 8352 32444
rect 7935 31776 7972 31804
rect 7935 31668 7963 31776
rect 8024 31680 8076 31686
rect 7935 31640 7972 31668
rect 7746 28792 7802 28801
rect 7656 28756 7708 28762
rect 7746 28727 7802 28736
rect 7656 28698 7708 28704
rect 7576 28614 7788 28642
rect 7564 26920 7616 26926
rect 7564 26862 7616 26868
rect 7576 26586 7604 26862
rect 7564 26580 7616 26586
rect 7564 26522 7616 26528
rect 7564 25356 7616 25362
rect 7564 25298 7616 25304
rect 7576 24954 7604 25298
rect 7656 25152 7708 25158
rect 7656 25094 7708 25100
rect 7564 24948 7616 24954
rect 7564 24890 7616 24896
rect 7470 24712 7526 24721
rect 7470 24647 7526 24656
rect 7484 24342 7512 24647
rect 7576 24410 7604 24890
rect 7668 24886 7696 25094
rect 7656 24880 7708 24886
rect 7656 24822 7708 24828
rect 7564 24404 7616 24410
rect 7564 24346 7616 24352
rect 7472 24336 7524 24342
rect 7472 24278 7524 24284
rect 7484 23866 7512 24278
rect 7472 23860 7524 23866
rect 7472 23802 7524 23808
rect 7564 23520 7616 23526
rect 7564 23462 7616 23468
rect 7472 23316 7524 23322
rect 7472 23258 7524 23264
rect 7484 23225 7512 23258
rect 7470 23216 7526 23225
rect 7470 23151 7526 23160
rect 7472 22976 7524 22982
rect 7576 22964 7604 23462
rect 7524 22936 7604 22964
rect 7472 22918 7524 22924
rect 7104 22102 7156 22108
rect 6920 22024 6972 22030
rect 6920 21966 6972 21972
rect 6736 21480 6788 21486
rect 6736 21422 6788 21428
rect 6748 21146 6776 21422
rect 7116 21418 7144 22102
rect 7300 22086 7420 22114
rect 7484 22556 7512 22918
rect 7564 22568 7616 22574
rect 7484 22528 7564 22556
rect 7300 22080 7328 22086
rect 7208 22052 7328 22080
rect 7104 21412 7156 21418
rect 7104 21354 7156 21360
rect 6736 21140 6788 21146
rect 6736 21082 6788 21088
rect 6748 19009 6776 21082
rect 7104 21004 7156 21010
rect 7104 20946 7156 20952
rect 6920 20936 6972 20942
rect 6920 20878 6972 20884
rect 6932 20618 6960 20878
rect 6840 20602 6960 20618
rect 6828 20596 6960 20602
rect 6880 20590 6960 20596
rect 6828 20538 6880 20544
rect 6828 20392 6880 20398
rect 6828 20334 6880 20340
rect 6840 19174 6868 20334
rect 7010 19816 7066 19825
rect 7010 19751 7012 19760
rect 7064 19751 7066 19760
rect 7012 19722 7064 19728
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6734 19000 6790 19009
rect 6734 18935 6790 18944
rect 6828 18760 6880 18766
rect 7116 18737 7144 20946
rect 7208 19310 7236 22052
rect 7484 21690 7512 22528
rect 7564 22510 7616 22516
rect 7564 22228 7616 22234
rect 7564 22170 7616 22176
rect 7576 21962 7604 22170
rect 7564 21956 7616 21962
rect 7564 21898 7616 21904
rect 7472 21684 7524 21690
rect 7472 21626 7524 21632
rect 7564 21412 7616 21418
rect 7564 21354 7616 21360
rect 7472 21344 7524 21350
rect 7472 21286 7524 21292
rect 7484 21010 7512 21286
rect 7472 21004 7524 21010
rect 7472 20946 7524 20952
rect 7380 20800 7432 20806
rect 7380 20742 7432 20748
rect 7288 20256 7340 20262
rect 7288 20198 7340 20204
rect 7300 19922 7328 20198
rect 7392 20058 7420 20742
rect 7380 20052 7432 20058
rect 7380 19994 7432 20000
rect 7576 19961 7604 21354
rect 7654 21040 7710 21049
rect 7654 20975 7710 20984
rect 7668 20942 7696 20975
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 7562 19952 7618 19961
rect 7288 19916 7340 19922
rect 7562 19887 7618 19896
rect 7288 19858 7340 19864
rect 7300 19825 7328 19858
rect 7472 19848 7524 19854
rect 7286 19816 7342 19825
rect 7472 19790 7524 19796
rect 7286 19751 7342 19760
rect 7484 19718 7512 19790
rect 7472 19712 7524 19718
rect 7472 19654 7524 19660
rect 7196 19304 7248 19310
rect 7196 19246 7248 19252
rect 7286 19000 7342 19009
rect 7286 18935 7342 18944
rect 7194 18864 7250 18873
rect 7194 18799 7250 18808
rect 6828 18702 6880 18708
rect 7102 18728 7158 18737
rect 6736 18624 6788 18630
rect 6736 18566 6788 18572
rect 6748 18426 6776 18566
rect 6736 18420 6788 18426
rect 6736 18362 6788 18368
rect 6736 18216 6788 18222
rect 6736 18158 6788 18164
rect 6748 17542 6776 18158
rect 6840 17882 6868 18702
rect 7102 18663 7158 18672
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6736 17536 6788 17542
rect 6736 17478 6788 17484
rect 6734 16552 6790 16561
rect 6734 16487 6790 16496
rect 7012 16516 7064 16522
rect 6748 13462 6776 16487
rect 7012 16458 7064 16464
rect 7024 16114 7052 16458
rect 7012 16108 7064 16114
rect 7012 16050 7064 16056
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6828 15428 6880 15434
rect 6828 15370 6880 15376
rect 6840 15162 6868 15370
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6932 15094 6960 15506
rect 7116 15502 7144 15846
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 6920 15088 6972 15094
rect 6920 15030 6972 15036
rect 6828 14272 6880 14278
rect 7024 14226 7052 15438
rect 7208 15144 7236 18799
rect 7300 17338 7328 18935
rect 7380 18828 7432 18834
rect 7380 18770 7432 18776
rect 7392 17542 7420 18770
rect 7484 17610 7512 19654
rect 7472 17604 7524 17610
rect 7472 17546 7524 17552
rect 7380 17536 7432 17542
rect 7576 17490 7604 19887
rect 7380 17478 7432 17484
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 6880 14220 7052 14226
rect 6828 14214 7052 14220
rect 6840 14198 7052 14214
rect 7116 15116 7236 15144
rect 6736 13456 6788 13462
rect 6736 13398 6788 13404
rect 6736 12776 6788 12782
rect 6736 12718 6788 12724
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6748 11257 6776 12718
rect 6840 12442 6868 12718
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6828 12232 6880 12238
rect 6826 12200 6828 12209
rect 6880 12200 6882 12209
rect 6826 12135 6882 12144
rect 6840 11354 6868 12135
rect 6932 11898 6960 14198
rect 7116 12918 7144 15116
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7208 14618 7236 14962
rect 7196 14612 7248 14618
rect 7248 14572 7328 14600
rect 7196 14554 7248 14560
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 7116 12714 7144 12854
rect 7104 12708 7156 12714
rect 7156 12668 7236 12696
rect 7104 12650 7156 12656
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 7024 11558 7052 12310
rect 7208 12186 7236 12668
rect 7116 12158 7236 12186
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6734 11248 6790 11257
rect 6734 11183 6790 11192
rect 7010 11112 7066 11121
rect 7010 11047 7066 11056
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6932 9518 6960 10406
rect 6644 9512 6696 9518
rect 6182 9480 6238 9489
rect 6644 9454 6696 9460
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6182 9415 6238 9424
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6289 9276 6585 9296
rect 6345 9274 6369 9276
rect 6425 9274 6449 9276
rect 6505 9274 6529 9276
rect 6367 9222 6369 9274
rect 6431 9222 6443 9274
rect 6505 9222 6507 9274
rect 6345 9220 6369 9222
rect 6425 9220 6449 9222
rect 6505 9220 6529 9222
rect 6289 9200 6585 9220
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6184 8560 6236 8566
rect 6184 8502 6236 8508
rect 6196 7886 6224 8502
rect 6472 8498 6500 8774
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6289 8188 6585 8208
rect 6345 8186 6369 8188
rect 6425 8186 6449 8188
rect 6505 8186 6529 8188
rect 6367 8134 6369 8186
rect 6431 8134 6443 8186
rect 6505 8134 6507 8186
rect 6345 8132 6369 8134
rect 6425 8132 6449 8134
rect 6505 8132 6529 8134
rect 6289 8112 6585 8132
rect 6656 8022 6684 9318
rect 6932 9178 6960 9454
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6932 8106 6960 8774
rect 6840 8090 6960 8106
rect 6828 8084 6960 8090
rect 6880 8078 6960 8084
rect 6828 8026 6880 8032
rect 6644 8016 6696 8022
rect 6644 7958 6696 7964
rect 6736 8016 6788 8022
rect 6736 7958 6788 7964
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6196 7546 6224 7822
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6289 7100 6585 7120
rect 6345 7098 6369 7100
rect 6425 7098 6449 7100
rect 6505 7098 6529 7100
rect 6367 7046 6369 7098
rect 6431 7046 6443 7098
rect 6505 7046 6507 7098
rect 6345 7044 6369 7046
rect 6425 7044 6449 7046
rect 6505 7044 6529 7046
rect 6289 7024 6585 7044
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 6184 6248 6236 6254
rect 6184 6190 6236 6196
rect 6012 6072 6132 6100
rect 6000 5840 6052 5846
rect 6000 5782 6052 5788
rect 5908 3664 5960 3670
rect 5908 3606 5960 3612
rect 5920 2514 5948 3606
rect 6012 2689 6040 5782
rect 6104 4146 6132 6072
rect 6196 5794 6224 6190
rect 6288 6186 6316 6802
rect 6276 6180 6328 6186
rect 6276 6122 6328 6128
rect 6289 6012 6585 6032
rect 6345 6010 6369 6012
rect 6425 6010 6449 6012
rect 6505 6010 6529 6012
rect 6367 5958 6369 6010
rect 6431 5958 6443 6010
rect 6505 5958 6507 6010
rect 6345 5956 6369 5958
rect 6425 5956 6449 5958
rect 6505 5956 6529 5958
rect 6289 5936 6585 5956
rect 6274 5808 6330 5817
rect 6196 5766 6274 5794
rect 6748 5794 6776 7958
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6826 6896 6882 6905
rect 6826 6831 6882 6840
rect 6840 6458 6868 6831
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6840 5846 6868 6054
rect 6274 5743 6330 5752
rect 6656 5766 6776 5794
rect 6828 5840 6880 5846
rect 6828 5782 6880 5788
rect 6182 5672 6238 5681
rect 6288 5642 6316 5743
rect 6182 5607 6238 5616
rect 6276 5636 6328 5642
rect 6196 4690 6224 5607
rect 6276 5578 6328 5584
rect 6289 4924 6585 4944
rect 6345 4922 6369 4924
rect 6425 4922 6449 4924
rect 6505 4922 6529 4924
rect 6367 4870 6369 4922
rect 6431 4870 6443 4922
rect 6505 4870 6507 4922
rect 6345 4868 6369 4870
rect 6425 4868 6449 4870
rect 6505 4868 6529 4870
rect 6289 4848 6585 4868
rect 6274 4720 6330 4729
rect 6184 4684 6236 4690
rect 6274 4655 6330 4664
rect 6460 4684 6512 4690
rect 6184 4626 6236 4632
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 6288 4078 6316 4655
rect 6460 4626 6512 4632
rect 6276 4072 6328 4078
rect 6182 4040 6238 4049
rect 6276 4014 6328 4020
rect 6472 4010 6500 4626
rect 6182 3975 6238 3984
rect 6460 4004 6512 4010
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6104 3398 6132 3878
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 5998 2680 6054 2689
rect 5998 2615 6054 2624
rect 5908 2508 5960 2514
rect 5908 2450 5960 2456
rect 6196 480 6224 3975
rect 6460 3946 6512 3952
rect 6289 3836 6585 3856
rect 6345 3834 6369 3836
rect 6425 3834 6449 3836
rect 6505 3834 6529 3836
rect 6367 3782 6369 3834
rect 6431 3782 6443 3834
rect 6505 3782 6507 3834
rect 6345 3780 6369 3782
rect 6425 3780 6449 3782
rect 6505 3780 6529 3782
rect 6289 3760 6585 3780
rect 6656 3618 6684 5766
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6564 3590 6684 3618
rect 6564 3194 6592 3590
rect 6642 3496 6698 3505
rect 6748 3466 6776 5646
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6840 4758 6868 4966
rect 6828 4752 6880 4758
rect 6828 4694 6880 4700
rect 6932 4706 6960 7686
rect 7024 6390 7052 11047
rect 7116 10130 7144 12158
rect 7196 12096 7248 12102
rect 7300 12084 7328 14572
rect 7248 12056 7328 12084
rect 7196 12038 7248 12044
rect 7300 11762 7328 12056
rect 7392 11801 7420 17478
rect 7484 17462 7604 17490
rect 7378 11792 7434 11801
rect 7288 11756 7340 11762
rect 7208 11716 7288 11744
rect 7208 11286 7236 11716
rect 7378 11727 7434 11736
rect 7288 11698 7340 11704
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 7300 11354 7328 11562
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7196 11280 7248 11286
rect 7196 11222 7248 11228
rect 7392 10266 7420 11630
rect 7484 11354 7512 17462
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 7576 14482 7604 16934
rect 7668 16658 7696 20878
rect 7656 16652 7708 16658
rect 7656 16594 7708 16600
rect 7656 15972 7708 15978
rect 7656 15914 7708 15920
rect 7668 15026 7696 15914
rect 7656 15020 7708 15026
rect 7656 14962 7708 14968
rect 7656 14884 7708 14890
rect 7656 14826 7708 14832
rect 7668 14618 7696 14826
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7576 14074 7604 14418
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 7656 13184 7708 13190
rect 7576 13144 7656 13172
rect 7576 11694 7604 13144
rect 7656 13126 7708 13132
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7484 10810 7512 11290
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7576 10470 7604 11154
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7196 10192 7248 10198
rect 7196 10134 7248 10140
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 7208 9654 7236 10134
rect 7104 9648 7156 9654
rect 7104 9590 7156 9596
rect 7196 9648 7248 9654
rect 7196 9590 7248 9596
rect 7116 9042 7144 9590
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7116 8634 7144 8978
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 6932 4678 7052 4706
rect 7024 4434 7052 4678
rect 6932 4406 7052 4434
rect 6826 3768 6882 3777
rect 6826 3703 6882 3712
rect 6642 3431 6698 3440
rect 6736 3460 6788 3466
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6564 2990 6592 3130
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 6289 2748 6585 2768
rect 6345 2746 6369 2748
rect 6425 2746 6449 2748
rect 6505 2746 6529 2748
rect 6367 2694 6369 2746
rect 6431 2694 6443 2746
rect 6505 2694 6507 2746
rect 6345 2692 6369 2694
rect 6425 2692 6449 2694
rect 6505 2692 6529 2694
rect 6289 2672 6585 2692
rect 6656 1714 6684 3431
rect 6736 3402 6788 3408
rect 6840 3126 6868 3703
rect 6828 3120 6880 3126
rect 6828 3062 6880 3068
rect 6564 1686 6684 1714
rect 6564 480 6592 1686
rect 6932 480 6960 4406
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 7024 3641 7052 3878
rect 7116 3777 7144 8570
rect 7194 7984 7250 7993
rect 7194 7919 7196 7928
rect 7248 7919 7250 7928
rect 7196 7890 7248 7896
rect 7208 7546 7236 7890
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 7300 6322 7328 6666
rect 7484 6322 7512 6802
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7576 6202 7604 10406
rect 7668 10198 7696 12786
rect 7760 11218 7788 28614
rect 7944 24750 7972 31640
rect 8024 31622 8076 31628
rect 8036 31346 8064 31622
rect 8024 31340 8076 31346
rect 8024 31282 8076 31288
rect 8116 31272 8168 31278
rect 8116 31214 8168 31220
rect 8128 30938 8156 31214
rect 8116 30932 8168 30938
rect 8116 30874 8168 30880
rect 8024 30864 8076 30870
rect 8496 30841 8524 34983
rect 8588 34513 8616 39520
rect 8956 37210 8984 39520
rect 8680 37182 8984 37210
rect 8574 34504 8630 34513
rect 8574 34439 8630 34448
rect 8680 32881 8708 37182
rect 8956 37020 9252 37040
rect 9012 37018 9036 37020
rect 9092 37018 9116 37020
rect 9172 37018 9196 37020
rect 9034 36966 9036 37018
rect 9098 36966 9110 37018
rect 9172 36966 9174 37018
rect 9012 36964 9036 36966
rect 9092 36964 9116 36966
rect 9172 36964 9196 36966
rect 8956 36944 9252 36964
rect 8956 35932 9252 35952
rect 9012 35930 9036 35932
rect 9092 35930 9116 35932
rect 9172 35930 9196 35932
rect 9034 35878 9036 35930
rect 9098 35878 9110 35930
rect 9172 35878 9174 35930
rect 9012 35876 9036 35878
rect 9092 35876 9116 35878
rect 9172 35876 9196 35878
rect 8956 35856 9252 35876
rect 8852 35488 8904 35494
rect 8852 35430 8904 35436
rect 8864 35193 8892 35430
rect 8850 35184 8906 35193
rect 8850 35119 8906 35128
rect 9312 35148 9364 35154
rect 9312 35090 9364 35096
rect 8956 34844 9252 34864
rect 9012 34842 9036 34844
rect 9092 34842 9116 34844
rect 9172 34842 9196 34844
rect 9034 34790 9036 34842
rect 9098 34790 9110 34842
rect 9172 34790 9174 34842
rect 9012 34788 9036 34790
rect 9092 34788 9116 34790
rect 9172 34788 9196 34790
rect 8956 34768 9252 34788
rect 8760 34468 8812 34474
rect 8760 34410 8812 34416
rect 8772 34202 8800 34410
rect 9324 34406 9352 35090
rect 9312 34400 9364 34406
rect 9312 34342 9364 34348
rect 8760 34196 8812 34202
rect 8760 34138 8812 34144
rect 9416 33946 9444 39520
rect 9784 35290 9812 39520
rect 9864 35760 9916 35766
rect 9862 35728 9864 35737
rect 9916 35728 9918 35737
rect 10152 35714 10180 39520
rect 10612 35714 10640 39520
rect 10980 39494 11100 39520
rect 9862 35663 9918 35672
rect 9968 35686 10180 35714
rect 10428 35686 10640 35714
rect 9772 35284 9824 35290
rect 9772 35226 9824 35232
rect 9772 35080 9824 35086
rect 9772 35022 9824 35028
rect 9784 34746 9812 35022
rect 9864 35012 9916 35018
rect 9864 34954 9916 34960
rect 9772 34740 9824 34746
rect 9772 34682 9824 34688
rect 9784 34649 9812 34682
rect 9876 34678 9904 34954
rect 9864 34672 9916 34678
rect 9770 34640 9826 34649
rect 9864 34614 9916 34620
rect 9770 34575 9826 34584
rect 9876 34202 9904 34614
rect 9864 34196 9916 34202
rect 9864 34138 9916 34144
rect 9416 33918 9536 33946
rect 9404 33856 9456 33862
rect 9404 33798 9456 33804
rect 8956 33756 9252 33776
rect 9012 33754 9036 33756
rect 9092 33754 9116 33756
rect 9172 33754 9196 33756
rect 9034 33702 9036 33754
rect 9098 33702 9110 33754
rect 9172 33702 9174 33754
rect 9012 33700 9036 33702
rect 9092 33700 9116 33702
rect 9172 33700 9196 33702
rect 8956 33680 9252 33700
rect 9312 33584 9364 33590
rect 9310 33552 9312 33561
rect 9364 33552 9366 33561
rect 9310 33487 9366 33496
rect 8758 33416 8814 33425
rect 9416 33386 9444 33798
rect 8758 33351 8814 33360
rect 9404 33380 9456 33386
rect 8666 32872 8722 32881
rect 8666 32807 8722 32816
rect 8576 32564 8628 32570
rect 8576 32506 8628 32512
rect 8588 32026 8616 32506
rect 8576 32020 8628 32026
rect 8576 31962 8628 31968
rect 8024 30806 8076 30812
rect 8482 30832 8538 30841
rect 8036 24857 8064 30806
rect 8482 30767 8538 30776
rect 8576 29504 8628 29510
rect 8576 29446 8628 29452
rect 8588 29170 8616 29446
rect 8576 29164 8628 29170
rect 8576 29106 8628 29112
rect 8300 29096 8352 29102
rect 8300 29038 8352 29044
rect 8116 28960 8168 28966
rect 8116 28902 8168 28908
rect 8128 26926 8156 28902
rect 8312 27554 8340 29038
rect 8392 28620 8444 28626
rect 8392 28562 8444 28568
rect 8404 27674 8432 28562
rect 8484 28552 8536 28558
rect 8484 28494 8536 28500
rect 8496 27946 8524 28494
rect 8588 28218 8616 29106
rect 8576 28212 8628 28218
rect 8576 28154 8628 28160
rect 8484 27940 8536 27946
rect 8484 27882 8536 27888
rect 8392 27668 8444 27674
rect 8392 27610 8444 27616
rect 8220 27538 8340 27554
rect 8208 27532 8340 27538
rect 8260 27526 8340 27532
rect 8208 27474 8260 27480
rect 8208 27328 8260 27334
rect 8208 27270 8260 27276
rect 8220 27130 8248 27270
rect 8208 27124 8260 27130
rect 8208 27066 8260 27072
rect 8116 26920 8168 26926
rect 8116 26862 8168 26868
rect 8312 25294 8340 27526
rect 8392 27328 8444 27334
rect 8392 27270 8444 27276
rect 8668 27328 8720 27334
rect 8668 27270 8720 27276
rect 8404 26994 8432 27270
rect 8392 26988 8444 26994
rect 8392 26930 8444 26936
rect 8576 26240 8628 26246
rect 8576 26182 8628 26188
rect 8588 25838 8616 26182
rect 8576 25832 8628 25838
rect 8576 25774 8628 25780
rect 8300 25288 8352 25294
rect 8300 25230 8352 25236
rect 8022 24848 8078 24857
rect 8312 24818 8340 25230
rect 8022 24783 8078 24792
rect 8300 24812 8352 24818
rect 8300 24754 8352 24760
rect 7932 24744 7984 24750
rect 7932 24686 7984 24692
rect 7944 24313 7972 24686
rect 8024 24608 8076 24614
rect 8024 24550 8076 24556
rect 7930 24304 7986 24313
rect 7930 24239 7986 24248
rect 8036 23866 8064 24550
rect 8392 24064 8444 24070
rect 8392 24006 8444 24012
rect 8024 23860 8076 23866
rect 8024 23802 8076 23808
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 8208 23180 8260 23186
rect 8208 23122 8260 23128
rect 7852 22234 7880 23122
rect 8024 23112 8076 23118
rect 8024 23054 8076 23060
rect 8036 22778 8064 23054
rect 8024 22772 8076 22778
rect 8024 22714 8076 22720
rect 8220 22438 8248 23122
rect 8404 22982 8432 24006
rect 8588 23338 8616 25774
rect 8496 23310 8616 23338
rect 8392 22976 8444 22982
rect 8392 22918 8444 22924
rect 8404 22658 8432 22918
rect 8496 22778 8524 23310
rect 8484 22772 8536 22778
rect 8484 22714 8536 22720
rect 8404 22630 8524 22658
rect 8208 22432 8260 22438
rect 8208 22374 8260 22380
rect 7840 22228 7892 22234
rect 7840 22170 7892 22176
rect 8220 22137 8248 22374
rect 8206 22128 8262 22137
rect 8206 22063 8262 22072
rect 8496 21894 8524 22630
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 8496 21486 8524 21830
rect 8484 21480 8536 21486
rect 8484 21422 8536 21428
rect 8496 21010 8524 21422
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 8484 21004 8536 21010
rect 8484 20946 8536 20952
rect 8024 20936 8076 20942
rect 8024 20878 8076 20884
rect 8220 20890 8248 20946
rect 8680 20890 8708 27270
rect 8772 25401 8800 33351
rect 9404 33322 9456 33328
rect 9312 33108 9364 33114
rect 9312 33050 9364 33056
rect 8852 32836 8904 32842
rect 8852 32778 8904 32784
rect 8864 32366 8892 32778
rect 8956 32668 9252 32688
rect 9012 32666 9036 32668
rect 9092 32666 9116 32668
rect 9172 32666 9196 32668
rect 9034 32614 9036 32666
rect 9098 32614 9110 32666
rect 9172 32614 9174 32666
rect 9012 32612 9036 32614
rect 9092 32612 9116 32614
rect 9172 32612 9196 32614
rect 8956 32592 9252 32612
rect 9324 32434 9352 33050
rect 9312 32428 9364 32434
rect 9312 32370 9364 32376
rect 8852 32360 8904 32366
rect 8852 32302 8904 32308
rect 8852 32224 8904 32230
rect 8852 32166 8904 32172
rect 8864 31686 8892 32166
rect 8852 31680 8904 31686
rect 8852 31622 8904 31628
rect 8864 31482 8892 31622
rect 8956 31580 9252 31600
rect 9012 31578 9036 31580
rect 9092 31578 9116 31580
rect 9172 31578 9196 31580
rect 9034 31526 9036 31578
rect 9098 31526 9110 31578
rect 9172 31526 9174 31578
rect 9012 31524 9036 31526
rect 9092 31524 9116 31526
rect 9172 31524 9196 31526
rect 8956 31504 9252 31524
rect 9416 31482 9444 33322
rect 9508 32745 9536 33918
rect 9680 33856 9732 33862
rect 9680 33798 9732 33804
rect 9692 33454 9720 33798
rect 9772 33516 9824 33522
rect 9772 33458 9824 33464
rect 9680 33448 9732 33454
rect 9680 33390 9732 33396
rect 9588 33312 9640 33318
rect 9640 33260 9720 33266
rect 9588 33254 9720 33260
rect 9600 33238 9720 33254
rect 9692 32978 9720 33238
rect 9680 32972 9732 32978
rect 9680 32914 9732 32920
rect 9678 32872 9734 32881
rect 9678 32807 9734 32816
rect 9494 32736 9550 32745
rect 9494 32671 9550 32680
rect 9692 32570 9720 32807
rect 9680 32564 9732 32570
rect 9680 32506 9732 32512
rect 9678 32328 9734 32337
rect 9678 32263 9680 32272
rect 9732 32263 9734 32272
rect 9680 32234 9732 32240
rect 9496 32020 9548 32026
rect 9496 31962 9548 31968
rect 8852 31476 8904 31482
rect 8852 31418 8904 31424
rect 9404 31476 9456 31482
rect 9404 31418 9456 31424
rect 9310 31376 9366 31385
rect 9310 31311 9366 31320
rect 9324 30938 9352 31311
rect 9508 31278 9536 31962
rect 9588 31680 9640 31686
rect 9588 31622 9640 31628
rect 9600 31414 9628 31622
rect 9588 31408 9640 31414
rect 9588 31350 9640 31356
rect 9496 31272 9548 31278
rect 9496 31214 9548 31220
rect 9680 31204 9732 31210
rect 9680 31146 9732 31152
rect 9588 31136 9640 31142
rect 9586 31104 9588 31113
rect 9640 31104 9642 31113
rect 9586 31039 9642 31048
rect 9312 30932 9364 30938
rect 9312 30874 9364 30880
rect 8956 30492 9252 30512
rect 9012 30490 9036 30492
rect 9092 30490 9116 30492
rect 9172 30490 9196 30492
rect 9034 30438 9036 30490
rect 9098 30438 9110 30490
rect 9172 30438 9174 30490
rect 9012 30436 9036 30438
rect 9092 30436 9116 30438
rect 9172 30436 9196 30438
rect 8956 30416 9252 30436
rect 9324 29782 9352 30874
rect 9312 29776 9364 29782
rect 9312 29718 9364 29724
rect 8956 29404 9252 29424
rect 9012 29402 9036 29404
rect 9092 29402 9116 29404
rect 9172 29402 9196 29404
rect 9034 29350 9036 29402
rect 9098 29350 9110 29402
rect 9172 29350 9174 29402
rect 9012 29348 9036 29350
rect 9092 29348 9116 29350
rect 9172 29348 9196 29350
rect 8956 29328 9252 29348
rect 9324 29306 9352 29718
rect 9312 29300 9364 29306
rect 9312 29242 9364 29248
rect 9588 29164 9640 29170
rect 9588 29106 9640 29112
rect 9600 28762 9628 29106
rect 9692 29050 9720 31146
rect 9784 31090 9812 33458
rect 9864 33312 9916 33318
rect 9864 33254 9916 33260
rect 9876 31385 9904 33254
rect 9862 31376 9918 31385
rect 9862 31311 9864 31320
rect 9916 31311 9918 31320
rect 9864 31282 9916 31288
rect 9876 31251 9904 31282
rect 9968 31210 9996 35686
rect 10048 35488 10100 35494
rect 10048 35430 10100 35436
rect 9956 31204 10008 31210
rect 9956 31146 10008 31152
rect 9784 31062 9996 31090
rect 9968 29510 9996 31062
rect 9956 29504 10008 29510
rect 9956 29446 10008 29452
rect 9968 29306 9996 29446
rect 9956 29300 10008 29306
rect 9956 29242 10008 29248
rect 9692 29022 9904 29050
rect 9680 28960 9732 28966
rect 9680 28902 9732 28908
rect 9588 28756 9640 28762
rect 9588 28698 9640 28704
rect 9692 28694 9720 28902
rect 9680 28688 9732 28694
rect 9586 28656 9642 28665
rect 9680 28630 9732 28636
rect 9586 28591 9642 28600
rect 9404 28552 9456 28558
rect 8850 28520 8906 28529
rect 9404 28494 9456 28500
rect 8850 28455 8906 28464
rect 8864 28150 8892 28455
rect 8956 28316 9252 28336
rect 9012 28314 9036 28316
rect 9092 28314 9116 28316
rect 9172 28314 9196 28316
rect 9034 28262 9036 28314
rect 9098 28262 9110 28314
rect 9172 28262 9174 28314
rect 9012 28260 9036 28262
rect 9092 28260 9116 28262
rect 9172 28260 9196 28262
rect 8956 28240 9252 28260
rect 8852 28144 8904 28150
rect 8852 28086 8904 28092
rect 8864 27878 8892 28086
rect 9416 28014 9444 28494
rect 9494 28112 9550 28121
rect 9494 28047 9550 28056
rect 9404 28008 9456 28014
rect 9404 27950 9456 27956
rect 8852 27872 8904 27878
rect 8852 27814 8904 27820
rect 9312 27872 9364 27878
rect 9312 27814 9364 27820
rect 9324 27713 9352 27814
rect 9310 27704 9366 27713
rect 9310 27639 9366 27648
rect 8956 27228 9252 27248
rect 9012 27226 9036 27228
rect 9092 27226 9116 27228
rect 9172 27226 9196 27228
rect 9034 27174 9036 27226
rect 9098 27174 9110 27226
rect 9172 27174 9174 27226
rect 9012 27172 9036 27174
rect 9092 27172 9116 27174
rect 9172 27172 9196 27174
rect 8956 27152 9252 27172
rect 9416 26314 9444 27950
rect 9508 27878 9536 28047
rect 9600 27946 9628 28591
rect 9692 28558 9720 28630
rect 9680 28552 9732 28558
rect 9680 28494 9732 28500
rect 9588 27940 9640 27946
rect 9588 27882 9640 27888
rect 9496 27872 9548 27878
rect 9496 27814 9548 27820
rect 9508 27334 9536 27814
rect 9496 27328 9548 27334
rect 9496 27270 9548 27276
rect 9600 27146 9628 27882
rect 9508 27118 9628 27146
rect 9404 26308 9456 26314
rect 9404 26250 9456 26256
rect 8956 26140 9252 26160
rect 9012 26138 9036 26140
rect 9092 26138 9116 26140
rect 9172 26138 9196 26140
rect 9034 26086 9036 26138
rect 9098 26086 9110 26138
rect 9172 26086 9174 26138
rect 9012 26084 9036 26086
rect 9092 26084 9116 26086
rect 9172 26084 9196 26086
rect 8956 26064 9252 26084
rect 9416 25906 9444 26250
rect 9312 25900 9364 25906
rect 9312 25842 9364 25848
rect 9404 25900 9456 25906
rect 9404 25842 9456 25848
rect 8852 25696 8904 25702
rect 8852 25638 8904 25644
rect 8864 25498 8892 25638
rect 9324 25498 9352 25842
rect 8852 25492 8904 25498
rect 8852 25434 8904 25440
rect 9312 25492 9364 25498
rect 9312 25434 9364 25440
rect 8758 25392 8814 25401
rect 8758 25327 8814 25336
rect 8772 24818 8800 25327
rect 8956 25052 9252 25072
rect 9012 25050 9036 25052
rect 9092 25050 9116 25052
rect 9172 25050 9196 25052
rect 9034 24998 9036 25050
rect 9098 24998 9110 25050
rect 9172 24998 9174 25050
rect 9012 24996 9036 24998
rect 9092 24996 9116 24998
rect 9172 24996 9196 24998
rect 8956 24976 9252 24996
rect 9402 24984 9458 24993
rect 9402 24919 9458 24928
rect 8760 24812 8812 24818
rect 8760 24754 8812 24760
rect 9128 24744 9180 24750
rect 9128 24686 9180 24692
rect 9220 24744 9272 24750
rect 9220 24686 9272 24692
rect 9140 24138 9168 24686
rect 9232 24410 9260 24686
rect 9312 24676 9364 24682
rect 9312 24618 9364 24624
rect 9220 24404 9272 24410
rect 9220 24346 9272 24352
rect 9128 24132 9180 24138
rect 9128 24074 9180 24080
rect 8956 23964 9252 23984
rect 9012 23962 9036 23964
rect 9092 23962 9116 23964
rect 9172 23962 9196 23964
rect 9034 23910 9036 23962
rect 9098 23910 9110 23962
rect 9172 23910 9174 23962
rect 9012 23908 9036 23910
rect 9092 23908 9116 23910
rect 9172 23908 9196 23910
rect 8956 23888 9252 23908
rect 8852 23792 8904 23798
rect 8850 23760 8852 23769
rect 8904 23760 8906 23769
rect 8850 23695 8906 23704
rect 8956 22876 9252 22896
rect 9012 22874 9036 22876
rect 9092 22874 9116 22876
rect 9172 22874 9196 22876
rect 9034 22822 9036 22874
rect 9098 22822 9110 22874
rect 9172 22822 9174 22874
rect 9012 22820 9036 22822
rect 9092 22820 9116 22822
rect 9172 22820 9196 22822
rect 8956 22800 9252 22820
rect 8956 21788 9252 21808
rect 9012 21786 9036 21788
rect 9092 21786 9116 21788
rect 9172 21786 9196 21788
rect 9034 21734 9036 21786
rect 9098 21734 9110 21786
rect 9172 21734 9174 21786
rect 9012 21732 9036 21734
rect 9092 21732 9116 21734
rect 9172 21732 9196 21734
rect 8956 21712 9252 21732
rect 8852 21412 8904 21418
rect 8852 21354 8904 21360
rect 8864 21146 8892 21354
rect 8852 21140 8904 21146
rect 8852 21082 8904 21088
rect 8760 21072 8812 21078
rect 8760 21014 8812 21020
rect 8036 20534 8064 20878
rect 8220 20862 8340 20890
rect 8312 20602 8340 20862
rect 8404 20862 8708 20890
rect 8300 20596 8352 20602
rect 8300 20538 8352 20544
rect 8024 20528 8076 20534
rect 8024 20470 8076 20476
rect 7840 20052 7892 20058
rect 7840 19994 7892 20000
rect 7852 17882 7880 19994
rect 8036 19378 8064 20470
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 8312 19854 8340 20198
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 8220 19446 8248 19790
rect 8208 19440 8260 19446
rect 8208 19382 8260 19388
rect 8024 19372 8076 19378
rect 8024 19314 8076 19320
rect 7932 19304 7984 19310
rect 7932 19246 7984 19252
rect 7840 17876 7892 17882
rect 7840 17818 7892 17824
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 7852 15162 7880 16390
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 7852 14958 7880 15098
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 7944 14618 7972 19246
rect 8036 18970 8064 19314
rect 8116 19168 8168 19174
rect 8116 19110 8168 19116
rect 8024 18964 8076 18970
rect 8024 18906 8076 18912
rect 8036 18358 8064 18906
rect 8024 18352 8076 18358
rect 8024 18294 8076 18300
rect 8022 18184 8078 18193
rect 8022 18119 8078 18128
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 7944 14074 7972 14554
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 8036 13954 8064 18119
rect 8128 15201 8156 19110
rect 8220 18970 8248 19382
rect 8208 18964 8260 18970
rect 8208 18906 8260 18912
rect 8312 18426 8340 19790
rect 8404 19258 8432 20862
rect 8772 19718 8800 21014
rect 8864 20058 8892 21082
rect 8956 20700 9252 20720
rect 9012 20698 9036 20700
rect 9092 20698 9116 20700
rect 9172 20698 9196 20700
rect 9034 20646 9036 20698
rect 9098 20646 9110 20698
rect 9172 20646 9174 20698
rect 9012 20644 9036 20646
rect 9092 20644 9116 20646
rect 9172 20644 9196 20646
rect 8956 20624 9252 20644
rect 8852 20052 8904 20058
rect 8852 19994 8904 20000
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 8666 19408 8722 19417
rect 8666 19343 8722 19352
rect 8680 19258 8708 19343
rect 8772 19310 8800 19654
rect 8864 19378 8892 19994
rect 8956 19612 9252 19632
rect 9012 19610 9036 19612
rect 9092 19610 9116 19612
rect 9172 19610 9196 19612
rect 9034 19558 9036 19610
rect 9098 19558 9110 19610
rect 9172 19558 9174 19610
rect 9012 19556 9036 19558
rect 9092 19556 9116 19558
rect 9172 19556 9196 19558
rect 8956 19536 9252 19556
rect 8852 19372 8904 19378
rect 8852 19314 8904 19320
rect 8404 19230 8708 19258
rect 8760 19304 8812 19310
rect 8760 19246 8812 19252
rect 8850 19272 8906 19281
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 8390 19000 8446 19009
rect 8390 18935 8446 18944
rect 8404 18698 8432 18935
rect 8392 18692 8444 18698
rect 8392 18634 8444 18640
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 8390 18184 8446 18193
rect 8390 18119 8446 18128
rect 8404 17814 8432 18119
rect 8496 17882 8524 19110
rect 8576 18352 8628 18358
rect 8576 18294 8628 18300
rect 8484 17876 8536 17882
rect 8484 17818 8536 17824
rect 8392 17808 8444 17814
rect 8392 17750 8444 17756
rect 8404 17270 8432 17750
rect 8496 17338 8524 17818
rect 8588 17678 8616 18294
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8392 17264 8444 17270
rect 8392 17206 8444 17212
rect 8588 17202 8616 17614
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8680 17082 8708 19230
rect 8496 17054 8708 17082
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8220 15706 8248 16594
rect 8300 16584 8352 16590
rect 8300 16526 8352 16532
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8312 15881 8340 16526
rect 8298 15872 8354 15881
rect 8298 15807 8354 15816
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8404 15366 8432 16526
rect 8208 15360 8260 15366
rect 8208 15302 8260 15308
rect 8392 15360 8444 15366
rect 8392 15302 8444 15308
rect 8114 15192 8170 15201
rect 8114 15127 8170 15136
rect 8114 14920 8170 14929
rect 8114 14855 8170 14864
rect 8128 14482 8156 14855
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 8128 14006 8156 14418
rect 8220 14414 8248 15302
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 7944 13926 8064 13954
rect 8116 14000 8168 14006
rect 8116 13942 8168 13948
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 7852 12986 7880 13330
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7944 11642 7972 13926
rect 8128 13841 8156 13942
rect 8220 13870 8248 14350
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 8208 13864 8260 13870
rect 8114 13832 8170 13841
rect 8208 13806 8260 13812
rect 8114 13767 8170 13776
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8128 12986 8156 13126
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 8220 12374 8248 13806
rect 8312 13530 8340 14214
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8496 13410 8524 17054
rect 8666 15192 8722 15201
rect 8666 15127 8722 15136
rect 8312 13382 8524 13410
rect 8576 13388 8628 13394
rect 8312 12617 8340 13382
rect 8576 13330 8628 13336
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 8404 12986 8432 13194
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 8298 12608 8354 12617
rect 8298 12543 8354 12552
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 8496 12209 8524 12786
rect 8588 12782 8616 13330
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8588 12374 8616 12718
rect 8680 12714 8708 15127
rect 8772 14226 8800 19246
rect 8850 19207 8852 19216
rect 8904 19207 8906 19216
rect 8852 19178 8904 19184
rect 9324 18850 9352 24618
rect 9416 23662 9444 24919
rect 9404 23656 9456 23662
rect 9404 23598 9456 23604
rect 9416 23322 9444 23598
rect 9404 23316 9456 23322
rect 9404 23258 9456 23264
rect 9416 23089 9444 23258
rect 9402 23080 9458 23089
rect 9402 23015 9458 23024
rect 9404 21344 9456 21350
rect 9404 21286 9456 21292
rect 9416 20602 9444 21286
rect 9404 20596 9456 20602
rect 9404 20538 9456 20544
rect 9324 18822 9444 18850
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 8956 18524 9252 18544
rect 9012 18522 9036 18524
rect 9092 18522 9116 18524
rect 9172 18522 9196 18524
rect 9034 18470 9036 18522
rect 9098 18470 9110 18522
rect 9172 18470 9174 18522
rect 9012 18468 9036 18470
rect 9092 18468 9116 18470
rect 9172 18468 9196 18470
rect 8956 18448 9252 18468
rect 9324 18358 9352 18702
rect 9312 18352 9364 18358
rect 9312 18294 9364 18300
rect 8956 17436 9252 17456
rect 9012 17434 9036 17436
rect 9092 17434 9116 17436
rect 9172 17434 9196 17436
rect 9034 17382 9036 17434
rect 9098 17382 9110 17434
rect 9172 17382 9174 17434
rect 9012 17380 9036 17382
rect 9092 17380 9116 17382
rect 9172 17380 9196 17382
rect 8956 17360 9252 17380
rect 9312 16516 9364 16522
rect 9312 16458 9364 16464
rect 8956 16348 9252 16368
rect 9012 16346 9036 16348
rect 9092 16346 9116 16348
rect 9172 16346 9196 16348
rect 9034 16294 9036 16346
rect 9098 16294 9110 16346
rect 9172 16294 9174 16346
rect 9012 16292 9036 16294
rect 9092 16292 9116 16294
rect 9172 16292 9196 16294
rect 8956 16272 9252 16292
rect 9218 16144 9274 16153
rect 9324 16130 9352 16458
rect 9274 16102 9352 16130
rect 9218 16079 9220 16088
rect 9272 16079 9274 16088
rect 9220 16050 9272 16056
rect 8852 15904 8904 15910
rect 8850 15872 8852 15881
rect 8904 15872 8906 15881
rect 8850 15807 8906 15816
rect 9232 15706 9260 16050
rect 9312 16040 9364 16046
rect 9416 15994 9444 18822
rect 9364 15988 9444 15994
rect 9312 15982 9444 15988
rect 9324 15966 9444 15982
rect 9220 15700 9272 15706
rect 9220 15642 9272 15648
rect 9232 15450 9260 15642
rect 9232 15422 9352 15450
rect 8956 15260 9252 15280
rect 9012 15258 9036 15260
rect 9092 15258 9116 15260
rect 9172 15258 9196 15260
rect 9034 15206 9036 15258
rect 9098 15206 9110 15258
rect 9172 15206 9174 15258
rect 9012 15204 9036 15206
rect 9092 15204 9116 15206
rect 9172 15204 9196 15206
rect 8956 15184 9252 15204
rect 8772 14198 8892 14226
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 8668 12708 8720 12714
rect 8668 12650 8720 12656
rect 8666 12608 8722 12617
rect 8666 12543 8722 12552
rect 8576 12368 8628 12374
rect 8576 12310 8628 12316
rect 8576 12232 8628 12238
rect 8482 12200 8538 12209
rect 8538 12180 8576 12186
rect 8538 12174 8628 12180
rect 8538 12158 8616 12174
rect 8482 12135 8538 12144
rect 8496 12075 8524 12135
rect 8588 11694 8616 12158
rect 8300 11688 8352 11694
rect 7944 11614 8064 11642
rect 8300 11630 8352 11636
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 7840 11552 7892 11558
rect 7892 11500 7972 11506
rect 7840 11494 7972 11500
rect 7852 11478 7972 11494
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 7852 10674 7880 11154
rect 7944 11150 7972 11478
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 7944 10810 7972 11086
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7760 9722 7788 10066
rect 7944 10062 7972 10746
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7748 9716 7800 9722
rect 7484 6174 7604 6202
rect 7668 9676 7748 9704
rect 7378 5672 7434 5681
rect 7378 5607 7434 5616
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7300 5234 7328 5510
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 7208 4729 7236 5102
rect 7194 4720 7250 4729
rect 7194 4655 7250 4664
rect 7102 3768 7158 3777
rect 7102 3703 7104 3712
rect 7156 3703 7158 3712
rect 7104 3674 7156 3680
rect 7010 3632 7066 3641
rect 7010 3567 7066 3576
rect 7010 2952 7066 2961
rect 7010 2887 7066 2896
rect 7024 2854 7052 2887
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7116 1465 7144 2246
rect 7102 1456 7158 1465
rect 7102 1391 7158 1400
rect 7392 480 7420 5607
rect 7484 5001 7512 6174
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7576 5710 7604 6054
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7470 4992 7526 5001
rect 7470 4927 7526 4936
rect 7576 4826 7604 5646
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7668 4298 7696 9676
rect 7748 9658 7800 9664
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 7746 9480 7802 9489
rect 7746 9415 7802 9424
rect 7760 9178 7788 9415
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7760 8090 7788 9114
rect 7944 8974 7972 9522
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 7944 8634 7972 8910
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7840 7268 7892 7274
rect 7840 7210 7892 7216
rect 7852 6798 7880 7210
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7760 6662 7788 6734
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7576 4270 7696 4298
rect 7760 4282 7788 6598
rect 7852 6118 7880 6734
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7944 5914 7972 6802
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 8036 5846 8064 11614
rect 8312 11218 8340 11630
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8392 11280 8444 11286
rect 8392 11222 8444 11228
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 8404 10538 8432 11222
rect 8392 10532 8444 10538
rect 8392 10474 8444 10480
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 8128 9586 8156 10406
rect 8404 10198 8432 10474
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8300 10056 8352 10062
rect 8496 10033 8524 11290
rect 8680 11121 8708 12543
rect 8666 11112 8722 11121
rect 8666 11047 8722 11056
rect 8772 10554 8800 14010
rect 8864 13682 8892 14198
rect 8956 14172 9252 14192
rect 9012 14170 9036 14172
rect 9092 14170 9116 14172
rect 9172 14170 9196 14172
rect 9034 14118 9036 14170
rect 9098 14118 9110 14170
rect 9172 14118 9174 14170
rect 9012 14116 9036 14118
rect 9092 14116 9116 14118
rect 9172 14116 9196 14118
rect 8956 14096 9252 14116
rect 8864 13654 8984 13682
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8864 12850 8892 13466
rect 8956 13297 8984 13654
rect 9324 13530 9352 15422
rect 9416 15094 9444 15966
rect 9404 15088 9456 15094
rect 9404 15030 9456 15036
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 8942 13288 8998 13297
rect 8942 13223 8998 13232
rect 9310 13288 9366 13297
rect 9310 13223 9366 13232
rect 8956 13084 9252 13104
rect 9012 13082 9036 13084
rect 9092 13082 9116 13084
rect 9172 13082 9196 13084
rect 9034 13030 9036 13082
rect 9098 13030 9110 13082
rect 9172 13030 9174 13082
rect 9012 13028 9036 13030
rect 9092 13028 9116 13030
rect 9172 13028 9196 13030
rect 8956 13008 9252 13028
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 8852 12708 8904 12714
rect 8852 12650 8904 12656
rect 8588 10526 8800 10554
rect 8300 9998 8352 10004
rect 8482 10024 8538 10033
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 8312 9178 8340 9998
rect 8482 9959 8538 9968
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8404 8838 8432 9522
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8208 8560 8260 8566
rect 8206 8528 8208 8537
rect 8260 8528 8262 8537
rect 8206 8463 8262 8472
rect 8404 8362 8432 8774
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8404 7886 8432 8298
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 8128 7342 8156 7686
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 8128 7206 8156 7278
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8024 5840 8076 5846
rect 8024 5782 8076 5788
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 7838 4584 7894 4593
rect 7838 4519 7894 4528
rect 7748 4276 7800 4282
rect 7576 3670 7604 4270
rect 7748 4218 7800 4224
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7564 3664 7616 3670
rect 7564 3606 7616 3612
rect 7668 3602 7696 4082
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7668 3194 7696 3538
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 7852 2258 7880 4519
rect 7944 4486 7972 5646
rect 8036 5370 8064 5782
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 7944 4146 7972 4422
rect 8036 4321 8064 5306
rect 8022 4312 8078 4321
rect 8022 4247 8078 4256
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 7944 4010 7972 4082
rect 7932 4004 7984 4010
rect 7932 3946 7984 3952
rect 7932 3664 7984 3670
rect 7932 3606 7984 3612
rect 7944 3194 7972 3606
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 8128 2990 8156 7142
rect 8496 6746 8524 9862
rect 8588 7313 8616 10526
rect 8758 10432 8814 10441
rect 8758 10367 8814 10376
rect 8668 9444 8720 9450
rect 8668 9386 8720 9392
rect 8680 7546 8708 9386
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8574 7304 8630 7313
rect 8574 7239 8630 7248
rect 8680 6934 8708 7482
rect 8668 6928 8720 6934
rect 8668 6870 8720 6876
rect 8496 6718 8708 6746
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8312 5914 8340 6598
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8220 3942 8248 5510
rect 8312 5370 8340 5850
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8312 4214 8340 4966
rect 8300 4208 8352 4214
rect 8300 4150 8352 4156
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 8220 2650 8248 3878
rect 8312 3097 8340 4150
rect 8404 4078 8432 6054
rect 8392 4072 8444 4078
rect 8496 4049 8524 6054
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8588 5166 8616 5850
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 8588 4865 8616 5102
rect 8574 4856 8630 4865
rect 8574 4791 8630 4800
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8588 4185 8616 4422
rect 8574 4176 8630 4185
rect 8574 4111 8630 4120
rect 8392 4014 8444 4020
rect 8482 4040 8538 4049
rect 8404 3738 8432 4014
rect 8482 3975 8538 3984
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8392 3460 8444 3466
rect 8392 3402 8444 3408
rect 8298 3088 8354 3097
rect 8298 3023 8354 3032
rect 8404 2922 8432 3402
rect 8300 2916 8352 2922
rect 8300 2858 8352 2864
rect 8392 2916 8444 2922
rect 8392 2858 8444 2864
rect 8576 2916 8628 2922
rect 8576 2858 8628 2864
rect 8312 2825 8340 2858
rect 8298 2816 8354 2825
rect 8298 2751 8354 2760
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 8024 2508 8076 2514
rect 8024 2450 8076 2456
rect 8036 2281 8064 2450
rect 8404 2378 8432 2858
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 7760 2230 7880 2258
rect 8022 2272 8078 2281
rect 7760 480 7788 2230
rect 8078 2230 8248 2258
rect 8022 2207 8078 2216
rect 8220 480 8248 2230
rect 8588 480 8616 2858
rect 8680 2650 8708 6718
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 8772 2582 8800 10367
rect 8864 4690 8892 12650
rect 9048 12442 9076 12718
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 8956 11996 9252 12016
rect 9012 11994 9036 11996
rect 9092 11994 9116 11996
rect 9172 11994 9196 11996
rect 9034 11942 9036 11994
rect 9098 11942 9110 11994
rect 9172 11942 9174 11994
rect 9012 11940 9036 11942
rect 9092 11940 9116 11942
rect 9172 11940 9196 11942
rect 8956 11920 9252 11940
rect 9324 11150 9352 13223
rect 9416 11354 9444 15030
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9402 11248 9458 11257
rect 9402 11183 9404 11192
rect 9456 11183 9458 11192
rect 9404 11154 9456 11160
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 8956 10908 9252 10928
rect 9012 10906 9036 10908
rect 9092 10906 9116 10908
rect 9172 10906 9196 10908
rect 9034 10854 9036 10906
rect 9098 10854 9110 10906
rect 9172 10854 9174 10906
rect 9012 10852 9036 10854
rect 9092 10852 9116 10854
rect 9172 10852 9196 10854
rect 8956 10832 9252 10852
rect 9312 9988 9364 9994
rect 9312 9930 9364 9936
rect 8956 9820 9252 9840
rect 9012 9818 9036 9820
rect 9092 9818 9116 9820
rect 9172 9818 9196 9820
rect 9034 9766 9036 9818
rect 9098 9766 9110 9818
rect 9172 9766 9174 9818
rect 9012 9764 9036 9766
rect 9092 9764 9116 9766
rect 9172 9764 9196 9766
rect 8956 9744 9252 9764
rect 8956 8732 9252 8752
rect 9012 8730 9036 8732
rect 9092 8730 9116 8732
rect 9172 8730 9196 8732
rect 9034 8678 9036 8730
rect 9098 8678 9110 8730
rect 9172 8678 9174 8730
rect 9012 8676 9036 8678
rect 9092 8676 9116 8678
rect 9172 8676 9196 8678
rect 8956 8656 9252 8676
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 9048 7886 9076 8366
rect 9324 8265 9352 9930
rect 9416 9926 9444 11154
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9404 9716 9456 9722
rect 9404 9658 9456 9664
rect 9310 8256 9366 8265
rect 9310 8191 9366 8200
rect 9310 8120 9366 8129
rect 9310 8055 9366 8064
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 8956 7644 9252 7664
rect 9012 7642 9036 7644
rect 9092 7642 9116 7644
rect 9172 7642 9196 7644
rect 9034 7590 9036 7642
rect 9098 7590 9110 7642
rect 9172 7590 9174 7642
rect 9012 7588 9036 7590
rect 9092 7588 9116 7590
rect 9172 7588 9196 7590
rect 8956 7568 9252 7588
rect 8956 6556 9252 6576
rect 9012 6554 9036 6556
rect 9092 6554 9116 6556
rect 9172 6554 9196 6556
rect 9034 6502 9036 6554
rect 9098 6502 9110 6554
rect 9172 6502 9174 6554
rect 9012 6500 9036 6502
rect 9092 6500 9116 6502
rect 9172 6500 9196 6502
rect 8956 6480 9252 6500
rect 9324 6440 9352 8055
rect 9048 6412 9352 6440
rect 9048 5914 9076 6412
rect 9416 6361 9444 9658
rect 9508 6458 9536 27118
rect 9588 26240 9640 26246
rect 9588 26182 9640 26188
rect 9600 25770 9628 26182
rect 9772 25900 9824 25906
rect 9772 25842 9824 25848
rect 9588 25764 9640 25770
rect 9640 25724 9720 25752
rect 9588 25706 9640 25712
rect 9692 24410 9720 25724
rect 9784 24954 9812 25842
rect 9876 24993 9904 29022
rect 9954 27432 10010 27441
rect 9954 27367 10010 27376
rect 9968 26364 9996 27367
rect 10060 26466 10088 35430
rect 10140 34944 10192 34950
rect 10140 34886 10192 34892
rect 10232 34944 10284 34950
rect 10232 34886 10284 34892
rect 10152 31890 10180 34886
rect 10244 34474 10272 34886
rect 10232 34468 10284 34474
rect 10232 34410 10284 34416
rect 10244 32910 10272 34410
rect 10322 34096 10378 34105
rect 10322 34031 10378 34040
rect 10232 32904 10284 32910
rect 10232 32846 10284 32852
rect 10336 32314 10364 34031
rect 10244 32286 10364 32314
rect 10244 32065 10272 32286
rect 10324 32224 10376 32230
rect 10324 32166 10376 32172
rect 10230 32056 10286 32065
rect 10336 32026 10364 32166
rect 10230 31991 10286 32000
rect 10324 32020 10376 32026
rect 10324 31962 10376 31968
rect 10232 31952 10284 31958
rect 10232 31894 10284 31900
rect 10140 31884 10192 31890
rect 10140 31826 10192 31832
rect 10152 30938 10180 31826
rect 10244 31142 10272 31894
rect 10324 31816 10376 31822
rect 10324 31758 10376 31764
rect 10336 31482 10364 31758
rect 10324 31476 10376 31482
rect 10324 31418 10376 31424
rect 10232 31136 10284 31142
rect 10232 31078 10284 31084
rect 10244 30977 10272 31078
rect 10230 30968 10286 30977
rect 10140 30932 10192 30938
rect 10230 30903 10286 30912
rect 10140 30874 10192 30880
rect 10428 30818 10456 35686
rect 10600 35284 10652 35290
rect 10600 35226 10652 35232
rect 10506 34504 10562 34513
rect 10506 34439 10562 34448
rect 10520 33153 10548 34439
rect 10506 33144 10562 33153
rect 10506 33079 10562 33088
rect 10508 32972 10560 32978
rect 10508 32914 10560 32920
rect 10520 32434 10548 32914
rect 10508 32428 10560 32434
rect 10508 32370 10560 32376
rect 10520 32026 10548 32370
rect 10508 32020 10560 32026
rect 10508 31962 10560 31968
rect 10506 31920 10562 31929
rect 10506 31855 10562 31864
rect 10244 30790 10456 30818
rect 10244 30297 10272 30790
rect 10520 30682 10548 31855
rect 10428 30654 10548 30682
rect 10324 30388 10376 30394
rect 10324 30330 10376 30336
rect 10230 30288 10286 30297
rect 10230 30223 10286 30232
rect 10232 29708 10284 29714
rect 10232 29650 10284 29656
rect 10244 28694 10272 29650
rect 10232 28688 10284 28694
rect 10232 28630 10284 28636
rect 10244 27334 10272 28630
rect 10232 27328 10284 27334
rect 10232 27270 10284 27276
rect 10140 26784 10192 26790
rect 10140 26726 10192 26732
rect 10152 26586 10180 26726
rect 10140 26580 10192 26586
rect 10140 26522 10192 26528
rect 10060 26438 10180 26466
rect 9968 26336 10088 26364
rect 9956 25696 10008 25702
rect 9956 25638 10008 25644
rect 9968 25430 9996 25638
rect 9956 25424 10008 25430
rect 9954 25392 9956 25401
rect 10008 25392 10010 25401
rect 9954 25327 10010 25336
rect 9862 24984 9918 24993
rect 9772 24948 9824 24954
rect 9862 24919 9918 24928
rect 9772 24890 9824 24896
rect 9784 24614 9812 24890
rect 9772 24608 9824 24614
rect 9772 24550 9824 24556
rect 9680 24404 9732 24410
rect 9680 24346 9732 24352
rect 9956 24200 10008 24206
rect 9956 24142 10008 24148
rect 9864 23724 9916 23730
rect 9864 23666 9916 23672
rect 9876 23322 9904 23666
rect 9968 23526 9996 24142
rect 9956 23520 10008 23526
rect 9956 23462 10008 23468
rect 9864 23316 9916 23322
rect 9864 23258 9916 23264
rect 9968 23202 9996 23462
rect 9876 23174 9996 23202
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9600 20448 9628 20742
rect 9772 20596 9824 20602
rect 9772 20538 9824 20544
rect 9784 20482 9812 20538
rect 9692 20454 9812 20482
rect 9692 20448 9720 20454
rect 9600 20420 9720 20448
rect 9876 20398 9904 23174
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9968 21078 9996 21830
rect 9956 21072 10008 21078
rect 9956 21014 10008 21020
rect 9968 20466 9996 21014
rect 9956 20460 10008 20466
rect 9956 20402 10008 20408
rect 9864 20392 9916 20398
rect 9678 20360 9734 20369
rect 9864 20334 9916 20340
rect 9678 20295 9734 20304
rect 9772 20324 9824 20330
rect 9692 20262 9720 20295
rect 9772 20266 9824 20272
rect 9680 20256 9732 20262
rect 9680 20198 9732 20204
rect 9678 19816 9734 19825
rect 9678 19751 9734 19760
rect 9692 18970 9720 19751
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9784 18850 9812 20266
rect 9956 19848 10008 19854
rect 9956 19790 10008 19796
rect 9692 18822 9812 18850
rect 9864 18828 9916 18834
rect 9692 17785 9720 18822
rect 9864 18770 9916 18776
rect 9772 18216 9824 18222
rect 9772 18158 9824 18164
rect 9678 17776 9734 17785
rect 9678 17711 9734 17720
rect 9692 16998 9720 17711
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9692 14618 9720 16934
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9692 13682 9720 13874
rect 9600 13654 9720 13682
rect 9600 12782 9628 13654
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9692 13433 9720 13466
rect 9678 13424 9734 13433
rect 9678 13359 9734 13368
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9600 12209 9628 12718
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9692 12238 9720 12582
rect 9680 12232 9732 12238
rect 9586 12200 9642 12209
rect 9680 12174 9732 12180
rect 9586 12135 9642 12144
rect 9600 11354 9628 12135
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9588 11348 9640 11354
rect 9588 11290 9640 11296
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9600 10266 9628 10950
rect 9692 10713 9720 12038
rect 9784 11354 9812 18158
rect 9876 18086 9904 18770
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9678 10704 9734 10713
rect 9678 10639 9734 10648
rect 9692 10606 9720 10639
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9680 10464 9732 10470
rect 9678 10432 9680 10441
rect 9784 10452 9812 11086
rect 9732 10432 9812 10452
rect 9734 10424 9812 10432
rect 9678 10367 9734 10376
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9692 9364 9720 9522
rect 9600 9336 9720 9364
rect 9600 8945 9628 9336
rect 9586 8936 9642 8945
rect 9586 8871 9642 8880
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9402 6352 9458 6361
rect 9600 6338 9628 8871
rect 9876 7857 9904 18022
rect 9968 17105 9996 19790
rect 10060 18834 10088 26336
rect 10152 19122 10180 26438
rect 10244 26042 10272 27270
rect 10336 26518 10364 30330
rect 10324 26512 10376 26518
rect 10324 26454 10376 26460
rect 10428 26450 10456 30654
rect 10508 30592 10560 30598
rect 10508 30534 10560 30540
rect 10416 26444 10468 26450
rect 10416 26386 10468 26392
rect 10232 26036 10284 26042
rect 10232 25978 10284 25984
rect 10244 25362 10272 25978
rect 10428 25838 10456 26386
rect 10520 25838 10548 30534
rect 10416 25832 10468 25838
rect 10416 25774 10468 25780
rect 10508 25832 10560 25838
rect 10508 25774 10560 25780
rect 10232 25356 10284 25362
rect 10232 25298 10284 25304
rect 10324 25288 10376 25294
rect 10324 25230 10376 25236
rect 10336 24818 10364 25230
rect 10324 24812 10376 24818
rect 10324 24754 10376 24760
rect 10336 24206 10364 24754
rect 10428 24274 10456 25774
rect 10520 25498 10548 25774
rect 10612 25770 10640 35226
rect 10784 34060 10836 34066
rect 10784 34002 10836 34008
rect 10692 33924 10744 33930
rect 10692 33866 10744 33872
rect 10704 33318 10732 33866
rect 10796 33862 10824 34002
rect 10876 33992 10928 33998
rect 10876 33934 10928 33940
rect 10784 33856 10836 33862
rect 10784 33798 10836 33804
rect 10692 33312 10744 33318
rect 10692 33254 10744 33260
rect 10690 33144 10746 33153
rect 10796 33114 10824 33798
rect 10888 33590 10916 33934
rect 10876 33584 10928 33590
rect 10876 33526 10928 33532
rect 10876 33312 10928 33318
rect 10876 33254 10928 33260
rect 10888 33114 10916 33254
rect 10690 33079 10746 33088
rect 10784 33108 10836 33114
rect 10704 32994 10732 33079
rect 10784 33050 10836 33056
rect 10876 33108 10928 33114
rect 10876 33050 10928 33056
rect 10704 32966 10824 32994
rect 10690 32736 10746 32745
rect 10690 32671 10746 32680
rect 10704 30394 10732 32671
rect 10796 30598 10824 32966
rect 11072 31668 11100 39494
rect 11152 37732 11204 37738
rect 11152 37674 11204 37680
rect 10980 31640 11100 31668
rect 10784 30592 10836 30598
rect 10784 30534 10836 30540
rect 10692 30388 10744 30394
rect 10692 30330 10744 30336
rect 10784 30320 10836 30326
rect 10782 30288 10784 30297
rect 10836 30288 10838 30297
rect 10692 30252 10744 30258
rect 10782 30223 10838 30232
rect 10692 30194 10744 30200
rect 10704 28150 10732 30194
rect 10782 29744 10838 29753
rect 10782 29679 10838 29688
rect 10796 28218 10824 29679
rect 10980 29306 11008 31640
rect 11164 31113 11192 37674
rect 11244 33448 11296 33454
rect 11244 33390 11296 33396
rect 11256 33289 11284 33390
rect 11242 33280 11298 33289
rect 11242 33215 11298 33224
rect 11150 31104 11206 31113
rect 11150 31039 11206 31048
rect 11164 30433 11192 31039
rect 11244 30592 11296 30598
rect 11244 30534 11296 30540
rect 11150 30424 11206 30433
rect 11150 30359 11206 30368
rect 11256 30190 11284 30534
rect 11244 30184 11296 30190
rect 11244 30126 11296 30132
rect 11152 30048 11204 30054
rect 11152 29990 11204 29996
rect 10968 29300 11020 29306
rect 10968 29242 11020 29248
rect 11058 29064 11114 29073
rect 11058 28999 11114 29008
rect 10968 28960 11020 28966
rect 10968 28902 11020 28908
rect 10784 28212 10836 28218
rect 10784 28154 10836 28160
rect 10692 28144 10744 28150
rect 10692 28086 10744 28092
rect 10692 27328 10744 27334
rect 10692 27270 10744 27276
rect 10704 26790 10732 27270
rect 10692 26784 10744 26790
rect 10692 26726 10744 26732
rect 10704 26042 10732 26726
rect 10784 26512 10836 26518
rect 10784 26454 10836 26460
rect 10796 26042 10824 26454
rect 10692 26036 10744 26042
rect 10692 25978 10744 25984
rect 10784 26036 10836 26042
rect 10784 25978 10836 25984
rect 10600 25764 10652 25770
rect 10600 25706 10652 25712
rect 10508 25492 10560 25498
rect 10508 25434 10560 25440
rect 10520 24954 10548 25434
rect 10508 24948 10560 24954
rect 10508 24890 10560 24896
rect 10692 24948 10744 24954
rect 10692 24890 10744 24896
rect 10598 24304 10654 24313
rect 10416 24268 10468 24274
rect 10598 24239 10654 24248
rect 10416 24210 10468 24216
rect 10324 24200 10376 24206
rect 10324 24142 10376 24148
rect 10336 23730 10364 24142
rect 10508 23860 10560 23866
rect 10508 23802 10560 23808
rect 10324 23724 10376 23730
rect 10324 23666 10376 23672
rect 10232 22432 10284 22438
rect 10232 22374 10284 22380
rect 10244 22030 10272 22374
rect 10324 22092 10376 22098
rect 10324 22034 10376 22040
rect 10232 22024 10284 22030
rect 10232 21966 10284 21972
rect 10244 21350 10272 21966
rect 10336 21690 10364 22034
rect 10324 21684 10376 21690
rect 10324 21626 10376 21632
rect 10232 21344 10284 21350
rect 10232 21286 10284 21292
rect 10244 21010 10272 21286
rect 10232 21004 10284 21010
rect 10232 20946 10284 20952
rect 10232 20596 10284 20602
rect 10232 20538 10284 20544
rect 10244 20398 10272 20538
rect 10232 20392 10284 20398
rect 10232 20334 10284 20340
rect 10336 20346 10364 21626
rect 10244 19786 10272 20334
rect 10336 20318 10456 20346
rect 10324 20256 10376 20262
rect 10324 20198 10376 20204
rect 10336 20058 10364 20198
rect 10324 20052 10376 20058
rect 10324 19994 10376 20000
rect 10232 19780 10284 19786
rect 10232 19722 10284 19728
rect 10336 19514 10364 19994
rect 10324 19508 10376 19514
rect 10324 19450 10376 19456
rect 10428 19446 10456 20318
rect 10520 19854 10548 23802
rect 10508 19848 10560 19854
rect 10508 19790 10560 19796
rect 10508 19712 10560 19718
rect 10508 19654 10560 19660
rect 10416 19440 10468 19446
rect 10416 19382 10468 19388
rect 10416 19304 10468 19310
rect 10416 19246 10468 19252
rect 10152 19094 10364 19122
rect 10140 18964 10192 18970
rect 10140 18906 10192 18912
rect 10048 18828 10100 18834
rect 10048 18770 10100 18776
rect 10152 18426 10180 18906
rect 10232 18896 10284 18902
rect 10232 18838 10284 18844
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 10244 18306 10272 18838
rect 10152 18278 10272 18306
rect 9954 17096 10010 17105
rect 10010 17054 10088 17082
rect 9954 17031 10010 17040
rect 10060 16998 10088 17054
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 9968 15706 9996 16934
rect 10060 16794 10088 16934
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 9968 15162 9996 15438
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 10152 14958 10180 18278
rect 10336 18222 10364 19094
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10232 18148 10284 18154
rect 10232 18090 10284 18096
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 10152 14618 10180 14894
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 9968 10198 9996 14554
rect 10140 13728 10192 13734
rect 10060 13676 10140 13682
rect 10060 13670 10192 13676
rect 10060 13654 10180 13670
rect 10060 13394 10088 13654
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 10060 12442 10088 13330
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10152 12986 10180 13262
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 10244 12481 10272 18090
rect 10324 18080 10376 18086
rect 10324 18022 10376 18028
rect 10336 17882 10364 18022
rect 10324 17876 10376 17882
rect 10324 17818 10376 17824
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 10336 16726 10364 17614
rect 10428 17610 10456 19246
rect 10520 19174 10548 19654
rect 10508 19168 10560 19174
rect 10508 19110 10560 19116
rect 10416 17604 10468 17610
rect 10416 17546 10468 17552
rect 10324 16720 10376 16726
rect 10324 16662 10376 16668
rect 10336 16454 10364 16662
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10336 15434 10364 16390
rect 10324 15428 10376 15434
rect 10324 15370 10376 15376
rect 10336 14550 10364 15370
rect 10520 15366 10548 19110
rect 10612 18834 10640 24239
rect 10704 18902 10732 24890
rect 10796 24342 10824 25978
rect 10980 25974 11008 28902
rect 11072 26382 11100 28999
rect 11164 28762 11192 29990
rect 11256 29306 11284 30126
rect 11244 29300 11296 29306
rect 11244 29242 11296 29248
rect 11244 29164 11296 29170
rect 11244 29106 11296 29112
rect 11256 29073 11284 29106
rect 11242 29064 11298 29073
rect 11242 28999 11298 29008
rect 11152 28756 11204 28762
rect 11152 28698 11204 28704
rect 11348 28257 11376 39520
rect 11808 37738 11836 39520
rect 11796 37732 11848 37738
rect 11796 37674 11848 37680
rect 11622 37564 11918 37584
rect 11678 37562 11702 37564
rect 11758 37562 11782 37564
rect 11838 37562 11862 37564
rect 11700 37510 11702 37562
rect 11764 37510 11776 37562
rect 11838 37510 11840 37562
rect 11678 37508 11702 37510
rect 11758 37508 11782 37510
rect 11838 37508 11862 37510
rect 11622 37488 11918 37508
rect 11622 36476 11918 36496
rect 11678 36474 11702 36476
rect 11758 36474 11782 36476
rect 11838 36474 11862 36476
rect 11700 36422 11702 36474
rect 11764 36422 11776 36474
rect 11838 36422 11840 36474
rect 11678 36420 11702 36422
rect 11758 36420 11782 36422
rect 11838 36420 11862 36422
rect 11622 36400 11918 36420
rect 12176 35714 12204 39520
rect 12176 35686 12480 35714
rect 11622 35388 11918 35408
rect 11678 35386 11702 35388
rect 11758 35386 11782 35388
rect 11838 35386 11862 35388
rect 11700 35334 11702 35386
rect 11764 35334 11776 35386
rect 11838 35334 11840 35386
rect 11678 35332 11702 35334
rect 11758 35332 11782 35334
rect 11838 35332 11862 35334
rect 11622 35312 11918 35332
rect 12164 34400 12216 34406
rect 12164 34342 12216 34348
rect 11622 34300 11918 34320
rect 11678 34298 11702 34300
rect 11758 34298 11782 34300
rect 11838 34298 11862 34300
rect 11700 34246 11702 34298
rect 11764 34246 11776 34298
rect 11838 34246 11840 34298
rect 11678 34244 11702 34246
rect 11758 34244 11782 34246
rect 11838 34244 11862 34246
rect 11622 34224 11918 34244
rect 11428 33992 11480 33998
rect 11428 33934 11480 33940
rect 11440 33318 11468 33934
rect 12176 33810 12204 34342
rect 12452 34134 12480 35686
rect 12440 34128 12492 34134
rect 12254 34096 12310 34105
rect 12440 34070 12492 34076
rect 12254 34031 12310 34040
rect 12348 34060 12400 34066
rect 12268 33998 12296 34031
rect 12348 34002 12400 34008
rect 12256 33992 12308 33998
rect 12256 33934 12308 33940
rect 12256 33856 12308 33862
rect 12176 33804 12256 33810
rect 12176 33798 12308 33804
rect 12176 33782 12296 33798
rect 11428 33312 11480 33318
rect 11428 33254 11480 33260
rect 11334 28248 11390 28257
rect 11334 28183 11390 28192
rect 11440 28098 11468 33254
rect 11622 33212 11918 33232
rect 11678 33210 11702 33212
rect 11758 33210 11782 33212
rect 11838 33210 11862 33212
rect 11700 33158 11702 33210
rect 11764 33158 11776 33210
rect 11838 33158 11840 33210
rect 11678 33156 11702 33158
rect 11758 33156 11782 33158
rect 11838 33156 11862 33158
rect 11622 33136 11918 33156
rect 12268 32978 12296 33782
rect 12360 33386 12388 34002
rect 12438 33960 12494 33969
rect 12438 33895 12494 33904
rect 12348 33380 12400 33386
rect 12348 33322 12400 33328
rect 12360 33114 12388 33322
rect 12348 33108 12400 33114
rect 12452 33096 12480 33895
rect 12544 33266 12572 39520
rect 13004 35057 13032 39520
rect 12990 35048 13046 35057
rect 12990 34983 13046 34992
rect 12716 34128 12768 34134
rect 12716 34070 12768 34076
rect 12728 33386 12756 34070
rect 12900 33516 12952 33522
rect 12900 33458 12952 33464
rect 12716 33380 12768 33386
rect 12716 33322 12768 33328
rect 12544 33238 12664 33266
rect 12452 33068 12572 33096
rect 12348 33050 12400 33056
rect 12256 32972 12308 32978
rect 12256 32914 12308 32920
rect 11520 32768 11572 32774
rect 11520 32710 11572 32716
rect 11532 31686 11560 32710
rect 12268 32570 12296 32914
rect 12256 32564 12308 32570
rect 12256 32506 12308 32512
rect 11622 32124 11918 32144
rect 11678 32122 11702 32124
rect 11758 32122 11782 32124
rect 11838 32122 11862 32124
rect 11700 32070 11702 32122
rect 11764 32070 11776 32122
rect 11838 32070 11840 32122
rect 11678 32068 11702 32070
rect 11758 32068 11782 32070
rect 11838 32068 11862 32070
rect 11622 32048 11918 32068
rect 11520 31680 11572 31686
rect 11520 31622 11572 31628
rect 11532 30598 11560 31622
rect 11622 31036 11918 31056
rect 11678 31034 11702 31036
rect 11758 31034 11782 31036
rect 11838 31034 11862 31036
rect 11700 30982 11702 31034
rect 11764 30982 11776 31034
rect 11838 30982 11840 31034
rect 11678 30980 11702 30982
rect 11758 30980 11782 30982
rect 11838 30980 11862 30982
rect 11622 30960 11918 30980
rect 11980 30796 12032 30802
rect 11980 30738 12032 30744
rect 11520 30592 11572 30598
rect 11520 30534 11572 30540
rect 11532 29646 11560 30534
rect 11992 30054 12020 30738
rect 12440 30592 12492 30598
rect 12440 30534 12492 30540
rect 12254 30424 12310 30433
rect 12254 30359 12310 30368
rect 11980 30048 12032 30054
rect 11980 29990 12032 29996
rect 11622 29948 11918 29968
rect 11678 29946 11702 29948
rect 11758 29946 11782 29948
rect 11838 29946 11862 29948
rect 11700 29894 11702 29946
rect 11764 29894 11776 29946
rect 11838 29894 11840 29946
rect 11678 29892 11702 29894
rect 11758 29892 11782 29894
rect 11838 29892 11862 29894
rect 11622 29872 11918 29892
rect 11520 29640 11572 29646
rect 11520 29582 11572 29588
rect 11886 29608 11942 29617
rect 11886 29543 11942 29552
rect 11900 29238 11928 29543
rect 11888 29232 11940 29238
rect 11888 29174 11940 29180
rect 11992 29170 12020 29990
rect 11980 29164 12032 29170
rect 11980 29106 12032 29112
rect 11520 29028 11572 29034
rect 11520 28970 11572 28976
rect 11532 28665 11560 28970
rect 11622 28860 11918 28880
rect 11678 28858 11702 28860
rect 11758 28858 11782 28860
rect 11838 28858 11862 28860
rect 11700 28806 11702 28858
rect 11764 28806 11776 28858
rect 11838 28806 11840 28858
rect 11678 28804 11702 28806
rect 11758 28804 11782 28806
rect 11838 28804 11862 28806
rect 11622 28784 11918 28804
rect 11518 28656 11574 28665
rect 11518 28591 11574 28600
rect 11992 28558 12020 29106
rect 12164 29028 12216 29034
rect 12164 28970 12216 28976
rect 12070 28792 12126 28801
rect 12070 28727 12072 28736
rect 12124 28727 12126 28736
rect 12072 28698 12124 28704
rect 11980 28552 12032 28558
rect 11980 28494 12032 28500
rect 12084 28218 12112 28698
rect 12072 28212 12124 28218
rect 12072 28154 12124 28160
rect 11348 28070 11468 28098
rect 12072 28076 12124 28082
rect 11244 27872 11296 27878
rect 11244 27814 11296 27820
rect 11150 27704 11206 27713
rect 11256 27674 11284 27814
rect 11150 27639 11206 27648
rect 11244 27668 11296 27674
rect 11164 26450 11192 27639
rect 11244 27610 11296 27616
rect 11256 27130 11284 27610
rect 11244 27124 11296 27130
rect 11244 27066 11296 27072
rect 11152 26444 11204 26450
rect 11152 26386 11204 26392
rect 11060 26376 11112 26382
rect 11060 26318 11112 26324
rect 10968 25968 11020 25974
rect 10968 25910 11020 25916
rect 11072 25906 11100 26318
rect 11152 25968 11204 25974
rect 11152 25910 11204 25916
rect 11060 25900 11112 25906
rect 11060 25842 11112 25848
rect 10968 25764 11020 25770
rect 10968 25706 11020 25712
rect 10784 24336 10836 24342
rect 10784 24278 10836 24284
rect 10796 23866 10824 24278
rect 10784 23860 10836 23866
rect 10784 23802 10836 23808
rect 10784 23724 10836 23730
rect 10784 23666 10836 23672
rect 10692 18896 10744 18902
rect 10692 18838 10744 18844
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10600 18692 10652 18698
rect 10600 18634 10652 18640
rect 10612 18290 10640 18634
rect 10692 18624 10744 18630
rect 10796 18612 10824 23666
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 10888 19990 10916 20402
rect 10876 19984 10928 19990
rect 10876 19926 10928 19932
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10888 19310 10916 19654
rect 10876 19304 10928 19310
rect 10876 19246 10928 19252
rect 10876 18828 10928 18834
rect 10876 18770 10928 18776
rect 10744 18584 10824 18612
rect 10692 18566 10744 18572
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 10612 17542 10640 18226
rect 10704 18154 10732 18566
rect 10692 18148 10744 18154
rect 10692 18090 10744 18096
rect 10784 17876 10836 17882
rect 10784 17818 10836 17824
rect 10600 17536 10652 17542
rect 10600 17478 10652 17484
rect 10612 17202 10640 17478
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10612 16658 10640 17138
rect 10796 16794 10824 17818
rect 10888 17746 10916 18770
rect 10876 17740 10928 17746
rect 10876 17682 10928 17688
rect 10888 17338 10916 17682
rect 10876 17332 10928 17338
rect 10876 17274 10928 17280
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10600 16652 10652 16658
rect 10600 16594 10652 16600
rect 10612 15910 10640 16594
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10782 15872 10838 15881
rect 10508 15360 10560 15366
rect 10508 15302 10560 15308
rect 10612 15026 10640 15846
rect 10782 15807 10838 15816
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10324 14544 10376 14550
rect 10324 14486 10376 14492
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10336 12646 10364 13262
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10230 12472 10286 12481
rect 10048 12436 10100 12442
rect 10230 12407 10286 12416
rect 10048 12378 10100 12384
rect 10416 12368 10468 12374
rect 10046 12336 10102 12345
rect 10046 12271 10102 12280
rect 10230 12336 10286 12345
rect 10416 12310 10468 12316
rect 10230 12271 10286 12280
rect 10060 11762 10088 12271
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 10060 11529 10088 11698
rect 10140 11552 10192 11558
rect 10046 11520 10102 11529
rect 10140 11494 10192 11500
rect 10046 11455 10102 11464
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9956 10056 10008 10062
rect 9956 9998 10008 10004
rect 9968 9110 9996 9998
rect 9956 9104 10008 9110
rect 9956 9046 10008 9052
rect 9954 8392 10010 8401
rect 9954 8327 10010 8336
rect 9862 7848 9918 7857
rect 9862 7783 9918 7792
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9692 6730 9720 7142
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9402 6287 9458 6296
rect 9508 6310 9628 6338
rect 9692 6322 9720 6666
rect 9784 6458 9812 6802
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9680 6316 9732 6322
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 9310 5808 9366 5817
rect 9310 5743 9366 5752
rect 8956 5468 9252 5488
rect 9012 5466 9036 5468
rect 9092 5466 9116 5468
rect 9172 5466 9196 5468
rect 9034 5414 9036 5466
rect 9098 5414 9110 5466
rect 9172 5414 9174 5466
rect 9012 5412 9036 5414
rect 9092 5412 9116 5414
rect 9172 5412 9196 5414
rect 8956 5392 9252 5412
rect 9324 5234 9352 5743
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9324 4826 9352 5170
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 8864 4282 8892 4626
rect 8956 4380 9252 4400
rect 9012 4378 9036 4380
rect 9092 4378 9116 4380
rect 9172 4378 9196 4380
rect 9034 4326 9036 4378
rect 9098 4326 9110 4378
rect 9172 4326 9174 4378
rect 9012 4324 9036 4326
rect 9092 4324 9116 4326
rect 9172 4324 9196 4326
rect 8956 4304 9252 4324
rect 8852 4276 8904 4282
rect 8852 4218 8904 4224
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8864 3194 8892 4082
rect 9324 3738 9352 4762
rect 9416 4146 9444 6122
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 8956 3292 9252 3312
rect 9012 3290 9036 3292
rect 9092 3290 9116 3292
rect 9172 3290 9196 3292
rect 9034 3238 9036 3290
rect 9098 3238 9110 3290
rect 9172 3238 9174 3290
rect 9012 3236 9036 3238
rect 9092 3236 9116 3238
rect 9172 3236 9196 3238
rect 8956 3216 9252 3236
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8760 2576 8812 2582
rect 8760 2518 8812 2524
rect 8864 1986 8892 2926
rect 9508 2854 9536 6310
rect 9680 6258 9732 6264
rect 9772 5840 9824 5846
rect 9772 5782 9824 5788
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9600 4808 9628 5510
rect 9784 5370 9812 5782
rect 9876 5681 9904 6598
rect 9862 5672 9918 5681
rect 9862 5607 9918 5616
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9680 4820 9732 4826
rect 9600 4780 9680 4808
rect 9680 4762 9732 4768
rect 9784 4690 9812 5306
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9600 4010 9628 4422
rect 9784 4282 9812 4626
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9588 4004 9640 4010
rect 9588 3946 9640 3952
rect 9770 3088 9826 3097
rect 9770 3023 9826 3032
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9494 2680 9550 2689
rect 9494 2615 9550 2624
rect 9508 2582 9536 2615
rect 9496 2576 9548 2582
rect 9496 2518 9548 2524
rect 9692 2514 9720 2790
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 8956 2204 9252 2224
rect 9012 2202 9036 2204
rect 9092 2202 9116 2204
rect 9172 2202 9196 2204
rect 9034 2150 9036 2202
rect 9098 2150 9110 2202
rect 9172 2150 9174 2202
rect 9012 2148 9036 2150
rect 9092 2148 9116 2150
rect 9172 2148 9196 2150
rect 8956 2128 9252 2148
rect 8864 1958 8984 1986
rect 8956 480 8984 1958
rect 9416 480 9444 2450
rect 9784 480 9812 3023
rect 9876 610 9904 5306
rect 9968 4554 9996 8327
rect 9956 4548 10008 4554
rect 9956 4490 10008 4496
rect 10060 3670 10088 11290
rect 10152 11286 10180 11494
rect 10140 11280 10192 11286
rect 10140 11222 10192 11228
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10152 9586 10180 10066
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10138 7440 10194 7449
rect 10138 7375 10194 7384
rect 10152 5370 10180 7375
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 10152 4282 10180 4558
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 10048 3664 10100 3670
rect 10048 3606 10100 3612
rect 10060 3194 10088 3606
rect 10152 3194 10180 4014
rect 10244 3534 10272 12271
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 10336 11694 10364 12106
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10336 10062 10364 11494
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10322 8256 10378 8265
rect 10322 8191 10378 8200
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 10048 3188 10100 3194
rect 9968 3148 10048 3176
rect 9968 678 9996 3148
rect 10048 3130 10100 3136
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10244 3097 10272 3470
rect 10230 3088 10286 3097
rect 10230 3023 10286 3032
rect 10336 2972 10364 8191
rect 10428 8129 10456 12310
rect 10520 12102 10548 14554
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10508 11824 10560 11830
rect 10508 11766 10560 11772
rect 10520 10470 10548 11766
rect 10612 10810 10640 12922
rect 10690 12880 10746 12889
rect 10690 12815 10746 12824
rect 10600 10804 10652 10810
rect 10600 10746 10652 10752
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10520 10198 10548 10406
rect 10612 10266 10640 10406
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10508 10192 10560 10198
rect 10704 10146 10732 12815
rect 10508 10134 10560 10140
rect 10612 10118 10732 10146
rect 10506 10024 10562 10033
rect 10506 9959 10562 9968
rect 10520 9586 10548 9959
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10414 8120 10470 8129
rect 10414 8055 10470 8064
rect 10520 4078 10548 9522
rect 10612 5370 10640 10118
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10704 9382 10732 9998
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10704 9178 10732 9318
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10796 6866 10824 15807
rect 10980 12374 11008 25706
rect 11072 25498 11100 25842
rect 11060 25492 11112 25498
rect 11060 25434 11112 25440
rect 11164 24018 11192 25910
rect 11244 25696 11296 25702
rect 11244 25638 11296 25644
rect 11256 24410 11284 25638
rect 11244 24404 11296 24410
rect 11244 24346 11296 24352
rect 11072 23990 11192 24018
rect 11072 23730 11100 23990
rect 11152 23860 11204 23866
rect 11152 23802 11204 23808
rect 11060 23724 11112 23730
rect 11060 23666 11112 23672
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 11072 15162 11100 15642
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 10968 12368 11020 12374
rect 10968 12310 11020 12316
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10888 11830 10916 12242
rect 10966 12200 11022 12209
rect 10966 12135 11022 12144
rect 10980 12102 11008 12135
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 10876 11824 10928 11830
rect 10876 11766 10928 11772
rect 10888 8838 10916 11766
rect 10980 10674 11008 12038
rect 11072 11354 11100 13806
rect 11164 11626 11192 23802
rect 11244 21140 11296 21146
rect 11244 21082 11296 21088
rect 11256 18698 11284 21082
rect 11348 21049 11376 28070
rect 12072 28018 12124 28024
rect 11428 27940 11480 27946
rect 11428 27882 11480 27888
rect 11440 27334 11468 27882
rect 11622 27772 11918 27792
rect 11678 27770 11702 27772
rect 11758 27770 11782 27772
rect 11838 27770 11862 27772
rect 11700 27718 11702 27770
rect 11764 27718 11776 27770
rect 11838 27718 11840 27770
rect 11678 27716 11702 27718
rect 11758 27716 11782 27718
rect 11838 27716 11862 27718
rect 11622 27696 11918 27716
rect 12084 27674 12112 28018
rect 12072 27668 12124 27674
rect 12072 27610 12124 27616
rect 11428 27328 11480 27334
rect 11428 27270 11480 27276
rect 11440 26586 11468 27270
rect 11622 26684 11918 26704
rect 11678 26682 11702 26684
rect 11758 26682 11782 26684
rect 11838 26682 11862 26684
rect 11700 26630 11702 26682
rect 11764 26630 11776 26682
rect 11838 26630 11840 26682
rect 11678 26628 11702 26630
rect 11758 26628 11782 26630
rect 11838 26628 11862 26630
rect 11622 26608 11918 26628
rect 11428 26580 11480 26586
rect 11428 26522 11480 26528
rect 11980 26444 12032 26450
rect 11980 26386 12032 26392
rect 11992 26042 12020 26386
rect 11980 26036 12032 26042
rect 11980 25978 12032 25984
rect 11622 25596 11918 25616
rect 11678 25594 11702 25596
rect 11758 25594 11782 25596
rect 11838 25594 11862 25596
rect 11700 25542 11702 25594
rect 11764 25542 11776 25594
rect 11838 25542 11840 25594
rect 11678 25540 11702 25542
rect 11758 25540 11782 25542
rect 11838 25540 11862 25542
rect 11622 25520 11918 25540
rect 11428 25424 11480 25430
rect 11428 25366 11480 25372
rect 11440 24970 11468 25366
rect 11888 25356 11940 25362
rect 11888 25298 11940 25304
rect 11440 24954 11560 24970
rect 11900 24954 11928 25298
rect 11992 24993 12020 25978
rect 11978 24984 12034 24993
rect 11428 24948 11560 24954
rect 11480 24942 11560 24948
rect 11428 24890 11480 24896
rect 11426 24848 11482 24857
rect 11426 24783 11482 24792
rect 11440 24342 11468 24783
rect 11428 24336 11480 24342
rect 11428 24278 11480 24284
rect 11440 23866 11468 24278
rect 11532 24206 11560 24942
rect 11888 24948 11940 24954
rect 11978 24919 12034 24928
rect 11888 24890 11940 24896
rect 11622 24508 11918 24528
rect 11678 24506 11702 24508
rect 11758 24506 11782 24508
rect 11838 24506 11862 24508
rect 11700 24454 11702 24506
rect 11764 24454 11776 24506
rect 11838 24454 11840 24506
rect 11678 24452 11702 24454
rect 11758 24452 11782 24454
rect 11838 24452 11862 24454
rect 11622 24432 11918 24452
rect 11520 24200 11572 24206
rect 11520 24142 11572 24148
rect 11532 23866 11560 24142
rect 11428 23860 11480 23866
rect 11428 23802 11480 23808
rect 11520 23860 11572 23866
rect 11520 23802 11572 23808
rect 11428 23724 11480 23730
rect 11428 23666 11480 23672
rect 11334 21040 11390 21049
rect 11334 20975 11390 20984
rect 11336 20256 11388 20262
rect 11336 20198 11388 20204
rect 11348 19174 11376 20198
rect 11336 19168 11388 19174
rect 11336 19110 11388 19116
rect 11336 18828 11388 18834
rect 11336 18770 11388 18776
rect 11244 18692 11296 18698
rect 11244 18634 11296 18640
rect 11348 18086 11376 18770
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 11348 16561 11376 18022
rect 11334 16552 11390 16561
rect 11334 16487 11390 16496
rect 11336 16448 11388 16454
rect 11336 16390 11388 16396
rect 11348 16250 11376 16390
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 11348 16153 11376 16186
rect 11334 16144 11390 16153
rect 11334 16079 11390 16088
rect 11244 13796 11296 13802
rect 11244 13738 11296 13744
rect 11256 13530 11284 13738
rect 11244 13524 11296 13530
rect 11244 13466 11296 13472
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 11348 12306 11376 12922
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 11242 11792 11298 11801
rect 11348 11762 11376 12242
rect 11242 11727 11298 11736
rect 11336 11756 11388 11762
rect 11152 11620 11204 11626
rect 11152 11562 11204 11568
rect 11150 11520 11206 11529
rect 11150 11455 11206 11464
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 11164 11286 11192 11455
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10968 10532 11020 10538
rect 10968 10474 11020 10480
rect 10980 9994 11008 10474
rect 10968 9988 11020 9994
rect 10968 9930 11020 9936
rect 11164 9722 11192 11222
rect 11256 10033 11284 11727
rect 11336 11698 11388 11704
rect 11440 11506 11468 23666
rect 11622 23420 11918 23440
rect 11678 23418 11702 23420
rect 11758 23418 11782 23420
rect 11838 23418 11862 23420
rect 11700 23366 11702 23418
rect 11764 23366 11776 23418
rect 11838 23366 11840 23418
rect 11678 23364 11702 23366
rect 11758 23364 11782 23366
rect 11838 23364 11862 23366
rect 11622 23344 11918 23364
rect 11622 22332 11918 22352
rect 11678 22330 11702 22332
rect 11758 22330 11782 22332
rect 11838 22330 11862 22332
rect 11700 22278 11702 22330
rect 11764 22278 11776 22330
rect 11838 22278 11840 22330
rect 11678 22276 11702 22278
rect 11758 22276 11782 22278
rect 11838 22276 11862 22278
rect 11622 22256 11918 22276
rect 11980 21344 12032 21350
rect 11980 21286 12032 21292
rect 11622 21244 11918 21264
rect 11678 21242 11702 21244
rect 11758 21242 11782 21244
rect 11838 21242 11862 21244
rect 11700 21190 11702 21242
rect 11764 21190 11776 21242
rect 11838 21190 11840 21242
rect 11678 21188 11702 21190
rect 11758 21188 11782 21190
rect 11838 21188 11862 21190
rect 11622 21168 11918 21188
rect 11992 21010 12020 21286
rect 12072 21072 12124 21078
rect 12072 21014 12124 21020
rect 11980 21004 12032 21010
rect 11980 20946 12032 20952
rect 11622 20156 11918 20176
rect 11678 20154 11702 20156
rect 11758 20154 11782 20156
rect 11838 20154 11862 20156
rect 11700 20102 11702 20154
rect 11764 20102 11776 20154
rect 11838 20102 11840 20154
rect 11678 20100 11702 20102
rect 11758 20100 11782 20102
rect 11838 20100 11862 20102
rect 11622 20080 11918 20100
rect 11888 19984 11940 19990
rect 11794 19952 11850 19961
rect 11992 19972 12020 20946
rect 12084 20398 12112 21014
rect 12072 20392 12124 20398
rect 12072 20334 12124 20340
rect 12176 19990 12204 28970
rect 12268 24410 12296 30359
rect 12452 30326 12480 30534
rect 12440 30320 12492 30326
rect 12440 30262 12492 30268
rect 12452 29714 12480 30262
rect 12544 30054 12572 33068
rect 12532 30048 12584 30054
rect 12532 29990 12584 29996
rect 12440 29708 12492 29714
rect 12440 29650 12492 29656
rect 12348 29640 12400 29646
rect 12348 29582 12400 29588
rect 12360 29238 12388 29582
rect 12348 29232 12400 29238
rect 12348 29174 12400 29180
rect 12348 28620 12400 28626
rect 12348 28562 12400 28568
rect 12360 28082 12388 28562
rect 12440 28552 12492 28558
rect 12440 28494 12492 28500
rect 12348 28076 12400 28082
rect 12348 28018 12400 28024
rect 12452 27674 12480 28494
rect 12636 28121 12664 33238
rect 12728 33114 12756 33322
rect 12912 33114 12940 33458
rect 13176 33380 13228 33386
rect 13176 33322 13228 33328
rect 12716 33108 12768 33114
rect 12716 33050 12768 33056
rect 12900 33108 12952 33114
rect 12900 33050 12952 33056
rect 12806 33008 12862 33017
rect 12806 32943 12862 32952
rect 12716 32904 12768 32910
rect 12716 32846 12768 32852
rect 12728 31521 12756 32846
rect 12714 31512 12770 31521
rect 12714 31447 12770 31456
rect 12622 28112 12678 28121
rect 12622 28047 12678 28056
rect 12440 27668 12492 27674
rect 12440 27610 12492 27616
rect 12452 26994 12480 27610
rect 12440 26988 12492 26994
rect 12440 26930 12492 26936
rect 12452 26382 12480 26930
rect 12440 26376 12492 26382
rect 12440 26318 12492 26324
rect 12452 26042 12480 26318
rect 12440 26036 12492 26042
rect 12440 25978 12492 25984
rect 12452 25498 12480 25978
rect 12440 25492 12492 25498
rect 12440 25434 12492 25440
rect 12256 24404 12308 24410
rect 12256 24346 12308 24352
rect 12268 23798 12296 24346
rect 12256 23792 12308 23798
rect 12256 23734 12308 23740
rect 12532 20800 12584 20806
rect 12532 20742 12584 20748
rect 12440 20528 12492 20534
rect 12440 20470 12492 20476
rect 12256 20460 12308 20466
rect 12256 20402 12308 20408
rect 11940 19944 12020 19972
rect 12164 19984 12216 19990
rect 11888 19926 11940 19932
rect 12164 19926 12216 19932
rect 11794 19887 11796 19896
rect 11848 19887 11850 19896
rect 11796 19858 11848 19864
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 12070 19816 12126 19825
rect 11520 19780 11572 19786
rect 11520 19722 11572 19728
rect 11532 19514 11560 19722
rect 11520 19508 11572 19514
rect 11520 19450 11572 19456
rect 11624 19446 11652 19790
rect 12070 19751 12126 19760
rect 11612 19440 11664 19446
rect 11612 19382 11664 19388
rect 11520 19168 11572 19174
rect 11520 19110 11572 19116
rect 11980 19168 12032 19174
rect 11980 19110 12032 19116
rect 11532 17678 11560 19110
rect 11622 19068 11918 19088
rect 11678 19066 11702 19068
rect 11758 19066 11782 19068
rect 11838 19066 11862 19068
rect 11700 19014 11702 19066
rect 11764 19014 11776 19066
rect 11838 19014 11840 19066
rect 11678 19012 11702 19014
rect 11758 19012 11782 19014
rect 11838 19012 11862 19014
rect 11622 18992 11918 19012
rect 11992 18873 12020 19110
rect 12084 18902 12112 19751
rect 12164 19712 12216 19718
rect 12164 19654 12216 19660
rect 12072 18896 12124 18902
rect 11978 18864 12034 18873
rect 12072 18838 12124 18844
rect 11978 18799 12034 18808
rect 11704 18760 11756 18766
rect 11702 18728 11704 18737
rect 12072 18760 12124 18766
rect 11756 18728 11758 18737
rect 12072 18702 12124 18708
rect 11702 18663 11758 18672
rect 11716 18426 11744 18663
rect 12084 18426 12112 18702
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 11622 17980 11918 18000
rect 11678 17978 11702 17980
rect 11758 17978 11782 17980
rect 11838 17978 11862 17980
rect 11700 17926 11702 17978
rect 11764 17926 11776 17978
rect 11838 17926 11840 17978
rect 11678 17924 11702 17926
rect 11758 17924 11782 17926
rect 11838 17924 11862 17926
rect 11622 17904 11918 17924
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 11622 16892 11918 16912
rect 11678 16890 11702 16892
rect 11758 16890 11782 16892
rect 11838 16890 11862 16892
rect 11700 16838 11702 16890
rect 11764 16838 11776 16890
rect 11838 16838 11840 16890
rect 11678 16836 11702 16838
rect 11758 16836 11782 16838
rect 11838 16836 11862 16838
rect 11622 16816 11918 16836
rect 11622 15804 11918 15824
rect 11678 15802 11702 15804
rect 11758 15802 11782 15804
rect 11838 15802 11862 15804
rect 11700 15750 11702 15802
rect 11764 15750 11776 15802
rect 11838 15750 11840 15802
rect 11678 15748 11702 15750
rect 11758 15748 11782 15750
rect 11838 15748 11862 15750
rect 11622 15728 11918 15748
rect 11622 14716 11918 14736
rect 11678 14714 11702 14716
rect 11758 14714 11782 14716
rect 11838 14714 11862 14716
rect 11700 14662 11702 14714
rect 11764 14662 11776 14714
rect 11838 14662 11840 14714
rect 11678 14660 11702 14662
rect 11758 14660 11782 14662
rect 11838 14660 11862 14662
rect 11622 14640 11918 14660
rect 11622 13628 11918 13648
rect 11678 13626 11702 13628
rect 11758 13626 11782 13628
rect 11838 13626 11862 13628
rect 11700 13574 11702 13626
rect 11764 13574 11776 13626
rect 11838 13574 11840 13626
rect 11678 13572 11702 13574
rect 11758 13572 11782 13574
rect 11838 13572 11862 13574
rect 11622 13552 11918 13572
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11624 12850 11652 13330
rect 11716 12918 11744 13330
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 11808 12986 11836 13262
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11704 12912 11756 12918
rect 11704 12854 11756 12860
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11622 12540 11918 12560
rect 11678 12538 11702 12540
rect 11758 12538 11782 12540
rect 11838 12538 11862 12540
rect 11700 12486 11702 12538
rect 11764 12486 11776 12538
rect 11838 12486 11840 12538
rect 11678 12484 11702 12486
rect 11758 12484 11782 12486
rect 11838 12484 11862 12486
rect 11622 12464 11918 12484
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11348 11478 11468 11506
rect 11348 11150 11376 11478
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 11348 10470 11376 11086
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11242 10024 11298 10033
rect 11242 9959 11298 9968
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 11256 9586 11284 9862
rect 11244 9580 11296 9586
rect 11164 9540 11244 9568
rect 11164 9110 11192 9540
rect 11244 9522 11296 9528
rect 11348 9466 11376 10406
rect 11428 9988 11480 9994
rect 11428 9930 11480 9936
rect 11256 9438 11376 9466
rect 11440 9450 11468 9930
rect 11428 9444 11480 9450
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 11152 9104 11204 9110
rect 11152 9046 11204 9052
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10980 8634 11008 9046
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 10612 5166 10640 5306
rect 10600 5160 10652 5166
rect 10598 5128 10600 5137
rect 10652 5128 10654 5137
rect 10598 5063 10654 5072
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 10600 5024 10652 5030
rect 10600 4966 10652 4972
rect 10612 4826 10640 4966
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10612 4010 10640 4762
rect 10704 4486 10732 5034
rect 10692 4480 10744 4486
rect 10888 4468 10916 8026
rect 10980 6848 11008 8434
rect 11164 8294 11192 8774
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11164 7886 11192 8230
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11164 7002 11192 7822
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 11060 6860 11112 6866
rect 10980 6820 11060 6848
rect 11060 6802 11112 6808
rect 11072 6458 11100 6802
rect 11060 6452 11112 6458
rect 10692 4422 10744 4428
rect 10796 4440 10916 4468
rect 10980 6412 11060 6440
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10520 3641 10548 3878
rect 10704 3738 10732 4422
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10506 3632 10562 3641
rect 10506 3567 10562 3576
rect 10046 2952 10102 2961
rect 10046 2887 10102 2896
rect 10244 2944 10364 2972
rect 10060 2650 10088 2887
rect 10244 2666 10272 2944
rect 10796 2922 10824 4440
rect 10980 3738 11008 6412
rect 11060 6394 11112 6400
rect 11150 5944 11206 5953
rect 11060 5908 11112 5914
rect 11150 5879 11152 5888
rect 11060 5850 11112 5856
rect 11204 5879 11206 5888
rect 11152 5850 11204 5856
rect 11072 5817 11100 5850
rect 11058 5808 11114 5817
rect 11058 5743 11114 5752
rect 11150 4992 11206 5001
rect 11150 4927 11206 4936
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 10980 3534 11008 3674
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10980 3058 11008 3470
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 11164 2922 11192 4927
rect 10784 2916 10836 2922
rect 10784 2858 10836 2864
rect 11060 2916 11112 2922
rect 11060 2858 11112 2864
rect 11152 2916 11204 2922
rect 11152 2858 11204 2864
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 10152 2638 10272 2666
rect 11072 2650 11100 2858
rect 11150 2816 11206 2825
rect 11150 2751 11206 2760
rect 11060 2644 11112 2650
rect 9956 672 10008 678
rect 9956 614 10008 620
rect 9864 604 9916 610
rect 9864 546 9916 552
rect 10152 480 10180 2638
rect 11060 2586 11112 2592
rect 11164 2582 11192 2751
rect 11152 2576 11204 2582
rect 11256 2553 11284 9438
rect 11428 9386 11480 9392
rect 11440 8090 11468 9386
rect 11532 9058 11560 11562
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11622 11452 11918 11472
rect 11678 11450 11702 11452
rect 11758 11450 11782 11452
rect 11838 11450 11862 11452
rect 11700 11398 11702 11450
rect 11764 11398 11776 11450
rect 11838 11398 11840 11450
rect 11678 11396 11702 11398
rect 11758 11396 11782 11398
rect 11838 11396 11862 11398
rect 11622 11376 11918 11396
rect 11992 11150 12020 11494
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11992 10470 12020 11086
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11622 10364 11918 10384
rect 11678 10362 11702 10364
rect 11758 10362 11782 10364
rect 11838 10362 11862 10364
rect 11700 10310 11702 10362
rect 11764 10310 11776 10362
rect 11838 10310 11840 10362
rect 11678 10308 11702 10310
rect 11758 10308 11782 10310
rect 11838 10308 11862 10310
rect 11622 10288 11918 10308
rect 11622 9276 11918 9296
rect 11678 9274 11702 9276
rect 11758 9274 11782 9276
rect 11838 9274 11862 9276
rect 11700 9222 11702 9274
rect 11764 9222 11776 9274
rect 11838 9222 11840 9274
rect 11678 9220 11702 9222
rect 11758 9220 11782 9222
rect 11838 9220 11862 9222
rect 11622 9200 11918 9220
rect 11992 9178 12020 10406
rect 12176 9654 12204 19654
rect 12268 13394 12296 20402
rect 12452 20058 12480 20470
rect 12440 20052 12492 20058
rect 12440 19994 12492 20000
rect 12544 19938 12572 20742
rect 12452 19910 12572 19938
rect 12624 19916 12676 19922
rect 12348 19848 12400 19854
rect 12452 19836 12480 19910
rect 12624 19858 12676 19864
rect 12400 19808 12480 19836
rect 12532 19848 12584 19854
rect 12348 19790 12400 19796
rect 12532 19790 12584 19796
rect 12544 19378 12572 19790
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 12636 19174 12664 19858
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12624 19168 12676 19174
rect 12624 19110 12676 19116
rect 12452 18193 12480 19110
rect 12438 18184 12494 18193
rect 12438 18119 12494 18128
rect 12348 17332 12400 17338
rect 12348 17274 12400 17280
rect 12360 16946 12388 17274
rect 12438 16960 12494 16969
rect 12360 16918 12438 16946
rect 12438 16895 12494 16904
rect 12636 16794 12664 19110
rect 12440 16788 12492 16794
rect 12440 16730 12492 16736
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 12164 9648 12216 9654
rect 12164 9590 12216 9596
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11532 9030 12020 9058
rect 11622 8188 11918 8208
rect 11678 8186 11702 8188
rect 11758 8186 11782 8188
rect 11838 8186 11862 8188
rect 11700 8134 11702 8186
rect 11764 8134 11776 8186
rect 11838 8134 11840 8186
rect 11678 8132 11702 8134
rect 11758 8132 11782 8134
rect 11838 8132 11862 8134
rect 11622 8112 11918 8132
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 11440 7546 11468 7890
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 11440 7002 11468 7482
rect 11622 7100 11918 7120
rect 11678 7098 11702 7100
rect 11758 7098 11782 7100
rect 11838 7098 11862 7100
rect 11700 7046 11702 7098
rect 11764 7046 11776 7098
rect 11838 7046 11840 7098
rect 11678 7044 11702 7046
rect 11758 7044 11782 7046
rect 11838 7044 11862 7046
rect 11622 7024 11918 7044
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11348 5846 11376 6054
rect 11336 5840 11388 5846
rect 11336 5782 11388 5788
rect 11440 5234 11468 6938
rect 11622 6012 11918 6032
rect 11678 6010 11702 6012
rect 11758 6010 11782 6012
rect 11838 6010 11862 6012
rect 11700 5958 11702 6010
rect 11764 5958 11776 6010
rect 11838 5958 11840 6010
rect 11678 5956 11702 5958
rect 11758 5956 11782 5958
rect 11838 5956 11862 5958
rect 11622 5936 11918 5956
rect 11428 5228 11480 5234
rect 11348 5188 11428 5216
rect 11348 4078 11376 5188
rect 11428 5170 11480 5176
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11532 4826 11560 4966
rect 11622 4924 11918 4944
rect 11678 4922 11702 4924
rect 11758 4922 11782 4924
rect 11838 4922 11862 4924
rect 11700 4870 11702 4922
rect 11764 4870 11776 4922
rect 11838 4870 11840 4922
rect 11678 4868 11702 4870
rect 11758 4868 11782 4870
rect 11838 4868 11862 4870
rect 11622 4848 11918 4868
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11336 4072 11388 4078
rect 11336 4014 11388 4020
rect 11440 4010 11468 4626
rect 11428 4004 11480 4010
rect 11428 3946 11480 3952
rect 11334 3904 11390 3913
rect 11334 3839 11390 3848
rect 11152 2518 11204 2524
rect 11242 2544 11298 2553
rect 11242 2479 11298 2488
rect 10600 604 10652 610
rect 10600 546 10652 552
rect 10968 604 11020 610
rect 10968 546 11020 552
rect 10612 480 10640 546
rect 10980 480 11008 546
rect 11348 480 11376 3839
rect 11440 3602 11468 3946
rect 11532 3738 11560 4762
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11808 4214 11836 4558
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 11622 3836 11918 3856
rect 11678 3834 11702 3836
rect 11758 3834 11782 3836
rect 11838 3834 11862 3836
rect 11700 3782 11702 3834
rect 11764 3782 11776 3834
rect 11838 3782 11840 3834
rect 11678 3780 11702 3782
rect 11758 3780 11782 3782
rect 11838 3780 11862 3782
rect 11622 3760 11918 3780
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11428 3596 11480 3602
rect 11428 3538 11480 3544
rect 11428 3052 11480 3058
rect 11428 2994 11480 3000
rect 11440 2650 11468 2994
rect 11622 2748 11918 2768
rect 11678 2746 11702 2748
rect 11758 2746 11782 2748
rect 11838 2746 11862 2748
rect 11700 2694 11702 2746
rect 11764 2694 11776 2746
rect 11838 2694 11840 2746
rect 11678 2692 11702 2694
rect 11758 2692 11782 2694
rect 11838 2692 11862 2694
rect 11622 2672 11918 2692
rect 11428 2644 11480 2650
rect 11428 2586 11480 2592
rect 11440 2446 11468 2586
rect 11992 2530 12020 9030
rect 12268 7993 12296 13330
rect 12452 11218 12480 16730
rect 12622 16688 12678 16697
rect 12622 16623 12678 16632
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12360 10742 12388 11154
rect 12348 10736 12400 10742
rect 12348 10678 12400 10684
rect 12360 10169 12388 10678
rect 12346 10160 12402 10169
rect 12346 10095 12402 10104
rect 12254 7984 12310 7993
rect 12254 7919 12310 7928
rect 12440 7744 12492 7750
rect 12440 7686 12492 7692
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 12084 6934 12112 7142
rect 12072 6928 12124 6934
rect 12072 6870 12124 6876
rect 12084 6118 12112 6870
rect 12162 6624 12218 6633
rect 12162 6559 12218 6568
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 12084 5778 12112 6054
rect 12072 5772 12124 5778
rect 12072 5714 12124 5720
rect 12084 5370 12112 5714
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 12176 4826 12204 6559
rect 12452 5114 12480 7686
rect 12636 5896 12664 16623
rect 12268 5086 12480 5114
rect 12544 5868 12664 5896
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 12268 4622 12296 5086
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12256 4616 12308 4622
rect 12256 4558 12308 4564
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 12268 3534 12296 4082
rect 12360 3738 12388 4966
rect 12438 4584 12494 4593
rect 12438 4519 12440 4528
rect 12492 4519 12494 4528
rect 12440 4490 12492 4496
rect 12348 3732 12400 3738
rect 12348 3674 12400 3680
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 12256 3528 12308 3534
rect 12256 3470 12308 3476
rect 12176 3194 12204 3470
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 12268 3074 12296 3470
rect 12084 3046 12296 3074
rect 12360 3058 12388 3674
rect 12438 3632 12494 3641
rect 12438 3567 12494 3576
rect 12452 3194 12480 3567
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12348 3052 12400 3058
rect 12084 2650 12112 3046
rect 12348 2994 12400 3000
rect 12164 2916 12216 2922
rect 12164 2858 12216 2864
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 11808 2502 12020 2530
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 11808 480 11836 2502
rect 12176 480 12204 2858
rect 12544 480 12572 5868
rect 12728 5273 12756 31447
rect 12820 27130 12848 32943
rect 12900 30592 12952 30598
rect 12900 30534 12952 30540
rect 12912 30297 12940 30534
rect 12898 30288 12954 30297
rect 12898 30223 12954 30232
rect 12912 30190 12940 30223
rect 12900 30184 12952 30190
rect 12900 30126 12952 30132
rect 12900 30048 12952 30054
rect 12900 29990 12952 29996
rect 12912 29753 12940 29990
rect 12898 29744 12954 29753
rect 12898 29679 12954 29688
rect 12992 29708 13044 29714
rect 12992 29650 13044 29656
rect 13004 28762 13032 29650
rect 13082 28792 13138 28801
rect 12992 28756 13044 28762
rect 13082 28727 13138 28736
rect 12992 28698 13044 28704
rect 12808 27124 12860 27130
rect 12808 27066 12860 27072
rect 13096 27010 13124 28727
rect 12820 26982 13124 27010
rect 12714 5264 12770 5273
rect 12714 5199 12770 5208
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12636 4146 12664 4762
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12728 3738 12756 5199
rect 12820 4690 12848 26982
rect 12900 26920 12952 26926
rect 12900 26862 12952 26868
rect 12912 20466 12940 26862
rect 12992 26580 13044 26586
rect 12992 26522 13044 26528
rect 13004 25702 13032 26522
rect 12992 25696 13044 25702
rect 12992 25638 13044 25644
rect 12990 23216 13046 23225
rect 12990 23151 13046 23160
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 13004 19922 13032 23151
rect 13188 20482 13216 33322
rect 13372 27033 13400 39520
rect 13648 39494 13768 39520
rect 13358 27024 13414 27033
rect 13358 26959 13414 26968
rect 13648 25106 13676 39494
rect 13728 30252 13780 30258
rect 13728 30194 13780 30200
rect 13740 30025 13768 30194
rect 13726 30016 13782 30025
rect 13726 29951 13782 29960
rect 13740 29850 13768 29951
rect 13728 29844 13780 29850
rect 13728 29786 13780 29792
rect 14200 29102 14228 39520
rect 14568 37210 14596 39520
rect 14568 37182 14688 37210
rect 14289 37020 14585 37040
rect 14345 37018 14369 37020
rect 14425 37018 14449 37020
rect 14505 37018 14529 37020
rect 14367 36966 14369 37018
rect 14431 36966 14443 37018
rect 14505 36966 14507 37018
rect 14345 36964 14369 36966
rect 14425 36964 14449 36966
rect 14505 36964 14529 36966
rect 14289 36944 14585 36964
rect 14289 35932 14585 35952
rect 14345 35930 14369 35932
rect 14425 35930 14449 35932
rect 14505 35930 14529 35932
rect 14367 35878 14369 35930
rect 14431 35878 14443 35930
rect 14505 35878 14507 35930
rect 14345 35876 14369 35878
rect 14425 35876 14449 35878
rect 14505 35876 14529 35878
rect 14289 35856 14585 35876
rect 14289 34844 14585 34864
rect 14345 34842 14369 34844
rect 14425 34842 14449 34844
rect 14505 34842 14529 34844
rect 14367 34790 14369 34842
rect 14431 34790 14443 34842
rect 14505 34790 14507 34842
rect 14345 34788 14369 34790
rect 14425 34788 14449 34790
rect 14505 34788 14529 34790
rect 14289 34768 14585 34788
rect 14289 33756 14585 33776
rect 14345 33754 14369 33756
rect 14425 33754 14449 33756
rect 14505 33754 14529 33756
rect 14367 33702 14369 33754
rect 14431 33702 14443 33754
rect 14505 33702 14507 33754
rect 14345 33700 14369 33702
rect 14425 33700 14449 33702
rect 14505 33700 14529 33702
rect 14289 33680 14585 33700
rect 14660 32910 14688 37182
rect 14936 33017 14964 39520
rect 15396 34105 15424 39520
rect 15382 34096 15438 34105
rect 15382 34031 15438 34040
rect 14922 33008 14978 33017
rect 14922 32943 14978 32952
rect 14648 32904 14700 32910
rect 14648 32846 14700 32852
rect 14289 32668 14585 32688
rect 14345 32666 14369 32668
rect 14425 32666 14449 32668
rect 14505 32666 14529 32668
rect 14367 32614 14369 32666
rect 14431 32614 14443 32666
rect 14505 32614 14507 32666
rect 14345 32612 14369 32614
rect 14425 32612 14449 32614
rect 14505 32612 14529 32614
rect 14289 32592 14585 32612
rect 14289 31580 14585 31600
rect 14345 31578 14369 31580
rect 14425 31578 14449 31580
rect 14505 31578 14529 31580
rect 14367 31526 14369 31578
rect 14431 31526 14443 31578
rect 14505 31526 14507 31578
rect 14345 31524 14369 31526
rect 14425 31524 14449 31526
rect 14505 31524 14529 31526
rect 14289 31504 14585 31524
rect 14289 30492 14585 30512
rect 14345 30490 14369 30492
rect 14425 30490 14449 30492
rect 14505 30490 14529 30492
rect 14367 30438 14369 30490
rect 14431 30438 14443 30490
rect 14505 30438 14507 30490
rect 14345 30436 14369 30438
rect 14425 30436 14449 30438
rect 14505 30436 14529 30438
rect 14289 30416 14585 30436
rect 14289 29404 14585 29424
rect 14345 29402 14369 29404
rect 14425 29402 14449 29404
rect 14505 29402 14529 29404
rect 14367 29350 14369 29402
rect 14431 29350 14443 29402
rect 14505 29350 14507 29402
rect 14345 29348 14369 29350
rect 14425 29348 14449 29350
rect 14505 29348 14529 29350
rect 14289 29328 14585 29348
rect 14188 29096 14240 29102
rect 14188 29038 14240 29044
rect 15764 28801 15792 39520
rect 15750 28792 15806 28801
rect 15750 28727 15806 28736
rect 14289 28316 14585 28336
rect 14345 28314 14369 28316
rect 14425 28314 14449 28316
rect 14505 28314 14529 28316
rect 14367 28262 14369 28314
rect 14431 28262 14443 28314
rect 14505 28262 14507 28314
rect 14345 28260 14369 28262
rect 14425 28260 14449 28262
rect 14505 28260 14529 28262
rect 14289 28240 14585 28260
rect 14289 27228 14585 27248
rect 14345 27226 14369 27228
rect 14425 27226 14449 27228
rect 14505 27226 14529 27228
rect 14367 27174 14369 27226
rect 14431 27174 14443 27226
rect 14505 27174 14507 27226
rect 14345 27172 14369 27174
rect 14425 27172 14449 27174
rect 14505 27172 14529 27174
rect 14289 27152 14585 27172
rect 14289 26140 14585 26160
rect 14345 26138 14369 26140
rect 14425 26138 14449 26140
rect 14505 26138 14529 26140
rect 14367 26086 14369 26138
rect 14431 26086 14443 26138
rect 14505 26086 14507 26138
rect 14345 26084 14369 26086
rect 14425 26084 14449 26086
rect 14505 26084 14529 26086
rect 14289 26064 14585 26084
rect 13556 25078 13676 25106
rect 13556 22681 13584 25078
rect 14289 25052 14585 25072
rect 14345 25050 14369 25052
rect 14425 25050 14449 25052
rect 14505 25050 14529 25052
rect 14367 24998 14369 25050
rect 14431 24998 14443 25050
rect 14505 24998 14507 25050
rect 14345 24996 14369 24998
rect 14425 24996 14449 24998
rect 14505 24996 14529 24998
rect 13634 24984 13690 24993
rect 14289 24976 14585 24996
rect 13634 24919 13690 24928
rect 13542 22672 13598 22681
rect 13542 22607 13598 22616
rect 13188 20454 13308 20482
rect 13176 20392 13228 20398
rect 13176 20334 13228 20340
rect 12992 19916 13044 19922
rect 12992 19858 13044 19864
rect 13188 19854 13216 20334
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 13176 19848 13228 19854
rect 13176 19790 13228 19796
rect 13096 19417 13124 19790
rect 13082 19408 13138 19417
rect 12992 19372 13044 19378
rect 13082 19343 13138 19352
rect 12992 19314 13044 19320
rect 13004 18970 13032 19314
rect 12992 18964 13044 18970
rect 12992 18906 13044 18912
rect 13004 18766 13032 18906
rect 13096 18902 13124 19343
rect 13084 18896 13136 18902
rect 13084 18838 13136 18844
rect 12992 18760 13044 18766
rect 12992 18702 13044 18708
rect 13280 14929 13308 20454
rect 13266 14920 13322 14929
rect 13266 14855 13322 14864
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 12898 7848 12954 7857
rect 12898 7783 12954 7792
rect 12808 4684 12860 4690
rect 12808 4626 12860 4632
rect 12820 4282 12848 4626
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 12820 3670 12848 4218
rect 12808 3664 12860 3670
rect 12808 3606 12860 3612
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 12912 3482 12940 7783
rect 13004 3942 13032 9590
rect 13358 5128 13414 5137
rect 13358 5063 13414 5072
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13268 3596 13320 3602
rect 13268 3538 13320 3544
rect 12622 3088 12678 3097
rect 12622 3023 12678 3032
rect 12636 2514 12664 3023
rect 12728 2990 12756 3470
rect 12912 3454 13032 3482
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12806 2952 12862 2961
rect 12806 2887 12808 2896
rect 12860 2887 12862 2896
rect 12808 2858 12860 2864
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 12806 2408 12862 2417
rect 12806 2343 12808 2352
rect 12860 2343 12862 2352
rect 12808 2314 12860 2320
rect 13004 480 13032 3454
rect 13084 3392 13136 3398
rect 13084 3334 13136 3340
rect 13096 3126 13124 3334
rect 13280 3194 13308 3538
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 13084 3120 13136 3126
rect 13084 3062 13136 3068
rect 13372 480 13400 5063
rect 13648 3505 13676 24919
rect 14289 23964 14585 23984
rect 14345 23962 14369 23964
rect 14425 23962 14449 23964
rect 14505 23962 14529 23964
rect 14367 23910 14369 23962
rect 14431 23910 14443 23962
rect 14505 23910 14507 23962
rect 14345 23908 14369 23910
rect 14425 23908 14449 23910
rect 14505 23908 14529 23910
rect 14289 23888 14585 23908
rect 14289 22876 14585 22896
rect 14345 22874 14369 22876
rect 14425 22874 14449 22876
rect 14505 22874 14529 22876
rect 14367 22822 14369 22874
rect 14431 22822 14443 22874
rect 14505 22822 14507 22874
rect 14345 22820 14369 22822
rect 14425 22820 14449 22822
rect 14505 22820 14529 22822
rect 14289 22800 14585 22820
rect 14289 21788 14585 21808
rect 14345 21786 14369 21788
rect 14425 21786 14449 21788
rect 14505 21786 14529 21788
rect 14367 21734 14369 21786
rect 14431 21734 14443 21786
rect 14505 21734 14507 21786
rect 14345 21732 14369 21734
rect 14425 21732 14449 21734
rect 14505 21732 14529 21734
rect 14289 21712 14585 21732
rect 14289 20700 14585 20720
rect 14345 20698 14369 20700
rect 14425 20698 14449 20700
rect 14505 20698 14529 20700
rect 14367 20646 14369 20698
rect 14431 20646 14443 20698
rect 14505 20646 14507 20698
rect 14345 20644 14369 20646
rect 14425 20644 14449 20646
rect 14505 20644 14529 20646
rect 14289 20624 14585 20644
rect 14289 19612 14585 19632
rect 14345 19610 14369 19612
rect 14425 19610 14449 19612
rect 14505 19610 14529 19612
rect 14367 19558 14369 19610
rect 14431 19558 14443 19610
rect 14505 19558 14507 19610
rect 14345 19556 14369 19558
rect 14425 19556 14449 19558
rect 14505 19556 14529 19558
rect 14289 19536 14585 19556
rect 14289 18524 14585 18544
rect 14345 18522 14369 18524
rect 14425 18522 14449 18524
rect 14505 18522 14529 18524
rect 14367 18470 14369 18522
rect 14431 18470 14443 18522
rect 14505 18470 14507 18522
rect 14345 18468 14369 18470
rect 14425 18468 14449 18470
rect 14505 18468 14529 18470
rect 14289 18448 14585 18468
rect 14289 17436 14585 17456
rect 14345 17434 14369 17436
rect 14425 17434 14449 17436
rect 14505 17434 14529 17436
rect 14367 17382 14369 17434
rect 14431 17382 14443 17434
rect 14505 17382 14507 17434
rect 14345 17380 14369 17382
rect 14425 17380 14449 17382
rect 14505 17380 14529 17382
rect 14289 17360 14585 17380
rect 14289 16348 14585 16368
rect 14345 16346 14369 16348
rect 14425 16346 14449 16348
rect 14505 16346 14529 16348
rect 14367 16294 14369 16346
rect 14431 16294 14443 16346
rect 14505 16294 14507 16346
rect 14345 16292 14369 16294
rect 14425 16292 14449 16294
rect 14505 16292 14529 16294
rect 14289 16272 14585 16292
rect 14289 15260 14585 15280
rect 14345 15258 14369 15260
rect 14425 15258 14449 15260
rect 14505 15258 14529 15260
rect 14367 15206 14369 15258
rect 14431 15206 14443 15258
rect 14505 15206 14507 15258
rect 14345 15204 14369 15206
rect 14425 15204 14449 15206
rect 14505 15204 14529 15206
rect 14289 15184 14585 15204
rect 14289 14172 14585 14192
rect 14345 14170 14369 14172
rect 14425 14170 14449 14172
rect 14505 14170 14529 14172
rect 14367 14118 14369 14170
rect 14431 14118 14443 14170
rect 14505 14118 14507 14170
rect 14345 14116 14369 14118
rect 14425 14116 14449 14118
rect 14505 14116 14529 14118
rect 14289 14096 14585 14116
rect 14289 13084 14585 13104
rect 14345 13082 14369 13084
rect 14425 13082 14449 13084
rect 14505 13082 14529 13084
rect 14367 13030 14369 13082
rect 14431 13030 14443 13082
rect 14505 13030 14507 13082
rect 14345 13028 14369 13030
rect 14425 13028 14449 13030
rect 14505 13028 14529 13030
rect 14289 13008 14585 13028
rect 14289 11996 14585 12016
rect 14345 11994 14369 11996
rect 14425 11994 14449 11996
rect 14505 11994 14529 11996
rect 14367 11942 14369 11994
rect 14431 11942 14443 11994
rect 14505 11942 14507 11994
rect 14345 11940 14369 11942
rect 14425 11940 14449 11942
rect 14505 11940 14529 11942
rect 14289 11920 14585 11940
rect 14289 10908 14585 10928
rect 14345 10906 14369 10908
rect 14425 10906 14449 10908
rect 14505 10906 14529 10908
rect 14367 10854 14369 10906
rect 14431 10854 14443 10906
rect 14505 10854 14507 10906
rect 14345 10852 14369 10854
rect 14425 10852 14449 10854
rect 14505 10852 14529 10854
rect 14289 10832 14585 10852
rect 14830 10160 14886 10169
rect 14830 10095 14886 10104
rect 14289 9820 14585 9840
rect 14345 9818 14369 9820
rect 14425 9818 14449 9820
rect 14505 9818 14529 9820
rect 14367 9766 14369 9818
rect 14431 9766 14443 9818
rect 14505 9766 14507 9818
rect 14345 9764 14369 9766
rect 14425 9764 14449 9766
rect 14505 9764 14529 9766
rect 14289 9744 14585 9764
rect 14289 8732 14585 8752
rect 14345 8730 14369 8732
rect 14425 8730 14449 8732
rect 14505 8730 14529 8732
rect 14367 8678 14369 8730
rect 14431 8678 14443 8730
rect 14505 8678 14507 8730
rect 14345 8676 14369 8678
rect 14425 8676 14449 8678
rect 14505 8676 14529 8678
rect 14289 8656 14585 8676
rect 14289 7644 14585 7664
rect 14345 7642 14369 7644
rect 14425 7642 14449 7644
rect 14505 7642 14529 7644
rect 14367 7590 14369 7642
rect 14431 7590 14443 7642
rect 14505 7590 14507 7642
rect 14345 7588 14369 7590
rect 14425 7588 14449 7590
rect 14505 7588 14529 7590
rect 14289 7568 14585 7588
rect 14289 6556 14585 6576
rect 14345 6554 14369 6556
rect 14425 6554 14449 6556
rect 14505 6554 14529 6556
rect 14367 6502 14369 6554
rect 14431 6502 14443 6554
rect 14505 6502 14507 6554
rect 14345 6500 14369 6502
rect 14425 6500 14449 6502
rect 14505 6500 14529 6502
rect 14289 6480 14585 6500
rect 14289 5468 14585 5488
rect 14345 5466 14369 5468
rect 14425 5466 14449 5468
rect 14505 5466 14529 5468
rect 14367 5414 14369 5466
rect 14431 5414 14443 5466
rect 14505 5414 14507 5466
rect 14345 5412 14369 5414
rect 14425 5412 14449 5414
rect 14505 5412 14529 5414
rect 14289 5392 14585 5412
rect 14646 4720 14702 4729
rect 14646 4655 14702 4664
rect 14289 4380 14585 4400
rect 14345 4378 14369 4380
rect 14425 4378 14449 4380
rect 14505 4378 14529 4380
rect 14367 4326 14369 4378
rect 14431 4326 14443 4378
rect 14505 4326 14507 4378
rect 14345 4324 14369 4326
rect 14425 4324 14449 4326
rect 14505 4324 14529 4326
rect 14289 4304 14585 4324
rect 13726 4040 13782 4049
rect 13726 3975 13782 3984
rect 13450 3496 13506 3505
rect 13450 3431 13452 3440
rect 13504 3431 13506 3440
rect 13634 3496 13690 3505
rect 13634 3431 13690 3440
rect 13452 3402 13504 3408
rect 13740 480 13768 3975
rect 14186 3496 14242 3505
rect 14186 3431 14242 3440
rect 14200 480 14228 3431
rect 14289 3292 14585 3312
rect 14345 3290 14369 3292
rect 14425 3290 14449 3292
rect 14505 3290 14529 3292
rect 14367 3238 14369 3290
rect 14431 3238 14443 3290
rect 14505 3238 14507 3290
rect 14345 3236 14369 3238
rect 14425 3236 14449 3238
rect 14505 3236 14529 3238
rect 14289 3216 14585 3236
rect 14289 2204 14585 2224
rect 14345 2202 14369 2204
rect 14425 2202 14449 2204
rect 14505 2202 14529 2204
rect 14367 2150 14369 2202
rect 14431 2150 14443 2202
rect 14505 2150 14507 2202
rect 14345 2148 14369 2150
rect 14425 2148 14449 2150
rect 14505 2148 14529 2150
rect 14289 2128 14585 2148
rect 14660 1986 14688 4655
rect 14844 3482 14872 10095
rect 15382 7304 15438 7313
rect 15382 7239 15438 7248
rect 14844 3454 14964 3482
rect 14568 1958 14688 1986
rect 14568 480 14596 1958
rect 14936 480 14964 3454
rect 15396 480 15424 7239
rect 15752 3936 15804 3942
rect 15752 3878 15804 3884
rect 15764 480 15792 3878
rect 202 0 258 480
rect 570 0 626 480
rect 938 0 994 480
rect 1398 0 1454 480
rect 1766 0 1822 480
rect 2134 0 2190 480
rect 2594 0 2650 480
rect 2962 0 3018 480
rect 3330 0 3386 480
rect 3790 0 3846 480
rect 4158 0 4214 480
rect 4526 0 4582 480
rect 4986 0 5042 480
rect 5354 0 5410 480
rect 5722 0 5778 480
rect 6182 0 6238 480
rect 6550 0 6606 480
rect 6918 0 6974 480
rect 7378 0 7434 480
rect 7746 0 7802 480
rect 8206 0 8262 480
rect 8574 0 8630 480
rect 8942 0 8998 480
rect 9402 0 9458 480
rect 9770 0 9826 480
rect 10138 0 10194 480
rect 10598 0 10654 480
rect 10966 0 11022 480
rect 11334 0 11390 480
rect 11794 0 11850 480
rect 12162 0 12218 480
rect 12530 0 12586 480
rect 12990 0 13046 480
rect 13358 0 13414 480
rect 13726 0 13782 480
rect 14186 0 14242 480
rect 14554 0 14610 480
rect 14922 0 14978 480
rect 15382 0 15438 480
rect 15750 0 15806 480
<< via2 >>
rect 202 34720 258 34776
rect 1582 38664 1638 38720
rect 1490 36352 1546 36408
rect 2962 35672 3018 35728
rect 2594 35264 2650 35320
rect 2134 34992 2190 35048
rect 3238 34740 3294 34776
rect 3238 34720 3240 34740
rect 3240 34720 3292 34740
rect 3292 34720 3294 34740
rect 1950 34176 2006 34232
rect 1674 34040 1730 34096
rect 3622 37018 3678 37020
rect 3702 37018 3758 37020
rect 3782 37018 3838 37020
rect 3862 37018 3918 37020
rect 3622 36966 3648 37018
rect 3648 36966 3678 37018
rect 3702 36966 3712 37018
rect 3712 36966 3758 37018
rect 3782 36966 3828 37018
rect 3828 36966 3838 37018
rect 3862 36966 3892 37018
rect 3892 36966 3918 37018
rect 3622 36964 3678 36966
rect 3702 36964 3758 36966
rect 3782 36964 3838 36966
rect 3862 36964 3918 36966
rect 3622 35930 3678 35932
rect 3702 35930 3758 35932
rect 3782 35930 3838 35932
rect 3862 35930 3918 35932
rect 3622 35878 3648 35930
rect 3648 35878 3678 35930
rect 3702 35878 3712 35930
rect 3712 35878 3758 35930
rect 3782 35878 3828 35930
rect 3828 35878 3838 35930
rect 3862 35878 3892 35930
rect 3892 35878 3918 35930
rect 3622 35876 3678 35878
rect 3702 35876 3758 35878
rect 3782 35876 3838 35878
rect 3862 35876 3918 35878
rect 3622 34842 3678 34844
rect 3702 34842 3758 34844
rect 3782 34842 3838 34844
rect 3862 34842 3918 34844
rect 3622 34790 3648 34842
rect 3648 34790 3678 34842
rect 3702 34790 3712 34842
rect 3712 34790 3758 34842
rect 3782 34790 3828 34842
rect 3828 34790 3838 34842
rect 3862 34790 3892 34842
rect 3892 34790 3918 34842
rect 3622 34788 3678 34790
rect 3702 34788 3758 34790
rect 3782 34788 3838 34790
rect 3862 34788 3918 34790
rect 3698 34620 3700 34640
rect 3700 34620 3752 34640
rect 3752 34620 3754 34640
rect 3698 34584 3754 34620
rect 2502 34040 2558 34096
rect 2042 33904 2098 33960
rect 2410 33532 2412 33552
rect 2412 33532 2464 33552
rect 2464 33532 2466 33552
rect 2410 33496 2466 33532
rect 1398 32972 1454 33008
rect 1398 32952 1400 32972
rect 1400 32952 1452 32972
rect 1452 32952 1454 32972
rect 1674 31592 1730 31648
rect 3622 33754 3678 33756
rect 3702 33754 3758 33756
rect 3782 33754 3838 33756
rect 3862 33754 3918 33756
rect 3622 33702 3648 33754
rect 3648 33702 3678 33754
rect 3702 33702 3712 33754
rect 3712 33702 3758 33754
rect 3782 33702 3828 33754
rect 3828 33702 3838 33754
rect 3862 33702 3892 33754
rect 3892 33702 3918 33754
rect 3622 33700 3678 33702
rect 3702 33700 3758 33702
rect 3782 33700 3838 33702
rect 3862 33700 3918 33702
rect 1950 30776 2006 30832
rect 2134 30116 2190 30152
rect 2134 30096 2136 30116
rect 2136 30096 2188 30116
rect 2188 30096 2190 30116
rect 2410 30252 2466 30288
rect 2410 30232 2412 30252
rect 2412 30232 2464 30252
rect 2464 30232 2466 30252
rect 2226 29996 2228 30016
rect 2228 29996 2280 30016
rect 2280 29996 2282 30016
rect 2226 29960 2282 29996
rect 1582 28872 1638 28928
rect 3622 32666 3678 32668
rect 3702 32666 3758 32668
rect 3782 32666 3838 32668
rect 3862 32666 3918 32668
rect 3622 32614 3648 32666
rect 3648 32614 3678 32666
rect 3702 32614 3712 32666
rect 3712 32614 3758 32666
rect 3782 32614 3828 32666
rect 3828 32614 3838 32666
rect 3862 32614 3892 32666
rect 3892 32614 3918 32666
rect 3622 32612 3678 32614
rect 3702 32612 3758 32614
rect 3782 32612 3838 32614
rect 3862 32612 3918 32614
rect 3622 31578 3678 31580
rect 3702 31578 3758 31580
rect 3782 31578 3838 31580
rect 3862 31578 3918 31580
rect 3622 31526 3648 31578
rect 3648 31526 3678 31578
rect 3702 31526 3712 31578
rect 3712 31526 3758 31578
rect 3782 31526 3828 31578
rect 3828 31526 3838 31578
rect 3862 31526 3892 31578
rect 3892 31526 3918 31578
rect 3622 31524 3678 31526
rect 3702 31524 3758 31526
rect 3782 31524 3838 31526
rect 3862 31524 3918 31526
rect 3622 30490 3678 30492
rect 3702 30490 3758 30492
rect 3782 30490 3838 30492
rect 3862 30490 3918 30492
rect 3622 30438 3648 30490
rect 3648 30438 3678 30490
rect 3702 30438 3712 30490
rect 3712 30438 3758 30490
rect 3782 30438 3828 30490
rect 3828 30438 3838 30490
rect 3862 30438 3892 30490
rect 3892 30438 3918 30490
rect 3622 30436 3678 30438
rect 3702 30436 3758 30438
rect 3782 30436 3838 30438
rect 3862 30436 3918 30438
rect 2226 27512 2282 27568
rect 1582 24520 1638 24576
rect 1674 22208 1730 22264
rect 1398 20304 1454 20360
rect 1674 20204 1676 20224
rect 1676 20204 1728 20224
rect 1728 20204 1730 20224
rect 1674 20168 1730 20204
rect 1674 19896 1730 19952
rect 3622 29402 3678 29404
rect 3702 29402 3758 29404
rect 3782 29402 3838 29404
rect 3862 29402 3918 29404
rect 3622 29350 3648 29402
rect 3648 29350 3678 29402
rect 3702 29350 3712 29402
rect 3712 29350 3758 29402
rect 3782 29350 3828 29402
rect 3828 29350 3838 29402
rect 3862 29350 3892 29402
rect 3892 29350 3918 29402
rect 3622 29348 3678 29350
rect 3702 29348 3758 29350
rect 3782 29348 3838 29350
rect 3862 29348 3918 29350
rect 3698 29008 3754 29064
rect 3622 28314 3678 28316
rect 3702 28314 3758 28316
rect 3782 28314 3838 28316
rect 3862 28314 3918 28316
rect 3622 28262 3648 28314
rect 3648 28262 3678 28314
rect 3702 28262 3712 28314
rect 3712 28262 3758 28314
rect 3782 28262 3828 28314
rect 3828 28262 3838 28314
rect 3862 28262 3892 28314
rect 3892 28262 3918 28314
rect 3622 28260 3678 28262
rect 3702 28260 3758 28262
rect 3782 28260 3838 28262
rect 3862 28260 3918 28262
rect 3622 27226 3678 27228
rect 3702 27226 3758 27228
rect 3782 27226 3838 27228
rect 3862 27226 3918 27228
rect 3622 27174 3648 27226
rect 3648 27174 3678 27226
rect 3702 27174 3712 27226
rect 3712 27174 3758 27226
rect 3782 27174 3828 27226
rect 3828 27174 3838 27226
rect 3862 27174 3892 27226
rect 3892 27174 3918 27226
rect 3622 27172 3678 27174
rect 3702 27172 3758 27174
rect 3782 27172 3838 27174
rect 3862 27172 3918 27174
rect 3622 26138 3678 26140
rect 3702 26138 3758 26140
rect 3782 26138 3838 26140
rect 3862 26138 3918 26140
rect 3622 26086 3648 26138
rect 3648 26086 3678 26138
rect 3702 26086 3712 26138
rect 3712 26086 3758 26138
rect 3782 26086 3828 26138
rect 3828 26086 3838 26138
rect 3862 26086 3892 26138
rect 3892 26086 3918 26138
rect 3622 26084 3678 26086
rect 3702 26084 3758 26086
rect 3782 26084 3838 26086
rect 3862 26084 3918 26086
rect 3622 25050 3678 25052
rect 3702 25050 3758 25052
rect 3782 25050 3838 25052
rect 3862 25050 3918 25052
rect 3622 24998 3648 25050
rect 3648 24998 3678 25050
rect 3702 24998 3712 25050
rect 3712 24998 3758 25050
rect 3782 24998 3828 25050
rect 3828 24998 3838 25050
rect 3862 24998 3892 25050
rect 3892 24998 3918 25050
rect 3622 24996 3678 24998
rect 3702 24996 3758 24998
rect 3782 24996 3838 24998
rect 3862 24996 3918 24998
rect 3622 23962 3678 23964
rect 3702 23962 3758 23964
rect 3782 23962 3838 23964
rect 3862 23962 3918 23964
rect 3622 23910 3648 23962
rect 3648 23910 3678 23962
rect 3702 23910 3712 23962
rect 3712 23910 3758 23962
rect 3782 23910 3828 23962
rect 3828 23910 3838 23962
rect 3862 23910 3892 23962
rect 3892 23910 3918 23962
rect 3622 23908 3678 23910
rect 3702 23908 3758 23910
rect 3782 23908 3838 23910
rect 3862 23908 3918 23910
rect 3622 22874 3678 22876
rect 3702 22874 3758 22876
rect 3782 22874 3838 22876
rect 3862 22874 3918 22876
rect 3622 22822 3648 22874
rect 3648 22822 3678 22874
rect 3702 22822 3712 22874
rect 3712 22822 3758 22874
rect 3782 22822 3828 22874
rect 3828 22822 3838 22874
rect 3862 22822 3892 22874
rect 3892 22822 3918 22874
rect 3622 22820 3678 22822
rect 3702 22820 3758 22822
rect 3782 22820 3838 22822
rect 3862 22820 3918 22822
rect 3622 21786 3678 21788
rect 3702 21786 3758 21788
rect 3782 21786 3838 21788
rect 3862 21786 3918 21788
rect 3622 21734 3648 21786
rect 3648 21734 3678 21786
rect 3702 21734 3712 21786
rect 3712 21734 3758 21786
rect 3782 21734 3828 21786
rect 3828 21734 3838 21786
rect 3862 21734 3892 21786
rect 3892 21734 3918 21786
rect 3622 21732 3678 21734
rect 3702 21732 3758 21734
rect 3782 21732 3838 21734
rect 3862 21732 3918 21734
rect 4250 35284 4306 35320
rect 4250 35264 4252 35284
rect 4252 35264 4304 35284
rect 4304 35264 4306 35284
rect 4342 34992 4398 35048
rect 4158 32272 4214 32328
rect 4894 34040 4950 34096
rect 4894 33768 4950 33824
rect 4066 30504 4122 30560
rect 4158 29960 4214 30016
rect 4802 30368 4858 30424
rect 4710 30268 4712 30288
rect 4712 30268 4764 30288
rect 4764 30268 4766 30288
rect 4710 30232 4766 30268
rect 6289 37562 6345 37564
rect 6369 37562 6425 37564
rect 6449 37562 6505 37564
rect 6529 37562 6585 37564
rect 6289 37510 6315 37562
rect 6315 37510 6345 37562
rect 6369 37510 6379 37562
rect 6379 37510 6425 37562
rect 6449 37510 6495 37562
rect 6495 37510 6505 37562
rect 6529 37510 6559 37562
rect 6559 37510 6585 37562
rect 6289 37508 6345 37510
rect 6369 37508 6425 37510
rect 6449 37508 6505 37510
rect 6529 37508 6585 37510
rect 6289 36474 6345 36476
rect 6369 36474 6425 36476
rect 6449 36474 6505 36476
rect 6529 36474 6585 36476
rect 6289 36422 6315 36474
rect 6315 36422 6345 36474
rect 6369 36422 6379 36474
rect 6379 36422 6425 36474
rect 6449 36422 6495 36474
rect 6495 36422 6505 36474
rect 6529 36422 6559 36474
rect 6559 36422 6585 36474
rect 6289 36420 6345 36422
rect 6369 36420 6425 36422
rect 6449 36420 6505 36422
rect 6529 36420 6585 36422
rect 5170 34040 5226 34096
rect 4618 27376 4674 27432
rect 4342 26968 4398 27024
rect 4158 23704 4214 23760
rect 3622 20698 3678 20700
rect 3702 20698 3758 20700
rect 3782 20698 3838 20700
rect 3862 20698 3918 20700
rect 3622 20646 3648 20698
rect 3648 20646 3678 20698
rect 3702 20646 3712 20698
rect 3712 20646 3758 20698
rect 3782 20646 3828 20698
rect 3828 20646 3838 20698
rect 3862 20646 3892 20698
rect 3892 20646 3918 20698
rect 3622 20644 3678 20646
rect 3702 20644 3758 20646
rect 3782 20644 3838 20646
rect 3862 20644 3918 20646
rect 3622 19610 3678 19612
rect 3702 19610 3758 19612
rect 3782 19610 3838 19612
rect 3862 19610 3918 19612
rect 3622 19558 3648 19610
rect 3648 19558 3678 19610
rect 3702 19558 3712 19610
rect 3712 19558 3758 19610
rect 3782 19558 3828 19610
rect 3828 19558 3838 19610
rect 3862 19558 3892 19610
rect 3892 19558 3918 19610
rect 3622 19556 3678 19558
rect 3702 19556 3758 19558
rect 3782 19556 3838 19558
rect 3862 19556 3918 19558
rect 3622 18522 3678 18524
rect 3702 18522 3758 18524
rect 3782 18522 3838 18524
rect 3862 18522 3918 18524
rect 3622 18470 3648 18522
rect 3648 18470 3678 18522
rect 3702 18470 3712 18522
rect 3712 18470 3758 18522
rect 3782 18470 3828 18522
rect 3828 18470 3838 18522
rect 3862 18470 3892 18522
rect 3892 18470 3918 18522
rect 3622 18468 3678 18470
rect 3702 18468 3758 18470
rect 3782 18468 3838 18470
rect 3862 18468 3918 18470
rect 4802 23568 4858 23624
rect 3054 17992 3110 18048
rect 3330 17992 3386 18048
rect 2778 17740 2834 17776
rect 2778 17720 2780 17740
rect 2780 17720 2832 17740
rect 2832 17720 2834 17740
rect 1582 17584 1638 17640
rect 2226 15852 2228 15872
rect 2228 15852 2280 15872
rect 2280 15852 2282 15872
rect 2226 15816 2282 15852
rect 1674 15136 1730 15192
rect 3622 17434 3678 17436
rect 3702 17434 3758 17436
rect 3782 17434 3838 17436
rect 3862 17434 3918 17436
rect 3622 17382 3648 17434
rect 3648 17382 3678 17434
rect 3702 17382 3712 17434
rect 3712 17382 3758 17434
rect 3782 17382 3828 17434
rect 3828 17382 3838 17434
rect 3862 17382 3892 17434
rect 3892 17382 3918 17434
rect 3622 17380 3678 17382
rect 3702 17380 3758 17382
rect 3782 17380 3838 17382
rect 3862 17380 3918 17382
rect 3974 17040 4030 17096
rect 3622 16346 3678 16348
rect 3702 16346 3758 16348
rect 3782 16346 3838 16348
rect 3862 16346 3918 16348
rect 3622 16294 3648 16346
rect 3648 16294 3678 16346
rect 3702 16294 3712 16346
rect 3712 16294 3758 16346
rect 3782 16294 3828 16346
rect 3828 16294 3838 16346
rect 3862 16294 3892 16346
rect 3892 16294 3918 16346
rect 3622 16292 3678 16294
rect 3702 16292 3758 16294
rect 3782 16292 3838 16294
rect 3862 16292 3918 16294
rect 3622 15258 3678 15260
rect 3702 15258 3758 15260
rect 3782 15258 3838 15260
rect 3862 15258 3918 15260
rect 3622 15206 3648 15258
rect 3648 15206 3678 15258
rect 3702 15206 3712 15258
rect 3712 15206 3758 15258
rect 3782 15206 3828 15258
rect 3828 15206 3838 15258
rect 3862 15206 3892 15258
rect 3892 15206 3918 15258
rect 3622 15204 3678 15206
rect 3702 15204 3758 15206
rect 3782 15204 3838 15206
rect 3862 15204 3918 15206
rect 2318 13776 2374 13832
rect 1398 13388 1454 13424
rect 1398 13368 1400 13388
rect 1400 13368 1452 13388
rect 1452 13368 1454 13388
rect 1582 12824 1638 12880
rect 1582 10512 1638 10568
rect 1582 8064 1638 8120
rect 1674 7384 1730 7440
rect 1490 6840 1546 6896
rect 1398 6704 1454 6760
rect 570 4256 626 4312
rect 938 3576 994 3632
rect 1582 5752 1638 5808
rect 2686 12844 2742 12880
rect 2686 12824 2688 12844
rect 2688 12824 2740 12844
rect 2740 12824 2742 12844
rect 3622 14170 3678 14172
rect 3702 14170 3758 14172
rect 3782 14170 3838 14172
rect 3862 14170 3918 14172
rect 3622 14118 3648 14170
rect 3648 14118 3678 14170
rect 3702 14118 3712 14170
rect 3712 14118 3758 14170
rect 3782 14118 3828 14170
rect 3828 14118 3838 14170
rect 3862 14118 3892 14170
rect 3892 14118 3918 14170
rect 3622 14116 3678 14118
rect 3702 14116 3758 14118
rect 3782 14116 3838 14118
rect 3862 14116 3918 14118
rect 3622 13082 3678 13084
rect 3702 13082 3758 13084
rect 3782 13082 3838 13084
rect 3862 13082 3918 13084
rect 3622 13030 3648 13082
rect 3648 13030 3678 13082
rect 3702 13030 3712 13082
rect 3712 13030 3758 13082
rect 3782 13030 3828 13082
rect 3828 13030 3838 13082
rect 3862 13030 3892 13082
rect 3892 13030 3918 13082
rect 3622 13028 3678 13030
rect 3702 13028 3758 13030
rect 3782 13028 3838 13030
rect 3862 13028 3918 13030
rect 2686 8880 2742 8936
rect 2778 8336 2834 8392
rect 2870 6704 2926 6760
rect 2594 6024 2650 6080
rect 1582 3440 1638 3496
rect 1766 2760 1822 2816
rect 2870 4256 2926 4312
rect 2594 2896 2650 2952
rect 3622 11994 3678 11996
rect 3702 11994 3758 11996
rect 3782 11994 3838 11996
rect 3862 11994 3918 11996
rect 3622 11942 3648 11994
rect 3648 11942 3678 11994
rect 3702 11942 3712 11994
rect 3712 11942 3758 11994
rect 3782 11942 3828 11994
rect 3828 11942 3838 11994
rect 3862 11942 3892 11994
rect 3892 11942 3918 11994
rect 3622 11940 3678 11942
rect 3702 11940 3758 11942
rect 3782 11940 3838 11942
rect 3862 11940 3918 11942
rect 3622 10906 3678 10908
rect 3702 10906 3758 10908
rect 3782 10906 3838 10908
rect 3862 10906 3918 10908
rect 3622 10854 3648 10906
rect 3648 10854 3678 10906
rect 3702 10854 3712 10906
rect 3712 10854 3758 10906
rect 3782 10854 3828 10906
rect 3828 10854 3838 10906
rect 3862 10854 3892 10906
rect 3892 10854 3918 10906
rect 3622 10852 3678 10854
rect 3702 10852 3758 10854
rect 3782 10852 3838 10854
rect 3862 10852 3918 10854
rect 3622 9818 3678 9820
rect 3702 9818 3758 9820
rect 3782 9818 3838 9820
rect 3862 9818 3918 9820
rect 3622 9766 3648 9818
rect 3648 9766 3678 9818
rect 3702 9766 3712 9818
rect 3712 9766 3758 9818
rect 3782 9766 3828 9818
rect 3828 9766 3838 9818
rect 3862 9766 3892 9818
rect 3892 9766 3918 9818
rect 3622 9764 3678 9766
rect 3702 9764 3758 9766
rect 3782 9764 3838 9766
rect 3862 9764 3918 9766
rect 4250 9968 4306 10024
rect 3622 8730 3678 8732
rect 3702 8730 3758 8732
rect 3782 8730 3838 8732
rect 3862 8730 3918 8732
rect 3622 8678 3648 8730
rect 3648 8678 3678 8730
rect 3702 8678 3712 8730
rect 3712 8678 3758 8730
rect 3782 8678 3828 8730
rect 3828 8678 3838 8730
rect 3862 8678 3892 8730
rect 3892 8678 3918 8730
rect 3622 8676 3678 8678
rect 3702 8676 3758 8678
rect 3782 8676 3838 8678
rect 3862 8676 3918 8678
rect 3622 7642 3678 7644
rect 3702 7642 3758 7644
rect 3782 7642 3838 7644
rect 3862 7642 3918 7644
rect 3622 7590 3648 7642
rect 3648 7590 3678 7642
rect 3702 7590 3712 7642
rect 3712 7590 3758 7642
rect 3782 7590 3828 7642
rect 3828 7590 3838 7642
rect 3862 7590 3892 7642
rect 3892 7590 3918 7642
rect 3622 7588 3678 7590
rect 3702 7588 3758 7590
rect 3782 7588 3838 7590
rect 3862 7588 3918 7590
rect 3622 6554 3678 6556
rect 3702 6554 3758 6556
rect 3782 6554 3838 6556
rect 3862 6554 3918 6556
rect 3622 6502 3648 6554
rect 3648 6502 3678 6554
rect 3702 6502 3712 6554
rect 3712 6502 3758 6554
rect 3782 6502 3828 6554
rect 3828 6502 3838 6554
rect 3862 6502 3892 6554
rect 3892 6502 3918 6554
rect 3622 6500 3678 6502
rect 3702 6500 3758 6502
rect 3782 6500 3838 6502
rect 3862 6500 3918 6502
rect 4066 5752 4122 5808
rect 3622 5466 3678 5468
rect 3702 5466 3758 5468
rect 3782 5466 3838 5468
rect 3862 5466 3918 5468
rect 3622 5414 3648 5466
rect 3648 5414 3678 5466
rect 3702 5414 3712 5466
rect 3712 5414 3758 5466
rect 3782 5414 3828 5466
rect 3828 5414 3838 5466
rect 3862 5414 3892 5466
rect 3892 5414 3918 5466
rect 3622 5412 3678 5414
rect 3702 5412 3758 5414
rect 3782 5412 3838 5414
rect 3862 5412 3918 5414
rect 3882 4972 3884 4992
rect 3884 4972 3936 4992
rect 3936 4972 3938 4992
rect 3882 4936 3938 4972
rect 3622 4378 3678 4380
rect 3702 4378 3758 4380
rect 3782 4378 3838 4380
rect 3862 4378 3918 4380
rect 3622 4326 3648 4378
rect 3648 4326 3678 4378
rect 3702 4326 3712 4378
rect 3712 4326 3758 4378
rect 3782 4326 3828 4378
rect 3828 4326 3838 4378
rect 3862 4326 3892 4378
rect 3892 4326 3918 4378
rect 3622 4324 3678 4326
rect 3702 4324 3758 4326
rect 3782 4324 3838 4326
rect 3862 4324 3918 4326
rect 3622 3290 3678 3292
rect 3702 3290 3758 3292
rect 3782 3290 3838 3292
rect 3862 3290 3918 3292
rect 3622 3238 3648 3290
rect 3648 3238 3678 3290
rect 3702 3238 3712 3290
rect 3712 3238 3758 3290
rect 3782 3238 3828 3290
rect 3828 3238 3838 3290
rect 3862 3238 3892 3290
rect 3892 3238 3918 3290
rect 3622 3236 3678 3238
rect 3702 3236 3758 3238
rect 3782 3236 3838 3238
rect 3862 3236 3918 3238
rect 4066 2624 4122 2680
rect 2962 2352 3018 2408
rect 2778 1128 2834 1184
rect 3622 2202 3678 2204
rect 3702 2202 3758 2204
rect 3782 2202 3838 2204
rect 3862 2202 3918 2204
rect 3622 2150 3648 2202
rect 3648 2150 3678 2202
rect 3702 2150 3712 2202
rect 3712 2150 3758 2202
rect 3782 2150 3828 2202
rect 3828 2150 3838 2202
rect 3862 2150 3892 2202
rect 3892 2150 3918 2202
rect 3622 2148 3678 2150
rect 3702 2148 3758 2150
rect 3782 2148 3838 2150
rect 3862 2148 3918 2150
rect 3330 1400 3386 1456
rect 4802 22072 4858 22128
rect 5262 31204 5318 31240
rect 5262 31184 5264 31204
rect 5264 31184 5316 31204
rect 5316 31184 5318 31204
rect 5262 30776 5318 30832
rect 5814 34584 5870 34640
rect 5722 32952 5778 33008
rect 5906 34448 5962 34504
rect 5998 34196 6054 34232
rect 5998 34176 6000 34196
rect 6000 34176 6052 34196
rect 6052 34176 6054 34196
rect 6289 35386 6345 35388
rect 6369 35386 6425 35388
rect 6449 35386 6505 35388
rect 6529 35386 6585 35388
rect 6289 35334 6315 35386
rect 6315 35334 6345 35386
rect 6369 35334 6379 35386
rect 6379 35334 6425 35386
rect 6449 35334 6495 35386
rect 6495 35334 6505 35386
rect 6529 35334 6559 35386
rect 6559 35334 6585 35386
rect 6289 35332 6345 35334
rect 6369 35332 6425 35334
rect 6449 35332 6505 35334
rect 6529 35332 6585 35334
rect 6289 34298 6345 34300
rect 6369 34298 6425 34300
rect 6449 34298 6505 34300
rect 6529 34298 6585 34300
rect 6289 34246 6315 34298
rect 6315 34246 6345 34298
rect 6369 34246 6379 34298
rect 6379 34246 6425 34298
rect 6449 34246 6495 34298
rect 6495 34246 6505 34298
rect 6529 34246 6559 34298
rect 6559 34246 6585 34298
rect 6289 34244 6345 34246
rect 6369 34244 6425 34246
rect 6449 34244 6505 34246
rect 6529 34244 6585 34246
rect 6550 33768 6606 33824
rect 5998 33360 6054 33416
rect 5906 32816 5962 32872
rect 5538 30776 5594 30832
rect 5538 28600 5594 28656
rect 5998 30504 6054 30560
rect 5906 29008 5962 29064
rect 5354 24656 5410 24712
rect 5262 23160 5318 23216
rect 5262 23024 5318 23080
rect 4710 19216 4766 19272
rect 5078 19216 5134 19272
rect 4618 12860 4620 12880
rect 4620 12860 4672 12880
rect 4672 12860 4674 12880
rect 4618 12824 4674 12860
rect 4618 12300 4674 12336
rect 4618 12280 4620 12300
rect 4620 12280 4672 12300
rect 4672 12280 4674 12300
rect 4526 10648 4582 10704
rect 5722 18808 5778 18864
rect 6289 33210 6345 33212
rect 6369 33210 6425 33212
rect 6449 33210 6505 33212
rect 6529 33210 6585 33212
rect 6289 33158 6315 33210
rect 6315 33158 6345 33210
rect 6369 33158 6379 33210
rect 6379 33158 6425 33210
rect 6449 33158 6495 33210
rect 6495 33158 6505 33210
rect 6529 33158 6559 33210
rect 6559 33158 6585 33210
rect 6289 33156 6345 33158
rect 6369 33156 6425 33158
rect 6449 33156 6505 33158
rect 6529 33156 6585 33158
rect 6289 32122 6345 32124
rect 6369 32122 6425 32124
rect 6449 32122 6505 32124
rect 6529 32122 6585 32124
rect 6289 32070 6315 32122
rect 6315 32070 6345 32122
rect 6369 32070 6379 32122
rect 6379 32070 6425 32122
rect 6449 32070 6495 32122
rect 6495 32070 6505 32122
rect 6529 32070 6559 32122
rect 6559 32070 6585 32122
rect 6289 32068 6345 32070
rect 6369 32068 6425 32070
rect 6449 32068 6505 32070
rect 6529 32068 6585 32070
rect 6289 31034 6345 31036
rect 6369 31034 6425 31036
rect 6449 31034 6505 31036
rect 6529 31034 6585 31036
rect 6289 30982 6315 31034
rect 6315 30982 6345 31034
rect 6369 30982 6379 31034
rect 6379 30982 6425 31034
rect 6449 30982 6495 31034
rect 6495 30982 6505 31034
rect 6529 30982 6559 31034
rect 6559 30982 6585 31034
rect 6289 30980 6345 30982
rect 6369 30980 6425 30982
rect 6449 30980 6505 30982
rect 6529 30980 6585 30982
rect 6642 30232 6698 30288
rect 6289 29946 6345 29948
rect 6369 29946 6425 29948
rect 6449 29946 6505 29948
rect 6529 29946 6585 29948
rect 6289 29894 6315 29946
rect 6315 29894 6345 29946
rect 6369 29894 6379 29946
rect 6379 29894 6425 29946
rect 6449 29894 6495 29946
rect 6495 29894 6505 29946
rect 6529 29894 6559 29946
rect 6559 29894 6585 29946
rect 6289 29892 6345 29894
rect 6369 29892 6425 29894
rect 6449 29892 6505 29894
rect 6529 29892 6585 29894
rect 6289 28858 6345 28860
rect 6369 28858 6425 28860
rect 6449 28858 6505 28860
rect 6529 28858 6585 28860
rect 6289 28806 6315 28858
rect 6315 28806 6345 28858
rect 6369 28806 6379 28858
rect 6379 28806 6425 28858
rect 6449 28806 6495 28858
rect 6495 28806 6505 28858
rect 6529 28806 6559 28858
rect 6559 28806 6585 28858
rect 6289 28804 6345 28806
rect 6369 28804 6425 28806
rect 6449 28804 6505 28806
rect 6529 28804 6585 28806
rect 6289 27770 6345 27772
rect 6369 27770 6425 27772
rect 6449 27770 6505 27772
rect 6529 27770 6585 27772
rect 6289 27718 6315 27770
rect 6315 27718 6345 27770
rect 6369 27718 6379 27770
rect 6379 27718 6425 27770
rect 6449 27718 6495 27770
rect 6495 27718 6505 27770
rect 6529 27718 6559 27770
rect 6559 27718 6585 27770
rect 6289 27716 6345 27718
rect 6369 27716 6425 27718
rect 6449 27716 6505 27718
rect 6529 27716 6585 27718
rect 7010 34040 7066 34096
rect 7194 34040 7250 34096
rect 7378 33224 7434 33280
rect 6826 30096 6882 30152
rect 6734 28464 6790 28520
rect 6642 26968 6698 27024
rect 6289 26682 6345 26684
rect 6369 26682 6425 26684
rect 6449 26682 6505 26684
rect 6529 26682 6585 26684
rect 6289 26630 6315 26682
rect 6315 26630 6345 26682
rect 6369 26630 6379 26682
rect 6379 26630 6425 26682
rect 6449 26630 6495 26682
rect 6495 26630 6505 26682
rect 6529 26630 6559 26682
rect 6559 26630 6585 26682
rect 6289 26628 6345 26630
rect 6369 26628 6425 26630
rect 6449 26628 6505 26630
rect 6529 26628 6585 26630
rect 6289 25594 6345 25596
rect 6369 25594 6425 25596
rect 6449 25594 6505 25596
rect 6529 25594 6585 25596
rect 6289 25542 6315 25594
rect 6315 25542 6345 25594
rect 6369 25542 6379 25594
rect 6379 25542 6425 25594
rect 6449 25542 6495 25594
rect 6495 25542 6505 25594
rect 6529 25542 6559 25594
rect 6559 25542 6585 25594
rect 6289 25540 6345 25542
rect 6369 25540 6425 25542
rect 6449 25540 6505 25542
rect 6529 25540 6585 25542
rect 6289 24506 6345 24508
rect 6369 24506 6425 24508
rect 6449 24506 6505 24508
rect 6529 24506 6585 24508
rect 6289 24454 6315 24506
rect 6315 24454 6345 24506
rect 6369 24454 6379 24506
rect 6379 24454 6425 24506
rect 6449 24454 6495 24506
rect 6495 24454 6505 24506
rect 6529 24454 6559 24506
rect 6559 24454 6585 24506
rect 6289 24452 6345 24454
rect 6369 24452 6425 24454
rect 6449 24452 6505 24454
rect 6529 24452 6585 24454
rect 5538 15816 5594 15872
rect 5262 13232 5318 13288
rect 5078 10648 5134 10704
rect 4342 6060 4344 6080
rect 4344 6060 4396 6080
rect 4396 6060 4398 6080
rect 4342 6024 4398 6060
rect 4434 5616 4490 5672
rect 4986 7420 4988 7440
rect 4988 7420 5040 7440
rect 5040 7420 5042 7440
rect 4986 7384 5042 7420
rect 5446 13812 5448 13832
rect 5448 13812 5500 13832
rect 5500 13812 5502 13832
rect 5446 13776 5502 13812
rect 5446 12824 5502 12880
rect 6090 20168 6146 20224
rect 5906 16768 5962 16824
rect 6289 23418 6345 23420
rect 6369 23418 6425 23420
rect 6449 23418 6505 23420
rect 6529 23418 6585 23420
rect 6289 23366 6315 23418
rect 6315 23366 6345 23418
rect 6369 23366 6379 23418
rect 6379 23366 6425 23418
rect 6449 23366 6495 23418
rect 6495 23366 6505 23418
rect 6529 23366 6559 23418
rect 6559 23366 6585 23418
rect 6289 23364 6345 23366
rect 6369 23364 6425 23366
rect 6449 23364 6505 23366
rect 6529 23364 6585 23366
rect 6918 23568 6974 23624
rect 7194 30368 7250 30424
rect 7194 27512 7250 27568
rect 7102 23296 7158 23352
rect 6289 22330 6345 22332
rect 6369 22330 6425 22332
rect 6449 22330 6505 22332
rect 6529 22330 6585 22332
rect 6289 22278 6315 22330
rect 6315 22278 6345 22330
rect 6369 22278 6379 22330
rect 6379 22278 6425 22330
rect 6449 22278 6495 22330
rect 6495 22278 6505 22330
rect 6529 22278 6559 22330
rect 6559 22278 6585 22330
rect 6289 22276 6345 22278
rect 6369 22276 6425 22278
rect 6449 22276 6505 22278
rect 6529 22276 6585 22278
rect 6289 21242 6345 21244
rect 6369 21242 6425 21244
rect 6449 21242 6505 21244
rect 6529 21242 6585 21244
rect 6289 21190 6315 21242
rect 6315 21190 6345 21242
rect 6369 21190 6379 21242
rect 6379 21190 6425 21242
rect 6449 21190 6495 21242
rect 6495 21190 6505 21242
rect 6529 21190 6559 21242
rect 6559 21190 6585 21242
rect 6289 21188 6345 21190
rect 6369 21188 6425 21190
rect 6449 21188 6505 21190
rect 6529 21188 6585 21190
rect 6289 20154 6345 20156
rect 6369 20154 6425 20156
rect 6449 20154 6505 20156
rect 6529 20154 6585 20156
rect 6289 20102 6315 20154
rect 6315 20102 6345 20154
rect 6369 20102 6379 20154
rect 6379 20102 6425 20154
rect 6449 20102 6495 20154
rect 6495 20102 6505 20154
rect 6529 20102 6559 20154
rect 6559 20102 6585 20154
rect 6289 20100 6345 20102
rect 6369 20100 6425 20102
rect 6449 20100 6505 20102
rect 6529 20100 6585 20102
rect 6458 19760 6514 19816
rect 6289 19066 6345 19068
rect 6369 19066 6425 19068
rect 6449 19066 6505 19068
rect 6529 19066 6585 19068
rect 6289 19014 6315 19066
rect 6315 19014 6345 19066
rect 6369 19014 6379 19066
rect 6379 19014 6425 19066
rect 6449 19014 6495 19066
rect 6495 19014 6505 19066
rect 6529 19014 6559 19066
rect 6559 19014 6585 19066
rect 6289 19012 6345 19014
rect 6369 19012 6425 19014
rect 6449 19012 6505 19014
rect 6529 19012 6585 19014
rect 6289 17978 6345 17980
rect 6369 17978 6425 17980
rect 6449 17978 6505 17980
rect 6529 17978 6585 17980
rect 6289 17926 6315 17978
rect 6315 17926 6345 17978
rect 6369 17926 6379 17978
rect 6379 17926 6425 17978
rect 6449 17926 6495 17978
rect 6495 17926 6505 17978
rect 6529 17926 6559 17978
rect 6559 17926 6585 17978
rect 6289 17924 6345 17926
rect 6369 17924 6425 17926
rect 6449 17924 6505 17926
rect 6529 17924 6585 17926
rect 6289 16890 6345 16892
rect 6369 16890 6425 16892
rect 6449 16890 6505 16892
rect 6529 16890 6585 16892
rect 6289 16838 6315 16890
rect 6315 16838 6345 16890
rect 6369 16838 6379 16890
rect 6379 16838 6425 16890
rect 6449 16838 6495 16890
rect 6495 16838 6505 16890
rect 6529 16838 6559 16890
rect 6559 16838 6585 16890
rect 6289 16836 6345 16838
rect 6369 16836 6425 16838
rect 6449 16836 6505 16838
rect 6529 16836 6585 16838
rect 6289 15802 6345 15804
rect 6369 15802 6425 15804
rect 6449 15802 6505 15804
rect 6529 15802 6585 15804
rect 6289 15750 6315 15802
rect 6315 15750 6345 15802
rect 6369 15750 6379 15802
rect 6379 15750 6425 15802
rect 6449 15750 6495 15802
rect 6495 15750 6505 15802
rect 6529 15750 6559 15802
rect 6559 15750 6585 15802
rect 6289 15748 6345 15750
rect 6369 15748 6425 15750
rect 6449 15748 6505 15750
rect 6529 15748 6585 15750
rect 6289 14714 6345 14716
rect 6369 14714 6425 14716
rect 6449 14714 6505 14716
rect 6529 14714 6585 14716
rect 6289 14662 6315 14714
rect 6315 14662 6345 14714
rect 6369 14662 6379 14714
rect 6379 14662 6425 14714
rect 6449 14662 6495 14714
rect 6495 14662 6505 14714
rect 6529 14662 6559 14714
rect 6559 14662 6585 14714
rect 6289 14660 6345 14662
rect 6369 14660 6425 14662
rect 6449 14660 6505 14662
rect 6529 14660 6585 14662
rect 5446 8472 5502 8528
rect 6090 13776 6146 13832
rect 6289 13626 6345 13628
rect 6369 13626 6425 13628
rect 6449 13626 6505 13628
rect 6529 13626 6585 13628
rect 6289 13574 6315 13626
rect 6315 13574 6345 13626
rect 6369 13574 6379 13626
rect 6379 13574 6425 13626
rect 6449 13574 6495 13626
rect 6495 13574 6505 13626
rect 6529 13574 6559 13626
rect 6559 13574 6585 13626
rect 6289 13572 6345 13574
rect 6369 13572 6425 13574
rect 6449 13572 6505 13574
rect 6529 13572 6585 13574
rect 5906 12144 5962 12200
rect 4802 5516 4804 5536
rect 4804 5516 4856 5536
rect 4856 5516 4858 5536
rect 4802 5480 4858 5516
rect 5078 4120 5134 4176
rect 4526 2216 4582 2272
rect 5630 6704 5686 6760
rect 5446 5208 5502 5264
rect 5630 2760 5686 2816
rect 5630 2508 5686 2544
rect 5630 2488 5632 2508
rect 5632 2488 5684 2508
rect 5684 2488 5686 2508
rect 5906 7384 5962 7440
rect 5814 5616 5870 5672
rect 6289 12538 6345 12540
rect 6369 12538 6425 12540
rect 6449 12538 6505 12540
rect 6529 12538 6585 12540
rect 6289 12486 6315 12538
rect 6315 12486 6345 12538
rect 6369 12486 6379 12538
rect 6379 12486 6425 12538
rect 6449 12486 6495 12538
rect 6495 12486 6505 12538
rect 6529 12486 6559 12538
rect 6559 12486 6585 12538
rect 6289 12484 6345 12486
rect 6369 12484 6425 12486
rect 6449 12484 6505 12486
rect 6529 12484 6585 12486
rect 6289 11450 6345 11452
rect 6369 11450 6425 11452
rect 6449 11450 6505 11452
rect 6529 11450 6585 11452
rect 6289 11398 6315 11450
rect 6315 11398 6345 11450
rect 6369 11398 6379 11450
rect 6379 11398 6425 11450
rect 6449 11398 6495 11450
rect 6495 11398 6505 11450
rect 6529 11398 6559 11450
rect 6559 11398 6585 11450
rect 6289 11396 6345 11398
rect 6369 11396 6425 11398
rect 6449 11396 6505 11398
rect 6529 11396 6585 11398
rect 6289 10362 6345 10364
rect 6369 10362 6425 10364
rect 6449 10362 6505 10364
rect 6529 10362 6585 10364
rect 6289 10310 6315 10362
rect 6315 10310 6345 10362
rect 6369 10310 6379 10362
rect 6379 10310 6425 10362
rect 6449 10310 6495 10362
rect 6495 10310 6505 10362
rect 6529 10310 6559 10362
rect 6559 10310 6585 10362
rect 6289 10308 6345 10310
rect 6369 10308 6425 10310
rect 6449 10308 6505 10310
rect 6529 10308 6585 10310
rect 7286 22616 7342 22672
rect 7562 32272 7618 32328
rect 7746 32408 7802 32464
rect 8482 34992 8538 35048
rect 8206 32972 8262 33008
rect 8206 32952 8208 32972
rect 8208 32952 8260 32972
rect 8260 32952 8262 32972
rect 7746 28736 7802 28792
rect 7470 24656 7526 24712
rect 7470 23160 7526 23216
rect 7010 19780 7066 19816
rect 7010 19760 7012 19780
rect 7012 19760 7064 19780
rect 7064 19760 7066 19780
rect 6734 18944 6790 19000
rect 7654 20984 7710 21040
rect 7562 19896 7618 19952
rect 7286 19760 7342 19816
rect 7286 18944 7342 19000
rect 7194 18808 7250 18864
rect 7102 18672 7158 18728
rect 6734 16496 6790 16552
rect 6826 12180 6828 12200
rect 6828 12180 6880 12200
rect 6880 12180 6882 12200
rect 6826 12144 6882 12180
rect 6734 11192 6790 11248
rect 7010 11056 7066 11112
rect 6182 9424 6238 9480
rect 6289 9274 6345 9276
rect 6369 9274 6425 9276
rect 6449 9274 6505 9276
rect 6529 9274 6585 9276
rect 6289 9222 6315 9274
rect 6315 9222 6345 9274
rect 6369 9222 6379 9274
rect 6379 9222 6425 9274
rect 6449 9222 6495 9274
rect 6495 9222 6505 9274
rect 6529 9222 6559 9274
rect 6559 9222 6585 9274
rect 6289 9220 6345 9222
rect 6369 9220 6425 9222
rect 6449 9220 6505 9222
rect 6529 9220 6585 9222
rect 6289 8186 6345 8188
rect 6369 8186 6425 8188
rect 6449 8186 6505 8188
rect 6529 8186 6585 8188
rect 6289 8134 6315 8186
rect 6315 8134 6345 8186
rect 6369 8134 6379 8186
rect 6379 8134 6425 8186
rect 6449 8134 6495 8186
rect 6495 8134 6505 8186
rect 6529 8134 6559 8186
rect 6559 8134 6585 8186
rect 6289 8132 6345 8134
rect 6369 8132 6425 8134
rect 6449 8132 6505 8134
rect 6529 8132 6585 8134
rect 6289 7098 6345 7100
rect 6369 7098 6425 7100
rect 6449 7098 6505 7100
rect 6529 7098 6585 7100
rect 6289 7046 6315 7098
rect 6315 7046 6345 7098
rect 6369 7046 6379 7098
rect 6379 7046 6425 7098
rect 6449 7046 6495 7098
rect 6495 7046 6505 7098
rect 6529 7046 6559 7098
rect 6559 7046 6585 7098
rect 6289 7044 6345 7046
rect 6369 7044 6425 7046
rect 6449 7044 6505 7046
rect 6529 7044 6585 7046
rect 6289 6010 6345 6012
rect 6369 6010 6425 6012
rect 6449 6010 6505 6012
rect 6529 6010 6585 6012
rect 6289 5958 6315 6010
rect 6315 5958 6345 6010
rect 6369 5958 6379 6010
rect 6379 5958 6425 6010
rect 6449 5958 6495 6010
rect 6495 5958 6505 6010
rect 6529 5958 6559 6010
rect 6559 5958 6585 6010
rect 6289 5956 6345 5958
rect 6369 5956 6425 5958
rect 6449 5956 6505 5958
rect 6529 5956 6585 5958
rect 6274 5752 6330 5808
rect 6826 6840 6882 6896
rect 6182 5616 6238 5672
rect 6289 4922 6345 4924
rect 6369 4922 6425 4924
rect 6449 4922 6505 4924
rect 6529 4922 6585 4924
rect 6289 4870 6315 4922
rect 6315 4870 6345 4922
rect 6369 4870 6379 4922
rect 6379 4870 6425 4922
rect 6449 4870 6495 4922
rect 6495 4870 6505 4922
rect 6529 4870 6559 4922
rect 6559 4870 6585 4922
rect 6289 4868 6345 4870
rect 6369 4868 6425 4870
rect 6449 4868 6505 4870
rect 6529 4868 6585 4870
rect 6274 4664 6330 4720
rect 6182 3984 6238 4040
rect 5998 2624 6054 2680
rect 6289 3834 6345 3836
rect 6369 3834 6425 3836
rect 6449 3834 6505 3836
rect 6529 3834 6585 3836
rect 6289 3782 6315 3834
rect 6315 3782 6345 3834
rect 6369 3782 6379 3834
rect 6379 3782 6425 3834
rect 6449 3782 6495 3834
rect 6495 3782 6505 3834
rect 6529 3782 6559 3834
rect 6559 3782 6585 3834
rect 6289 3780 6345 3782
rect 6369 3780 6425 3782
rect 6449 3780 6505 3782
rect 6529 3780 6585 3782
rect 6642 3440 6698 3496
rect 7378 11736 7434 11792
rect 6826 3712 6882 3768
rect 6289 2746 6345 2748
rect 6369 2746 6425 2748
rect 6449 2746 6505 2748
rect 6529 2746 6585 2748
rect 6289 2694 6315 2746
rect 6315 2694 6345 2746
rect 6369 2694 6379 2746
rect 6379 2694 6425 2746
rect 6449 2694 6495 2746
rect 6495 2694 6505 2746
rect 6529 2694 6559 2746
rect 6559 2694 6585 2746
rect 6289 2692 6345 2694
rect 6369 2692 6425 2694
rect 6449 2692 6505 2694
rect 6529 2692 6585 2694
rect 7194 7948 7250 7984
rect 7194 7928 7196 7948
rect 7196 7928 7248 7948
rect 7248 7928 7250 7948
rect 8574 34448 8630 34504
rect 8956 37018 9012 37020
rect 9036 37018 9092 37020
rect 9116 37018 9172 37020
rect 9196 37018 9252 37020
rect 8956 36966 8982 37018
rect 8982 36966 9012 37018
rect 9036 36966 9046 37018
rect 9046 36966 9092 37018
rect 9116 36966 9162 37018
rect 9162 36966 9172 37018
rect 9196 36966 9226 37018
rect 9226 36966 9252 37018
rect 8956 36964 9012 36966
rect 9036 36964 9092 36966
rect 9116 36964 9172 36966
rect 9196 36964 9252 36966
rect 8956 35930 9012 35932
rect 9036 35930 9092 35932
rect 9116 35930 9172 35932
rect 9196 35930 9252 35932
rect 8956 35878 8982 35930
rect 8982 35878 9012 35930
rect 9036 35878 9046 35930
rect 9046 35878 9092 35930
rect 9116 35878 9162 35930
rect 9162 35878 9172 35930
rect 9196 35878 9226 35930
rect 9226 35878 9252 35930
rect 8956 35876 9012 35878
rect 9036 35876 9092 35878
rect 9116 35876 9172 35878
rect 9196 35876 9252 35878
rect 8850 35128 8906 35184
rect 8956 34842 9012 34844
rect 9036 34842 9092 34844
rect 9116 34842 9172 34844
rect 9196 34842 9252 34844
rect 8956 34790 8982 34842
rect 8982 34790 9012 34842
rect 9036 34790 9046 34842
rect 9046 34790 9092 34842
rect 9116 34790 9162 34842
rect 9162 34790 9172 34842
rect 9196 34790 9226 34842
rect 9226 34790 9252 34842
rect 8956 34788 9012 34790
rect 9036 34788 9092 34790
rect 9116 34788 9172 34790
rect 9196 34788 9252 34790
rect 9862 35708 9864 35728
rect 9864 35708 9916 35728
rect 9916 35708 9918 35728
rect 9862 35672 9918 35708
rect 9770 34584 9826 34640
rect 8956 33754 9012 33756
rect 9036 33754 9092 33756
rect 9116 33754 9172 33756
rect 9196 33754 9252 33756
rect 8956 33702 8982 33754
rect 8982 33702 9012 33754
rect 9036 33702 9046 33754
rect 9046 33702 9092 33754
rect 9116 33702 9162 33754
rect 9162 33702 9172 33754
rect 9196 33702 9226 33754
rect 9226 33702 9252 33754
rect 8956 33700 9012 33702
rect 9036 33700 9092 33702
rect 9116 33700 9172 33702
rect 9196 33700 9252 33702
rect 9310 33532 9312 33552
rect 9312 33532 9364 33552
rect 9364 33532 9366 33552
rect 9310 33496 9366 33532
rect 8758 33360 8814 33416
rect 8666 32816 8722 32872
rect 8482 30776 8538 30832
rect 8022 24792 8078 24848
rect 7930 24248 7986 24304
rect 8206 22072 8262 22128
rect 8956 32666 9012 32668
rect 9036 32666 9092 32668
rect 9116 32666 9172 32668
rect 9196 32666 9252 32668
rect 8956 32614 8982 32666
rect 8982 32614 9012 32666
rect 9036 32614 9046 32666
rect 9046 32614 9092 32666
rect 9116 32614 9162 32666
rect 9162 32614 9172 32666
rect 9196 32614 9226 32666
rect 9226 32614 9252 32666
rect 8956 32612 9012 32614
rect 9036 32612 9092 32614
rect 9116 32612 9172 32614
rect 9196 32612 9252 32614
rect 8956 31578 9012 31580
rect 9036 31578 9092 31580
rect 9116 31578 9172 31580
rect 9196 31578 9252 31580
rect 8956 31526 8982 31578
rect 8982 31526 9012 31578
rect 9036 31526 9046 31578
rect 9046 31526 9092 31578
rect 9116 31526 9162 31578
rect 9162 31526 9172 31578
rect 9196 31526 9226 31578
rect 9226 31526 9252 31578
rect 8956 31524 9012 31526
rect 9036 31524 9092 31526
rect 9116 31524 9172 31526
rect 9196 31524 9252 31526
rect 9678 32816 9734 32872
rect 9494 32680 9550 32736
rect 9678 32292 9734 32328
rect 9678 32272 9680 32292
rect 9680 32272 9732 32292
rect 9732 32272 9734 32292
rect 9310 31320 9366 31376
rect 9586 31084 9588 31104
rect 9588 31084 9640 31104
rect 9640 31084 9642 31104
rect 9586 31048 9642 31084
rect 8956 30490 9012 30492
rect 9036 30490 9092 30492
rect 9116 30490 9172 30492
rect 9196 30490 9252 30492
rect 8956 30438 8982 30490
rect 8982 30438 9012 30490
rect 9036 30438 9046 30490
rect 9046 30438 9092 30490
rect 9116 30438 9162 30490
rect 9162 30438 9172 30490
rect 9196 30438 9226 30490
rect 9226 30438 9252 30490
rect 8956 30436 9012 30438
rect 9036 30436 9092 30438
rect 9116 30436 9172 30438
rect 9196 30436 9252 30438
rect 8956 29402 9012 29404
rect 9036 29402 9092 29404
rect 9116 29402 9172 29404
rect 9196 29402 9252 29404
rect 8956 29350 8982 29402
rect 8982 29350 9012 29402
rect 9036 29350 9046 29402
rect 9046 29350 9092 29402
rect 9116 29350 9162 29402
rect 9162 29350 9172 29402
rect 9196 29350 9226 29402
rect 9226 29350 9252 29402
rect 8956 29348 9012 29350
rect 9036 29348 9092 29350
rect 9116 29348 9172 29350
rect 9196 29348 9252 29350
rect 9862 31340 9918 31376
rect 9862 31320 9864 31340
rect 9864 31320 9916 31340
rect 9916 31320 9918 31340
rect 9586 28600 9642 28656
rect 8850 28464 8906 28520
rect 8956 28314 9012 28316
rect 9036 28314 9092 28316
rect 9116 28314 9172 28316
rect 9196 28314 9252 28316
rect 8956 28262 8982 28314
rect 8982 28262 9012 28314
rect 9036 28262 9046 28314
rect 9046 28262 9092 28314
rect 9116 28262 9162 28314
rect 9162 28262 9172 28314
rect 9196 28262 9226 28314
rect 9226 28262 9252 28314
rect 8956 28260 9012 28262
rect 9036 28260 9092 28262
rect 9116 28260 9172 28262
rect 9196 28260 9252 28262
rect 9494 28056 9550 28112
rect 9310 27648 9366 27704
rect 8956 27226 9012 27228
rect 9036 27226 9092 27228
rect 9116 27226 9172 27228
rect 9196 27226 9252 27228
rect 8956 27174 8982 27226
rect 8982 27174 9012 27226
rect 9036 27174 9046 27226
rect 9046 27174 9092 27226
rect 9116 27174 9162 27226
rect 9162 27174 9172 27226
rect 9196 27174 9226 27226
rect 9226 27174 9252 27226
rect 8956 27172 9012 27174
rect 9036 27172 9092 27174
rect 9116 27172 9172 27174
rect 9196 27172 9252 27174
rect 8956 26138 9012 26140
rect 9036 26138 9092 26140
rect 9116 26138 9172 26140
rect 9196 26138 9252 26140
rect 8956 26086 8982 26138
rect 8982 26086 9012 26138
rect 9036 26086 9046 26138
rect 9046 26086 9092 26138
rect 9116 26086 9162 26138
rect 9162 26086 9172 26138
rect 9196 26086 9226 26138
rect 9226 26086 9252 26138
rect 8956 26084 9012 26086
rect 9036 26084 9092 26086
rect 9116 26084 9172 26086
rect 9196 26084 9252 26086
rect 8758 25336 8814 25392
rect 8956 25050 9012 25052
rect 9036 25050 9092 25052
rect 9116 25050 9172 25052
rect 9196 25050 9252 25052
rect 8956 24998 8982 25050
rect 8982 24998 9012 25050
rect 9036 24998 9046 25050
rect 9046 24998 9092 25050
rect 9116 24998 9162 25050
rect 9162 24998 9172 25050
rect 9196 24998 9226 25050
rect 9226 24998 9252 25050
rect 8956 24996 9012 24998
rect 9036 24996 9092 24998
rect 9116 24996 9172 24998
rect 9196 24996 9252 24998
rect 9402 24928 9458 24984
rect 8956 23962 9012 23964
rect 9036 23962 9092 23964
rect 9116 23962 9172 23964
rect 9196 23962 9252 23964
rect 8956 23910 8982 23962
rect 8982 23910 9012 23962
rect 9036 23910 9046 23962
rect 9046 23910 9092 23962
rect 9116 23910 9162 23962
rect 9162 23910 9172 23962
rect 9196 23910 9226 23962
rect 9226 23910 9252 23962
rect 8956 23908 9012 23910
rect 9036 23908 9092 23910
rect 9116 23908 9172 23910
rect 9196 23908 9252 23910
rect 8850 23740 8852 23760
rect 8852 23740 8904 23760
rect 8904 23740 8906 23760
rect 8850 23704 8906 23740
rect 8956 22874 9012 22876
rect 9036 22874 9092 22876
rect 9116 22874 9172 22876
rect 9196 22874 9252 22876
rect 8956 22822 8982 22874
rect 8982 22822 9012 22874
rect 9036 22822 9046 22874
rect 9046 22822 9092 22874
rect 9116 22822 9162 22874
rect 9162 22822 9172 22874
rect 9196 22822 9226 22874
rect 9226 22822 9252 22874
rect 8956 22820 9012 22822
rect 9036 22820 9092 22822
rect 9116 22820 9172 22822
rect 9196 22820 9252 22822
rect 8956 21786 9012 21788
rect 9036 21786 9092 21788
rect 9116 21786 9172 21788
rect 9196 21786 9252 21788
rect 8956 21734 8982 21786
rect 8982 21734 9012 21786
rect 9036 21734 9046 21786
rect 9046 21734 9092 21786
rect 9116 21734 9162 21786
rect 9162 21734 9172 21786
rect 9196 21734 9226 21786
rect 9226 21734 9252 21786
rect 8956 21732 9012 21734
rect 9036 21732 9092 21734
rect 9116 21732 9172 21734
rect 9196 21732 9252 21734
rect 8022 18128 8078 18184
rect 8956 20698 9012 20700
rect 9036 20698 9092 20700
rect 9116 20698 9172 20700
rect 9196 20698 9252 20700
rect 8956 20646 8982 20698
rect 8982 20646 9012 20698
rect 9036 20646 9046 20698
rect 9046 20646 9092 20698
rect 9116 20646 9162 20698
rect 9162 20646 9172 20698
rect 9196 20646 9226 20698
rect 9226 20646 9252 20698
rect 8956 20644 9012 20646
rect 9036 20644 9092 20646
rect 9116 20644 9172 20646
rect 9196 20644 9252 20646
rect 8666 19352 8722 19408
rect 8956 19610 9012 19612
rect 9036 19610 9092 19612
rect 9116 19610 9172 19612
rect 9196 19610 9252 19612
rect 8956 19558 8982 19610
rect 8982 19558 9012 19610
rect 9036 19558 9046 19610
rect 9046 19558 9092 19610
rect 9116 19558 9162 19610
rect 9162 19558 9172 19610
rect 9196 19558 9226 19610
rect 9226 19558 9252 19610
rect 8956 19556 9012 19558
rect 9036 19556 9092 19558
rect 9116 19556 9172 19558
rect 9196 19556 9252 19558
rect 8390 18944 8446 19000
rect 8390 18128 8446 18184
rect 8298 15816 8354 15872
rect 8114 15136 8170 15192
rect 8114 14864 8170 14920
rect 8114 13776 8170 13832
rect 8666 15136 8722 15192
rect 8298 12552 8354 12608
rect 8850 19236 8906 19272
rect 8850 19216 8852 19236
rect 8852 19216 8904 19236
rect 8904 19216 8906 19236
rect 9402 23024 9458 23080
rect 8956 18522 9012 18524
rect 9036 18522 9092 18524
rect 9116 18522 9172 18524
rect 9196 18522 9252 18524
rect 8956 18470 8982 18522
rect 8982 18470 9012 18522
rect 9036 18470 9046 18522
rect 9046 18470 9092 18522
rect 9116 18470 9162 18522
rect 9162 18470 9172 18522
rect 9196 18470 9226 18522
rect 9226 18470 9252 18522
rect 8956 18468 9012 18470
rect 9036 18468 9092 18470
rect 9116 18468 9172 18470
rect 9196 18468 9252 18470
rect 8956 17434 9012 17436
rect 9036 17434 9092 17436
rect 9116 17434 9172 17436
rect 9196 17434 9252 17436
rect 8956 17382 8982 17434
rect 8982 17382 9012 17434
rect 9036 17382 9046 17434
rect 9046 17382 9092 17434
rect 9116 17382 9162 17434
rect 9162 17382 9172 17434
rect 9196 17382 9226 17434
rect 9226 17382 9252 17434
rect 8956 17380 9012 17382
rect 9036 17380 9092 17382
rect 9116 17380 9172 17382
rect 9196 17380 9252 17382
rect 8956 16346 9012 16348
rect 9036 16346 9092 16348
rect 9116 16346 9172 16348
rect 9196 16346 9252 16348
rect 8956 16294 8982 16346
rect 8982 16294 9012 16346
rect 9036 16294 9046 16346
rect 9046 16294 9092 16346
rect 9116 16294 9162 16346
rect 9162 16294 9172 16346
rect 9196 16294 9226 16346
rect 9226 16294 9252 16346
rect 8956 16292 9012 16294
rect 9036 16292 9092 16294
rect 9116 16292 9172 16294
rect 9196 16292 9252 16294
rect 9218 16108 9274 16144
rect 9218 16088 9220 16108
rect 9220 16088 9272 16108
rect 9272 16088 9274 16108
rect 8850 15852 8852 15872
rect 8852 15852 8904 15872
rect 8904 15852 8906 15872
rect 8850 15816 8906 15852
rect 8956 15258 9012 15260
rect 9036 15258 9092 15260
rect 9116 15258 9172 15260
rect 9196 15258 9252 15260
rect 8956 15206 8982 15258
rect 8982 15206 9012 15258
rect 9036 15206 9046 15258
rect 9046 15206 9092 15258
rect 9116 15206 9162 15258
rect 9162 15206 9172 15258
rect 9196 15206 9226 15258
rect 9226 15206 9252 15258
rect 8956 15204 9012 15206
rect 9036 15204 9092 15206
rect 9116 15204 9172 15206
rect 9196 15204 9252 15206
rect 8666 12552 8722 12608
rect 8482 12144 8538 12200
rect 7378 5616 7434 5672
rect 7194 4664 7250 4720
rect 7102 3732 7158 3768
rect 7102 3712 7104 3732
rect 7104 3712 7156 3732
rect 7156 3712 7158 3732
rect 7010 3576 7066 3632
rect 7010 2896 7066 2952
rect 7102 1400 7158 1456
rect 7470 4936 7526 4992
rect 7746 9424 7802 9480
rect 8666 11056 8722 11112
rect 8956 14170 9012 14172
rect 9036 14170 9092 14172
rect 9116 14170 9172 14172
rect 9196 14170 9252 14172
rect 8956 14118 8982 14170
rect 8982 14118 9012 14170
rect 9036 14118 9046 14170
rect 9046 14118 9092 14170
rect 9116 14118 9162 14170
rect 9162 14118 9172 14170
rect 9196 14118 9226 14170
rect 9226 14118 9252 14170
rect 8956 14116 9012 14118
rect 9036 14116 9092 14118
rect 9116 14116 9172 14118
rect 9196 14116 9252 14118
rect 8942 13232 8998 13288
rect 9310 13232 9366 13288
rect 8956 13082 9012 13084
rect 9036 13082 9092 13084
rect 9116 13082 9172 13084
rect 9196 13082 9252 13084
rect 8956 13030 8982 13082
rect 8982 13030 9012 13082
rect 9036 13030 9046 13082
rect 9046 13030 9092 13082
rect 9116 13030 9162 13082
rect 9162 13030 9172 13082
rect 9196 13030 9226 13082
rect 9226 13030 9252 13082
rect 8956 13028 9012 13030
rect 9036 13028 9092 13030
rect 9116 13028 9172 13030
rect 9196 13028 9252 13030
rect 8482 9968 8538 10024
rect 8206 8508 8208 8528
rect 8208 8508 8260 8528
rect 8260 8508 8262 8528
rect 8206 8472 8262 8508
rect 7838 4528 7894 4584
rect 8022 4256 8078 4312
rect 8758 10376 8814 10432
rect 8574 7248 8630 7304
rect 8574 4800 8630 4856
rect 8574 4120 8630 4176
rect 8482 3984 8538 4040
rect 8298 3032 8354 3088
rect 8298 2760 8354 2816
rect 8022 2216 8078 2272
rect 8956 11994 9012 11996
rect 9036 11994 9092 11996
rect 9116 11994 9172 11996
rect 9196 11994 9252 11996
rect 8956 11942 8982 11994
rect 8982 11942 9012 11994
rect 9036 11942 9046 11994
rect 9046 11942 9092 11994
rect 9116 11942 9162 11994
rect 9162 11942 9172 11994
rect 9196 11942 9226 11994
rect 9226 11942 9252 11994
rect 8956 11940 9012 11942
rect 9036 11940 9092 11942
rect 9116 11940 9172 11942
rect 9196 11940 9252 11942
rect 9402 11212 9458 11248
rect 9402 11192 9404 11212
rect 9404 11192 9456 11212
rect 9456 11192 9458 11212
rect 8956 10906 9012 10908
rect 9036 10906 9092 10908
rect 9116 10906 9172 10908
rect 9196 10906 9252 10908
rect 8956 10854 8982 10906
rect 8982 10854 9012 10906
rect 9036 10854 9046 10906
rect 9046 10854 9092 10906
rect 9116 10854 9162 10906
rect 9162 10854 9172 10906
rect 9196 10854 9226 10906
rect 9226 10854 9252 10906
rect 8956 10852 9012 10854
rect 9036 10852 9092 10854
rect 9116 10852 9172 10854
rect 9196 10852 9252 10854
rect 8956 9818 9012 9820
rect 9036 9818 9092 9820
rect 9116 9818 9172 9820
rect 9196 9818 9252 9820
rect 8956 9766 8982 9818
rect 8982 9766 9012 9818
rect 9036 9766 9046 9818
rect 9046 9766 9092 9818
rect 9116 9766 9162 9818
rect 9162 9766 9172 9818
rect 9196 9766 9226 9818
rect 9226 9766 9252 9818
rect 8956 9764 9012 9766
rect 9036 9764 9092 9766
rect 9116 9764 9172 9766
rect 9196 9764 9252 9766
rect 8956 8730 9012 8732
rect 9036 8730 9092 8732
rect 9116 8730 9172 8732
rect 9196 8730 9252 8732
rect 8956 8678 8982 8730
rect 8982 8678 9012 8730
rect 9036 8678 9046 8730
rect 9046 8678 9092 8730
rect 9116 8678 9162 8730
rect 9162 8678 9172 8730
rect 9196 8678 9226 8730
rect 9226 8678 9252 8730
rect 8956 8676 9012 8678
rect 9036 8676 9092 8678
rect 9116 8676 9172 8678
rect 9196 8676 9252 8678
rect 9310 8200 9366 8256
rect 9310 8064 9366 8120
rect 8956 7642 9012 7644
rect 9036 7642 9092 7644
rect 9116 7642 9172 7644
rect 9196 7642 9252 7644
rect 8956 7590 8982 7642
rect 8982 7590 9012 7642
rect 9036 7590 9046 7642
rect 9046 7590 9092 7642
rect 9116 7590 9162 7642
rect 9162 7590 9172 7642
rect 9196 7590 9226 7642
rect 9226 7590 9252 7642
rect 8956 7588 9012 7590
rect 9036 7588 9092 7590
rect 9116 7588 9172 7590
rect 9196 7588 9252 7590
rect 8956 6554 9012 6556
rect 9036 6554 9092 6556
rect 9116 6554 9172 6556
rect 9196 6554 9252 6556
rect 8956 6502 8982 6554
rect 8982 6502 9012 6554
rect 9036 6502 9046 6554
rect 9046 6502 9092 6554
rect 9116 6502 9162 6554
rect 9162 6502 9172 6554
rect 9196 6502 9226 6554
rect 9226 6502 9252 6554
rect 8956 6500 9012 6502
rect 9036 6500 9092 6502
rect 9116 6500 9172 6502
rect 9196 6500 9252 6502
rect 9954 27376 10010 27432
rect 10322 34040 10378 34096
rect 10230 32000 10286 32056
rect 10230 30912 10286 30968
rect 10506 34448 10562 34504
rect 10506 33088 10562 33144
rect 10506 31864 10562 31920
rect 10230 30232 10286 30288
rect 9954 25372 9956 25392
rect 9956 25372 10008 25392
rect 10008 25372 10010 25392
rect 9954 25336 10010 25372
rect 9862 24928 9918 24984
rect 9678 20304 9734 20360
rect 9678 19760 9734 19816
rect 9678 17720 9734 17776
rect 9678 13368 9734 13424
rect 9586 12144 9642 12200
rect 9678 10648 9734 10704
rect 9678 10412 9680 10432
rect 9680 10412 9732 10432
rect 9732 10412 9734 10432
rect 9678 10376 9734 10412
rect 9586 8880 9642 8936
rect 9402 6296 9458 6352
rect 10690 33088 10746 33144
rect 10690 32680 10746 32736
rect 10782 30268 10784 30288
rect 10784 30268 10836 30288
rect 10836 30268 10838 30288
rect 10782 30232 10838 30268
rect 10782 29688 10838 29744
rect 11242 33224 11298 33280
rect 11150 31048 11206 31104
rect 11150 30368 11206 30424
rect 11058 29008 11114 29064
rect 10598 24248 10654 24304
rect 9954 17040 10010 17096
rect 11242 29008 11298 29064
rect 11622 37562 11678 37564
rect 11702 37562 11758 37564
rect 11782 37562 11838 37564
rect 11862 37562 11918 37564
rect 11622 37510 11648 37562
rect 11648 37510 11678 37562
rect 11702 37510 11712 37562
rect 11712 37510 11758 37562
rect 11782 37510 11828 37562
rect 11828 37510 11838 37562
rect 11862 37510 11892 37562
rect 11892 37510 11918 37562
rect 11622 37508 11678 37510
rect 11702 37508 11758 37510
rect 11782 37508 11838 37510
rect 11862 37508 11918 37510
rect 11622 36474 11678 36476
rect 11702 36474 11758 36476
rect 11782 36474 11838 36476
rect 11862 36474 11918 36476
rect 11622 36422 11648 36474
rect 11648 36422 11678 36474
rect 11702 36422 11712 36474
rect 11712 36422 11758 36474
rect 11782 36422 11828 36474
rect 11828 36422 11838 36474
rect 11862 36422 11892 36474
rect 11892 36422 11918 36474
rect 11622 36420 11678 36422
rect 11702 36420 11758 36422
rect 11782 36420 11838 36422
rect 11862 36420 11918 36422
rect 11622 35386 11678 35388
rect 11702 35386 11758 35388
rect 11782 35386 11838 35388
rect 11862 35386 11918 35388
rect 11622 35334 11648 35386
rect 11648 35334 11678 35386
rect 11702 35334 11712 35386
rect 11712 35334 11758 35386
rect 11782 35334 11828 35386
rect 11828 35334 11838 35386
rect 11862 35334 11892 35386
rect 11892 35334 11918 35386
rect 11622 35332 11678 35334
rect 11702 35332 11758 35334
rect 11782 35332 11838 35334
rect 11862 35332 11918 35334
rect 11622 34298 11678 34300
rect 11702 34298 11758 34300
rect 11782 34298 11838 34300
rect 11862 34298 11918 34300
rect 11622 34246 11648 34298
rect 11648 34246 11678 34298
rect 11702 34246 11712 34298
rect 11712 34246 11758 34298
rect 11782 34246 11828 34298
rect 11828 34246 11838 34298
rect 11862 34246 11892 34298
rect 11892 34246 11918 34298
rect 11622 34244 11678 34246
rect 11702 34244 11758 34246
rect 11782 34244 11838 34246
rect 11862 34244 11918 34246
rect 12254 34040 12310 34096
rect 11334 28192 11390 28248
rect 11622 33210 11678 33212
rect 11702 33210 11758 33212
rect 11782 33210 11838 33212
rect 11862 33210 11918 33212
rect 11622 33158 11648 33210
rect 11648 33158 11678 33210
rect 11702 33158 11712 33210
rect 11712 33158 11758 33210
rect 11782 33158 11828 33210
rect 11828 33158 11838 33210
rect 11862 33158 11892 33210
rect 11892 33158 11918 33210
rect 11622 33156 11678 33158
rect 11702 33156 11758 33158
rect 11782 33156 11838 33158
rect 11862 33156 11918 33158
rect 12438 33904 12494 33960
rect 12990 34992 13046 35048
rect 11622 32122 11678 32124
rect 11702 32122 11758 32124
rect 11782 32122 11838 32124
rect 11862 32122 11918 32124
rect 11622 32070 11648 32122
rect 11648 32070 11678 32122
rect 11702 32070 11712 32122
rect 11712 32070 11758 32122
rect 11782 32070 11828 32122
rect 11828 32070 11838 32122
rect 11862 32070 11892 32122
rect 11892 32070 11918 32122
rect 11622 32068 11678 32070
rect 11702 32068 11758 32070
rect 11782 32068 11838 32070
rect 11862 32068 11918 32070
rect 11622 31034 11678 31036
rect 11702 31034 11758 31036
rect 11782 31034 11838 31036
rect 11862 31034 11918 31036
rect 11622 30982 11648 31034
rect 11648 30982 11678 31034
rect 11702 30982 11712 31034
rect 11712 30982 11758 31034
rect 11782 30982 11828 31034
rect 11828 30982 11838 31034
rect 11862 30982 11892 31034
rect 11892 30982 11918 31034
rect 11622 30980 11678 30982
rect 11702 30980 11758 30982
rect 11782 30980 11838 30982
rect 11862 30980 11918 30982
rect 12254 30368 12310 30424
rect 11622 29946 11678 29948
rect 11702 29946 11758 29948
rect 11782 29946 11838 29948
rect 11862 29946 11918 29948
rect 11622 29894 11648 29946
rect 11648 29894 11678 29946
rect 11702 29894 11712 29946
rect 11712 29894 11758 29946
rect 11782 29894 11828 29946
rect 11828 29894 11838 29946
rect 11862 29894 11892 29946
rect 11892 29894 11918 29946
rect 11622 29892 11678 29894
rect 11702 29892 11758 29894
rect 11782 29892 11838 29894
rect 11862 29892 11918 29894
rect 11886 29552 11942 29608
rect 11622 28858 11678 28860
rect 11702 28858 11758 28860
rect 11782 28858 11838 28860
rect 11862 28858 11918 28860
rect 11622 28806 11648 28858
rect 11648 28806 11678 28858
rect 11702 28806 11712 28858
rect 11712 28806 11758 28858
rect 11782 28806 11828 28858
rect 11828 28806 11838 28858
rect 11862 28806 11892 28858
rect 11892 28806 11918 28858
rect 11622 28804 11678 28806
rect 11702 28804 11758 28806
rect 11782 28804 11838 28806
rect 11862 28804 11918 28806
rect 11518 28600 11574 28656
rect 12070 28756 12126 28792
rect 12070 28736 12072 28756
rect 12072 28736 12124 28756
rect 12124 28736 12126 28756
rect 11150 27648 11206 27704
rect 10782 15816 10838 15872
rect 10230 12416 10286 12472
rect 10046 12280 10102 12336
rect 10230 12280 10286 12336
rect 10046 11464 10102 11520
rect 9954 8336 10010 8392
rect 9862 7792 9918 7848
rect 9310 5752 9366 5808
rect 8956 5466 9012 5468
rect 9036 5466 9092 5468
rect 9116 5466 9172 5468
rect 9196 5466 9252 5468
rect 8956 5414 8982 5466
rect 8982 5414 9012 5466
rect 9036 5414 9046 5466
rect 9046 5414 9092 5466
rect 9116 5414 9162 5466
rect 9162 5414 9172 5466
rect 9196 5414 9226 5466
rect 9226 5414 9252 5466
rect 8956 5412 9012 5414
rect 9036 5412 9092 5414
rect 9116 5412 9172 5414
rect 9196 5412 9252 5414
rect 8956 4378 9012 4380
rect 9036 4378 9092 4380
rect 9116 4378 9172 4380
rect 9196 4378 9252 4380
rect 8956 4326 8982 4378
rect 8982 4326 9012 4378
rect 9036 4326 9046 4378
rect 9046 4326 9092 4378
rect 9116 4326 9162 4378
rect 9162 4326 9172 4378
rect 9196 4326 9226 4378
rect 9226 4326 9252 4378
rect 8956 4324 9012 4326
rect 9036 4324 9092 4326
rect 9116 4324 9172 4326
rect 9196 4324 9252 4326
rect 8956 3290 9012 3292
rect 9036 3290 9092 3292
rect 9116 3290 9172 3292
rect 9196 3290 9252 3292
rect 8956 3238 8982 3290
rect 8982 3238 9012 3290
rect 9036 3238 9046 3290
rect 9046 3238 9092 3290
rect 9116 3238 9162 3290
rect 9162 3238 9172 3290
rect 9196 3238 9226 3290
rect 9226 3238 9252 3290
rect 8956 3236 9012 3238
rect 9036 3236 9092 3238
rect 9116 3236 9172 3238
rect 9196 3236 9252 3238
rect 9862 5616 9918 5672
rect 9770 3032 9826 3088
rect 9494 2624 9550 2680
rect 8956 2202 9012 2204
rect 9036 2202 9092 2204
rect 9116 2202 9172 2204
rect 9196 2202 9252 2204
rect 8956 2150 8982 2202
rect 8982 2150 9012 2202
rect 9036 2150 9046 2202
rect 9046 2150 9092 2202
rect 9116 2150 9162 2202
rect 9162 2150 9172 2202
rect 9196 2150 9226 2202
rect 9226 2150 9252 2202
rect 8956 2148 9012 2150
rect 9036 2148 9092 2150
rect 9116 2148 9172 2150
rect 9196 2148 9252 2150
rect 10138 7384 10194 7440
rect 10322 8200 10378 8256
rect 10230 3032 10286 3088
rect 10690 12824 10746 12880
rect 10506 9968 10562 10024
rect 10414 8064 10470 8120
rect 10966 12144 11022 12200
rect 11622 27770 11678 27772
rect 11702 27770 11758 27772
rect 11782 27770 11838 27772
rect 11862 27770 11918 27772
rect 11622 27718 11648 27770
rect 11648 27718 11678 27770
rect 11702 27718 11712 27770
rect 11712 27718 11758 27770
rect 11782 27718 11828 27770
rect 11828 27718 11838 27770
rect 11862 27718 11892 27770
rect 11892 27718 11918 27770
rect 11622 27716 11678 27718
rect 11702 27716 11758 27718
rect 11782 27716 11838 27718
rect 11862 27716 11918 27718
rect 11622 26682 11678 26684
rect 11702 26682 11758 26684
rect 11782 26682 11838 26684
rect 11862 26682 11918 26684
rect 11622 26630 11648 26682
rect 11648 26630 11678 26682
rect 11702 26630 11712 26682
rect 11712 26630 11758 26682
rect 11782 26630 11828 26682
rect 11828 26630 11838 26682
rect 11862 26630 11892 26682
rect 11892 26630 11918 26682
rect 11622 26628 11678 26630
rect 11702 26628 11758 26630
rect 11782 26628 11838 26630
rect 11862 26628 11918 26630
rect 11622 25594 11678 25596
rect 11702 25594 11758 25596
rect 11782 25594 11838 25596
rect 11862 25594 11918 25596
rect 11622 25542 11648 25594
rect 11648 25542 11678 25594
rect 11702 25542 11712 25594
rect 11712 25542 11758 25594
rect 11782 25542 11828 25594
rect 11828 25542 11838 25594
rect 11862 25542 11892 25594
rect 11892 25542 11918 25594
rect 11622 25540 11678 25542
rect 11702 25540 11758 25542
rect 11782 25540 11838 25542
rect 11862 25540 11918 25542
rect 11426 24792 11482 24848
rect 11978 24928 12034 24984
rect 11622 24506 11678 24508
rect 11702 24506 11758 24508
rect 11782 24506 11838 24508
rect 11862 24506 11918 24508
rect 11622 24454 11648 24506
rect 11648 24454 11678 24506
rect 11702 24454 11712 24506
rect 11712 24454 11758 24506
rect 11782 24454 11828 24506
rect 11828 24454 11838 24506
rect 11862 24454 11892 24506
rect 11892 24454 11918 24506
rect 11622 24452 11678 24454
rect 11702 24452 11758 24454
rect 11782 24452 11838 24454
rect 11862 24452 11918 24454
rect 11334 20984 11390 21040
rect 11334 16496 11390 16552
rect 11334 16088 11390 16144
rect 11242 11736 11298 11792
rect 11150 11464 11206 11520
rect 11622 23418 11678 23420
rect 11702 23418 11758 23420
rect 11782 23418 11838 23420
rect 11862 23418 11918 23420
rect 11622 23366 11648 23418
rect 11648 23366 11678 23418
rect 11702 23366 11712 23418
rect 11712 23366 11758 23418
rect 11782 23366 11828 23418
rect 11828 23366 11838 23418
rect 11862 23366 11892 23418
rect 11892 23366 11918 23418
rect 11622 23364 11678 23366
rect 11702 23364 11758 23366
rect 11782 23364 11838 23366
rect 11862 23364 11918 23366
rect 11622 22330 11678 22332
rect 11702 22330 11758 22332
rect 11782 22330 11838 22332
rect 11862 22330 11918 22332
rect 11622 22278 11648 22330
rect 11648 22278 11678 22330
rect 11702 22278 11712 22330
rect 11712 22278 11758 22330
rect 11782 22278 11828 22330
rect 11828 22278 11838 22330
rect 11862 22278 11892 22330
rect 11892 22278 11918 22330
rect 11622 22276 11678 22278
rect 11702 22276 11758 22278
rect 11782 22276 11838 22278
rect 11862 22276 11918 22278
rect 11622 21242 11678 21244
rect 11702 21242 11758 21244
rect 11782 21242 11838 21244
rect 11862 21242 11918 21244
rect 11622 21190 11648 21242
rect 11648 21190 11678 21242
rect 11702 21190 11712 21242
rect 11712 21190 11758 21242
rect 11782 21190 11828 21242
rect 11828 21190 11838 21242
rect 11862 21190 11892 21242
rect 11892 21190 11918 21242
rect 11622 21188 11678 21190
rect 11702 21188 11758 21190
rect 11782 21188 11838 21190
rect 11862 21188 11918 21190
rect 11622 20154 11678 20156
rect 11702 20154 11758 20156
rect 11782 20154 11838 20156
rect 11862 20154 11918 20156
rect 11622 20102 11648 20154
rect 11648 20102 11678 20154
rect 11702 20102 11712 20154
rect 11712 20102 11758 20154
rect 11782 20102 11828 20154
rect 11828 20102 11838 20154
rect 11862 20102 11892 20154
rect 11892 20102 11918 20154
rect 11622 20100 11678 20102
rect 11702 20100 11758 20102
rect 11782 20100 11838 20102
rect 11862 20100 11918 20102
rect 11794 19916 11850 19952
rect 12806 32952 12862 33008
rect 12714 31456 12770 31512
rect 12622 28056 12678 28112
rect 11794 19896 11796 19916
rect 11796 19896 11848 19916
rect 11848 19896 11850 19916
rect 12070 19760 12126 19816
rect 11622 19066 11678 19068
rect 11702 19066 11758 19068
rect 11782 19066 11838 19068
rect 11862 19066 11918 19068
rect 11622 19014 11648 19066
rect 11648 19014 11678 19066
rect 11702 19014 11712 19066
rect 11712 19014 11758 19066
rect 11782 19014 11828 19066
rect 11828 19014 11838 19066
rect 11862 19014 11892 19066
rect 11892 19014 11918 19066
rect 11622 19012 11678 19014
rect 11702 19012 11758 19014
rect 11782 19012 11838 19014
rect 11862 19012 11918 19014
rect 11978 18808 12034 18864
rect 11702 18708 11704 18728
rect 11704 18708 11756 18728
rect 11756 18708 11758 18728
rect 11702 18672 11758 18708
rect 11622 17978 11678 17980
rect 11702 17978 11758 17980
rect 11782 17978 11838 17980
rect 11862 17978 11918 17980
rect 11622 17926 11648 17978
rect 11648 17926 11678 17978
rect 11702 17926 11712 17978
rect 11712 17926 11758 17978
rect 11782 17926 11828 17978
rect 11828 17926 11838 17978
rect 11862 17926 11892 17978
rect 11892 17926 11918 17978
rect 11622 17924 11678 17926
rect 11702 17924 11758 17926
rect 11782 17924 11838 17926
rect 11862 17924 11918 17926
rect 11622 16890 11678 16892
rect 11702 16890 11758 16892
rect 11782 16890 11838 16892
rect 11862 16890 11918 16892
rect 11622 16838 11648 16890
rect 11648 16838 11678 16890
rect 11702 16838 11712 16890
rect 11712 16838 11758 16890
rect 11782 16838 11828 16890
rect 11828 16838 11838 16890
rect 11862 16838 11892 16890
rect 11892 16838 11918 16890
rect 11622 16836 11678 16838
rect 11702 16836 11758 16838
rect 11782 16836 11838 16838
rect 11862 16836 11918 16838
rect 11622 15802 11678 15804
rect 11702 15802 11758 15804
rect 11782 15802 11838 15804
rect 11862 15802 11918 15804
rect 11622 15750 11648 15802
rect 11648 15750 11678 15802
rect 11702 15750 11712 15802
rect 11712 15750 11758 15802
rect 11782 15750 11828 15802
rect 11828 15750 11838 15802
rect 11862 15750 11892 15802
rect 11892 15750 11918 15802
rect 11622 15748 11678 15750
rect 11702 15748 11758 15750
rect 11782 15748 11838 15750
rect 11862 15748 11918 15750
rect 11622 14714 11678 14716
rect 11702 14714 11758 14716
rect 11782 14714 11838 14716
rect 11862 14714 11918 14716
rect 11622 14662 11648 14714
rect 11648 14662 11678 14714
rect 11702 14662 11712 14714
rect 11712 14662 11758 14714
rect 11782 14662 11828 14714
rect 11828 14662 11838 14714
rect 11862 14662 11892 14714
rect 11892 14662 11918 14714
rect 11622 14660 11678 14662
rect 11702 14660 11758 14662
rect 11782 14660 11838 14662
rect 11862 14660 11918 14662
rect 11622 13626 11678 13628
rect 11702 13626 11758 13628
rect 11782 13626 11838 13628
rect 11862 13626 11918 13628
rect 11622 13574 11648 13626
rect 11648 13574 11678 13626
rect 11702 13574 11712 13626
rect 11712 13574 11758 13626
rect 11782 13574 11828 13626
rect 11828 13574 11838 13626
rect 11862 13574 11892 13626
rect 11892 13574 11918 13626
rect 11622 13572 11678 13574
rect 11702 13572 11758 13574
rect 11782 13572 11838 13574
rect 11862 13572 11918 13574
rect 11622 12538 11678 12540
rect 11702 12538 11758 12540
rect 11782 12538 11838 12540
rect 11862 12538 11918 12540
rect 11622 12486 11648 12538
rect 11648 12486 11678 12538
rect 11702 12486 11712 12538
rect 11712 12486 11758 12538
rect 11782 12486 11828 12538
rect 11828 12486 11838 12538
rect 11862 12486 11892 12538
rect 11892 12486 11918 12538
rect 11622 12484 11678 12486
rect 11702 12484 11758 12486
rect 11782 12484 11838 12486
rect 11862 12484 11918 12486
rect 11242 9968 11298 10024
rect 10598 5108 10600 5128
rect 10600 5108 10652 5128
rect 10652 5108 10654 5128
rect 10598 5072 10654 5108
rect 10506 3576 10562 3632
rect 10046 2896 10102 2952
rect 11150 5908 11206 5944
rect 11150 5888 11152 5908
rect 11152 5888 11204 5908
rect 11204 5888 11206 5908
rect 11058 5752 11114 5808
rect 11150 4936 11206 4992
rect 11150 2760 11206 2816
rect 11622 11450 11678 11452
rect 11702 11450 11758 11452
rect 11782 11450 11838 11452
rect 11862 11450 11918 11452
rect 11622 11398 11648 11450
rect 11648 11398 11678 11450
rect 11702 11398 11712 11450
rect 11712 11398 11758 11450
rect 11782 11398 11828 11450
rect 11828 11398 11838 11450
rect 11862 11398 11892 11450
rect 11892 11398 11918 11450
rect 11622 11396 11678 11398
rect 11702 11396 11758 11398
rect 11782 11396 11838 11398
rect 11862 11396 11918 11398
rect 11622 10362 11678 10364
rect 11702 10362 11758 10364
rect 11782 10362 11838 10364
rect 11862 10362 11918 10364
rect 11622 10310 11648 10362
rect 11648 10310 11678 10362
rect 11702 10310 11712 10362
rect 11712 10310 11758 10362
rect 11782 10310 11828 10362
rect 11828 10310 11838 10362
rect 11862 10310 11892 10362
rect 11892 10310 11918 10362
rect 11622 10308 11678 10310
rect 11702 10308 11758 10310
rect 11782 10308 11838 10310
rect 11862 10308 11918 10310
rect 11622 9274 11678 9276
rect 11702 9274 11758 9276
rect 11782 9274 11838 9276
rect 11862 9274 11918 9276
rect 11622 9222 11648 9274
rect 11648 9222 11678 9274
rect 11702 9222 11712 9274
rect 11712 9222 11758 9274
rect 11782 9222 11828 9274
rect 11828 9222 11838 9274
rect 11862 9222 11892 9274
rect 11892 9222 11918 9274
rect 11622 9220 11678 9222
rect 11702 9220 11758 9222
rect 11782 9220 11838 9222
rect 11862 9220 11918 9222
rect 12438 18128 12494 18184
rect 12438 16904 12494 16960
rect 11622 8186 11678 8188
rect 11702 8186 11758 8188
rect 11782 8186 11838 8188
rect 11862 8186 11918 8188
rect 11622 8134 11648 8186
rect 11648 8134 11678 8186
rect 11702 8134 11712 8186
rect 11712 8134 11758 8186
rect 11782 8134 11828 8186
rect 11828 8134 11838 8186
rect 11862 8134 11892 8186
rect 11892 8134 11918 8186
rect 11622 8132 11678 8134
rect 11702 8132 11758 8134
rect 11782 8132 11838 8134
rect 11862 8132 11918 8134
rect 11622 7098 11678 7100
rect 11702 7098 11758 7100
rect 11782 7098 11838 7100
rect 11862 7098 11918 7100
rect 11622 7046 11648 7098
rect 11648 7046 11678 7098
rect 11702 7046 11712 7098
rect 11712 7046 11758 7098
rect 11782 7046 11828 7098
rect 11828 7046 11838 7098
rect 11862 7046 11892 7098
rect 11892 7046 11918 7098
rect 11622 7044 11678 7046
rect 11702 7044 11758 7046
rect 11782 7044 11838 7046
rect 11862 7044 11918 7046
rect 11622 6010 11678 6012
rect 11702 6010 11758 6012
rect 11782 6010 11838 6012
rect 11862 6010 11918 6012
rect 11622 5958 11648 6010
rect 11648 5958 11678 6010
rect 11702 5958 11712 6010
rect 11712 5958 11758 6010
rect 11782 5958 11828 6010
rect 11828 5958 11838 6010
rect 11862 5958 11892 6010
rect 11892 5958 11918 6010
rect 11622 5956 11678 5958
rect 11702 5956 11758 5958
rect 11782 5956 11838 5958
rect 11862 5956 11918 5958
rect 11622 4922 11678 4924
rect 11702 4922 11758 4924
rect 11782 4922 11838 4924
rect 11862 4922 11918 4924
rect 11622 4870 11648 4922
rect 11648 4870 11678 4922
rect 11702 4870 11712 4922
rect 11712 4870 11758 4922
rect 11782 4870 11828 4922
rect 11828 4870 11838 4922
rect 11862 4870 11892 4922
rect 11892 4870 11918 4922
rect 11622 4868 11678 4870
rect 11702 4868 11758 4870
rect 11782 4868 11838 4870
rect 11862 4868 11918 4870
rect 11334 3848 11390 3904
rect 11242 2488 11298 2544
rect 11622 3834 11678 3836
rect 11702 3834 11758 3836
rect 11782 3834 11838 3836
rect 11862 3834 11918 3836
rect 11622 3782 11648 3834
rect 11648 3782 11678 3834
rect 11702 3782 11712 3834
rect 11712 3782 11758 3834
rect 11782 3782 11828 3834
rect 11828 3782 11838 3834
rect 11862 3782 11892 3834
rect 11892 3782 11918 3834
rect 11622 3780 11678 3782
rect 11702 3780 11758 3782
rect 11782 3780 11838 3782
rect 11862 3780 11918 3782
rect 11622 2746 11678 2748
rect 11702 2746 11758 2748
rect 11782 2746 11838 2748
rect 11862 2746 11918 2748
rect 11622 2694 11648 2746
rect 11648 2694 11678 2746
rect 11702 2694 11712 2746
rect 11712 2694 11758 2746
rect 11782 2694 11828 2746
rect 11828 2694 11838 2746
rect 11862 2694 11892 2746
rect 11892 2694 11918 2746
rect 11622 2692 11678 2694
rect 11702 2692 11758 2694
rect 11782 2692 11838 2694
rect 11862 2692 11918 2694
rect 12622 16632 12678 16688
rect 12346 10104 12402 10160
rect 12254 7928 12310 7984
rect 12162 6568 12218 6624
rect 12438 4548 12494 4584
rect 12438 4528 12440 4548
rect 12440 4528 12492 4548
rect 12492 4528 12494 4548
rect 12438 3576 12494 3632
rect 12898 30232 12954 30288
rect 12898 29688 12954 29744
rect 13082 28736 13138 28792
rect 12714 5208 12770 5264
rect 12990 23160 13046 23216
rect 13358 26968 13414 27024
rect 13726 29960 13782 30016
rect 14289 37018 14345 37020
rect 14369 37018 14425 37020
rect 14449 37018 14505 37020
rect 14529 37018 14585 37020
rect 14289 36966 14315 37018
rect 14315 36966 14345 37018
rect 14369 36966 14379 37018
rect 14379 36966 14425 37018
rect 14449 36966 14495 37018
rect 14495 36966 14505 37018
rect 14529 36966 14559 37018
rect 14559 36966 14585 37018
rect 14289 36964 14345 36966
rect 14369 36964 14425 36966
rect 14449 36964 14505 36966
rect 14529 36964 14585 36966
rect 14289 35930 14345 35932
rect 14369 35930 14425 35932
rect 14449 35930 14505 35932
rect 14529 35930 14585 35932
rect 14289 35878 14315 35930
rect 14315 35878 14345 35930
rect 14369 35878 14379 35930
rect 14379 35878 14425 35930
rect 14449 35878 14495 35930
rect 14495 35878 14505 35930
rect 14529 35878 14559 35930
rect 14559 35878 14585 35930
rect 14289 35876 14345 35878
rect 14369 35876 14425 35878
rect 14449 35876 14505 35878
rect 14529 35876 14585 35878
rect 14289 34842 14345 34844
rect 14369 34842 14425 34844
rect 14449 34842 14505 34844
rect 14529 34842 14585 34844
rect 14289 34790 14315 34842
rect 14315 34790 14345 34842
rect 14369 34790 14379 34842
rect 14379 34790 14425 34842
rect 14449 34790 14495 34842
rect 14495 34790 14505 34842
rect 14529 34790 14559 34842
rect 14559 34790 14585 34842
rect 14289 34788 14345 34790
rect 14369 34788 14425 34790
rect 14449 34788 14505 34790
rect 14529 34788 14585 34790
rect 14289 33754 14345 33756
rect 14369 33754 14425 33756
rect 14449 33754 14505 33756
rect 14529 33754 14585 33756
rect 14289 33702 14315 33754
rect 14315 33702 14345 33754
rect 14369 33702 14379 33754
rect 14379 33702 14425 33754
rect 14449 33702 14495 33754
rect 14495 33702 14505 33754
rect 14529 33702 14559 33754
rect 14559 33702 14585 33754
rect 14289 33700 14345 33702
rect 14369 33700 14425 33702
rect 14449 33700 14505 33702
rect 14529 33700 14585 33702
rect 15382 34040 15438 34096
rect 14922 32952 14978 33008
rect 14289 32666 14345 32668
rect 14369 32666 14425 32668
rect 14449 32666 14505 32668
rect 14529 32666 14585 32668
rect 14289 32614 14315 32666
rect 14315 32614 14345 32666
rect 14369 32614 14379 32666
rect 14379 32614 14425 32666
rect 14449 32614 14495 32666
rect 14495 32614 14505 32666
rect 14529 32614 14559 32666
rect 14559 32614 14585 32666
rect 14289 32612 14345 32614
rect 14369 32612 14425 32614
rect 14449 32612 14505 32614
rect 14529 32612 14585 32614
rect 14289 31578 14345 31580
rect 14369 31578 14425 31580
rect 14449 31578 14505 31580
rect 14529 31578 14585 31580
rect 14289 31526 14315 31578
rect 14315 31526 14345 31578
rect 14369 31526 14379 31578
rect 14379 31526 14425 31578
rect 14449 31526 14495 31578
rect 14495 31526 14505 31578
rect 14529 31526 14559 31578
rect 14559 31526 14585 31578
rect 14289 31524 14345 31526
rect 14369 31524 14425 31526
rect 14449 31524 14505 31526
rect 14529 31524 14585 31526
rect 14289 30490 14345 30492
rect 14369 30490 14425 30492
rect 14449 30490 14505 30492
rect 14529 30490 14585 30492
rect 14289 30438 14315 30490
rect 14315 30438 14345 30490
rect 14369 30438 14379 30490
rect 14379 30438 14425 30490
rect 14449 30438 14495 30490
rect 14495 30438 14505 30490
rect 14529 30438 14559 30490
rect 14559 30438 14585 30490
rect 14289 30436 14345 30438
rect 14369 30436 14425 30438
rect 14449 30436 14505 30438
rect 14529 30436 14585 30438
rect 14289 29402 14345 29404
rect 14369 29402 14425 29404
rect 14449 29402 14505 29404
rect 14529 29402 14585 29404
rect 14289 29350 14315 29402
rect 14315 29350 14345 29402
rect 14369 29350 14379 29402
rect 14379 29350 14425 29402
rect 14449 29350 14495 29402
rect 14495 29350 14505 29402
rect 14529 29350 14559 29402
rect 14559 29350 14585 29402
rect 14289 29348 14345 29350
rect 14369 29348 14425 29350
rect 14449 29348 14505 29350
rect 14529 29348 14585 29350
rect 15750 28736 15806 28792
rect 14289 28314 14345 28316
rect 14369 28314 14425 28316
rect 14449 28314 14505 28316
rect 14529 28314 14585 28316
rect 14289 28262 14315 28314
rect 14315 28262 14345 28314
rect 14369 28262 14379 28314
rect 14379 28262 14425 28314
rect 14449 28262 14495 28314
rect 14495 28262 14505 28314
rect 14529 28262 14559 28314
rect 14559 28262 14585 28314
rect 14289 28260 14345 28262
rect 14369 28260 14425 28262
rect 14449 28260 14505 28262
rect 14529 28260 14585 28262
rect 14289 27226 14345 27228
rect 14369 27226 14425 27228
rect 14449 27226 14505 27228
rect 14529 27226 14585 27228
rect 14289 27174 14315 27226
rect 14315 27174 14345 27226
rect 14369 27174 14379 27226
rect 14379 27174 14425 27226
rect 14449 27174 14495 27226
rect 14495 27174 14505 27226
rect 14529 27174 14559 27226
rect 14559 27174 14585 27226
rect 14289 27172 14345 27174
rect 14369 27172 14425 27174
rect 14449 27172 14505 27174
rect 14529 27172 14585 27174
rect 14289 26138 14345 26140
rect 14369 26138 14425 26140
rect 14449 26138 14505 26140
rect 14529 26138 14585 26140
rect 14289 26086 14315 26138
rect 14315 26086 14345 26138
rect 14369 26086 14379 26138
rect 14379 26086 14425 26138
rect 14449 26086 14495 26138
rect 14495 26086 14505 26138
rect 14529 26086 14559 26138
rect 14559 26086 14585 26138
rect 14289 26084 14345 26086
rect 14369 26084 14425 26086
rect 14449 26084 14505 26086
rect 14529 26084 14585 26086
rect 14289 25050 14345 25052
rect 14369 25050 14425 25052
rect 14449 25050 14505 25052
rect 14529 25050 14585 25052
rect 14289 24998 14315 25050
rect 14315 24998 14345 25050
rect 14369 24998 14379 25050
rect 14379 24998 14425 25050
rect 14449 24998 14495 25050
rect 14495 24998 14505 25050
rect 14529 24998 14559 25050
rect 14559 24998 14585 25050
rect 14289 24996 14345 24998
rect 14369 24996 14425 24998
rect 14449 24996 14505 24998
rect 14529 24996 14585 24998
rect 13634 24928 13690 24984
rect 13542 22616 13598 22672
rect 13082 19352 13138 19408
rect 13266 14864 13322 14920
rect 12898 7792 12954 7848
rect 13358 5072 13414 5128
rect 12622 3032 12678 3088
rect 12806 2916 12862 2952
rect 12806 2896 12808 2916
rect 12808 2896 12860 2916
rect 12860 2896 12862 2916
rect 12806 2372 12862 2408
rect 12806 2352 12808 2372
rect 12808 2352 12860 2372
rect 12860 2352 12862 2372
rect 14289 23962 14345 23964
rect 14369 23962 14425 23964
rect 14449 23962 14505 23964
rect 14529 23962 14585 23964
rect 14289 23910 14315 23962
rect 14315 23910 14345 23962
rect 14369 23910 14379 23962
rect 14379 23910 14425 23962
rect 14449 23910 14495 23962
rect 14495 23910 14505 23962
rect 14529 23910 14559 23962
rect 14559 23910 14585 23962
rect 14289 23908 14345 23910
rect 14369 23908 14425 23910
rect 14449 23908 14505 23910
rect 14529 23908 14585 23910
rect 14289 22874 14345 22876
rect 14369 22874 14425 22876
rect 14449 22874 14505 22876
rect 14529 22874 14585 22876
rect 14289 22822 14315 22874
rect 14315 22822 14345 22874
rect 14369 22822 14379 22874
rect 14379 22822 14425 22874
rect 14449 22822 14495 22874
rect 14495 22822 14505 22874
rect 14529 22822 14559 22874
rect 14559 22822 14585 22874
rect 14289 22820 14345 22822
rect 14369 22820 14425 22822
rect 14449 22820 14505 22822
rect 14529 22820 14585 22822
rect 14289 21786 14345 21788
rect 14369 21786 14425 21788
rect 14449 21786 14505 21788
rect 14529 21786 14585 21788
rect 14289 21734 14315 21786
rect 14315 21734 14345 21786
rect 14369 21734 14379 21786
rect 14379 21734 14425 21786
rect 14449 21734 14495 21786
rect 14495 21734 14505 21786
rect 14529 21734 14559 21786
rect 14559 21734 14585 21786
rect 14289 21732 14345 21734
rect 14369 21732 14425 21734
rect 14449 21732 14505 21734
rect 14529 21732 14585 21734
rect 14289 20698 14345 20700
rect 14369 20698 14425 20700
rect 14449 20698 14505 20700
rect 14529 20698 14585 20700
rect 14289 20646 14315 20698
rect 14315 20646 14345 20698
rect 14369 20646 14379 20698
rect 14379 20646 14425 20698
rect 14449 20646 14495 20698
rect 14495 20646 14505 20698
rect 14529 20646 14559 20698
rect 14559 20646 14585 20698
rect 14289 20644 14345 20646
rect 14369 20644 14425 20646
rect 14449 20644 14505 20646
rect 14529 20644 14585 20646
rect 14289 19610 14345 19612
rect 14369 19610 14425 19612
rect 14449 19610 14505 19612
rect 14529 19610 14585 19612
rect 14289 19558 14315 19610
rect 14315 19558 14345 19610
rect 14369 19558 14379 19610
rect 14379 19558 14425 19610
rect 14449 19558 14495 19610
rect 14495 19558 14505 19610
rect 14529 19558 14559 19610
rect 14559 19558 14585 19610
rect 14289 19556 14345 19558
rect 14369 19556 14425 19558
rect 14449 19556 14505 19558
rect 14529 19556 14585 19558
rect 14289 18522 14345 18524
rect 14369 18522 14425 18524
rect 14449 18522 14505 18524
rect 14529 18522 14585 18524
rect 14289 18470 14315 18522
rect 14315 18470 14345 18522
rect 14369 18470 14379 18522
rect 14379 18470 14425 18522
rect 14449 18470 14495 18522
rect 14495 18470 14505 18522
rect 14529 18470 14559 18522
rect 14559 18470 14585 18522
rect 14289 18468 14345 18470
rect 14369 18468 14425 18470
rect 14449 18468 14505 18470
rect 14529 18468 14585 18470
rect 14289 17434 14345 17436
rect 14369 17434 14425 17436
rect 14449 17434 14505 17436
rect 14529 17434 14585 17436
rect 14289 17382 14315 17434
rect 14315 17382 14345 17434
rect 14369 17382 14379 17434
rect 14379 17382 14425 17434
rect 14449 17382 14495 17434
rect 14495 17382 14505 17434
rect 14529 17382 14559 17434
rect 14559 17382 14585 17434
rect 14289 17380 14345 17382
rect 14369 17380 14425 17382
rect 14449 17380 14505 17382
rect 14529 17380 14585 17382
rect 14289 16346 14345 16348
rect 14369 16346 14425 16348
rect 14449 16346 14505 16348
rect 14529 16346 14585 16348
rect 14289 16294 14315 16346
rect 14315 16294 14345 16346
rect 14369 16294 14379 16346
rect 14379 16294 14425 16346
rect 14449 16294 14495 16346
rect 14495 16294 14505 16346
rect 14529 16294 14559 16346
rect 14559 16294 14585 16346
rect 14289 16292 14345 16294
rect 14369 16292 14425 16294
rect 14449 16292 14505 16294
rect 14529 16292 14585 16294
rect 14289 15258 14345 15260
rect 14369 15258 14425 15260
rect 14449 15258 14505 15260
rect 14529 15258 14585 15260
rect 14289 15206 14315 15258
rect 14315 15206 14345 15258
rect 14369 15206 14379 15258
rect 14379 15206 14425 15258
rect 14449 15206 14495 15258
rect 14495 15206 14505 15258
rect 14529 15206 14559 15258
rect 14559 15206 14585 15258
rect 14289 15204 14345 15206
rect 14369 15204 14425 15206
rect 14449 15204 14505 15206
rect 14529 15204 14585 15206
rect 14289 14170 14345 14172
rect 14369 14170 14425 14172
rect 14449 14170 14505 14172
rect 14529 14170 14585 14172
rect 14289 14118 14315 14170
rect 14315 14118 14345 14170
rect 14369 14118 14379 14170
rect 14379 14118 14425 14170
rect 14449 14118 14495 14170
rect 14495 14118 14505 14170
rect 14529 14118 14559 14170
rect 14559 14118 14585 14170
rect 14289 14116 14345 14118
rect 14369 14116 14425 14118
rect 14449 14116 14505 14118
rect 14529 14116 14585 14118
rect 14289 13082 14345 13084
rect 14369 13082 14425 13084
rect 14449 13082 14505 13084
rect 14529 13082 14585 13084
rect 14289 13030 14315 13082
rect 14315 13030 14345 13082
rect 14369 13030 14379 13082
rect 14379 13030 14425 13082
rect 14449 13030 14495 13082
rect 14495 13030 14505 13082
rect 14529 13030 14559 13082
rect 14559 13030 14585 13082
rect 14289 13028 14345 13030
rect 14369 13028 14425 13030
rect 14449 13028 14505 13030
rect 14529 13028 14585 13030
rect 14289 11994 14345 11996
rect 14369 11994 14425 11996
rect 14449 11994 14505 11996
rect 14529 11994 14585 11996
rect 14289 11942 14315 11994
rect 14315 11942 14345 11994
rect 14369 11942 14379 11994
rect 14379 11942 14425 11994
rect 14449 11942 14495 11994
rect 14495 11942 14505 11994
rect 14529 11942 14559 11994
rect 14559 11942 14585 11994
rect 14289 11940 14345 11942
rect 14369 11940 14425 11942
rect 14449 11940 14505 11942
rect 14529 11940 14585 11942
rect 14289 10906 14345 10908
rect 14369 10906 14425 10908
rect 14449 10906 14505 10908
rect 14529 10906 14585 10908
rect 14289 10854 14315 10906
rect 14315 10854 14345 10906
rect 14369 10854 14379 10906
rect 14379 10854 14425 10906
rect 14449 10854 14495 10906
rect 14495 10854 14505 10906
rect 14529 10854 14559 10906
rect 14559 10854 14585 10906
rect 14289 10852 14345 10854
rect 14369 10852 14425 10854
rect 14449 10852 14505 10854
rect 14529 10852 14585 10854
rect 14830 10104 14886 10160
rect 14289 9818 14345 9820
rect 14369 9818 14425 9820
rect 14449 9818 14505 9820
rect 14529 9818 14585 9820
rect 14289 9766 14315 9818
rect 14315 9766 14345 9818
rect 14369 9766 14379 9818
rect 14379 9766 14425 9818
rect 14449 9766 14495 9818
rect 14495 9766 14505 9818
rect 14529 9766 14559 9818
rect 14559 9766 14585 9818
rect 14289 9764 14345 9766
rect 14369 9764 14425 9766
rect 14449 9764 14505 9766
rect 14529 9764 14585 9766
rect 14289 8730 14345 8732
rect 14369 8730 14425 8732
rect 14449 8730 14505 8732
rect 14529 8730 14585 8732
rect 14289 8678 14315 8730
rect 14315 8678 14345 8730
rect 14369 8678 14379 8730
rect 14379 8678 14425 8730
rect 14449 8678 14495 8730
rect 14495 8678 14505 8730
rect 14529 8678 14559 8730
rect 14559 8678 14585 8730
rect 14289 8676 14345 8678
rect 14369 8676 14425 8678
rect 14449 8676 14505 8678
rect 14529 8676 14585 8678
rect 14289 7642 14345 7644
rect 14369 7642 14425 7644
rect 14449 7642 14505 7644
rect 14529 7642 14585 7644
rect 14289 7590 14315 7642
rect 14315 7590 14345 7642
rect 14369 7590 14379 7642
rect 14379 7590 14425 7642
rect 14449 7590 14495 7642
rect 14495 7590 14505 7642
rect 14529 7590 14559 7642
rect 14559 7590 14585 7642
rect 14289 7588 14345 7590
rect 14369 7588 14425 7590
rect 14449 7588 14505 7590
rect 14529 7588 14585 7590
rect 14289 6554 14345 6556
rect 14369 6554 14425 6556
rect 14449 6554 14505 6556
rect 14529 6554 14585 6556
rect 14289 6502 14315 6554
rect 14315 6502 14345 6554
rect 14369 6502 14379 6554
rect 14379 6502 14425 6554
rect 14449 6502 14495 6554
rect 14495 6502 14505 6554
rect 14529 6502 14559 6554
rect 14559 6502 14585 6554
rect 14289 6500 14345 6502
rect 14369 6500 14425 6502
rect 14449 6500 14505 6502
rect 14529 6500 14585 6502
rect 14289 5466 14345 5468
rect 14369 5466 14425 5468
rect 14449 5466 14505 5468
rect 14529 5466 14585 5468
rect 14289 5414 14315 5466
rect 14315 5414 14345 5466
rect 14369 5414 14379 5466
rect 14379 5414 14425 5466
rect 14449 5414 14495 5466
rect 14495 5414 14505 5466
rect 14529 5414 14559 5466
rect 14559 5414 14585 5466
rect 14289 5412 14345 5414
rect 14369 5412 14425 5414
rect 14449 5412 14505 5414
rect 14529 5412 14585 5414
rect 14646 4664 14702 4720
rect 14289 4378 14345 4380
rect 14369 4378 14425 4380
rect 14449 4378 14505 4380
rect 14529 4378 14585 4380
rect 14289 4326 14315 4378
rect 14315 4326 14345 4378
rect 14369 4326 14379 4378
rect 14379 4326 14425 4378
rect 14449 4326 14495 4378
rect 14495 4326 14505 4378
rect 14529 4326 14559 4378
rect 14559 4326 14585 4378
rect 14289 4324 14345 4326
rect 14369 4324 14425 4326
rect 14449 4324 14505 4326
rect 14529 4324 14585 4326
rect 13726 3984 13782 4040
rect 13450 3460 13506 3496
rect 13450 3440 13452 3460
rect 13452 3440 13504 3460
rect 13504 3440 13506 3460
rect 13634 3440 13690 3496
rect 14186 3440 14242 3496
rect 14289 3290 14345 3292
rect 14369 3290 14425 3292
rect 14449 3290 14505 3292
rect 14529 3290 14585 3292
rect 14289 3238 14315 3290
rect 14315 3238 14345 3290
rect 14369 3238 14379 3290
rect 14379 3238 14425 3290
rect 14449 3238 14495 3290
rect 14495 3238 14505 3290
rect 14529 3238 14559 3290
rect 14559 3238 14585 3290
rect 14289 3236 14345 3238
rect 14369 3236 14425 3238
rect 14449 3236 14505 3238
rect 14529 3236 14585 3238
rect 14289 2202 14345 2204
rect 14369 2202 14425 2204
rect 14449 2202 14505 2204
rect 14529 2202 14585 2204
rect 14289 2150 14315 2202
rect 14315 2150 14345 2202
rect 14369 2150 14379 2202
rect 14379 2150 14425 2202
rect 14449 2150 14495 2202
rect 14495 2150 14505 2202
rect 14529 2150 14559 2202
rect 14559 2150 14585 2202
rect 14289 2148 14345 2150
rect 14369 2148 14425 2150
rect 14449 2148 14505 2150
rect 14529 2148 14585 2150
rect 15382 7248 15438 7304
<< metal3 >>
rect 0 38722 480 38752
rect 1577 38722 1643 38725
rect 0 38720 1643 38722
rect 0 38664 1582 38720
rect 1638 38664 1643 38720
rect 0 38662 1643 38664
rect 0 38632 480 38662
rect 1577 38659 1643 38662
rect 6277 37568 6597 37569
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 37503 6597 37504
rect 11610 37568 11930 37569
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 37503 11930 37504
rect 3610 37024 3930 37025
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3930 37024
rect 3610 36959 3930 36960
rect 8944 37024 9264 37025
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 36959 9264 36960
rect 14277 37024 14597 37025
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 36959 14597 36960
rect 6277 36480 6597 36481
rect 0 36410 480 36440
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 36415 6597 36416
rect 11610 36480 11930 36481
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 36415 11930 36416
rect 1485 36410 1551 36413
rect 0 36408 1551 36410
rect 0 36352 1490 36408
rect 1546 36352 1551 36408
rect 0 36350 1551 36352
rect 0 36320 480 36350
rect 1485 36347 1551 36350
rect 3610 35936 3930 35937
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3930 35936
rect 3610 35871 3930 35872
rect 8944 35936 9264 35937
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 35871 9264 35872
rect 14277 35936 14597 35937
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 35871 14597 35872
rect 2957 35730 3023 35733
rect 9857 35730 9923 35733
rect 2957 35728 9923 35730
rect 2957 35672 2962 35728
rect 3018 35672 9862 35728
rect 9918 35672 9923 35728
rect 2957 35670 9923 35672
rect 2957 35667 3023 35670
rect 9857 35667 9923 35670
rect 6277 35392 6597 35393
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 35327 6597 35328
rect 11610 35392 11930 35393
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 35327 11930 35328
rect 2589 35322 2655 35325
rect 4245 35322 4311 35325
rect 2589 35320 4311 35322
rect 2589 35264 2594 35320
rect 2650 35264 4250 35320
rect 4306 35264 4311 35320
rect 2589 35262 4311 35264
rect 2589 35259 2655 35262
rect 4245 35259 4311 35262
rect 8845 35186 8911 35189
rect 11462 35186 11468 35188
rect 8845 35184 11468 35186
rect 8845 35128 8850 35184
rect 8906 35128 11468 35184
rect 8845 35126 11468 35128
rect 8845 35123 8911 35126
rect 11462 35124 11468 35126
rect 11532 35124 11538 35188
rect 2129 35050 2195 35053
rect 4337 35050 4403 35053
rect 2129 35048 4403 35050
rect 2129 34992 2134 35048
rect 2190 34992 4342 35048
rect 4398 34992 4403 35048
rect 2129 34990 4403 34992
rect 2129 34987 2195 34990
rect 4337 34987 4403 34990
rect 8477 35050 8543 35053
rect 12985 35050 13051 35053
rect 8477 35048 13051 35050
rect 8477 34992 8482 35048
rect 8538 34992 12990 35048
rect 13046 34992 13051 35048
rect 8477 34990 13051 34992
rect 8477 34987 8543 34990
rect 12985 34987 13051 34990
rect 3610 34848 3930 34849
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3930 34848
rect 3610 34783 3930 34784
rect 8944 34848 9264 34849
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 34783 9264 34784
rect 14277 34848 14597 34849
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 34783 14597 34784
rect 197 34778 263 34781
rect 3233 34778 3299 34781
rect 197 34776 3299 34778
rect 197 34720 202 34776
rect 258 34720 3238 34776
rect 3294 34720 3299 34776
rect 197 34718 3299 34720
rect 197 34715 263 34718
rect 3233 34715 3299 34718
rect 3693 34642 3759 34645
rect 5809 34642 5875 34645
rect 9765 34642 9831 34645
rect 3693 34640 9831 34642
rect 3693 34584 3698 34640
rect 3754 34584 5814 34640
rect 5870 34584 9770 34640
rect 9826 34584 9831 34640
rect 3693 34582 9831 34584
rect 3693 34579 3759 34582
rect 5809 34579 5875 34582
rect 9765 34579 9831 34582
rect 5901 34506 5967 34509
rect 8569 34506 8635 34509
rect 10501 34506 10567 34509
rect 5901 34504 10567 34506
rect 5901 34448 5906 34504
rect 5962 34448 8574 34504
rect 8630 34448 10506 34504
rect 10562 34448 10567 34504
rect 5901 34446 10567 34448
rect 5901 34443 5967 34446
rect 8569 34443 8635 34446
rect 10501 34443 10567 34446
rect 6277 34304 6597 34305
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 34239 6597 34240
rect 11610 34304 11930 34305
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 34239 11930 34240
rect 1945 34234 2011 34237
rect 5993 34234 6059 34237
rect 1945 34232 6059 34234
rect 1945 34176 1950 34232
rect 2006 34176 5998 34232
rect 6054 34176 6059 34232
rect 1945 34174 6059 34176
rect 1945 34171 2011 34174
rect 5993 34171 6059 34174
rect 0 34098 480 34128
rect 1669 34098 1735 34101
rect 0 34096 1735 34098
rect 0 34040 1674 34096
rect 1730 34040 1735 34096
rect 0 34038 1735 34040
rect 0 34008 480 34038
rect 1669 34035 1735 34038
rect 2497 34098 2563 34101
rect 4889 34098 4955 34101
rect 2497 34096 4955 34098
rect 2497 34040 2502 34096
rect 2558 34040 4894 34096
rect 4950 34040 4955 34096
rect 2497 34038 4955 34040
rect 2497 34035 2563 34038
rect 4889 34035 4955 34038
rect 5165 34098 5231 34101
rect 7005 34098 7071 34101
rect 5165 34096 7071 34098
rect 5165 34040 5170 34096
rect 5226 34040 7010 34096
rect 7066 34040 7071 34096
rect 5165 34038 7071 34040
rect 5165 34035 5231 34038
rect 7005 34035 7071 34038
rect 7189 34098 7255 34101
rect 10317 34098 10383 34101
rect 7189 34096 10383 34098
rect 7189 34040 7194 34096
rect 7250 34040 10322 34096
rect 10378 34040 10383 34096
rect 7189 34038 10383 34040
rect 7189 34035 7255 34038
rect 10317 34035 10383 34038
rect 12249 34098 12315 34101
rect 15377 34098 15443 34101
rect 12249 34096 15443 34098
rect 12249 34040 12254 34096
rect 12310 34040 15382 34096
rect 15438 34040 15443 34096
rect 12249 34038 15443 34040
rect 12249 34035 12315 34038
rect 15377 34035 15443 34038
rect 2037 33962 2103 33965
rect 12433 33962 12499 33965
rect 2037 33960 12499 33962
rect 2037 33904 2042 33960
rect 2098 33904 12438 33960
rect 12494 33904 12499 33960
rect 2037 33902 12499 33904
rect 2037 33899 2103 33902
rect 12433 33899 12499 33902
rect 4889 33826 4955 33829
rect 6545 33826 6611 33829
rect 4889 33824 6611 33826
rect 4889 33768 4894 33824
rect 4950 33768 6550 33824
rect 6606 33768 6611 33824
rect 4889 33766 6611 33768
rect 4889 33763 4955 33766
rect 6545 33763 6611 33766
rect 3610 33760 3930 33761
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3930 33760
rect 3610 33695 3930 33696
rect 8944 33760 9264 33761
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 33695 9264 33696
rect 14277 33760 14597 33761
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 33695 14597 33696
rect 2405 33554 2471 33557
rect 9305 33554 9371 33557
rect 2405 33552 9371 33554
rect 2405 33496 2410 33552
rect 2466 33496 9310 33552
rect 9366 33496 9371 33552
rect 2405 33494 9371 33496
rect 2405 33491 2471 33494
rect 9305 33491 9371 33494
rect 5993 33418 6059 33421
rect 8753 33418 8819 33421
rect 5993 33416 8819 33418
rect 5993 33360 5998 33416
rect 6054 33360 8758 33416
rect 8814 33360 8819 33416
rect 5993 33358 8819 33360
rect 5993 33355 6059 33358
rect 8753 33355 8819 33358
rect 7373 33282 7439 33285
rect 11237 33282 11303 33285
rect 7373 33280 11303 33282
rect 7373 33224 7378 33280
rect 7434 33224 11242 33280
rect 11298 33224 11303 33280
rect 7373 33222 11303 33224
rect 7373 33219 7439 33222
rect 11237 33219 11303 33222
rect 6277 33216 6597 33217
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 33151 6597 33152
rect 11610 33216 11930 33217
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 33151 11930 33152
rect 10501 33146 10567 33149
rect 10685 33146 10751 33149
rect 10501 33144 10751 33146
rect 10501 33088 10506 33144
rect 10562 33088 10690 33144
rect 10746 33088 10751 33144
rect 10501 33086 10751 33088
rect 10501 33083 10567 33086
rect 10685 33083 10751 33086
rect 1393 33010 1459 33013
rect 5717 33010 5783 33013
rect 1393 33008 5783 33010
rect 1393 32952 1398 33008
rect 1454 32952 5722 33008
rect 5778 32952 5783 33008
rect 1393 32950 5783 32952
rect 1393 32947 1459 32950
rect 5717 32947 5783 32950
rect 8201 33010 8267 33013
rect 12801 33010 12867 33013
rect 14917 33010 14983 33013
rect 8201 33008 14983 33010
rect 8201 32952 8206 33008
rect 8262 32952 12806 33008
rect 12862 32952 14922 33008
rect 14978 32952 14983 33008
rect 8201 32950 14983 32952
rect 8201 32947 8267 32950
rect 12801 32947 12867 32950
rect 14917 32947 14983 32950
rect 5901 32874 5967 32877
rect 8661 32874 8727 32877
rect 9673 32874 9739 32877
rect 5901 32872 9739 32874
rect 5901 32816 5906 32872
rect 5962 32816 8666 32872
rect 8722 32816 9678 32872
rect 9734 32816 9739 32872
rect 5901 32814 9739 32816
rect 5901 32811 5967 32814
rect 8661 32811 8727 32814
rect 9673 32811 9739 32814
rect 9489 32738 9555 32741
rect 10685 32738 10751 32741
rect 9446 32736 10751 32738
rect 9446 32680 9494 32736
rect 9550 32680 10690 32736
rect 10746 32680 10751 32736
rect 9446 32678 10751 32680
rect 9446 32675 9555 32678
rect 10685 32675 10751 32678
rect 3610 32672 3930 32673
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3930 32672
rect 3610 32607 3930 32608
rect 8944 32672 9264 32673
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 32607 9264 32608
rect 7741 32466 7807 32469
rect 9446 32466 9506 32675
rect 14277 32672 14597 32673
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 32607 14597 32608
rect 7741 32464 9506 32466
rect 7741 32408 7746 32464
rect 7802 32408 9506 32464
rect 7741 32406 9506 32408
rect 7741 32403 7807 32406
rect 4153 32330 4219 32333
rect 7557 32330 7623 32333
rect 9673 32330 9739 32333
rect 4153 32328 9739 32330
rect 4153 32272 4158 32328
rect 4214 32272 7562 32328
rect 7618 32272 9678 32328
rect 9734 32272 9739 32328
rect 4153 32270 9739 32272
rect 4153 32267 4219 32270
rect 7557 32267 7623 32270
rect 9673 32267 9739 32270
rect 6277 32128 6597 32129
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 32063 6597 32064
rect 11610 32128 11930 32129
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 32063 11930 32064
rect 10225 32058 10291 32061
rect 10225 32056 10426 32058
rect 10225 32000 10230 32056
rect 10286 32000 10426 32056
rect 10225 31998 10426 32000
rect 10225 31995 10291 31998
rect 10366 31922 10426 31998
rect 10501 31922 10567 31925
rect 10366 31920 10567 31922
rect 10366 31864 10506 31920
rect 10562 31864 10567 31920
rect 10366 31862 10567 31864
rect 10501 31859 10567 31862
rect 0 31650 480 31680
rect 1669 31650 1735 31653
rect 0 31648 1735 31650
rect 0 31592 1674 31648
rect 1730 31592 1735 31648
rect 0 31590 1735 31592
rect 0 31560 480 31590
rect 1669 31587 1735 31590
rect 3610 31584 3930 31585
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3930 31584
rect 3610 31519 3930 31520
rect 8944 31584 9264 31585
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 31519 9264 31520
rect 14277 31584 14597 31585
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 31519 14597 31520
rect 9622 31452 9628 31516
rect 9692 31514 9698 31516
rect 12709 31514 12775 31517
rect 9692 31512 12775 31514
rect 9692 31456 12714 31512
rect 12770 31456 12775 31512
rect 9692 31454 12775 31456
rect 9692 31452 9698 31454
rect 12709 31451 12775 31454
rect 9305 31378 9371 31381
rect 9857 31378 9923 31381
rect 9305 31376 9923 31378
rect 9305 31320 9310 31376
rect 9366 31320 9862 31376
rect 9918 31320 9923 31376
rect 9305 31318 9923 31320
rect 9305 31315 9371 31318
rect 9857 31315 9923 31318
rect 5257 31242 5323 31245
rect 9622 31242 9628 31244
rect 5257 31240 9628 31242
rect 5257 31184 5262 31240
rect 5318 31184 9628 31240
rect 5257 31182 9628 31184
rect 5257 31179 5323 31182
rect 9622 31180 9628 31182
rect 9692 31180 9698 31244
rect 9581 31106 9647 31109
rect 11145 31106 11211 31109
rect 9581 31104 11211 31106
rect 9581 31048 9586 31104
rect 9642 31048 11150 31104
rect 11206 31048 11211 31104
rect 9581 31046 11211 31048
rect 9581 31043 9647 31046
rect 11145 31043 11211 31046
rect 6277 31040 6597 31041
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 30975 6597 30976
rect 11610 31040 11930 31041
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 30975 11930 30976
rect 10225 30970 10291 30973
rect 10182 30968 10291 30970
rect 10182 30912 10230 30968
rect 10286 30912 10291 30968
rect 10182 30907 10291 30912
rect 1945 30834 2011 30837
rect 5257 30834 5323 30837
rect 5533 30834 5599 30837
rect 8477 30834 8543 30837
rect 1945 30832 5458 30834
rect 1945 30776 1950 30832
rect 2006 30776 5262 30832
rect 5318 30776 5458 30832
rect 1945 30774 5458 30776
rect 1945 30771 2011 30774
rect 5257 30771 5323 30774
rect 5398 30698 5458 30774
rect 5533 30832 8543 30834
rect 5533 30776 5538 30832
rect 5594 30776 8482 30832
rect 8538 30776 8543 30832
rect 5533 30774 8543 30776
rect 5533 30771 5599 30774
rect 8477 30771 8543 30774
rect 10182 30698 10242 30907
rect 5398 30638 10242 30698
rect 4061 30562 4127 30565
rect 5993 30562 6059 30565
rect 4061 30560 6059 30562
rect 4061 30504 4066 30560
rect 4122 30504 5998 30560
rect 6054 30504 6059 30560
rect 4061 30502 6059 30504
rect 4061 30499 4127 30502
rect 5993 30499 6059 30502
rect 3610 30496 3930 30497
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3930 30496
rect 3610 30431 3930 30432
rect 8944 30496 9264 30497
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 30431 9264 30432
rect 14277 30496 14597 30497
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 30431 14597 30432
rect 4797 30426 4863 30429
rect 7189 30426 7255 30429
rect 4797 30424 7255 30426
rect 4797 30368 4802 30424
rect 4858 30368 7194 30424
rect 7250 30368 7255 30424
rect 4797 30366 7255 30368
rect 4797 30363 4863 30366
rect 7189 30363 7255 30366
rect 11145 30426 11211 30429
rect 12249 30426 12315 30429
rect 11145 30424 12315 30426
rect 11145 30368 11150 30424
rect 11206 30368 12254 30424
rect 12310 30368 12315 30424
rect 11145 30366 12315 30368
rect 11145 30363 11211 30366
rect 12249 30363 12315 30366
rect 2405 30290 2471 30293
rect 4705 30290 4771 30293
rect 2405 30288 4771 30290
rect 2405 30232 2410 30288
rect 2466 30232 4710 30288
rect 4766 30232 4771 30288
rect 2405 30230 4771 30232
rect 2405 30227 2471 30230
rect 4705 30227 4771 30230
rect 6637 30290 6703 30293
rect 10225 30290 10291 30293
rect 6637 30288 10291 30290
rect 6637 30232 6642 30288
rect 6698 30232 10230 30288
rect 10286 30232 10291 30288
rect 6637 30230 10291 30232
rect 6637 30227 6703 30230
rect 10225 30227 10291 30230
rect 10777 30290 10843 30293
rect 12893 30290 12959 30293
rect 10777 30288 12959 30290
rect 10777 30232 10782 30288
rect 10838 30232 12898 30288
rect 12954 30232 12959 30288
rect 10777 30230 12959 30232
rect 10777 30227 10843 30230
rect 12893 30227 12959 30230
rect 2129 30154 2195 30157
rect 6821 30154 6887 30157
rect 2129 30152 6887 30154
rect 2129 30096 2134 30152
rect 2190 30096 6826 30152
rect 6882 30096 6887 30152
rect 2129 30094 6887 30096
rect 2129 30091 2195 30094
rect 6821 30091 6887 30094
rect 2221 30018 2287 30021
rect 4153 30018 4219 30021
rect 2221 30016 4219 30018
rect 2221 29960 2226 30016
rect 2282 29960 4158 30016
rect 4214 29960 4219 30016
rect 2221 29958 4219 29960
rect 2221 29955 2287 29958
rect 4153 29955 4219 29958
rect 13721 30018 13787 30021
rect 15520 30018 16000 30048
rect 13721 30016 16000 30018
rect 13721 29960 13726 30016
rect 13782 29960 16000 30016
rect 13721 29958 16000 29960
rect 13721 29955 13787 29958
rect 6277 29952 6597 29953
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 29887 6597 29888
rect 11610 29952 11930 29953
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 15520 29928 16000 29958
rect 11610 29887 11930 29888
rect 10777 29746 10843 29749
rect 12893 29746 12959 29749
rect 10777 29744 12959 29746
rect 10777 29688 10782 29744
rect 10838 29688 12898 29744
rect 12954 29688 12959 29744
rect 10777 29686 12959 29688
rect 10777 29683 10843 29686
rect 12893 29683 12959 29686
rect 11462 29548 11468 29612
rect 11532 29610 11538 29612
rect 11881 29610 11947 29613
rect 11532 29608 11947 29610
rect 11532 29552 11886 29608
rect 11942 29552 11947 29608
rect 11532 29550 11947 29552
rect 11532 29548 11538 29550
rect 11881 29547 11947 29550
rect 3610 29408 3930 29409
rect 0 29338 480 29368
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3930 29408
rect 3610 29343 3930 29344
rect 8944 29408 9264 29409
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 29343 9264 29344
rect 14277 29408 14597 29409
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 29343 14597 29344
rect 0 29278 1594 29338
rect 0 29248 480 29278
rect 1534 28933 1594 29278
rect 3693 29066 3759 29069
rect 5901 29066 5967 29069
rect 3693 29064 5967 29066
rect 3693 29008 3698 29064
rect 3754 29008 5906 29064
rect 5962 29008 5967 29064
rect 3693 29006 5967 29008
rect 3693 29003 3759 29006
rect 5901 29003 5967 29006
rect 11053 29066 11119 29069
rect 11237 29066 11303 29069
rect 11053 29064 11303 29066
rect 11053 29008 11058 29064
rect 11114 29008 11242 29064
rect 11298 29008 11303 29064
rect 11053 29006 11303 29008
rect 11053 29003 11119 29006
rect 11237 29003 11303 29006
rect 1534 28928 1643 28933
rect 1534 28872 1582 28928
rect 1638 28872 1643 28928
rect 1534 28870 1643 28872
rect 1577 28867 1643 28870
rect 6277 28864 6597 28865
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 28799 6597 28800
rect 11610 28864 11930 28865
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 28799 11930 28800
rect 7741 28794 7807 28797
rect 6686 28792 7807 28794
rect 6686 28736 7746 28792
rect 7802 28736 7807 28792
rect 6686 28734 7807 28736
rect 5533 28658 5599 28661
rect 6686 28658 6746 28734
rect 7741 28731 7807 28734
rect 12065 28794 12131 28797
rect 13077 28794 13143 28797
rect 15745 28794 15811 28797
rect 12065 28792 15811 28794
rect 12065 28736 12070 28792
rect 12126 28736 13082 28792
rect 13138 28736 15750 28792
rect 15806 28736 15811 28792
rect 12065 28734 15811 28736
rect 12065 28731 12131 28734
rect 13077 28731 13143 28734
rect 15745 28731 15811 28734
rect 5533 28656 6746 28658
rect 5533 28600 5538 28656
rect 5594 28600 6746 28656
rect 5533 28598 6746 28600
rect 9581 28658 9647 28661
rect 11513 28658 11579 28661
rect 9581 28656 11579 28658
rect 9581 28600 9586 28656
rect 9642 28600 11518 28656
rect 11574 28600 11579 28656
rect 9581 28598 11579 28600
rect 5533 28595 5599 28598
rect 9581 28595 9647 28598
rect 11513 28595 11579 28598
rect 6729 28522 6795 28525
rect 8845 28522 8911 28525
rect 6729 28520 8911 28522
rect 6729 28464 6734 28520
rect 6790 28464 8850 28520
rect 8906 28464 8911 28520
rect 6729 28462 8911 28464
rect 6729 28459 6795 28462
rect 8845 28459 8911 28462
rect 3610 28320 3930 28321
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3930 28320
rect 3610 28255 3930 28256
rect 8944 28320 9264 28321
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 28255 9264 28256
rect 14277 28320 14597 28321
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 28255 14597 28256
rect 11329 28250 11395 28253
rect 11462 28250 11468 28252
rect 11329 28248 11468 28250
rect 11329 28192 11334 28248
rect 11390 28192 11468 28248
rect 11329 28190 11468 28192
rect 11329 28187 11395 28190
rect 11462 28188 11468 28190
rect 11532 28188 11538 28252
rect 9489 28114 9555 28117
rect 12617 28114 12683 28117
rect 9489 28112 12683 28114
rect 9489 28056 9494 28112
rect 9550 28056 12622 28112
rect 12678 28056 12683 28112
rect 9489 28054 12683 28056
rect 9489 28051 9555 28054
rect 12617 28051 12683 28054
rect 6277 27776 6597 27777
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 27711 6597 27712
rect 11610 27776 11930 27777
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 27711 11930 27712
rect 9305 27706 9371 27709
rect 11145 27706 11211 27709
rect 9305 27704 11211 27706
rect 9305 27648 9310 27704
rect 9366 27648 11150 27704
rect 11206 27648 11211 27704
rect 9305 27646 11211 27648
rect 9305 27643 9371 27646
rect 11145 27643 11211 27646
rect 2221 27570 2287 27573
rect 7189 27570 7255 27573
rect 2221 27568 7255 27570
rect 2221 27512 2226 27568
rect 2282 27512 7194 27568
rect 7250 27512 7255 27568
rect 2221 27510 7255 27512
rect 2221 27507 2287 27510
rect 7189 27507 7255 27510
rect 4613 27434 4679 27437
rect 9949 27434 10015 27437
rect 4613 27432 10015 27434
rect 4613 27376 4618 27432
rect 4674 27376 9954 27432
rect 10010 27376 10015 27432
rect 4613 27374 10015 27376
rect 4613 27371 4679 27374
rect 9949 27371 10015 27374
rect 3610 27232 3930 27233
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3930 27232
rect 3610 27167 3930 27168
rect 8944 27232 9264 27233
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 27167 9264 27168
rect 14277 27232 14597 27233
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 27167 14597 27168
rect 0 27026 480 27056
rect 4337 27026 4403 27029
rect 0 27024 4403 27026
rect 0 26968 4342 27024
rect 4398 26968 4403 27024
rect 0 26966 4403 26968
rect 0 26936 480 26966
rect 4337 26963 4403 26966
rect 6637 27026 6703 27029
rect 13353 27026 13419 27029
rect 6637 27024 13419 27026
rect 6637 26968 6642 27024
rect 6698 26968 13358 27024
rect 13414 26968 13419 27024
rect 6637 26966 13419 26968
rect 6637 26963 6703 26966
rect 13353 26963 13419 26966
rect 6277 26688 6597 26689
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 26623 6597 26624
rect 11610 26688 11930 26689
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 26623 11930 26624
rect 3610 26144 3930 26145
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3930 26144
rect 3610 26079 3930 26080
rect 8944 26144 9264 26145
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 26079 9264 26080
rect 14277 26144 14597 26145
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 26079 14597 26080
rect 6277 25600 6597 25601
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 25535 6597 25536
rect 11610 25600 11930 25601
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 25535 11930 25536
rect 8753 25394 8819 25397
rect 9949 25394 10015 25397
rect 8753 25392 10015 25394
rect 8753 25336 8758 25392
rect 8814 25336 9954 25392
rect 10010 25336 10015 25392
rect 8753 25334 10015 25336
rect 8753 25331 8819 25334
rect 9949 25331 10015 25334
rect 3610 25056 3930 25057
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3930 25056
rect 3610 24991 3930 24992
rect 8944 25056 9264 25057
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 24991 9264 24992
rect 14277 25056 14597 25057
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 24991 14597 24992
rect 9397 24986 9463 24989
rect 9857 24986 9923 24989
rect 9397 24984 9923 24986
rect 9397 24928 9402 24984
rect 9458 24928 9862 24984
rect 9918 24928 9923 24984
rect 9397 24926 9923 24928
rect 9397 24923 9463 24926
rect 9857 24923 9923 24926
rect 11973 24986 12039 24989
rect 13629 24986 13695 24989
rect 11973 24984 13695 24986
rect 11973 24928 11978 24984
rect 12034 24928 13634 24984
rect 13690 24928 13695 24984
rect 11973 24926 13695 24928
rect 11973 24923 12039 24926
rect 13629 24923 13695 24926
rect 8017 24850 8083 24853
rect 11421 24850 11487 24853
rect 8017 24848 11487 24850
rect 8017 24792 8022 24848
rect 8078 24792 11426 24848
rect 11482 24792 11487 24848
rect 8017 24790 11487 24792
rect 8017 24787 8083 24790
rect 11421 24787 11487 24790
rect 5349 24714 5415 24717
rect 7465 24714 7531 24717
rect 5349 24712 7531 24714
rect 5349 24656 5354 24712
rect 5410 24656 7470 24712
rect 7526 24656 7531 24712
rect 5349 24654 7531 24656
rect 5349 24651 5415 24654
rect 7465 24651 7531 24654
rect 0 24578 480 24608
rect 1577 24578 1643 24581
rect 0 24576 1643 24578
rect 0 24520 1582 24576
rect 1638 24520 1643 24576
rect 0 24518 1643 24520
rect 0 24488 480 24518
rect 1577 24515 1643 24518
rect 6277 24512 6597 24513
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 24447 6597 24448
rect 11610 24512 11930 24513
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 24447 11930 24448
rect 7925 24306 7991 24309
rect 10593 24306 10659 24309
rect 7925 24304 10659 24306
rect 7925 24248 7930 24304
rect 7986 24248 10598 24304
rect 10654 24248 10659 24304
rect 7925 24246 10659 24248
rect 7925 24243 7991 24246
rect 10593 24243 10659 24246
rect 3610 23968 3930 23969
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3930 23968
rect 3610 23903 3930 23904
rect 8944 23968 9264 23969
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 23903 9264 23904
rect 14277 23968 14597 23969
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 23903 14597 23904
rect 4153 23762 4219 23765
rect 8845 23762 8911 23765
rect 4153 23760 8911 23762
rect 4153 23704 4158 23760
rect 4214 23704 8850 23760
rect 8906 23704 8911 23760
rect 4153 23702 8911 23704
rect 4153 23699 4219 23702
rect 8845 23699 8911 23702
rect 4797 23626 4863 23629
rect 6913 23626 6979 23629
rect 4797 23624 6979 23626
rect 4797 23568 4802 23624
rect 4858 23568 6918 23624
rect 6974 23568 6979 23624
rect 4797 23566 6979 23568
rect 4797 23563 4863 23566
rect 6913 23563 6979 23566
rect 6277 23424 6597 23425
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 23359 6597 23360
rect 11610 23424 11930 23425
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 23359 11930 23360
rect 7097 23354 7163 23357
rect 7097 23352 7666 23354
rect 7097 23296 7102 23352
rect 7158 23296 7666 23352
rect 7097 23294 7666 23296
rect 7097 23291 7163 23294
rect 5257 23218 5323 23221
rect 7465 23218 7531 23221
rect 5257 23216 7531 23218
rect 5257 23160 5262 23216
rect 5318 23160 7470 23216
rect 7526 23160 7531 23216
rect 5257 23158 7531 23160
rect 7606 23218 7666 23294
rect 12985 23218 13051 23221
rect 7606 23216 13051 23218
rect 7606 23160 12990 23216
rect 13046 23160 13051 23216
rect 7606 23158 13051 23160
rect 5257 23155 5323 23158
rect 7465 23155 7531 23158
rect 12985 23155 13051 23158
rect 5257 23082 5323 23085
rect 9397 23082 9463 23085
rect 5257 23080 9463 23082
rect 5257 23024 5262 23080
rect 5318 23024 9402 23080
rect 9458 23024 9463 23080
rect 5257 23022 9463 23024
rect 5257 23019 5323 23022
rect 9397 23019 9463 23022
rect 3610 22880 3930 22881
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3930 22880
rect 3610 22815 3930 22816
rect 8944 22880 9264 22881
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 22815 9264 22816
rect 14277 22880 14597 22881
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 22815 14597 22816
rect 7281 22674 7347 22677
rect 13537 22674 13603 22677
rect 7281 22672 13603 22674
rect 7281 22616 7286 22672
rect 7342 22616 13542 22672
rect 13598 22616 13603 22672
rect 7281 22614 13603 22616
rect 7281 22611 7347 22614
rect 13537 22611 13603 22614
rect 6277 22336 6597 22337
rect 0 22266 480 22296
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 22271 6597 22272
rect 11610 22336 11930 22337
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 22271 11930 22272
rect 1669 22266 1735 22269
rect 0 22264 1735 22266
rect 0 22208 1674 22264
rect 1730 22208 1735 22264
rect 0 22206 1735 22208
rect 0 22176 480 22206
rect 1669 22203 1735 22206
rect 4797 22130 4863 22133
rect 8201 22130 8267 22133
rect 4797 22128 8267 22130
rect 4797 22072 4802 22128
rect 4858 22072 8206 22128
rect 8262 22072 8267 22128
rect 4797 22070 8267 22072
rect 4797 22067 4863 22070
rect 8201 22067 8267 22070
rect 3610 21792 3930 21793
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3930 21792
rect 3610 21727 3930 21728
rect 8944 21792 9264 21793
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 21727 9264 21728
rect 14277 21792 14597 21793
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 21727 14597 21728
rect 6277 21248 6597 21249
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 21183 6597 21184
rect 11610 21248 11930 21249
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 21183 11930 21184
rect 7649 21042 7715 21045
rect 11329 21042 11395 21045
rect 7649 21040 11395 21042
rect 7649 20984 7654 21040
rect 7710 20984 11334 21040
rect 11390 20984 11395 21040
rect 7649 20982 11395 20984
rect 7649 20979 7715 20982
rect 11329 20979 11395 20982
rect 3610 20704 3930 20705
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3930 20704
rect 3610 20639 3930 20640
rect 8944 20704 9264 20705
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 20639 9264 20640
rect 14277 20704 14597 20705
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 20639 14597 20640
rect 1393 20362 1459 20365
rect 9673 20362 9739 20365
rect 1393 20360 9739 20362
rect 1393 20304 1398 20360
rect 1454 20304 9678 20360
rect 9734 20304 9739 20360
rect 1393 20302 9739 20304
rect 1393 20299 1459 20302
rect 9673 20299 9739 20302
rect 1669 20226 1735 20229
rect 6085 20226 6151 20229
rect 1669 20224 6151 20226
rect 1669 20168 1674 20224
rect 1730 20168 6090 20224
rect 6146 20168 6151 20224
rect 1669 20166 6151 20168
rect 1669 20163 1735 20166
rect 6085 20163 6151 20166
rect 6277 20160 6597 20161
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 20095 6597 20096
rect 11610 20160 11930 20161
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 20095 11930 20096
rect 0 19954 480 19984
rect 1669 19954 1735 19957
rect 0 19952 1735 19954
rect 0 19896 1674 19952
rect 1730 19896 1735 19952
rect 0 19894 1735 19896
rect 0 19864 480 19894
rect 1669 19891 1735 19894
rect 7557 19954 7623 19957
rect 11789 19954 11855 19957
rect 7557 19952 11855 19954
rect 7557 19896 7562 19952
rect 7618 19896 11794 19952
rect 11850 19896 11855 19952
rect 7557 19894 11855 19896
rect 7557 19891 7623 19894
rect 11789 19891 11855 19894
rect 6453 19818 6519 19821
rect 7005 19818 7071 19821
rect 6453 19816 7071 19818
rect 6453 19760 6458 19816
rect 6514 19760 7010 19816
rect 7066 19760 7071 19816
rect 6453 19758 7071 19760
rect 6453 19755 6519 19758
rect 7005 19755 7071 19758
rect 7281 19818 7347 19821
rect 9673 19818 9739 19821
rect 7281 19816 9739 19818
rect 7281 19760 7286 19816
rect 7342 19760 9678 19816
rect 9734 19760 9739 19816
rect 7281 19758 9739 19760
rect 7281 19755 7347 19758
rect 9673 19755 9739 19758
rect 11462 19756 11468 19820
rect 11532 19818 11538 19820
rect 12065 19818 12131 19821
rect 11532 19816 12131 19818
rect 11532 19760 12070 19816
rect 12126 19760 12131 19816
rect 11532 19758 12131 19760
rect 11532 19756 11538 19758
rect 12065 19755 12131 19758
rect 3610 19616 3930 19617
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3930 19616
rect 3610 19551 3930 19552
rect 8944 19616 9264 19617
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 19551 9264 19552
rect 14277 19616 14597 19617
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 19551 14597 19552
rect 8661 19410 8727 19413
rect 13077 19410 13143 19413
rect 8661 19408 13143 19410
rect 8661 19352 8666 19408
rect 8722 19352 13082 19408
rect 13138 19352 13143 19408
rect 8661 19350 13143 19352
rect 8661 19347 8727 19350
rect 13077 19347 13143 19350
rect 4705 19274 4771 19277
rect 5073 19274 5139 19277
rect 8845 19274 8911 19277
rect 4705 19272 8911 19274
rect 4705 19216 4710 19272
rect 4766 19216 5078 19272
rect 5134 19216 8850 19272
rect 8906 19216 8911 19272
rect 4705 19214 8911 19216
rect 4705 19211 4771 19214
rect 5073 19211 5139 19214
rect 8845 19211 8911 19214
rect 6277 19072 6597 19073
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 19007 6597 19008
rect 11610 19072 11930 19073
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 19007 11930 19008
rect 6729 19002 6795 19005
rect 7281 19002 7347 19005
rect 8385 19002 8451 19005
rect 6729 19000 8451 19002
rect 6729 18944 6734 19000
rect 6790 18944 7286 19000
rect 7342 18944 8390 19000
rect 8446 18944 8451 19000
rect 6729 18942 8451 18944
rect 6729 18939 6795 18942
rect 7281 18939 7347 18942
rect 8385 18939 8451 18942
rect 5717 18866 5783 18869
rect 7189 18866 7255 18869
rect 11973 18866 12039 18869
rect 5717 18864 12039 18866
rect 5717 18808 5722 18864
rect 5778 18808 7194 18864
rect 7250 18808 11978 18864
rect 12034 18808 12039 18864
rect 5717 18806 12039 18808
rect 5717 18803 5783 18806
rect 7189 18803 7255 18806
rect 11973 18803 12039 18806
rect 7097 18730 7163 18733
rect 11697 18730 11763 18733
rect 7097 18728 11763 18730
rect 7097 18672 7102 18728
rect 7158 18672 11702 18728
rect 11758 18672 11763 18728
rect 7097 18670 11763 18672
rect 7097 18667 7163 18670
rect 3610 18528 3930 18529
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3930 18528
rect 3610 18463 3930 18464
rect 7974 18189 8034 18670
rect 11697 18667 11763 18670
rect 8944 18528 9264 18529
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 18463 9264 18464
rect 14277 18528 14597 18529
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 18463 14597 18464
rect 7974 18184 8083 18189
rect 7974 18128 8022 18184
rect 8078 18128 8083 18184
rect 7974 18126 8083 18128
rect 8017 18123 8083 18126
rect 8385 18186 8451 18189
rect 12433 18186 12499 18189
rect 8385 18184 12499 18186
rect 8385 18128 8390 18184
rect 8446 18128 12438 18184
rect 12494 18128 12499 18184
rect 8385 18126 12499 18128
rect 8385 18123 8451 18126
rect 12433 18123 12499 18126
rect 3049 18050 3115 18053
rect 3325 18050 3391 18053
rect 3049 18048 3391 18050
rect 3049 17992 3054 18048
rect 3110 17992 3330 18048
rect 3386 17992 3391 18048
rect 3049 17990 3391 17992
rect 3049 17987 3115 17990
rect 3325 17987 3391 17990
rect 6277 17984 6597 17985
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 17919 6597 17920
rect 11610 17984 11930 17985
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 17919 11930 17920
rect 2773 17778 2839 17781
rect 9673 17778 9739 17781
rect 2773 17776 9739 17778
rect 2773 17720 2778 17776
rect 2834 17720 9678 17776
rect 9734 17720 9739 17776
rect 2773 17718 9739 17720
rect 2773 17715 2839 17718
rect 9673 17715 9739 17718
rect 0 17642 480 17672
rect 1577 17642 1643 17645
rect 0 17640 1643 17642
rect 0 17584 1582 17640
rect 1638 17584 1643 17640
rect 0 17582 1643 17584
rect 0 17552 480 17582
rect 1577 17579 1643 17582
rect 3610 17440 3930 17441
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3930 17440
rect 3610 17375 3930 17376
rect 8944 17440 9264 17441
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 17375 9264 17376
rect 14277 17440 14597 17441
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 17375 14597 17376
rect 3969 17098 4035 17101
rect 9622 17098 9628 17100
rect 3969 17096 9628 17098
rect 3969 17040 3974 17096
rect 4030 17040 9628 17096
rect 3969 17038 9628 17040
rect 3969 17035 4035 17038
rect 9622 17036 9628 17038
rect 9692 17098 9698 17100
rect 9949 17098 10015 17101
rect 9692 17096 10015 17098
rect 9692 17040 9954 17096
rect 10010 17040 10015 17096
rect 9692 17038 10015 17040
rect 9692 17036 9698 17038
rect 9949 17035 10015 17038
rect 12433 16962 12499 16965
rect 12433 16960 12634 16962
rect 12433 16904 12438 16960
rect 12494 16904 12634 16960
rect 12433 16902 12634 16904
rect 12433 16899 12499 16902
rect 6277 16896 6597 16897
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 16831 6597 16832
rect 11610 16896 11930 16897
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 16831 11930 16832
rect 5901 16828 5967 16829
rect 5901 16824 5948 16828
rect 6012 16826 6018 16828
rect 5901 16768 5906 16824
rect 5901 16764 5948 16768
rect 6012 16766 6058 16826
rect 6012 16764 6018 16766
rect 5901 16763 5967 16764
rect 12574 16693 12634 16902
rect 12574 16688 12683 16693
rect 12574 16632 12622 16688
rect 12678 16632 12683 16688
rect 12574 16630 12683 16632
rect 12617 16627 12683 16630
rect 6729 16554 6795 16557
rect 11329 16554 11395 16557
rect 6729 16552 11395 16554
rect 6729 16496 6734 16552
rect 6790 16496 11334 16552
rect 11390 16496 11395 16552
rect 6729 16494 11395 16496
rect 6729 16491 6795 16494
rect 11329 16491 11395 16494
rect 3610 16352 3930 16353
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3930 16352
rect 3610 16287 3930 16288
rect 8944 16352 9264 16353
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 16287 9264 16288
rect 14277 16352 14597 16353
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 16287 14597 16288
rect 9213 16146 9279 16149
rect 11329 16146 11395 16149
rect 9213 16144 11395 16146
rect 9213 16088 9218 16144
rect 9274 16088 11334 16144
rect 11390 16088 11395 16144
rect 9213 16086 11395 16088
rect 9213 16083 9279 16086
rect 11329 16083 11395 16086
rect 2221 15874 2287 15877
rect 5533 15874 5599 15877
rect 2221 15872 5599 15874
rect 2221 15816 2226 15872
rect 2282 15816 5538 15872
rect 5594 15816 5599 15872
rect 2221 15814 5599 15816
rect 2221 15811 2287 15814
rect 5533 15811 5599 15814
rect 8293 15874 8359 15877
rect 8845 15874 8911 15877
rect 10777 15874 10843 15877
rect 8293 15872 10843 15874
rect 8293 15816 8298 15872
rect 8354 15816 8850 15872
rect 8906 15816 10782 15872
rect 10838 15816 10843 15872
rect 8293 15814 10843 15816
rect 8293 15811 8359 15814
rect 8845 15811 8911 15814
rect 10777 15811 10843 15814
rect 6277 15808 6597 15809
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 15743 6597 15744
rect 11610 15808 11930 15809
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 15743 11930 15744
rect 3610 15264 3930 15265
rect 0 15194 480 15224
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3930 15264
rect 3610 15199 3930 15200
rect 8944 15264 9264 15265
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 15199 9264 15200
rect 14277 15264 14597 15265
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 15199 14597 15200
rect 1669 15194 1735 15197
rect 0 15192 1735 15194
rect 0 15136 1674 15192
rect 1730 15136 1735 15192
rect 0 15134 1735 15136
rect 0 15104 480 15134
rect 1669 15131 1735 15134
rect 8109 15194 8175 15197
rect 8661 15194 8727 15197
rect 8109 15192 8727 15194
rect 8109 15136 8114 15192
rect 8170 15136 8666 15192
rect 8722 15136 8727 15192
rect 8109 15134 8727 15136
rect 8109 15131 8175 15134
rect 8661 15131 8727 15134
rect 8109 14922 8175 14925
rect 13261 14922 13327 14925
rect 8109 14920 13327 14922
rect 8109 14864 8114 14920
rect 8170 14864 13266 14920
rect 13322 14864 13327 14920
rect 8109 14862 13327 14864
rect 8109 14859 8175 14862
rect 13261 14859 13327 14862
rect 6277 14720 6597 14721
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 14655 6597 14656
rect 11610 14720 11930 14721
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 14655 11930 14656
rect 3610 14176 3930 14177
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3930 14176
rect 3610 14111 3930 14112
rect 8944 14176 9264 14177
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 14111 9264 14112
rect 14277 14176 14597 14177
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 14111 14597 14112
rect 2313 13834 2379 13837
rect 5441 13834 5507 13837
rect 2313 13832 5507 13834
rect 2313 13776 2318 13832
rect 2374 13776 5446 13832
rect 5502 13776 5507 13832
rect 2313 13774 5507 13776
rect 2313 13771 2379 13774
rect 5441 13771 5507 13774
rect 6085 13834 6151 13837
rect 8109 13834 8175 13837
rect 6085 13832 8175 13834
rect 6085 13776 6090 13832
rect 6146 13776 8114 13832
rect 8170 13776 8175 13832
rect 6085 13774 8175 13776
rect 6085 13771 6151 13774
rect 8109 13771 8175 13774
rect 6277 13632 6597 13633
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 13567 6597 13568
rect 11610 13632 11930 13633
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 13567 11930 13568
rect 1393 13426 1459 13429
rect 9673 13426 9739 13429
rect 1393 13424 9739 13426
rect 1393 13368 1398 13424
rect 1454 13368 9678 13424
rect 9734 13368 9739 13424
rect 1393 13366 9739 13368
rect 1393 13363 1459 13366
rect 9673 13363 9739 13366
rect 5257 13290 5323 13293
rect 8937 13290 9003 13293
rect 9305 13290 9371 13293
rect 5257 13288 9371 13290
rect 5257 13232 5262 13288
rect 5318 13232 8942 13288
rect 8998 13232 9310 13288
rect 9366 13232 9371 13288
rect 5257 13230 9371 13232
rect 5257 13227 5323 13230
rect 8937 13227 9003 13230
rect 9305 13227 9371 13230
rect 3610 13088 3930 13089
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3930 13088
rect 3610 13023 3930 13024
rect 8944 13088 9264 13089
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 13023 9264 13024
rect 14277 13088 14597 13089
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 13023 14597 13024
rect 0 12882 480 12912
rect 1577 12882 1643 12885
rect 0 12880 1643 12882
rect 0 12824 1582 12880
rect 1638 12824 1643 12880
rect 0 12822 1643 12824
rect 0 12792 480 12822
rect 1577 12819 1643 12822
rect 2681 12882 2747 12885
rect 4613 12882 4679 12885
rect 2681 12880 4679 12882
rect 2681 12824 2686 12880
rect 2742 12824 4618 12880
rect 4674 12824 4679 12880
rect 2681 12822 4679 12824
rect 2681 12819 2747 12822
rect 4613 12819 4679 12822
rect 5441 12882 5507 12885
rect 10685 12882 10751 12885
rect 5441 12880 10751 12882
rect 5441 12824 5446 12880
rect 5502 12824 10690 12880
rect 10746 12824 10751 12880
rect 5441 12822 10751 12824
rect 5441 12819 5507 12822
rect 10685 12819 10751 12822
rect 8293 12610 8359 12613
rect 8661 12610 8727 12613
rect 8293 12608 8727 12610
rect 8293 12552 8298 12608
rect 8354 12552 8666 12608
rect 8722 12552 8727 12608
rect 8293 12550 8727 12552
rect 8293 12547 8359 12550
rect 8661 12547 8727 12550
rect 6277 12544 6597 12545
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 12479 6597 12480
rect 11610 12544 11930 12545
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 12479 11930 12480
rect 10225 12474 10291 12477
rect 10182 12472 10291 12474
rect 10182 12416 10230 12472
rect 10286 12416 10291 12472
rect 10182 12411 10291 12416
rect 10182 12341 10242 12411
rect 4613 12338 4679 12341
rect 9622 12338 9628 12340
rect 4613 12336 9628 12338
rect 4613 12280 4618 12336
rect 4674 12280 9628 12336
rect 4613 12278 9628 12280
rect 4613 12275 4679 12278
rect 9622 12276 9628 12278
rect 9692 12338 9698 12340
rect 10041 12338 10107 12341
rect 9692 12336 10107 12338
rect 9692 12280 10046 12336
rect 10102 12280 10107 12336
rect 9692 12278 10107 12280
rect 10182 12336 10291 12341
rect 10182 12280 10230 12336
rect 10286 12280 10291 12336
rect 10182 12278 10291 12280
rect 9692 12276 9698 12278
rect 10041 12275 10107 12278
rect 10225 12275 10291 12278
rect 5901 12204 5967 12205
rect 5901 12202 5948 12204
rect 5856 12200 5948 12202
rect 5856 12144 5906 12200
rect 5856 12142 5948 12144
rect 5901 12140 5948 12142
rect 6012 12140 6018 12204
rect 6821 12202 6887 12205
rect 8477 12202 8543 12205
rect 6821 12200 8543 12202
rect 6821 12144 6826 12200
rect 6882 12144 8482 12200
rect 8538 12144 8543 12200
rect 6821 12142 8543 12144
rect 5901 12139 5967 12140
rect 6821 12139 6887 12142
rect 8477 12139 8543 12142
rect 9581 12202 9647 12205
rect 10961 12202 11027 12205
rect 9581 12200 11027 12202
rect 9581 12144 9586 12200
rect 9642 12144 10966 12200
rect 11022 12144 11027 12200
rect 9581 12142 11027 12144
rect 9581 12139 9647 12142
rect 10961 12139 11027 12142
rect 3610 12000 3930 12001
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3930 12000
rect 3610 11935 3930 11936
rect 8944 12000 9264 12001
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 11935 9264 11936
rect 14277 12000 14597 12001
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 11935 14597 11936
rect 7373 11794 7439 11797
rect 11237 11794 11303 11797
rect 7373 11792 11303 11794
rect 7373 11736 7378 11792
rect 7434 11736 11242 11792
rect 11298 11736 11303 11792
rect 7373 11734 11303 11736
rect 7373 11731 7439 11734
rect 11237 11731 11303 11734
rect 10041 11522 10107 11525
rect 11145 11522 11211 11525
rect 10041 11520 11211 11522
rect 10041 11464 10046 11520
rect 10102 11464 11150 11520
rect 11206 11464 11211 11520
rect 10041 11462 11211 11464
rect 10041 11459 10107 11462
rect 11145 11459 11211 11462
rect 6277 11456 6597 11457
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 11391 6597 11392
rect 11610 11456 11930 11457
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 11391 11930 11392
rect 6729 11250 6795 11253
rect 9397 11250 9463 11253
rect 6729 11248 9463 11250
rect 6729 11192 6734 11248
rect 6790 11192 9402 11248
rect 9458 11192 9463 11248
rect 6729 11190 9463 11192
rect 6729 11187 6795 11190
rect 9397 11187 9463 11190
rect 7005 11114 7071 11117
rect 8661 11114 8727 11117
rect 7005 11112 8727 11114
rect 7005 11056 7010 11112
rect 7066 11056 8666 11112
rect 8722 11056 8727 11112
rect 7005 11054 8727 11056
rect 7005 11051 7071 11054
rect 8661 11051 8727 11054
rect 3610 10912 3930 10913
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3930 10912
rect 3610 10847 3930 10848
rect 8944 10912 9264 10913
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 10847 9264 10848
rect 14277 10912 14597 10913
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 10847 14597 10848
rect 4521 10706 4587 10709
rect 5073 10706 5139 10709
rect 9673 10706 9739 10709
rect 4521 10704 9739 10706
rect 4521 10648 4526 10704
rect 4582 10648 5078 10704
rect 5134 10648 9678 10704
rect 9734 10648 9739 10704
rect 4521 10646 9739 10648
rect 4521 10643 4587 10646
rect 5073 10643 5139 10646
rect 9673 10643 9739 10646
rect 0 10570 480 10600
rect 1577 10570 1643 10573
rect 0 10568 1643 10570
rect 0 10512 1582 10568
rect 1638 10512 1643 10568
rect 0 10510 1643 10512
rect 0 10480 480 10510
rect 1577 10507 1643 10510
rect 8753 10434 8819 10437
rect 9673 10434 9739 10437
rect 8753 10432 9739 10434
rect 8753 10376 8758 10432
rect 8814 10376 9678 10432
rect 9734 10376 9739 10432
rect 8753 10374 9739 10376
rect 8753 10371 8819 10374
rect 9673 10371 9739 10374
rect 6277 10368 6597 10369
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 10303 6597 10304
rect 11610 10368 11930 10369
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 10303 11930 10304
rect 12341 10162 12407 10165
rect 14825 10162 14891 10165
rect 12341 10160 14891 10162
rect 12341 10104 12346 10160
rect 12402 10104 14830 10160
rect 14886 10104 14891 10160
rect 12341 10102 14891 10104
rect 12341 10099 12407 10102
rect 14825 10099 14891 10102
rect 4245 10026 4311 10029
rect 8477 10026 8543 10029
rect 10501 10026 10567 10029
rect 4245 10024 10567 10026
rect 4245 9968 4250 10024
rect 4306 9968 8482 10024
rect 8538 9968 10506 10024
rect 10562 9968 10567 10024
rect 4245 9966 10567 9968
rect 4245 9963 4311 9966
rect 8477 9963 8543 9966
rect 10501 9963 10567 9966
rect 11237 10026 11303 10029
rect 15520 10026 16000 10056
rect 11237 10024 16000 10026
rect 11237 9968 11242 10024
rect 11298 9968 16000 10024
rect 11237 9966 16000 9968
rect 11237 9963 11303 9966
rect 15520 9936 16000 9966
rect 3610 9824 3930 9825
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3930 9824
rect 3610 9759 3930 9760
rect 8944 9824 9264 9825
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 9759 9264 9760
rect 14277 9824 14597 9825
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 9759 14597 9760
rect 6177 9482 6243 9485
rect 7741 9482 7807 9485
rect 6177 9480 7807 9482
rect 6177 9424 6182 9480
rect 6238 9424 7746 9480
rect 7802 9424 7807 9480
rect 6177 9422 7807 9424
rect 6177 9419 6243 9422
rect 7741 9419 7807 9422
rect 6277 9280 6597 9281
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 9215 6597 9216
rect 11610 9280 11930 9281
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 9215 11930 9216
rect 2681 8938 2747 8941
rect 9581 8938 9647 8941
rect 2681 8936 9647 8938
rect 2681 8880 2686 8936
rect 2742 8880 9586 8936
rect 9642 8880 9647 8936
rect 2681 8878 9647 8880
rect 2681 8875 2747 8878
rect 9581 8875 9647 8878
rect 3610 8736 3930 8737
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3930 8736
rect 3610 8671 3930 8672
rect 8944 8736 9264 8737
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 8671 9264 8672
rect 14277 8736 14597 8737
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 8671 14597 8672
rect 5441 8530 5507 8533
rect 8201 8530 8267 8533
rect 5441 8528 8267 8530
rect 5441 8472 5446 8528
rect 5502 8472 8206 8528
rect 8262 8472 8267 8528
rect 5441 8470 8267 8472
rect 5441 8467 5507 8470
rect 8201 8467 8267 8470
rect 2773 8394 2839 8397
rect 9949 8394 10015 8397
rect 2773 8392 10015 8394
rect 2773 8336 2778 8392
rect 2834 8336 9954 8392
rect 10010 8336 10015 8392
rect 2773 8334 10015 8336
rect 2773 8331 2839 8334
rect 9949 8331 10015 8334
rect 9305 8258 9371 8261
rect 10317 8258 10383 8261
rect 9305 8256 10383 8258
rect 9305 8200 9310 8256
rect 9366 8200 10322 8256
rect 10378 8200 10383 8256
rect 9305 8198 10383 8200
rect 9305 8195 9371 8198
rect 10317 8195 10383 8198
rect 6277 8192 6597 8193
rect 0 8122 480 8152
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 8127 6597 8128
rect 11610 8192 11930 8193
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 8127 11930 8128
rect 1577 8122 1643 8125
rect 0 8120 1643 8122
rect 0 8064 1582 8120
rect 1638 8064 1643 8120
rect 0 8062 1643 8064
rect 0 8032 480 8062
rect 1577 8059 1643 8062
rect 9305 8122 9371 8125
rect 10409 8122 10475 8125
rect 9305 8120 10475 8122
rect 9305 8064 9310 8120
rect 9366 8064 10414 8120
rect 10470 8064 10475 8120
rect 9305 8062 10475 8064
rect 9305 8059 9371 8062
rect 10409 8059 10475 8062
rect 7189 7986 7255 7989
rect 12249 7986 12315 7989
rect 7189 7984 12315 7986
rect 7189 7928 7194 7984
rect 7250 7928 12254 7984
rect 12310 7928 12315 7984
rect 7189 7926 12315 7928
rect 7189 7923 7255 7926
rect 12249 7923 12315 7926
rect 9857 7850 9923 7853
rect 12893 7850 12959 7853
rect 9857 7848 12959 7850
rect 9857 7792 9862 7848
rect 9918 7792 12898 7848
rect 12954 7792 12959 7848
rect 9857 7790 12959 7792
rect 9857 7787 9923 7790
rect 12893 7787 12959 7790
rect 3610 7648 3930 7649
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3930 7648
rect 3610 7583 3930 7584
rect 8944 7648 9264 7649
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 7583 9264 7584
rect 14277 7648 14597 7649
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 7583 14597 7584
rect 1669 7442 1735 7445
rect 4981 7442 5047 7445
rect 1669 7440 5047 7442
rect 1669 7384 1674 7440
rect 1730 7384 4986 7440
rect 5042 7384 5047 7440
rect 1669 7382 5047 7384
rect 1669 7379 1735 7382
rect 4981 7379 5047 7382
rect 5901 7442 5967 7445
rect 10133 7442 10199 7445
rect 5901 7440 10199 7442
rect 5901 7384 5906 7440
rect 5962 7384 10138 7440
rect 10194 7384 10199 7440
rect 5901 7382 10199 7384
rect 5901 7379 5967 7382
rect 10133 7379 10199 7382
rect 8569 7306 8635 7309
rect 15377 7306 15443 7309
rect 8569 7304 15443 7306
rect 8569 7248 8574 7304
rect 8630 7248 15382 7304
rect 15438 7248 15443 7304
rect 8569 7246 15443 7248
rect 8569 7243 8635 7246
rect 15377 7243 15443 7246
rect 6277 7104 6597 7105
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 7039 6597 7040
rect 11610 7104 11930 7105
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 7039 11930 7040
rect 1485 6898 1551 6901
rect 6821 6898 6887 6901
rect 1485 6896 6887 6898
rect 1485 6840 1490 6896
rect 1546 6840 6826 6896
rect 6882 6840 6887 6896
rect 1485 6838 6887 6840
rect 1485 6835 1551 6838
rect 6821 6835 6887 6838
rect 1393 6762 1459 6765
rect 2865 6762 2931 6765
rect 1393 6760 2931 6762
rect 1393 6704 1398 6760
rect 1454 6704 2870 6760
rect 2926 6704 2931 6760
rect 1393 6702 2931 6704
rect 1393 6699 1459 6702
rect 2865 6699 2931 6702
rect 5625 6762 5691 6765
rect 5625 6760 9506 6762
rect 5625 6704 5630 6760
rect 5686 6704 9506 6760
rect 5625 6702 9506 6704
rect 5625 6699 5691 6702
rect 9446 6626 9506 6702
rect 12157 6626 12223 6629
rect 9446 6624 12223 6626
rect 9446 6568 12162 6624
rect 12218 6568 12223 6624
rect 9446 6566 12223 6568
rect 12157 6563 12223 6566
rect 3610 6560 3930 6561
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3930 6560
rect 3610 6495 3930 6496
rect 8944 6560 9264 6561
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 6495 9264 6496
rect 14277 6560 14597 6561
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 6495 14597 6496
rect 9397 6356 9463 6357
rect 9397 6352 9444 6356
rect 9508 6354 9514 6356
rect 9397 6296 9402 6352
rect 9397 6292 9444 6296
rect 9508 6294 9554 6354
rect 9508 6292 9514 6294
rect 9397 6291 9463 6292
rect 2589 6082 2655 6085
rect 4337 6082 4403 6085
rect 2589 6080 4403 6082
rect 2589 6024 2594 6080
rect 2650 6024 4342 6080
rect 4398 6024 4403 6080
rect 2589 6022 4403 6024
rect 2589 6019 2655 6022
rect 4337 6019 4403 6022
rect 6277 6016 6597 6017
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 5951 6597 5952
rect 11610 6016 11930 6017
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 5951 11930 5952
rect 11145 5946 11211 5949
rect 6686 5944 11211 5946
rect 6686 5888 11150 5944
rect 11206 5888 11211 5944
rect 6686 5886 11211 5888
rect 0 5810 480 5840
rect 1577 5810 1643 5813
rect 0 5808 1643 5810
rect 0 5752 1582 5808
rect 1638 5752 1643 5808
rect 0 5750 1643 5752
rect 0 5720 480 5750
rect 1577 5747 1643 5750
rect 4061 5810 4127 5813
rect 6269 5810 6335 5813
rect 4061 5808 6335 5810
rect 4061 5752 4066 5808
rect 4122 5752 6274 5808
rect 6330 5752 6335 5808
rect 4061 5750 6335 5752
rect 4061 5747 4127 5750
rect 6269 5747 6335 5750
rect 4429 5674 4495 5677
rect 5809 5674 5875 5677
rect 6177 5674 6243 5677
rect 6686 5674 6746 5886
rect 11145 5883 11211 5886
rect 9305 5810 9371 5813
rect 11053 5810 11119 5813
rect 9305 5808 11119 5810
rect 9305 5752 9310 5808
rect 9366 5752 11058 5808
rect 11114 5752 11119 5808
rect 9305 5750 11119 5752
rect 9305 5747 9371 5750
rect 11053 5747 11119 5750
rect 4429 5672 5875 5674
rect 4429 5616 4434 5672
rect 4490 5616 5814 5672
rect 5870 5616 5875 5672
rect 4429 5614 5875 5616
rect 4429 5611 4495 5614
rect 5809 5611 5875 5614
rect 5950 5672 6746 5674
rect 5950 5616 6182 5672
rect 6238 5616 6746 5672
rect 5950 5614 6746 5616
rect 7373 5674 7439 5677
rect 9857 5674 9923 5677
rect 7373 5672 9923 5674
rect 7373 5616 7378 5672
rect 7434 5616 9862 5672
rect 9918 5616 9923 5672
rect 7373 5614 9923 5616
rect 4797 5538 4863 5541
rect 5950 5538 6010 5614
rect 6177 5611 6243 5614
rect 7373 5611 7439 5614
rect 9857 5611 9923 5614
rect 4797 5536 6010 5538
rect 4797 5480 4802 5536
rect 4858 5480 6010 5536
rect 4797 5478 6010 5480
rect 4797 5475 4863 5478
rect 3610 5472 3930 5473
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3930 5472
rect 3610 5407 3930 5408
rect 8944 5472 9264 5473
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 5407 9264 5408
rect 14277 5472 14597 5473
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 5407 14597 5408
rect 5441 5266 5507 5269
rect 12709 5266 12775 5269
rect 5441 5264 12775 5266
rect 5441 5208 5446 5264
rect 5502 5208 12714 5264
rect 12770 5208 12775 5264
rect 5441 5206 12775 5208
rect 5441 5203 5507 5206
rect 12709 5203 12775 5206
rect 10593 5130 10659 5133
rect 13353 5130 13419 5133
rect 5950 5070 7114 5130
rect 3877 4994 3943 4997
rect 5950 4994 6010 5070
rect 3877 4992 6010 4994
rect 3877 4936 3882 4992
rect 3938 4936 6010 4992
rect 3877 4934 6010 4936
rect 7054 4994 7114 5070
rect 10593 5128 13419 5130
rect 10593 5072 10598 5128
rect 10654 5072 13358 5128
rect 13414 5072 13419 5128
rect 10593 5070 13419 5072
rect 10593 5067 10659 5070
rect 13353 5067 13419 5070
rect 7465 4994 7531 4997
rect 11145 4994 11211 4997
rect 7054 4992 11211 4994
rect 7054 4936 7470 4992
rect 7526 4936 11150 4992
rect 11206 4936 11211 4992
rect 7054 4934 11211 4936
rect 3877 4931 3943 4934
rect 7465 4931 7531 4934
rect 11145 4931 11211 4934
rect 6277 4928 6597 4929
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 4863 6597 4864
rect 11610 4928 11930 4929
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 4863 11930 4864
rect 8569 4858 8635 4861
rect 6686 4856 8635 4858
rect 6686 4800 8574 4856
rect 8630 4800 8635 4856
rect 6686 4798 8635 4800
rect 6269 4722 6335 4725
rect 6686 4722 6746 4798
rect 8569 4795 8635 4798
rect 6269 4720 6746 4722
rect 6269 4664 6274 4720
rect 6330 4664 6746 4720
rect 6269 4662 6746 4664
rect 7189 4722 7255 4725
rect 14641 4722 14707 4725
rect 7189 4720 14707 4722
rect 7189 4664 7194 4720
rect 7250 4664 14646 4720
rect 14702 4664 14707 4720
rect 7189 4662 14707 4664
rect 6269 4659 6335 4662
rect 7189 4659 7255 4662
rect 14641 4659 14707 4662
rect 7833 4586 7899 4589
rect 12433 4586 12499 4589
rect 7833 4584 12499 4586
rect 7833 4528 7838 4584
rect 7894 4528 12438 4584
rect 12494 4528 12499 4584
rect 7833 4526 12499 4528
rect 7833 4523 7899 4526
rect 12433 4523 12499 4526
rect 3610 4384 3930 4385
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3930 4384
rect 3610 4319 3930 4320
rect 8944 4384 9264 4385
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 4319 9264 4320
rect 14277 4384 14597 4385
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 4319 14597 4320
rect 565 4314 631 4317
rect 2865 4314 2931 4317
rect 565 4312 2931 4314
rect 565 4256 570 4312
rect 626 4256 2870 4312
rect 2926 4256 2931 4312
rect 565 4254 2931 4256
rect 565 4251 631 4254
rect 2865 4251 2931 4254
rect 8017 4314 8083 4317
rect 8017 4312 8770 4314
rect 8017 4256 8022 4312
rect 8078 4256 8770 4312
rect 8017 4254 8770 4256
rect 8017 4251 8083 4254
rect 5073 4178 5139 4181
rect 8569 4178 8635 4181
rect 5073 4176 8635 4178
rect 5073 4120 5078 4176
rect 5134 4120 8574 4176
rect 8630 4120 8635 4176
rect 5073 4118 8635 4120
rect 8710 4178 8770 4254
rect 8710 4118 11346 4178
rect 5073 4115 5139 4118
rect 8569 4115 8635 4118
rect 6177 4042 6243 4045
rect 8477 4042 8543 4045
rect 6177 4040 8543 4042
rect 6177 3984 6182 4040
rect 6238 3984 8482 4040
rect 8538 3984 8543 4040
rect 6177 3982 8543 3984
rect 6177 3979 6243 3982
rect 8477 3979 8543 3982
rect 11286 3909 11346 4118
rect 13721 4042 13787 4045
rect 11470 4040 13787 4042
rect 11470 3984 13726 4040
rect 13782 3984 13787 4040
rect 11470 3982 13787 3984
rect 11286 3904 11395 3909
rect 11286 3848 11334 3904
rect 11390 3848 11395 3904
rect 11286 3846 11395 3848
rect 11329 3843 11395 3846
rect 6277 3840 6597 3841
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 3775 6597 3776
rect 6821 3770 6887 3773
rect 7097 3770 7163 3773
rect 11470 3770 11530 3982
rect 13721 3979 13787 3982
rect 11610 3840 11930 3841
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 3775 11930 3776
rect 6821 3768 11530 3770
rect 6821 3712 6826 3768
rect 6882 3712 7102 3768
rect 7158 3712 11530 3768
rect 6821 3710 11530 3712
rect 6821 3707 6887 3710
rect 7097 3707 7163 3710
rect 933 3634 999 3637
rect 7005 3634 7071 3637
rect 933 3632 7071 3634
rect 933 3576 938 3632
rect 994 3576 7010 3632
rect 7066 3576 7071 3632
rect 933 3574 7071 3576
rect 933 3571 999 3574
rect 7005 3571 7071 3574
rect 10501 3634 10567 3637
rect 12433 3634 12499 3637
rect 10501 3632 12499 3634
rect 10501 3576 10506 3632
rect 10562 3576 12438 3632
rect 12494 3576 12499 3632
rect 10501 3574 12499 3576
rect 10501 3571 10567 3574
rect 12433 3571 12499 3574
rect 0 3498 480 3528
rect 1577 3498 1643 3501
rect 0 3496 1643 3498
rect 0 3440 1582 3496
rect 1638 3440 1643 3496
rect 0 3438 1643 3440
rect 0 3408 480 3438
rect 1577 3435 1643 3438
rect 6637 3498 6703 3501
rect 13445 3498 13511 3501
rect 6637 3496 13511 3498
rect 6637 3440 6642 3496
rect 6698 3440 13450 3496
rect 13506 3440 13511 3496
rect 6637 3438 13511 3440
rect 6637 3435 6703 3438
rect 13445 3435 13511 3438
rect 13629 3498 13695 3501
rect 14181 3498 14247 3501
rect 13629 3496 14247 3498
rect 13629 3440 13634 3496
rect 13690 3440 14186 3496
rect 14242 3440 14247 3496
rect 13629 3438 14247 3440
rect 13629 3435 13695 3438
rect 14181 3435 14247 3438
rect 3610 3296 3930 3297
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3930 3296
rect 3610 3231 3930 3232
rect 8944 3296 9264 3297
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 3231 9264 3232
rect 14277 3296 14597 3297
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 3231 14597 3232
rect 8293 3090 8359 3093
rect 9765 3090 9831 3093
rect 8293 3088 9831 3090
rect 8293 3032 8298 3088
rect 8354 3032 9770 3088
rect 9826 3032 9831 3088
rect 8293 3030 9831 3032
rect 8293 3027 8359 3030
rect 9765 3027 9831 3030
rect 10225 3090 10291 3093
rect 12617 3090 12683 3093
rect 10225 3088 12683 3090
rect 10225 3032 10230 3088
rect 10286 3032 12622 3088
rect 12678 3032 12683 3088
rect 10225 3030 12683 3032
rect 10225 3027 10291 3030
rect 12617 3027 12683 3030
rect 2589 2954 2655 2957
rect 7005 2954 7071 2957
rect 2589 2952 7071 2954
rect 2589 2896 2594 2952
rect 2650 2896 7010 2952
rect 7066 2896 7071 2952
rect 2589 2894 7071 2896
rect 2589 2891 2655 2894
rect 7005 2891 7071 2894
rect 10041 2954 10107 2957
rect 12801 2954 12867 2957
rect 10041 2952 12867 2954
rect 10041 2896 10046 2952
rect 10102 2896 12806 2952
rect 12862 2896 12867 2952
rect 10041 2894 12867 2896
rect 10041 2891 10107 2894
rect 12801 2891 12867 2894
rect 1761 2818 1827 2821
rect 5625 2818 5691 2821
rect 1761 2816 5691 2818
rect 1761 2760 1766 2816
rect 1822 2760 5630 2816
rect 5686 2760 5691 2816
rect 1761 2758 5691 2760
rect 1761 2755 1827 2758
rect 5625 2755 5691 2758
rect 8293 2818 8359 2821
rect 11145 2818 11211 2821
rect 8293 2816 11211 2818
rect 8293 2760 8298 2816
rect 8354 2760 11150 2816
rect 11206 2760 11211 2816
rect 8293 2758 11211 2760
rect 8293 2755 8359 2758
rect 11145 2755 11211 2758
rect 6277 2752 6597 2753
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2687 6597 2688
rect 11610 2752 11930 2753
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2687 11930 2688
rect 4061 2682 4127 2685
rect 5993 2682 6059 2685
rect 9489 2684 9555 2685
rect 4061 2680 6059 2682
rect 4061 2624 4066 2680
rect 4122 2624 5998 2680
rect 6054 2624 6059 2680
rect 4061 2622 6059 2624
rect 4061 2619 4127 2622
rect 5993 2619 6059 2622
rect 9438 2620 9444 2684
rect 9508 2682 9555 2684
rect 9508 2680 9600 2682
rect 9550 2624 9600 2680
rect 9508 2622 9600 2624
rect 9508 2620 9555 2622
rect 9489 2619 9555 2620
rect 5625 2546 5691 2549
rect 11237 2546 11303 2549
rect 5625 2544 11303 2546
rect 5625 2488 5630 2544
rect 5686 2488 11242 2544
rect 11298 2488 11303 2544
rect 5625 2486 11303 2488
rect 5625 2483 5691 2486
rect 11237 2483 11303 2486
rect 2957 2410 3023 2413
rect 12801 2410 12867 2413
rect 2957 2408 12867 2410
rect 2957 2352 2962 2408
rect 3018 2352 12806 2408
rect 12862 2352 12867 2408
rect 2957 2350 12867 2352
rect 2957 2347 3023 2350
rect 12801 2347 12867 2350
rect 4521 2274 4587 2277
rect 8017 2274 8083 2277
rect 4521 2272 8083 2274
rect 4521 2216 4526 2272
rect 4582 2216 8022 2272
rect 8078 2216 8083 2272
rect 4521 2214 8083 2216
rect 4521 2211 4587 2214
rect 8017 2211 8083 2214
rect 3610 2208 3930 2209
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3930 2208
rect 3610 2143 3930 2144
rect 8944 2208 9264 2209
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2143 9264 2144
rect 14277 2208 14597 2209
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2143 14597 2144
rect 3325 1458 3391 1461
rect 7097 1458 7163 1461
rect 3325 1456 7163 1458
rect 3325 1400 3330 1456
rect 3386 1400 7102 1456
rect 7158 1400 7163 1456
rect 3325 1398 7163 1400
rect 3325 1395 3391 1398
rect 7097 1395 7163 1398
rect 0 1186 480 1216
rect 2773 1186 2839 1189
rect 0 1184 2839 1186
rect 0 1128 2778 1184
rect 2834 1128 2839 1184
rect 0 1126 2839 1128
rect 0 1096 480 1126
rect 2773 1123 2839 1126
<< via3 >>
rect 6285 37564 6349 37568
rect 6285 37508 6289 37564
rect 6289 37508 6345 37564
rect 6345 37508 6349 37564
rect 6285 37504 6349 37508
rect 6365 37564 6429 37568
rect 6365 37508 6369 37564
rect 6369 37508 6425 37564
rect 6425 37508 6429 37564
rect 6365 37504 6429 37508
rect 6445 37564 6509 37568
rect 6445 37508 6449 37564
rect 6449 37508 6505 37564
rect 6505 37508 6509 37564
rect 6445 37504 6509 37508
rect 6525 37564 6589 37568
rect 6525 37508 6529 37564
rect 6529 37508 6585 37564
rect 6585 37508 6589 37564
rect 6525 37504 6589 37508
rect 11618 37564 11682 37568
rect 11618 37508 11622 37564
rect 11622 37508 11678 37564
rect 11678 37508 11682 37564
rect 11618 37504 11682 37508
rect 11698 37564 11762 37568
rect 11698 37508 11702 37564
rect 11702 37508 11758 37564
rect 11758 37508 11762 37564
rect 11698 37504 11762 37508
rect 11778 37564 11842 37568
rect 11778 37508 11782 37564
rect 11782 37508 11838 37564
rect 11838 37508 11842 37564
rect 11778 37504 11842 37508
rect 11858 37564 11922 37568
rect 11858 37508 11862 37564
rect 11862 37508 11918 37564
rect 11918 37508 11922 37564
rect 11858 37504 11922 37508
rect 3618 37020 3682 37024
rect 3618 36964 3622 37020
rect 3622 36964 3678 37020
rect 3678 36964 3682 37020
rect 3618 36960 3682 36964
rect 3698 37020 3762 37024
rect 3698 36964 3702 37020
rect 3702 36964 3758 37020
rect 3758 36964 3762 37020
rect 3698 36960 3762 36964
rect 3778 37020 3842 37024
rect 3778 36964 3782 37020
rect 3782 36964 3838 37020
rect 3838 36964 3842 37020
rect 3778 36960 3842 36964
rect 3858 37020 3922 37024
rect 3858 36964 3862 37020
rect 3862 36964 3918 37020
rect 3918 36964 3922 37020
rect 3858 36960 3922 36964
rect 8952 37020 9016 37024
rect 8952 36964 8956 37020
rect 8956 36964 9012 37020
rect 9012 36964 9016 37020
rect 8952 36960 9016 36964
rect 9032 37020 9096 37024
rect 9032 36964 9036 37020
rect 9036 36964 9092 37020
rect 9092 36964 9096 37020
rect 9032 36960 9096 36964
rect 9112 37020 9176 37024
rect 9112 36964 9116 37020
rect 9116 36964 9172 37020
rect 9172 36964 9176 37020
rect 9112 36960 9176 36964
rect 9192 37020 9256 37024
rect 9192 36964 9196 37020
rect 9196 36964 9252 37020
rect 9252 36964 9256 37020
rect 9192 36960 9256 36964
rect 14285 37020 14349 37024
rect 14285 36964 14289 37020
rect 14289 36964 14345 37020
rect 14345 36964 14349 37020
rect 14285 36960 14349 36964
rect 14365 37020 14429 37024
rect 14365 36964 14369 37020
rect 14369 36964 14425 37020
rect 14425 36964 14429 37020
rect 14365 36960 14429 36964
rect 14445 37020 14509 37024
rect 14445 36964 14449 37020
rect 14449 36964 14505 37020
rect 14505 36964 14509 37020
rect 14445 36960 14509 36964
rect 14525 37020 14589 37024
rect 14525 36964 14529 37020
rect 14529 36964 14585 37020
rect 14585 36964 14589 37020
rect 14525 36960 14589 36964
rect 6285 36476 6349 36480
rect 6285 36420 6289 36476
rect 6289 36420 6345 36476
rect 6345 36420 6349 36476
rect 6285 36416 6349 36420
rect 6365 36476 6429 36480
rect 6365 36420 6369 36476
rect 6369 36420 6425 36476
rect 6425 36420 6429 36476
rect 6365 36416 6429 36420
rect 6445 36476 6509 36480
rect 6445 36420 6449 36476
rect 6449 36420 6505 36476
rect 6505 36420 6509 36476
rect 6445 36416 6509 36420
rect 6525 36476 6589 36480
rect 6525 36420 6529 36476
rect 6529 36420 6585 36476
rect 6585 36420 6589 36476
rect 6525 36416 6589 36420
rect 11618 36476 11682 36480
rect 11618 36420 11622 36476
rect 11622 36420 11678 36476
rect 11678 36420 11682 36476
rect 11618 36416 11682 36420
rect 11698 36476 11762 36480
rect 11698 36420 11702 36476
rect 11702 36420 11758 36476
rect 11758 36420 11762 36476
rect 11698 36416 11762 36420
rect 11778 36476 11842 36480
rect 11778 36420 11782 36476
rect 11782 36420 11838 36476
rect 11838 36420 11842 36476
rect 11778 36416 11842 36420
rect 11858 36476 11922 36480
rect 11858 36420 11862 36476
rect 11862 36420 11918 36476
rect 11918 36420 11922 36476
rect 11858 36416 11922 36420
rect 3618 35932 3682 35936
rect 3618 35876 3622 35932
rect 3622 35876 3678 35932
rect 3678 35876 3682 35932
rect 3618 35872 3682 35876
rect 3698 35932 3762 35936
rect 3698 35876 3702 35932
rect 3702 35876 3758 35932
rect 3758 35876 3762 35932
rect 3698 35872 3762 35876
rect 3778 35932 3842 35936
rect 3778 35876 3782 35932
rect 3782 35876 3838 35932
rect 3838 35876 3842 35932
rect 3778 35872 3842 35876
rect 3858 35932 3922 35936
rect 3858 35876 3862 35932
rect 3862 35876 3918 35932
rect 3918 35876 3922 35932
rect 3858 35872 3922 35876
rect 8952 35932 9016 35936
rect 8952 35876 8956 35932
rect 8956 35876 9012 35932
rect 9012 35876 9016 35932
rect 8952 35872 9016 35876
rect 9032 35932 9096 35936
rect 9032 35876 9036 35932
rect 9036 35876 9092 35932
rect 9092 35876 9096 35932
rect 9032 35872 9096 35876
rect 9112 35932 9176 35936
rect 9112 35876 9116 35932
rect 9116 35876 9172 35932
rect 9172 35876 9176 35932
rect 9112 35872 9176 35876
rect 9192 35932 9256 35936
rect 9192 35876 9196 35932
rect 9196 35876 9252 35932
rect 9252 35876 9256 35932
rect 9192 35872 9256 35876
rect 14285 35932 14349 35936
rect 14285 35876 14289 35932
rect 14289 35876 14345 35932
rect 14345 35876 14349 35932
rect 14285 35872 14349 35876
rect 14365 35932 14429 35936
rect 14365 35876 14369 35932
rect 14369 35876 14425 35932
rect 14425 35876 14429 35932
rect 14365 35872 14429 35876
rect 14445 35932 14509 35936
rect 14445 35876 14449 35932
rect 14449 35876 14505 35932
rect 14505 35876 14509 35932
rect 14445 35872 14509 35876
rect 14525 35932 14589 35936
rect 14525 35876 14529 35932
rect 14529 35876 14585 35932
rect 14585 35876 14589 35932
rect 14525 35872 14589 35876
rect 6285 35388 6349 35392
rect 6285 35332 6289 35388
rect 6289 35332 6345 35388
rect 6345 35332 6349 35388
rect 6285 35328 6349 35332
rect 6365 35388 6429 35392
rect 6365 35332 6369 35388
rect 6369 35332 6425 35388
rect 6425 35332 6429 35388
rect 6365 35328 6429 35332
rect 6445 35388 6509 35392
rect 6445 35332 6449 35388
rect 6449 35332 6505 35388
rect 6505 35332 6509 35388
rect 6445 35328 6509 35332
rect 6525 35388 6589 35392
rect 6525 35332 6529 35388
rect 6529 35332 6585 35388
rect 6585 35332 6589 35388
rect 6525 35328 6589 35332
rect 11618 35388 11682 35392
rect 11618 35332 11622 35388
rect 11622 35332 11678 35388
rect 11678 35332 11682 35388
rect 11618 35328 11682 35332
rect 11698 35388 11762 35392
rect 11698 35332 11702 35388
rect 11702 35332 11758 35388
rect 11758 35332 11762 35388
rect 11698 35328 11762 35332
rect 11778 35388 11842 35392
rect 11778 35332 11782 35388
rect 11782 35332 11838 35388
rect 11838 35332 11842 35388
rect 11778 35328 11842 35332
rect 11858 35388 11922 35392
rect 11858 35332 11862 35388
rect 11862 35332 11918 35388
rect 11918 35332 11922 35388
rect 11858 35328 11922 35332
rect 11468 35124 11532 35188
rect 3618 34844 3682 34848
rect 3618 34788 3622 34844
rect 3622 34788 3678 34844
rect 3678 34788 3682 34844
rect 3618 34784 3682 34788
rect 3698 34844 3762 34848
rect 3698 34788 3702 34844
rect 3702 34788 3758 34844
rect 3758 34788 3762 34844
rect 3698 34784 3762 34788
rect 3778 34844 3842 34848
rect 3778 34788 3782 34844
rect 3782 34788 3838 34844
rect 3838 34788 3842 34844
rect 3778 34784 3842 34788
rect 3858 34844 3922 34848
rect 3858 34788 3862 34844
rect 3862 34788 3918 34844
rect 3918 34788 3922 34844
rect 3858 34784 3922 34788
rect 8952 34844 9016 34848
rect 8952 34788 8956 34844
rect 8956 34788 9012 34844
rect 9012 34788 9016 34844
rect 8952 34784 9016 34788
rect 9032 34844 9096 34848
rect 9032 34788 9036 34844
rect 9036 34788 9092 34844
rect 9092 34788 9096 34844
rect 9032 34784 9096 34788
rect 9112 34844 9176 34848
rect 9112 34788 9116 34844
rect 9116 34788 9172 34844
rect 9172 34788 9176 34844
rect 9112 34784 9176 34788
rect 9192 34844 9256 34848
rect 9192 34788 9196 34844
rect 9196 34788 9252 34844
rect 9252 34788 9256 34844
rect 9192 34784 9256 34788
rect 14285 34844 14349 34848
rect 14285 34788 14289 34844
rect 14289 34788 14345 34844
rect 14345 34788 14349 34844
rect 14285 34784 14349 34788
rect 14365 34844 14429 34848
rect 14365 34788 14369 34844
rect 14369 34788 14425 34844
rect 14425 34788 14429 34844
rect 14365 34784 14429 34788
rect 14445 34844 14509 34848
rect 14445 34788 14449 34844
rect 14449 34788 14505 34844
rect 14505 34788 14509 34844
rect 14445 34784 14509 34788
rect 14525 34844 14589 34848
rect 14525 34788 14529 34844
rect 14529 34788 14585 34844
rect 14585 34788 14589 34844
rect 14525 34784 14589 34788
rect 6285 34300 6349 34304
rect 6285 34244 6289 34300
rect 6289 34244 6345 34300
rect 6345 34244 6349 34300
rect 6285 34240 6349 34244
rect 6365 34300 6429 34304
rect 6365 34244 6369 34300
rect 6369 34244 6425 34300
rect 6425 34244 6429 34300
rect 6365 34240 6429 34244
rect 6445 34300 6509 34304
rect 6445 34244 6449 34300
rect 6449 34244 6505 34300
rect 6505 34244 6509 34300
rect 6445 34240 6509 34244
rect 6525 34300 6589 34304
rect 6525 34244 6529 34300
rect 6529 34244 6585 34300
rect 6585 34244 6589 34300
rect 6525 34240 6589 34244
rect 11618 34300 11682 34304
rect 11618 34244 11622 34300
rect 11622 34244 11678 34300
rect 11678 34244 11682 34300
rect 11618 34240 11682 34244
rect 11698 34300 11762 34304
rect 11698 34244 11702 34300
rect 11702 34244 11758 34300
rect 11758 34244 11762 34300
rect 11698 34240 11762 34244
rect 11778 34300 11842 34304
rect 11778 34244 11782 34300
rect 11782 34244 11838 34300
rect 11838 34244 11842 34300
rect 11778 34240 11842 34244
rect 11858 34300 11922 34304
rect 11858 34244 11862 34300
rect 11862 34244 11918 34300
rect 11918 34244 11922 34300
rect 11858 34240 11922 34244
rect 3618 33756 3682 33760
rect 3618 33700 3622 33756
rect 3622 33700 3678 33756
rect 3678 33700 3682 33756
rect 3618 33696 3682 33700
rect 3698 33756 3762 33760
rect 3698 33700 3702 33756
rect 3702 33700 3758 33756
rect 3758 33700 3762 33756
rect 3698 33696 3762 33700
rect 3778 33756 3842 33760
rect 3778 33700 3782 33756
rect 3782 33700 3838 33756
rect 3838 33700 3842 33756
rect 3778 33696 3842 33700
rect 3858 33756 3922 33760
rect 3858 33700 3862 33756
rect 3862 33700 3918 33756
rect 3918 33700 3922 33756
rect 3858 33696 3922 33700
rect 8952 33756 9016 33760
rect 8952 33700 8956 33756
rect 8956 33700 9012 33756
rect 9012 33700 9016 33756
rect 8952 33696 9016 33700
rect 9032 33756 9096 33760
rect 9032 33700 9036 33756
rect 9036 33700 9092 33756
rect 9092 33700 9096 33756
rect 9032 33696 9096 33700
rect 9112 33756 9176 33760
rect 9112 33700 9116 33756
rect 9116 33700 9172 33756
rect 9172 33700 9176 33756
rect 9112 33696 9176 33700
rect 9192 33756 9256 33760
rect 9192 33700 9196 33756
rect 9196 33700 9252 33756
rect 9252 33700 9256 33756
rect 9192 33696 9256 33700
rect 14285 33756 14349 33760
rect 14285 33700 14289 33756
rect 14289 33700 14345 33756
rect 14345 33700 14349 33756
rect 14285 33696 14349 33700
rect 14365 33756 14429 33760
rect 14365 33700 14369 33756
rect 14369 33700 14425 33756
rect 14425 33700 14429 33756
rect 14365 33696 14429 33700
rect 14445 33756 14509 33760
rect 14445 33700 14449 33756
rect 14449 33700 14505 33756
rect 14505 33700 14509 33756
rect 14445 33696 14509 33700
rect 14525 33756 14589 33760
rect 14525 33700 14529 33756
rect 14529 33700 14585 33756
rect 14585 33700 14589 33756
rect 14525 33696 14589 33700
rect 6285 33212 6349 33216
rect 6285 33156 6289 33212
rect 6289 33156 6345 33212
rect 6345 33156 6349 33212
rect 6285 33152 6349 33156
rect 6365 33212 6429 33216
rect 6365 33156 6369 33212
rect 6369 33156 6425 33212
rect 6425 33156 6429 33212
rect 6365 33152 6429 33156
rect 6445 33212 6509 33216
rect 6445 33156 6449 33212
rect 6449 33156 6505 33212
rect 6505 33156 6509 33212
rect 6445 33152 6509 33156
rect 6525 33212 6589 33216
rect 6525 33156 6529 33212
rect 6529 33156 6585 33212
rect 6585 33156 6589 33212
rect 6525 33152 6589 33156
rect 11618 33212 11682 33216
rect 11618 33156 11622 33212
rect 11622 33156 11678 33212
rect 11678 33156 11682 33212
rect 11618 33152 11682 33156
rect 11698 33212 11762 33216
rect 11698 33156 11702 33212
rect 11702 33156 11758 33212
rect 11758 33156 11762 33212
rect 11698 33152 11762 33156
rect 11778 33212 11842 33216
rect 11778 33156 11782 33212
rect 11782 33156 11838 33212
rect 11838 33156 11842 33212
rect 11778 33152 11842 33156
rect 11858 33212 11922 33216
rect 11858 33156 11862 33212
rect 11862 33156 11918 33212
rect 11918 33156 11922 33212
rect 11858 33152 11922 33156
rect 3618 32668 3682 32672
rect 3618 32612 3622 32668
rect 3622 32612 3678 32668
rect 3678 32612 3682 32668
rect 3618 32608 3682 32612
rect 3698 32668 3762 32672
rect 3698 32612 3702 32668
rect 3702 32612 3758 32668
rect 3758 32612 3762 32668
rect 3698 32608 3762 32612
rect 3778 32668 3842 32672
rect 3778 32612 3782 32668
rect 3782 32612 3838 32668
rect 3838 32612 3842 32668
rect 3778 32608 3842 32612
rect 3858 32668 3922 32672
rect 3858 32612 3862 32668
rect 3862 32612 3918 32668
rect 3918 32612 3922 32668
rect 3858 32608 3922 32612
rect 8952 32668 9016 32672
rect 8952 32612 8956 32668
rect 8956 32612 9012 32668
rect 9012 32612 9016 32668
rect 8952 32608 9016 32612
rect 9032 32668 9096 32672
rect 9032 32612 9036 32668
rect 9036 32612 9092 32668
rect 9092 32612 9096 32668
rect 9032 32608 9096 32612
rect 9112 32668 9176 32672
rect 9112 32612 9116 32668
rect 9116 32612 9172 32668
rect 9172 32612 9176 32668
rect 9112 32608 9176 32612
rect 9192 32668 9256 32672
rect 9192 32612 9196 32668
rect 9196 32612 9252 32668
rect 9252 32612 9256 32668
rect 9192 32608 9256 32612
rect 14285 32668 14349 32672
rect 14285 32612 14289 32668
rect 14289 32612 14345 32668
rect 14345 32612 14349 32668
rect 14285 32608 14349 32612
rect 14365 32668 14429 32672
rect 14365 32612 14369 32668
rect 14369 32612 14425 32668
rect 14425 32612 14429 32668
rect 14365 32608 14429 32612
rect 14445 32668 14509 32672
rect 14445 32612 14449 32668
rect 14449 32612 14505 32668
rect 14505 32612 14509 32668
rect 14445 32608 14509 32612
rect 14525 32668 14589 32672
rect 14525 32612 14529 32668
rect 14529 32612 14585 32668
rect 14585 32612 14589 32668
rect 14525 32608 14589 32612
rect 6285 32124 6349 32128
rect 6285 32068 6289 32124
rect 6289 32068 6345 32124
rect 6345 32068 6349 32124
rect 6285 32064 6349 32068
rect 6365 32124 6429 32128
rect 6365 32068 6369 32124
rect 6369 32068 6425 32124
rect 6425 32068 6429 32124
rect 6365 32064 6429 32068
rect 6445 32124 6509 32128
rect 6445 32068 6449 32124
rect 6449 32068 6505 32124
rect 6505 32068 6509 32124
rect 6445 32064 6509 32068
rect 6525 32124 6589 32128
rect 6525 32068 6529 32124
rect 6529 32068 6585 32124
rect 6585 32068 6589 32124
rect 6525 32064 6589 32068
rect 11618 32124 11682 32128
rect 11618 32068 11622 32124
rect 11622 32068 11678 32124
rect 11678 32068 11682 32124
rect 11618 32064 11682 32068
rect 11698 32124 11762 32128
rect 11698 32068 11702 32124
rect 11702 32068 11758 32124
rect 11758 32068 11762 32124
rect 11698 32064 11762 32068
rect 11778 32124 11842 32128
rect 11778 32068 11782 32124
rect 11782 32068 11838 32124
rect 11838 32068 11842 32124
rect 11778 32064 11842 32068
rect 11858 32124 11922 32128
rect 11858 32068 11862 32124
rect 11862 32068 11918 32124
rect 11918 32068 11922 32124
rect 11858 32064 11922 32068
rect 3618 31580 3682 31584
rect 3618 31524 3622 31580
rect 3622 31524 3678 31580
rect 3678 31524 3682 31580
rect 3618 31520 3682 31524
rect 3698 31580 3762 31584
rect 3698 31524 3702 31580
rect 3702 31524 3758 31580
rect 3758 31524 3762 31580
rect 3698 31520 3762 31524
rect 3778 31580 3842 31584
rect 3778 31524 3782 31580
rect 3782 31524 3838 31580
rect 3838 31524 3842 31580
rect 3778 31520 3842 31524
rect 3858 31580 3922 31584
rect 3858 31524 3862 31580
rect 3862 31524 3918 31580
rect 3918 31524 3922 31580
rect 3858 31520 3922 31524
rect 8952 31580 9016 31584
rect 8952 31524 8956 31580
rect 8956 31524 9012 31580
rect 9012 31524 9016 31580
rect 8952 31520 9016 31524
rect 9032 31580 9096 31584
rect 9032 31524 9036 31580
rect 9036 31524 9092 31580
rect 9092 31524 9096 31580
rect 9032 31520 9096 31524
rect 9112 31580 9176 31584
rect 9112 31524 9116 31580
rect 9116 31524 9172 31580
rect 9172 31524 9176 31580
rect 9112 31520 9176 31524
rect 9192 31580 9256 31584
rect 9192 31524 9196 31580
rect 9196 31524 9252 31580
rect 9252 31524 9256 31580
rect 9192 31520 9256 31524
rect 14285 31580 14349 31584
rect 14285 31524 14289 31580
rect 14289 31524 14345 31580
rect 14345 31524 14349 31580
rect 14285 31520 14349 31524
rect 14365 31580 14429 31584
rect 14365 31524 14369 31580
rect 14369 31524 14425 31580
rect 14425 31524 14429 31580
rect 14365 31520 14429 31524
rect 14445 31580 14509 31584
rect 14445 31524 14449 31580
rect 14449 31524 14505 31580
rect 14505 31524 14509 31580
rect 14445 31520 14509 31524
rect 14525 31580 14589 31584
rect 14525 31524 14529 31580
rect 14529 31524 14585 31580
rect 14585 31524 14589 31580
rect 14525 31520 14589 31524
rect 9628 31452 9692 31516
rect 9628 31180 9692 31244
rect 6285 31036 6349 31040
rect 6285 30980 6289 31036
rect 6289 30980 6345 31036
rect 6345 30980 6349 31036
rect 6285 30976 6349 30980
rect 6365 31036 6429 31040
rect 6365 30980 6369 31036
rect 6369 30980 6425 31036
rect 6425 30980 6429 31036
rect 6365 30976 6429 30980
rect 6445 31036 6509 31040
rect 6445 30980 6449 31036
rect 6449 30980 6505 31036
rect 6505 30980 6509 31036
rect 6445 30976 6509 30980
rect 6525 31036 6589 31040
rect 6525 30980 6529 31036
rect 6529 30980 6585 31036
rect 6585 30980 6589 31036
rect 6525 30976 6589 30980
rect 11618 31036 11682 31040
rect 11618 30980 11622 31036
rect 11622 30980 11678 31036
rect 11678 30980 11682 31036
rect 11618 30976 11682 30980
rect 11698 31036 11762 31040
rect 11698 30980 11702 31036
rect 11702 30980 11758 31036
rect 11758 30980 11762 31036
rect 11698 30976 11762 30980
rect 11778 31036 11842 31040
rect 11778 30980 11782 31036
rect 11782 30980 11838 31036
rect 11838 30980 11842 31036
rect 11778 30976 11842 30980
rect 11858 31036 11922 31040
rect 11858 30980 11862 31036
rect 11862 30980 11918 31036
rect 11918 30980 11922 31036
rect 11858 30976 11922 30980
rect 3618 30492 3682 30496
rect 3618 30436 3622 30492
rect 3622 30436 3678 30492
rect 3678 30436 3682 30492
rect 3618 30432 3682 30436
rect 3698 30492 3762 30496
rect 3698 30436 3702 30492
rect 3702 30436 3758 30492
rect 3758 30436 3762 30492
rect 3698 30432 3762 30436
rect 3778 30492 3842 30496
rect 3778 30436 3782 30492
rect 3782 30436 3838 30492
rect 3838 30436 3842 30492
rect 3778 30432 3842 30436
rect 3858 30492 3922 30496
rect 3858 30436 3862 30492
rect 3862 30436 3918 30492
rect 3918 30436 3922 30492
rect 3858 30432 3922 30436
rect 8952 30492 9016 30496
rect 8952 30436 8956 30492
rect 8956 30436 9012 30492
rect 9012 30436 9016 30492
rect 8952 30432 9016 30436
rect 9032 30492 9096 30496
rect 9032 30436 9036 30492
rect 9036 30436 9092 30492
rect 9092 30436 9096 30492
rect 9032 30432 9096 30436
rect 9112 30492 9176 30496
rect 9112 30436 9116 30492
rect 9116 30436 9172 30492
rect 9172 30436 9176 30492
rect 9112 30432 9176 30436
rect 9192 30492 9256 30496
rect 9192 30436 9196 30492
rect 9196 30436 9252 30492
rect 9252 30436 9256 30492
rect 9192 30432 9256 30436
rect 14285 30492 14349 30496
rect 14285 30436 14289 30492
rect 14289 30436 14345 30492
rect 14345 30436 14349 30492
rect 14285 30432 14349 30436
rect 14365 30492 14429 30496
rect 14365 30436 14369 30492
rect 14369 30436 14425 30492
rect 14425 30436 14429 30492
rect 14365 30432 14429 30436
rect 14445 30492 14509 30496
rect 14445 30436 14449 30492
rect 14449 30436 14505 30492
rect 14505 30436 14509 30492
rect 14445 30432 14509 30436
rect 14525 30492 14589 30496
rect 14525 30436 14529 30492
rect 14529 30436 14585 30492
rect 14585 30436 14589 30492
rect 14525 30432 14589 30436
rect 6285 29948 6349 29952
rect 6285 29892 6289 29948
rect 6289 29892 6345 29948
rect 6345 29892 6349 29948
rect 6285 29888 6349 29892
rect 6365 29948 6429 29952
rect 6365 29892 6369 29948
rect 6369 29892 6425 29948
rect 6425 29892 6429 29948
rect 6365 29888 6429 29892
rect 6445 29948 6509 29952
rect 6445 29892 6449 29948
rect 6449 29892 6505 29948
rect 6505 29892 6509 29948
rect 6445 29888 6509 29892
rect 6525 29948 6589 29952
rect 6525 29892 6529 29948
rect 6529 29892 6585 29948
rect 6585 29892 6589 29948
rect 6525 29888 6589 29892
rect 11618 29948 11682 29952
rect 11618 29892 11622 29948
rect 11622 29892 11678 29948
rect 11678 29892 11682 29948
rect 11618 29888 11682 29892
rect 11698 29948 11762 29952
rect 11698 29892 11702 29948
rect 11702 29892 11758 29948
rect 11758 29892 11762 29948
rect 11698 29888 11762 29892
rect 11778 29948 11842 29952
rect 11778 29892 11782 29948
rect 11782 29892 11838 29948
rect 11838 29892 11842 29948
rect 11778 29888 11842 29892
rect 11858 29948 11922 29952
rect 11858 29892 11862 29948
rect 11862 29892 11918 29948
rect 11918 29892 11922 29948
rect 11858 29888 11922 29892
rect 11468 29548 11532 29612
rect 3618 29404 3682 29408
rect 3618 29348 3622 29404
rect 3622 29348 3678 29404
rect 3678 29348 3682 29404
rect 3618 29344 3682 29348
rect 3698 29404 3762 29408
rect 3698 29348 3702 29404
rect 3702 29348 3758 29404
rect 3758 29348 3762 29404
rect 3698 29344 3762 29348
rect 3778 29404 3842 29408
rect 3778 29348 3782 29404
rect 3782 29348 3838 29404
rect 3838 29348 3842 29404
rect 3778 29344 3842 29348
rect 3858 29404 3922 29408
rect 3858 29348 3862 29404
rect 3862 29348 3918 29404
rect 3918 29348 3922 29404
rect 3858 29344 3922 29348
rect 8952 29404 9016 29408
rect 8952 29348 8956 29404
rect 8956 29348 9012 29404
rect 9012 29348 9016 29404
rect 8952 29344 9016 29348
rect 9032 29404 9096 29408
rect 9032 29348 9036 29404
rect 9036 29348 9092 29404
rect 9092 29348 9096 29404
rect 9032 29344 9096 29348
rect 9112 29404 9176 29408
rect 9112 29348 9116 29404
rect 9116 29348 9172 29404
rect 9172 29348 9176 29404
rect 9112 29344 9176 29348
rect 9192 29404 9256 29408
rect 9192 29348 9196 29404
rect 9196 29348 9252 29404
rect 9252 29348 9256 29404
rect 9192 29344 9256 29348
rect 14285 29404 14349 29408
rect 14285 29348 14289 29404
rect 14289 29348 14345 29404
rect 14345 29348 14349 29404
rect 14285 29344 14349 29348
rect 14365 29404 14429 29408
rect 14365 29348 14369 29404
rect 14369 29348 14425 29404
rect 14425 29348 14429 29404
rect 14365 29344 14429 29348
rect 14445 29404 14509 29408
rect 14445 29348 14449 29404
rect 14449 29348 14505 29404
rect 14505 29348 14509 29404
rect 14445 29344 14509 29348
rect 14525 29404 14589 29408
rect 14525 29348 14529 29404
rect 14529 29348 14585 29404
rect 14585 29348 14589 29404
rect 14525 29344 14589 29348
rect 6285 28860 6349 28864
rect 6285 28804 6289 28860
rect 6289 28804 6345 28860
rect 6345 28804 6349 28860
rect 6285 28800 6349 28804
rect 6365 28860 6429 28864
rect 6365 28804 6369 28860
rect 6369 28804 6425 28860
rect 6425 28804 6429 28860
rect 6365 28800 6429 28804
rect 6445 28860 6509 28864
rect 6445 28804 6449 28860
rect 6449 28804 6505 28860
rect 6505 28804 6509 28860
rect 6445 28800 6509 28804
rect 6525 28860 6589 28864
rect 6525 28804 6529 28860
rect 6529 28804 6585 28860
rect 6585 28804 6589 28860
rect 6525 28800 6589 28804
rect 11618 28860 11682 28864
rect 11618 28804 11622 28860
rect 11622 28804 11678 28860
rect 11678 28804 11682 28860
rect 11618 28800 11682 28804
rect 11698 28860 11762 28864
rect 11698 28804 11702 28860
rect 11702 28804 11758 28860
rect 11758 28804 11762 28860
rect 11698 28800 11762 28804
rect 11778 28860 11842 28864
rect 11778 28804 11782 28860
rect 11782 28804 11838 28860
rect 11838 28804 11842 28860
rect 11778 28800 11842 28804
rect 11858 28860 11922 28864
rect 11858 28804 11862 28860
rect 11862 28804 11918 28860
rect 11918 28804 11922 28860
rect 11858 28800 11922 28804
rect 3618 28316 3682 28320
rect 3618 28260 3622 28316
rect 3622 28260 3678 28316
rect 3678 28260 3682 28316
rect 3618 28256 3682 28260
rect 3698 28316 3762 28320
rect 3698 28260 3702 28316
rect 3702 28260 3758 28316
rect 3758 28260 3762 28316
rect 3698 28256 3762 28260
rect 3778 28316 3842 28320
rect 3778 28260 3782 28316
rect 3782 28260 3838 28316
rect 3838 28260 3842 28316
rect 3778 28256 3842 28260
rect 3858 28316 3922 28320
rect 3858 28260 3862 28316
rect 3862 28260 3918 28316
rect 3918 28260 3922 28316
rect 3858 28256 3922 28260
rect 8952 28316 9016 28320
rect 8952 28260 8956 28316
rect 8956 28260 9012 28316
rect 9012 28260 9016 28316
rect 8952 28256 9016 28260
rect 9032 28316 9096 28320
rect 9032 28260 9036 28316
rect 9036 28260 9092 28316
rect 9092 28260 9096 28316
rect 9032 28256 9096 28260
rect 9112 28316 9176 28320
rect 9112 28260 9116 28316
rect 9116 28260 9172 28316
rect 9172 28260 9176 28316
rect 9112 28256 9176 28260
rect 9192 28316 9256 28320
rect 9192 28260 9196 28316
rect 9196 28260 9252 28316
rect 9252 28260 9256 28316
rect 9192 28256 9256 28260
rect 14285 28316 14349 28320
rect 14285 28260 14289 28316
rect 14289 28260 14345 28316
rect 14345 28260 14349 28316
rect 14285 28256 14349 28260
rect 14365 28316 14429 28320
rect 14365 28260 14369 28316
rect 14369 28260 14425 28316
rect 14425 28260 14429 28316
rect 14365 28256 14429 28260
rect 14445 28316 14509 28320
rect 14445 28260 14449 28316
rect 14449 28260 14505 28316
rect 14505 28260 14509 28316
rect 14445 28256 14509 28260
rect 14525 28316 14589 28320
rect 14525 28260 14529 28316
rect 14529 28260 14585 28316
rect 14585 28260 14589 28316
rect 14525 28256 14589 28260
rect 11468 28188 11532 28252
rect 6285 27772 6349 27776
rect 6285 27716 6289 27772
rect 6289 27716 6345 27772
rect 6345 27716 6349 27772
rect 6285 27712 6349 27716
rect 6365 27772 6429 27776
rect 6365 27716 6369 27772
rect 6369 27716 6425 27772
rect 6425 27716 6429 27772
rect 6365 27712 6429 27716
rect 6445 27772 6509 27776
rect 6445 27716 6449 27772
rect 6449 27716 6505 27772
rect 6505 27716 6509 27772
rect 6445 27712 6509 27716
rect 6525 27772 6589 27776
rect 6525 27716 6529 27772
rect 6529 27716 6585 27772
rect 6585 27716 6589 27772
rect 6525 27712 6589 27716
rect 11618 27772 11682 27776
rect 11618 27716 11622 27772
rect 11622 27716 11678 27772
rect 11678 27716 11682 27772
rect 11618 27712 11682 27716
rect 11698 27772 11762 27776
rect 11698 27716 11702 27772
rect 11702 27716 11758 27772
rect 11758 27716 11762 27772
rect 11698 27712 11762 27716
rect 11778 27772 11842 27776
rect 11778 27716 11782 27772
rect 11782 27716 11838 27772
rect 11838 27716 11842 27772
rect 11778 27712 11842 27716
rect 11858 27772 11922 27776
rect 11858 27716 11862 27772
rect 11862 27716 11918 27772
rect 11918 27716 11922 27772
rect 11858 27712 11922 27716
rect 3618 27228 3682 27232
rect 3618 27172 3622 27228
rect 3622 27172 3678 27228
rect 3678 27172 3682 27228
rect 3618 27168 3682 27172
rect 3698 27228 3762 27232
rect 3698 27172 3702 27228
rect 3702 27172 3758 27228
rect 3758 27172 3762 27228
rect 3698 27168 3762 27172
rect 3778 27228 3842 27232
rect 3778 27172 3782 27228
rect 3782 27172 3838 27228
rect 3838 27172 3842 27228
rect 3778 27168 3842 27172
rect 3858 27228 3922 27232
rect 3858 27172 3862 27228
rect 3862 27172 3918 27228
rect 3918 27172 3922 27228
rect 3858 27168 3922 27172
rect 8952 27228 9016 27232
rect 8952 27172 8956 27228
rect 8956 27172 9012 27228
rect 9012 27172 9016 27228
rect 8952 27168 9016 27172
rect 9032 27228 9096 27232
rect 9032 27172 9036 27228
rect 9036 27172 9092 27228
rect 9092 27172 9096 27228
rect 9032 27168 9096 27172
rect 9112 27228 9176 27232
rect 9112 27172 9116 27228
rect 9116 27172 9172 27228
rect 9172 27172 9176 27228
rect 9112 27168 9176 27172
rect 9192 27228 9256 27232
rect 9192 27172 9196 27228
rect 9196 27172 9252 27228
rect 9252 27172 9256 27228
rect 9192 27168 9256 27172
rect 14285 27228 14349 27232
rect 14285 27172 14289 27228
rect 14289 27172 14345 27228
rect 14345 27172 14349 27228
rect 14285 27168 14349 27172
rect 14365 27228 14429 27232
rect 14365 27172 14369 27228
rect 14369 27172 14425 27228
rect 14425 27172 14429 27228
rect 14365 27168 14429 27172
rect 14445 27228 14509 27232
rect 14445 27172 14449 27228
rect 14449 27172 14505 27228
rect 14505 27172 14509 27228
rect 14445 27168 14509 27172
rect 14525 27228 14589 27232
rect 14525 27172 14529 27228
rect 14529 27172 14585 27228
rect 14585 27172 14589 27228
rect 14525 27168 14589 27172
rect 6285 26684 6349 26688
rect 6285 26628 6289 26684
rect 6289 26628 6345 26684
rect 6345 26628 6349 26684
rect 6285 26624 6349 26628
rect 6365 26684 6429 26688
rect 6365 26628 6369 26684
rect 6369 26628 6425 26684
rect 6425 26628 6429 26684
rect 6365 26624 6429 26628
rect 6445 26684 6509 26688
rect 6445 26628 6449 26684
rect 6449 26628 6505 26684
rect 6505 26628 6509 26684
rect 6445 26624 6509 26628
rect 6525 26684 6589 26688
rect 6525 26628 6529 26684
rect 6529 26628 6585 26684
rect 6585 26628 6589 26684
rect 6525 26624 6589 26628
rect 11618 26684 11682 26688
rect 11618 26628 11622 26684
rect 11622 26628 11678 26684
rect 11678 26628 11682 26684
rect 11618 26624 11682 26628
rect 11698 26684 11762 26688
rect 11698 26628 11702 26684
rect 11702 26628 11758 26684
rect 11758 26628 11762 26684
rect 11698 26624 11762 26628
rect 11778 26684 11842 26688
rect 11778 26628 11782 26684
rect 11782 26628 11838 26684
rect 11838 26628 11842 26684
rect 11778 26624 11842 26628
rect 11858 26684 11922 26688
rect 11858 26628 11862 26684
rect 11862 26628 11918 26684
rect 11918 26628 11922 26684
rect 11858 26624 11922 26628
rect 3618 26140 3682 26144
rect 3618 26084 3622 26140
rect 3622 26084 3678 26140
rect 3678 26084 3682 26140
rect 3618 26080 3682 26084
rect 3698 26140 3762 26144
rect 3698 26084 3702 26140
rect 3702 26084 3758 26140
rect 3758 26084 3762 26140
rect 3698 26080 3762 26084
rect 3778 26140 3842 26144
rect 3778 26084 3782 26140
rect 3782 26084 3838 26140
rect 3838 26084 3842 26140
rect 3778 26080 3842 26084
rect 3858 26140 3922 26144
rect 3858 26084 3862 26140
rect 3862 26084 3918 26140
rect 3918 26084 3922 26140
rect 3858 26080 3922 26084
rect 8952 26140 9016 26144
rect 8952 26084 8956 26140
rect 8956 26084 9012 26140
rect 9012 26084 9016 26140
rect 8952 26080 9016 26084
rect 9032 26140 9096 26144
rect 9032 26084 9036 26140
rect 9036 26084 9092 26140
rect 9092 26084 9096 26140
rect 9032 26080 9096 26084
rect 9112 26140 9176 26144
rect 9112 26084 9116 26140
rect 9116 26084 9172 26140
rect 9172 26084 9176 26140
rect 9112 26080 9176 26084
rect 9192 26140 9256 26144
rect 9192 26084 9196 26140
rect 9196 26084 9252 26140
rect 9252 26084 9256 26140
rect 9192 26080 9256 26084
rect 14285 26140 14349 26144
rect 14285 26084 14289 26140
rect 14289 26084 14345 26140
rect 14345 26084 14349 26140
rect 14285 26080 14349 26084
rect 14365 26140 14429 26144
rect 14365 26084 14369 26140
rect 14369 26084 14425 26140
rect 14425 26084 14429 26140
rect 14365 26080 14429 26084
rect 14445 26140 14509 26144
rect 14445 26084 14449 26140
rect 14449 26084 14505 26140
rect 14505 26084 14509 26140
rect 14445 26080 14509 26084
rect 14525 26140 14589 26144
rect 14525 26084 14529 26140
rect 14529 26084 14585 26140
rect 14585 26084 14589 26140
rect 14525 26080 14589 26084
rect 6285 25596 6349 25600
rect 6285 25540 6289 25596
rect 6289 25540 6345 25596
rect 6345 25540 6349 25596
rect 6285 25536 6349 25540
rect 6365 25596 6429 25600
rect 6365 25540 6369 25596
rect 6369 25540 6425 25596
rect 6425 25540 6429 25596
rect 6365 25536 6429 25540
rect 6445 25596 6509 25600
rect 6445 25540 6449 25596
rect 6449 25540 6505 25596
rect 6505 25540 6509 25596
rect 6445 25536 6509 25540
rect 6525 25596 6589 25600
rect 6525 25540 6529 25596
rect 6529 25540 6585 25596
rect 6585 25540 6589 25596
rect 6525 25536 6589 25540
rect 11618 25596 11682 25600
rect 11618 25540 11622 25596
rect 11622 25540 11678 25596
rect 11678 25540 11682 25596
rect 11618 25536 11682 25540
rect 11698 25596 11762 25600
rect 11698 25540 11702 25596
rect 11702 25540 11758 25596
rect 11758 25540 11762 25596
rect 11698 25536 11762 25540
rect 11778 25596 11842 25600
rect 11778 25540 11782 25596
rect 11782 25540 11838 25596
rect 11838 25540 11842 25596
rect 11778 25536 11842 25540
rect 11858 25596 11922 25600
rect 11858 25540 11862 25596
rect 11862 25540 11918 25596
rect 11918 25540 11922 25596
rect 11858 25536 11922 25540
rect 3618 25052 3682 25056
rect 3618 24996 3622 25052
rect 3622 24996 3678 25052
rect 3678 24996 3682 25052
rect 3618 24992 3682 24996
rect 3698 25052 3762 25056
rect 3698 24996 3702 25052
rect 3702 24996 3758 25052
rect 3758 24996 3762 25052
rect 3698 24992 3762 24996
rect 3778 25052 3842 25056
rect 3778 24996 3782 25052
rect 3782 24996 3838 25052
rect 3838 24996 3842 25052
rect 3778 24992 3842 24996
rect 3858 25052 3922 25056
rect 3858 24996 3862 25052
rect 3862 24996 3918 25052
rect 3918 24996 3922 25052
rect 3858 24992 3922 24996
rect 8952 25052 9016 25056
rect 8952 24996 8956 25052
rect 8956 24996 9012 25052
rect 9012 24996 9016 25052
rect 8952 24992 9016 24996
rect 9032 25052 9096 25056
rect 9032 24996 9036 25052
rect 9036 24996 9092 25052
rect 9092 24996 9096 25052
rect 9032 24992 9096 24996
rect 9112 25052 9176 25056
rect 9112 24996 9116 25052
rect 9116 24996 9172 25052
rect 9172 24996 9176 25052
rect 9112 24992 9176 24996
rect 9192 25052 9256 25056
rect 9192 24996 9196 25052
rect 9196 24996 9252 25052
rect 9252 24996 9256 25052
rect 9192 24992 9256 24996
rect 14285 25052 14349 25056
rect 14285 24996 14289 25052
rect 14289 24996 14345 25052
rect 14345 24996 14349 25052
rect 14285 24992 14349 24996
rect 14365 25052 14429 25056
rect 14365 24996 14369 25052
rect 14369 24996 14425 25052
rect 14425 24996 14429 25052
rect 14365 24992 14429 24996
rect 14445 25052 14509 25056
rect 14445 24996 14449 25052
rect 14449 24996 14505 25052
rect 14505 24996 14509 25052
rect 14445 24992 14509 24996
rect 14525 25052 14589 25056
rect 14525 24996 14529 25052
rect 14529 24996 14585 25052
rect 14585 24996 14589 25052
rect 14525 24992 14589 24996
rect 6285 24508 6349 24512
rect 6285 24452 6289 24508
rect 6289 24452 6345 24508
rect 6345 24452 6349 24508
rect 6285 24448 6349 24452
rect 6365 24508 6429 24512
rect 6365 24452 6369 24508
rect 6369 24452 6425 24508
rect 6425 24452 6429 24508
rect 6365 24448 6429 24452
rect 6445 24508 6509 24512
rect 6445 24452 6449 24508
rect 6449 24452 6505 24508
rect 6505 24452 6509 24508
rect 6445 24448 6509 24452
rect 6525 24508 6589 24512
rect 6525 24452 6529 24508
rect 6529 24452 6585 24508
rect 6585 24452 6589 24508
rect 6525 24448 6589 24452
rect 11618 24508 11682 24512
rect 11618 24452 11622 24508
rect 11622 24452 11678 24508
rect 11678 24452 11682 24508
rect 11618 24448 11682 24452
rect 11698 24508 11762 24512
rect 11698 24452 11702 24508
rect 11702 24452 11758 24508
rect 11758 24452 11762 24508
rect 11698 24448 11762 24452
rect 11778 24508 11842 24512
rect 11778 24452 11782 24508
rect 11782 24452 11838 24508
rect 11838 24452 11842 24508
rect 11778 24448 11842 24452
rect 11858 24508 11922 24512
rect 11858 24452 11862 24508
rect 11862 24452 11918 24508
rect 11918 24452 11922 24508
rect 11858 24448 11922 24452
rect 3618 23964 3682 23968
rect 3618 23908 3622 23964
rect 3622 23908 3678 23964
rect 3678 23908 3682 23964
rect 3618 23904 3682 23908
rect 3698 23964 3762 23968
rect 3698 23908 3702 23964
rect 3702 23908 3758 23964
rect 3758 23908 3762 23964
rect 3698 23904 3762 23908
rect 3778 23964 3842 23968
rect 3778 23908 3782 23964
rect 3782 23908 3838 23964
rect 3838 23908 3842 23964
rect 3778 23904 3842 23908
rect 3858 23964 3922 23968
rect 3858 23908 3862 23964
rect 3862 23908 3918 23964
rect 3918 23908 3922 23964
rect 3858 23904 3922 23908
rect 8952 23964 9016 23968
rect 8952 23908 8956 23964
rect 8956 23908 9012 23964
rect 9012 23908 9016 23964
rect 8952 23904 9016 23908
rect 9032 23964 9096 23968
rect 9032 23908 9036 23964
rect 9036 23908 9092 23964
rect 9092 23908 9096 23964
rect 9032 23904 9096 23908
rect 9112 23964 9176 23968
rect 9112 23908 9116 23964
rect 9116 23908 9172 23964
rect 9172 23908 9176 23964
rect 9112 23904 9176 23908
rect 9192 23964 9256 23968
rect 9192 23908 9196 23964
rect 9196 23908 9252 23964
rect 9252 23908 9256 23964
rect 9192 23904 9256 23908
rect 14285 23964 14349 23968
rect 14285 23908 14289 23964
rect 14289 23908 14345 23964
rect 14345 23908 14349 23964
rect 14285 23904 14349 23908
rect 14365 23964 14429 23968
rect 14365 23908 14369 23964
rect 14369 23908 14425 23964
rect 14425 23908 14429 23964
rect 14365 23904 14429 23908
rect 14445 23964 14509 23968
rect 14445 23908 14449 23964
rect 14449 23908 14505 23964
rect 14505 23908 14509 23964
rect 14445 23904 14509 23908
rect 14525 23964 14589 23968
rect 14525 23908 14529 23964
rect 14529 23908 14585 23964
rect 14585 23908 14589 23964
rect 14525 23904 14589 23908
rect 6285 23420 6349 23424
rect 6285 23364 6289 23420
rect 6289 23364 6345 23420
rect 6345 23364 6349 23420
rect 6285 23360 6349 23364
rect 6365 23420 6429 23424
rect 6365 23364 6369 23420
rect 6369 23364 6425 23420
rect 6425 23364 6429 23420
rect 6365 23360 6429 23364
rect 6445 23420 6509 23424
rect 6445 23364 6449 23420
rect 6449 23364 6505 23420
rect 6505 23364 6509 23420
rect 6445 23360 6509 23364
rect 6525 23420 6589 23424
rect 6525 23364 6529 23420
rect 6529 23364 6585 23420
rect 6585 23364 6589 23420
rect 6525 23360 6589 23364
rect 11618 23420 11682 23424
rect 11618 23364 11622 23420
rect 11622 23364 11678 23420
rect 11678 23364 11682 23420
rect 11618 23360 11682 23364
rect 11698 23420 11762 23424
rect 11698 23364 11702 23420
rect 11702 23364 11758 23420
rect 11758 23364 11762 23420
rect 11698 23360 11762 23364
rect 11778 23420 11842 23424
rect 11778 23364 11782 23420
rect 11782 23364 11838 23420
rect 11838 23364 11842 23420
rect 11778 23360 11842 23364
rect 11858 23420 11922 23424
rect 11858 23364 11862 23420
rect 11862 23364 11918 23420
rect 11918 23364 11922 23420
rect 11858 23360 11922 23364
rect 3618 22876 3682 22880
rect 3618 22820 3622 22876
rect 3622 22820 3678 22876
rect 3678 22820 3682 22876
rect 3618 22816 3682 22820
rect 3698 22876 3762 22880
rect 3698 22820 3702 22876
rect 3702 22820 3758 22876
rect 3758 22820 3762 22876
rect 3698 22816 3762 22820
rect 3778 22876 3842 22880
rect 3778 22820 3782 22876
rect 3782 22820 3838 22876
rect 3838 22820 3842 22876
rect 3778 22816 3842 22820
rect 3858 22876 3922 22880
rect 3858 22820 3862 22876
rect 3862 22820 3918 22876
rect 3918 22820 3922 22876
rect 3858 22816 3922 22820
rect 8952 22876 9016 22880
rect 8952 22820 8956 22876
rect 8956 22820 9012 22876
rect 9012 22820 9016 22876
rect 8952 22816 9016 22820
rect 9032 22876 9096 22880
rect 9032 22820 9036 22876
rect 9036 22820 9092 22876
rect 9092 22820 9096 22876
rect 9032 22816 9096 22820
rect 9112 22876 9176 22880
rect 9112 22820 9116 22876
rect 9116 22820 9172 22876
rect 9172 22820 9176 22876
rect 9112 22816 9176 22820
rect 9192 22876 9256 22880
rect 9192 22820 9196 22876
rect 9196 22820 9252 22876
rect 9252 22820 9256 22876
rect 9192 22816 9256 22820
rect 14285 22876 14349 22880
rect 14285 22820 14289 22876
rect 14289 22820 14345 22876
rect 14345 22820 14349 22876
rect 14285 22816 14349 22820
rect 14365 22876 14429 22880
rect 14365 22820 14369 22876
rect 14369 22820 14425 22876
rect 14425 22820 14429 22876
rect 14365 22816 14429 22820
rect 14445 22876 14509 22880
rect 14445 22820 14449 22876
rect 14449 22820 14505 22876
rect 14505 22820 14509 22876
rect 14445 22816 14509 22820
rect 14525 22876 14589 22880
rect 14525 22820 14529 22876
rect 14529 22820 14585 22876
rect 14585 22820 14589 22876
rect 14525 22816 14589 22820
rect 6285 22332 6349 22336
rect 6285 22276 6289 22332
rect 6289 22276 6345 22332
rect 6345 22276 6349 22332
rect 6285 22272 6349 22276
rect 6365 22332 6429 22336
rect 6365 22276 6369 22332
rect 6369 22276 6425 22332
rect 6425 22276 6429 22332
rect 6365 22272 6429 22276
rect 6445 22332 6509 22336
rect 6445 22276 6449 22332
rect 6449 22276 6505 22332
rect 6505 22276 6509 22332
rect 6445 22272 6509 22276
rect 6525 22332 6589 22336
rect 6525 22276 6529 22332
rect 6529 22276 6585 22332
rect 6585 22276 6589 22332
rect 6525 22272 6589 22276
rect 11618 22332 11682 22336
rect 11618 22276 11622 22332
rect 11622 22276 11678 22332
rect 11678 22276 11682 22332
rect 11618 22272 11682 22276
rect 11698 22332 11762 22336
rect 11698 22276 11702 22332
rect 11702 22276 11758 22332
rect 11758 22276 11762 22332
rect 11698 22272 11762 22276
rect 11778 22332 11842 22336
rect 11778 22276 11782 22332
rect 11782 22276 11838 22332
rect 11838 22276 11842 22332
rect 11778 22272 11842 22276
rect 11858 22332 11922 22336
rect 11858 22276 11862 22332
rect 11862 22276 11918 22332
rect 11918 22276 11922 22332
rect 11858 22272 11922 22276
rect 3618 21788 3682 21792
rect 3618 21732 3622 21788
rect 3622 21732 3678 21788
rect 3678 21732 3682 21788
rect 3618 21728 3682 21732
rect 3698 21788 3762 21792
rect 3698 21732 3702 21788
rect 3702 21732 3758 21788
rect 3758 21732 3762 21788
rect 3698 21728 3762 21732
rect 3778 21788 3842 21792
rect 3778 21732 3782 21788
rect 3782 21732 3838 21788
rect 3838 21732 3842 21788
rect 3778 21728 3842 21732
rect 3858 21788 3922 21792
rect 3858 21732 3862 21788
rect 3862 21732 3918 21788
rect 3918 21732 3922 21788
rect 3858 21728 3922 21732
rect 8952 21788 9016 21792
rect 8952 21732 8956 21788
rect 8956 21732 9012 21788
rect 9012 21732 9016 21788
rect 8952 21728 9016 21732
rect 9032 21788 9096 21792
rect 9032 21732 9036 21788
rect 9036 21732 9092 21788
rect 9092 21732 9096 21788
rect 9032 21728 9096 21732
rect 9112 21788 9176 21792
rect 9112 21732 9116 21788
rect 9116 21732 9172 21788
rect 9172 21732 9176 21788
rect 9112 21728 9176 21732
rect 9192 21788 9256 21792
rect 9192 21732 9196 21788
rect 9196 21732 9252 21788
rect 9252 21732 9256 21788
rect 9192 21728 9256 21732
rect 14285 21788 14349 21792
rect 14285 21732 14289 21788
rect 14289 21732 14345 21788
rect 14345 21732 14349 21788
rect 14285 21728 14349 21732
rect 14365 21788 14429 21792
rect 14365 21732 14369 21788
rect 14369 21732 14425 21788
rect 14425 21732 14429 21788
rect 14365 21728 14429 21732
rect 14445 21788 14509 21792
rect 14445 21732 14449 21788
rect 14449 21732 14505 21788
rect 14505 21732 14509 21788
rect 14445 21728 14509 21732
rect 14525 21788 14589 21792
rect 14525 21732 14529 21788
rect 14529 21732 14585 21788
rect 14585 21732 14589 21788
rect 14525 21728 14589 21732
rect 6285 21244 6349 21248
rect 6285 21188 6289 21244
rect 6289 21188 6345 21244
rect 6345 21188 6349 21244
rect 6285 21184 6349 21188
rect 6365 21244 6429 21248
rect 6365 21188 6369 21244
rect 6369 21188 6425 21244
rect 6425 21188 6429 21244
rect 6365 21184 6429 21188
rect 6445 21244 6509 21248
rect 6445 21188 6449 21244
rect 6449 21188 6505 21244
rect 6505 21188 6509 21244
rect 6445 21184 6509 21188
rect 6525 21244 6589 21248
rect 6525 21188 6529 21244
rect 6529 21188 6585 21244
rect 6585 21188 6589 21244
rect 6525 21184 6589 21188
rect 11618 21244 11682 21248
rect 11618 21188 11622 21244
rect 11622 21188 11678 21244
rect 11678 21188 11682 21244
rect 11618 21184 11682 21188
rect 11698 21244 11762 21248
rect 11698 21188 11702 21244
rect 11702 21188 11758 21244
rect 11758 21188 11762 21244
rect 11698 21184 11762 21188
rect 11778 21244 11842 21248
rect 11778 21188 11782 21244
rect 11782 21188 11838 21244
rect 11838 21188 11842 21244
rect 11778 21184 11842 21188
rect 11858 21244 11922 21248
rect 11858 21188 11862 21244
rect 11862 21188 11918 21244
rect 11918 21188 11922 21244
rect 11858 21184 11922 21188
rect 3618 20700 3682 20704
rect 3618 20644 3622 20700
rect 3622 20644 3678 20700
rect 3678 20644 3682 20700
rect 3618 20640 3682 20644
rect 3698 20700 3762 20704
rect 3698 20644 3702 20700
rect 3702 20644 3758 20700
rect 3758 20644 3762 20700
rect 3698 20640 3762 20644
rect 3778 20700 3842 20704
rect 3778 20644 3782 20700
rect 3782 20644 3838 20700
rect 3838 20644 3842 20700
rect 3778 20640 3842 20644
rect 3858 20700 3922 20704
rect 3858 20644 3862 20700
rect 3862 20644 3918 20700
rect 3918 20644 3922 20700
rect 3858 20640 3922 20644
rect 8952 20700 9016 20704
rect 8952 20644 8956 20700
rect 8956 20644 9012 20700
rect 9012 20644 9016 20700
rect 8952 20640 9016 20644
rect 9032 20700 9096 20704
rect 9032 20644 9036 20700
rect 9036 20644 9092 20700
rect 9092 20644 9096 20700
rect 9032 20640 9096 20644
rect 9112 20700 9176 20704
rect 9112 20644 9116 20700
rect 9116 20644 9172 20700
rect 9172 20644 9176 20700
rect 9112 20640 9176 20644
rect 9192 20700 9256 20704
rect 9192 20644 9196 20700
rect 9196 20644 9252 20700
rect 9252 20644 9256 20700
rect 9192 20640 9256 20644
rect 14285 20700 14349 20704
rect 14285 20644 14289 20700
rect 14289 20644 14345 20700
rect 14345 20644 14349 20700
rect 14285 20640 14349 20644
rect 14365 20700 14429 20704
rect 14365 20644 14369 20700
rect 14369 20644 14425 20700
rect 14425 20644 14429 20700
rect 14365 20640 14429 20644
rect 14445 20700 14509 20704
rect 14445 20644 14449 20700
rect 14449 20644 14505 20700
rect 14505 20644 14509 20700
rect 14445 20640 14509 20644
rect 14525 20700 14589 20704
rect 14525 20644 14529 20700
rect 14529 20644 14585 20700
rect 14585 20644 14589 20700
rect 14525 20640 14589 20644
rect 6285 20156 6349 20160
rect 6285 20100 6289 20156
rect 6289 20100 6345 20156
rect 6345 20100 6349 20156
rect 6285 20096 6349 20100
rect 6365 20156 6429 20160
rect 6365 20100 6369 20156
rect 6369 20100 6425 20156
rect 6425 20100 6429 20156
rect 6365 20096 6429 20100
rect 6445 20156 6509 20160
rect 6445 20100 6449 20156
rect 6449 20100 6505 20156
rect 6505 20100 6509 20156
rect 6445 20096 6509 20100
rect 6525 20156 6589 20160
rect 6525 20100 6529 20156
rect 6529 20100 6585 20156
rect 6585 20100 6589 20156
rect 6525 20096 6589 20100
rect 11618 20156 11682 20160
rect 11618 20100 11622 20156
rect 11622 20100 11678 20156
rect 11678 20100 11682 20156
rect 11618 20096 11682 20100
rect 11698 20156 11762 20160
rect 11698 20100 11702 20156
rect 11702 20100 11758 20156
rect 11758 20100 11762 20156
rect 11698 20096 11762 20100
rect 11778 20156 11842 20160
rect 11778 20100 11782 20156
rect 11782 20100 11838 20156
rect 11838 20100 11842 20156
rect 11778 20096 11842 20100
rect 11858 20156 11922 20160
rect 11858 20100 11862 20156
rect 11862 20100 11918 20156
rect 11918 20100 11922 20156
rect 11858 20096 11922 20100
rect 11468 19756 11532 19820
rect 3618 19612 3682 19616
rect 3618 19556 3622 19612
rect 3622 19556 3678 19612
rect 3678 19556 3682 19612
rect 3618 19552 3682 19556
rect 3698 19612 3762 19616
rect 3698 19556 3702 19612
rect 3702 19556 3758 19612
rect 3758 19556 3762 19612
rect 3698 19552 3762 19556
rect 3778 19612 3842 19616
rect 3778 19556 3782 19612
rect 3782 19556 3838 19612
rect 3838 19556 3842 19612
rect 3778 19552 3842 19556
rect 3858 19612 3922 19616
rect 3858 19556 3862 19612
rect 3862 19556 3918 19612
rect 3918 19556 3922 19612
rect 3858 19552 3922 19556
rect 8952 19612 9016 19616
rect 8952 19556 8956 19612
rect 8956 19556 9012 19612
rect 9012 19556 9016 19612
rect 8952 19552 9016 19556
rect 9032 19612 9096 19616
rect 9032 19556 9036 19612
rect 9036 19556 9092 19612
rect 9092 19556 9096 19612
rect 9032 19552 9096 19556
rect 9112 19612 9176 19616
rect 9112 19556 9116 19612
rect 9116 19556 9172 19612
rect 9172 19556 9176 19612
rect 9112 19552 9176 19556
rect 9192 19612 9256 19616
rect 9192 19556 9196 19612
rect 9196 19556 9252 19612
rect 9252 19556 9256 19612
rect 9192 19552 9256 19556
rect 14285 19612 14349 19616
rect 14285 19556 14289 19612
rect 14289 19556 14345 19612
rect 14345 19556 14349 19612
rect 14285 19552 14349 19556
rect 14365 19612 14429 19616
rect 14365 19556 14369 19612
rect 14369 19556 14425 19612
rect 14425 19556 14429 19612
rect 14365 19552 14429 19556
rect 14445 19612 14509 19616
rect 14445 19556 14449 19612
rect 14449 19556 14505 19612
rect 14505 19556 14509 19612
rect 14445 19552 14509 19556
rect 14525 19612 14589 19616
rect 14525 19556 14529 19612
rect 14529 19556 14585 19612
rect 14585 19556 14589 19612
rect 14525 19552 14589 19556
rect 6285 19068 6349 19072
rect 6285 19012 6289 19068
rect 6289 19012 6345 19068
rect 6345 19012 6349 19068
rect 6285 19008 6349 19012
rect 6365 19068 6429 19072
rect 6365 19012 6369 19068
rect 6369 19012 6425 19068
rect 6425 19012 6429 19068
rect 6365 19008 6429 19012
rect 6445 19068 6509 19072
rect 6445 19012 6449 19068
rect 6449 19012 6505 19068
rect 6505 19012 6509 19068
rect 6445 19008 6509 19012
rect 6525 19068 6589 19072
rect 6525 19012 6529 19068
rect 6529 19012 6585 19068
rect 6585 19012 6589 19068
rect 6525 19008 6589 19012
rect 11618 19068 11682 19072
rect 11618 19012 11622 19068
rect 11622 19012 11678 19068
rect 11678 19012 11682 19068
rect 11618 19008 11682 19012
rect 11698 19068 11762 19072
rect 11698 19012 11702 19068
rect 11702 19012 11758 19068
rect 11758 19012 11762 19068
rect 11698 19008 11762 19012
rect 11778 19068 11842 19072
rect 11778 19012 11782 19068
rect 11782 19012 11838 19068
rect 11838 19012 11842 19068
rect 11778 19008 11842 19012
rect 11858 19068 11922 19072
rect 11858 19012 11862 19068
rect 11862 19012 11918 19068
rect 11918 19012 11922 19068
rect 11858 19008 11922 19012
rect 3618 18524 3682 18528
rect 3618 18468 3622 18524
rect 3622 18468 3678 18524
rect 3678 18468 3682 18524
rect 3618 18464 3682 18468
rect 3698 18524 3762 18528
rect 3698 18468 3702 18524
rect 3702 18468 3758 18524
rect 3758 18468 3762 18524
rect 3698 18464 3762 18468
rect 3778 18524 3842 18528
rect 3778 18468 3782 18524
rect 3782 18468 3838 18524
rect 3838 18468 3842 18524
rect 3778 18464 3842 18468
rect 3858 18524 3922 18528
rect 3858 18468 3862 18524
rect 3862 18468 3918 18524
rect 3918 18468 3922 18524
rect 3858 18464 3922 18468
rect 8952 18524 9016 18528
rect 8952 18468 8956 18524
rect 8956 18468 9012 18524
rect 9012 18468 9016 18524
rect 8952 18464 9016 18468
rect 9032 18524 9096 18528
rect 9032 18468 9036 18524
rect 9036 18468 9092 18524
rect 9092 18468 9096 18524
rect 9032 18464 9096 18468
rect 9112 18524 9176 18528
rect 9112 18468 9116 18524
rect 9116 18468 9172 18524
rect 9172 18468 9176 18524
rect 9112 18464 9176 18468
rect 9192 18524 9256 18528
rect 9192 18468 9196 18524
rect 9196 18468 9252 18524
rect 9252 18468 9256 18524
rect 9192 18464 9256 18468
rect 14285 18524 14349 18528
rect 14285 18468 14289 18524
rect 14289 18468 14345 18524
rect 14345 18468 14349 18524
rect 14285 18464 14349 18468
rect 14365 18524 14429 18528
rect 14365 18468 14369 18524
rect 14369 18468 14425 18524
rect 14425 18468 14429 18524
rect 14365 18464 14429 18468
rect 14445 18524 14509 18528
rect 14445 18468 14449 18524
rect 14449 18468 14505 18524
rect 14505 18468 14509 18524
rect 14445 18464 14509 18468
rect 14525 18524 14589 18528
rect 14525 18468 14529 18524
rect 14529 18468 14585 18524
rect 14585 18468 14589 18524
rect 14525 18464 14589 18468
rect 6285 17980 6349 17984
rect 6285 17924 6289 17980
rect 6289 17924 6345 17980
rect 6345 17924 6349 17980
rect 6285 17920 6349 17924
rect 6365 17980 6429 17984
rect 6365 17924 6369 17980
rect 6369 17924 6425 17980
rect 6425 17924 6429 17980
rect 6365 17920 6429 17924
rect 6445 17980 6509 17984
rect 6445 17924 6449 17980
rect 6449 17924 6505 17980
rect 6505 17924 6509 17980
rect 6445 17920 6509 17924
rect 6525 17980 6589 17984
rect 6525 17924 6529 17980
rect 6529 17924 6585 17980
rect 6585 17924 6589 17980
rect 6525 17920 6589 17924
rect 11618 17980 11682 17984
rect 11618 17924 11622 17980
rect 11622 17924 11678 17980
rect 11678 17924 11682 17980
rect 11618 17920 11682 17924
rect 11698 17980 11762 17984
rect 11698 17924 11702 17980
rect 11702 17924 11758 17980
rect 11758 17924 11762 17980
rect 11698 17920 11762 17924
rect 11778 17980 11842 17984
rect 11778 17924 11782 17980
rect 11782 17924 11838 17980
rect 11838 17924 11842 17980
rect 11778 17920 11842 17924
rect 11858 17980 11922 17984
rect 11858 17924 11862 17980
rect 11862 17924 11918 17980
rect 11918 17924 11922 17980
rect 11858 17920 11922 17924
rect 3618 17436 3682 17440
rect 3618 17380 3622 17436
rect 3622 17380 3678 17436
rect 3678 17380 3682 17436
rect 3618 17376 3682 17380
rect 3698 17436 3762 17440
rect 3698 17380 3702 17436
rect 3702 17380 3758 17436
rect 3758 17380 3762 17436
rect 3698 17376 3762 17380
rect 3778 17436 3842 17440
rect 3778 17380 3782 17436
rect 3782 17380 3838 17436
rect 3838 17380 3842 17436
rect 3778 17376 3842 17380
rect 3858 17436 3922 17440
rect 3858 17380 3862 17436
rect 3862 17380 3918 17436
rect 3918 17380 3922 17436
rect 3858 17376 3922 17380
rect 8952 17436 9016 17440
rect 8952 17380 8956 17436
rect 8956 17380 9012 17436
rect 9012 17380 9016 17436
rect 8952 17376 9016 17380
rect 9032 17436 9096 17440
rect 9032 17380 9036 17436
rect 9036 17380 9092 17436
rect 9092 17380 9096 17436
rect 9032 17376 9096 17380
rect 9112 17436 9176 17440
rect 9112 17380 9116 17436
rect 9116 17380 9172 17436
rect 9172 17380 9176 17436
rect 9112 17376 9176 17380
rect 9192 17436 9256 17440
rect 9192 17380 9196 17436
rect 9196 17380 9252 17436
rect 9252 17380 9256 17436
rect 9192 17376 9256 17380
rect 14285 17436 14349 17440
rect 14285 17380 14289 17436
rect 14289 17380 14345 17436
rect 14345 17380 14349 17436
rect 14285 17376 14349 17380
rect 14365 17436 14429 17440
rect 14365 17380 14369 17436
rect 14369 17380 14425 17436
rect 14425 17380 14429 17436
rect 14365 17376 14429 17380
rect 14445 17436 14509 17440
rect 14445 17380 14449 17436
rect 14449 17380 14505 17436
rect 14505 17380 14509 17436
rect 14445 17376 14509 17380
rect 14525 17436 14589 17440
rect 14525 17380 14529 17436
rect 14529 17380 14585 17436
rect 14585 17380 14589 17436
rect 14525 17376 14589 17380
rect 9628 17036 9692 17100
rect 6285 16892 6349 16896
rect 6285 16836 6289 16892
rect 6289 16836 6345 16892
rect 6345 16836 6349 16892
rect 6285 16832 6349 16836
rect 6365 16892 6429 16896
rect 6365 16836 6369 16892
rect 6369 16836 6425 16892
rect 6425 16836 6429 16892
rect 6365 16832 6429 16836
rect 6445 16892 6509 16896
rect 6445 16836 6449 16892
rect 6449 16836 6505 16892
rect 6505 16836 6509 16892
rect 6445 16832 6509 16836
rect 6525 16892 6589 16896
rect 6525 16836 6529 16892
rect 6529 16836 6585 16892
rect 6585 16836 6589 16892
rect 6525 16832 6589 16836
rect 11618 16892 11682 16896
rect 11618 16836 11622 16892
rect 11622 16836 11678 16892
rect 11678 16836 11682 16892
rect 11618 16832 11682 16836
rect 11698 16892 11762 16896
rect 11698 16836 11702 16892
rect 11702 16836 11758 16892
rect 11758 16836 11762 16892
rect 11698 16832 11762 16836
rect 11778 16892 11842 16896
rect 11778 16836 11782 16892
rect 11782 16836 11838 16892
rect 11838 16836 11842 16892
rect 11778 16832 11842 16836
rect 11858 16892 11922 16896
rect 11858 16836 11862 16892
rect 11862 16836 11918 16892
rect 11918 16836 11922 16892
rect 11858 16832 11922 16836
rect 5948 16824 6012 16828
rect 5948 16768 5962 16824
rect 5962 16768 6012 16824
rect 5948 16764 6012 16768
rect 3618 16348 3682 16352
rect 3618 16292 3622 16348
rect 3622 16292 3678 16348
rect 3678 16292 3682 16348
rect 3618 16288 3682 16292
rect 3698 16348 3762 16352
rect 3698 16292 3702 16348
rect 3702 16292 3758 16348
rect 3758 16292 3762 16348
rect 3698 16288 3762 16292
rect 3778 16348 3842 16352
rect 3778 16292 3782 16348
rect 3782 16292 3838 16348
rect 3838 16292 3842 16348
rect 3778 16288 3842 16292
rect 3858 16348 3922 16352
rect 3858 16292 3862 16348
rect 3862 16292 3918 16348
rect 3918 16292 3922 16348
rect 3858 16288 3922 16292
rect 8952 16348 9016 16352
rect 8952 16292 8956 16348
rect 8956 16292 9012 16348
rect 9012 16292 9016 16348
rect 8952 16288 9016 16292
rect 9032 16348 9096 16352
rect 9032 16292 9036 16348
rect 9036 16292 9092 16348
rect 9092 16292 9096 16348
rect 9032 16288 9096 16292
rect 9112 16348 9176 16352
rect 9112 16292 9116 16348
rect 9116 16292 9172 16348
rect 9172 16292 9176 16348
rect 9112 16288 9176 16292
rect 9192 16348 9256 16352
rect 9192 16292 9196 16348
rect 9196 16292 9252 16348
rect 9252 16292 9256 16348
rect 9192 16288 9256 16292
rect 14285 16348 14349 16352
rect 14285 16292 14289 16348
rect 14289 16292 14345 16348
rect 14345 16292 14349 16348
rect 14285 16288 14349 16292
rect 14365 16348 14429 16352
rect 14365 16292 14369 16348
rect 14369 16292 14425 16348
rect 14425 16292 14429 16348
rect 14365 16288 14429 16292
rect 14445 16348 14509 16352
rect 14445 16292 14449 16348
rect 14449 16292 14505 16348
rect 14505 16292 14509 16348
rect 14445 16288 14509 16292
rect 14525 16348 14589 16352
rect 14525 16292 14529 16348
rect 14529 16292 14585 16348
rect 14585 16292 14589 16348
rect 14525 16288 14589 16292
rect 6285 15804 6349 15808
rect 6285 15748 6289 15804
rect 6289 15748 6345 15804
rect 6345 15748 6349 15804
rect 6285 15744 6349 15748
rect 6365 15804 6429 15808
rect 6365 15748 6369 15804
rect 6369 15748 6425 15804
rect 6425 15748 6429 15804
rect 6365 15744 6429 15748
rect 6445 15804 6509 15808
rect 6445 15748 6449 15804
rect 6449 15748 6505 15804
rect 6505 15748 6509 15804
rect 6445 15744 6509 15748
rect 6525 15804 6589 15808
rect 6525 15748 6529 15804
rect 6529 15748 6585 15804
rect 6585 15748 6589 15804
rect 6525 15744 6589 15748
rect 11618 15804 11682 15808
rect 11618 15748 11622 15804
rect 11622 15748 11678 15804
rect 11678 15748 11682 15804
rect 11618 15744 11682 15748
rect 11698 15804 11762 15808
rect 11698 15748 11702 15804
rect 11702 15748 11758 15804
rect 11758 15748 11762 15804
rect 11698 15744 11762 15748
rect 11778 15804 11842 15808
rect 11778 15748 11782 15804
rect 11782 15748 11838 15804
rect 11838 15748 11842 15804
rect 11778 15744 11842 15748
rect 11858 15804 11922 15808
rect 11858 15748 11862 15804
rect 11862 15748 11918 15804
rect 11918 15748 11922 15804
rect 11858 15744 11922 15748
rect 3618 15260 3682 15264
rect 3618 15204 3622 15260
rect 3622 15204 3678 15260
rect 3678 15204 3682 15260
rect 3618 15200 3682 15204
rect 3698 15260 3762 15264
rect 3698 15204 3702 15260
rect 3702 15204 3758 15260
rect 3758 15204 3762 15260
rect 3698 15200 3762 15204
rect 3778 15260 3842 15264
rect 3778 15204 3782 15260
rect 3782 15204 3838 15260
rect 3838 15204 3842 15260
rect 3778 15200 3842 15204
rect 3858 15260 3922 15264
rect 3858 15204 3862 15260
rect 3862 15204 3918 15260
rect 3918 15204 3922 15260
rect 3858 15200 3922 15204
rect 8952 15260 9016 15264
rect 8952 15204 8956 15260
rect 8956 15204 9012 15260
rect 9012 15204 9016 15260
rect 8952 15200 9016 15204
rect 9032 15260 9096 15264
rect 9032 15204 9036 15260
rect 9036 15204 9092 15260
rect 9092 15204 9096 15260
rect 9032 15200 9096 15204
rect 9112 15260 9176 15264
rect 9112 15204 9116 15260
rect 9116 15204 9172 15260
rect 9172 15204 9176 15260
rect 9112 15200 9176 15204
rect 9192 15260 9256 15264
rect 9192 15204 9196 15260
rect 9196 15204 9252 15260
rect 9252 15204 9256 15260
rect 9192 15200 9256 15204
rect 14285 15260 14349 15264
rect 14285 15204 14289 15260
rect 14289 15204 14345 15260
rect 14345 15204 14349 15260
rect 14285 15200 14349 15204
rect 14365 15260 14429 15264
rect 14365 15204 14369 15260
rect 14369 15204 14425 15260
rect 14425 15204 14429 15260
rect 14365 15200 14429 15204
rect 14445 15260 14509 15264
rect 14445 15204 14449 15260
rect 14449 15204 14505 15260
rect 14505 15204 14509 15260
rect 14445 15200 14509 15204
rect 14525 15260 14589 15264
rect 14525 15204 14529 15260
rect 14529 15204 14585 15260
rect 14585 15204 14589 15260
rect 14525 15200 14589 15204
rect 6285 14716 6349 14720
rect 6285 14660 6289 14716
rect 6289 14660 6345 14716
rect 6345 14660 6349 14716
rect 6285 14656 6349 14660
rect 6365 14716 6429 14720
rect 6365 14660 6369 14716
rect 6369 14660 6425 14716
rect 6425 14660 6429 14716
rect 6365 14656 6429 14660
rect 6445 14716 6509 14720
rect 6445 14660 6449 14716
rect 6449 14660 6505 14716
rect 6505 14660 6509 14716
rect 6445 14656 6509 14660
rect 6525 14716 6589 14720
rect 6525 14660 6529 14716
rect 6529 14660 6585 14716
rect 6585 14660 6589 14716
rect 6525 14656 6589 14660
rect 11618 14716 11682 14720
rect 11618 14660 11622 14716
rect 11622 14660 11678 14716
rect 11678 14660 11682 14716
rect 11618 14656 11682 14660
rect 11698 14716 11762 14720
rect 11698 14660 11702 14716
rect 11702 14660 11758 14716
rect 11758 14660 11762 14716
rect 11698 14656 11762 14660
rect 11778 14716 11842 14720
rect 11778 14660 11782 14716
rect 11782 14660 11838 14716
rect 11838 14660 11842 14716
rect 11778 14656 11842 14660
rect 11858 14716 11922 14720
rect 11858 14660 11862 14716
rect 11862 14660 11918 14716
rect 11918 14660 11922 14716
rect 11858 14656 11922 14660
rect 3618 14172 3682 14176
rect 3618 14116 3622 14172
rect 3622 14116 3678 14172
rect 3678 14116 3682 14172
rect 3618 14112 3682 14116
rect 3698 14172 3762 14176
rect 3698 14116 3702 14172
rect 3702 14116 3758 14172
rect 3758 14116 3762 14172
rect 3698 14112 3762 14116
rect 3778 14172 3842 14176
rect 3778 14116 3782 14172
rect 3782 14116 3838 14172
rect 3838 14116 3842 14172
rect 3778 14112 3842 14116
rect 3858 14172 3922 14176
rect 3858 14116 3862 14172
rect 3862 14116 3918 14172
rect 3918 14116 3922 14172
rect 3858 14112 3922 14116
rect 8952 14172 9016 14176
rect 8952 14116 8956 14172
rect 8956 14116 9012 14172
rect 9012 14116 9016 14172
rect 8952 14112 9016 14116
rect 9032 14172 9096 14176
rect 9032 14116 9036 14172
rect 9036 14116 9092 14172
rect 9092 14116 9096 14172
rect 9032 14112 9096 14116
rect 9112 14172 9176 14176
rect 9112 14116 9116 14172
rect 9116 14116 9172 14172
rect 9172 14116 9176 14172
rect 9112 14112 9176 14116
rect 9192 14172 9256 14176
rect 9192 14116 9196 14172
rect 9196 14116 9252 14172
rect 9252 14116 9256 14172
rect 9192 14112 9256 14116
rect 14285 14172 14349 14176
rect 14285 14116 14289 14172
rect 14289 14116 14345 14172
rect 14345 14116 14349 14172
rect 14285 14112 14349 14116
rect 14365 14172 14429 14176
rect 14365 14116 14369 14172
rect 14369 14116 14425 14172
rect 14425 14116 14429 14172
rect 14365 14112 14429 14116
rect 14445 14172 14509 14176
rect 14445 14116 14449 14172
rect 14449 14116 14505 14172
rect 14505 14116 14509 14172
rect 14445 14112 14509 14116
rect 14525 14172 14589 14176
rect 14525 14116 14529 14172
rect 14529 14116 14585 14172
rect 14585 14116 14589 14172
rect 14525 14112 14589 14116
rect 6285 13628 6349 13632
rect 6285 13572 6289 13628
rect 6289 13572 6345 13628
rect 6345 13572 6349 13628
rect 6285 13568 6349 13572
rect 6365 13628 6429 13632
rect 6365 13572 6369 13628
rect 6369 13572 6425 13628
rect 6425 13572 6429 13628
rect 6365 13568 6429 13572
rect 6445 13628 6509 13632
rect 6445 13572 6449 13628
rect 6449 13572 6505 13628
rect 6505 13572 6509 13628
rect 6445 13568 6509 13572
rect 6525 13628 6589 13632
rect 6525 13572 6529 13628
rect 6529 13572 6585 13628
rect 6585 13572 6589 13628
rect 6525 13568 6589 13572
rect 11618 13628 11682 13632
rect 11618 13572 11622 13628
rect 11622 13572 11678 13628
rect 11678 13572 11682 13628
rect 11618 13568 11682 13572
rect 11698 13628 11762 13632
rect 11698 13572 11702 13628
rect 11702 13572 11758 13628
rect 11758 13572 11762 13628
rect 11698 13568 11762 13572
rect 11778 13628 11842 13632
rect 11778 13572 11782 13628
rect 11782 13572 11838 13628
rect 11838 13572 11842 13628
rect 11778 13568 11842 13572
rect 11858 13628 11922 13632
rect 11858 13572 11862 13628
rect 11862 13572 11918 13628
rect 11918 13572 11922 13628
rect 11858 13568 11922 13572
rect 3618 13084 3682 13088
rect 3618 13028 3622 13084
rect 3622 13028 3678 13084
rect 3678 13028 3682 13084
rect 3618 13024 3682 13028
rect 3698 13084 3762 13088
rect 3698 13028 3702 13084
rect 3702 13028 3758 13084
rect 3758 13028 3762 13084
rect 3698 13024 3762 13028
rect 3778 13084 3842 13088
rect 3778 13028 3782 13084
rect 3782 13028 3838 13084
rect 3838 13028 3842 13084
rect 3778 13024 3842 13028
rect 3858 13084 3922 13088
rect 3858 13028 3862 13084
rect 3862 13028 3918 13084
rect 3918 13028 3922 13084
rect 3858 13024 3922 13028
rect 8952 13084 9016 13088
rect 8952 13028 8956 13084
rect 8956 13028 9012 13084
rect 9012 13028 9016 13084
rect 8952 13024 9016 13028
rect 9032 13084 9096 13088
rect 9032 13028 9036 13084
rect 9036 13028 9092 13084
rect 9092 13028 9096 13084
rect 9032 13024 9096 13028
rect 9112 13084 9176 13088
rect 9112 13028 9116 13084
rect 9116 13028 9172 13084
rect 9172 13028 9176 13084
rect 9112 13024 9176 13028
rect 9192 13084 9256 13088
rect 9192 13028 9196 13084
rect 9196 13028 9252 13084
rect 9252 13028 9256 13084
rect 9192 13024 9256 13028
rect 14285 13084 14349 13088
rect 14285 13028 14289 13084
rect 14289 13028 14345 13084
rect 14345 13028 14349 13084
rect 14285 13024 14349 13028
rect 14365 13084 14429 13088
rect 14365 13028 14369 13084
rect 14369 13028 14425 13084
rect 14425 13028 14429 13084
rect 14365 13024 14429 13028
rect 14445 13084 14509 13088
rect 14445 13028 14449 13084
rect 14449 13028 14505 13084
rect 14505 13028 14509 13084
rect 14445 13024 14509 13028
rect 14525 13084 14589 13088
rect 14525 13028 14529 13084
rect 14529 13028 14585 13084
rect 14585 13028 14589 13084
rect 14525 13024 14589 13028
rect 6285 12540 6349 12544
rect 6285 12484 6289 12540
rect 6289 12484 6345 12540
rect 6345 12484 6349 12540
rect 6285 12480 6349 12484
rect 6365 12540 6429 12544
rect 6365 12484 6369 12540
rect 6369 12484 6425 12540
rect 6425 12484 6429 12540
rect 6365 12480 6429 12484
rect 6445 12540 6509 12544
rect 6445 12484 6449 12540
rect 6449 12484 6505 12540
rect 6505 12484 6509 12540
rect 6445 12480 6509 12484
rect 6525 12540 6589 12544
rect 6525 12484 6529 12540
rect 6529 12484 6585 12540
rect 6585 12484 6589 12540
rect 6525 12480 6589 12484
rect 11618 12540 11682 12544
rect 11618 12484 11622 12540
rect 11622 12484 11678 12540
rect 11678 12484 11682 12540
rect 11618 12480 11682 12484
rect 11698 12540 11762 12544
rect 11698 12484 11702 12540
rect 11702 12484 11758 12540
rect 11758 12484 11762 12540
rect 11698 12480 11762 12484
rect 11778 12540 11842 12544
rect 11778 12484 11782 12540
rect 11782 12484 11838 12540
rect 11838 12484 11842 12540
rect 11778 12480 11842 12484
rect 11858 12540 11922 12544
rect 11858 12484 11862 12540
rect 11862 12484 11918 12540
rect 11918 12484 11922 12540
rect 11858 12480 11922 12484
rect 9628 12276 9692 12340
rect 5948 12200 6012 12204
rect 5948 12144 5962 12200
rect 5962 12144 6012 12200
rect 5948 12140 6012 12144
rect 3618 11996 3682 12000
rect 3618 11940 3622 11996
rect 3622 11940 3678 11996
rect 3678 11940 3682 11996
rect 3618 11936 3682 11940
rect 3698 11996 3762 12000
rect 3698 11940 3702 11996
rect 3702 11940 3758 11996
rect 3758 11940 3762 11996
rect 3698 11936 3762 11940
rect 3778 11996 3842 12000
rect 3778 11940 3782 11996
rect 3782 11940 3838 11996
rect 3838 11940 3842 11996
rect 3778 11936 3842 11940
rect 3858 11996 3922 12000
rect 3858 11940 3862 11996
rect 3862 11940 3918 11996
rect 3918 11940 3922 11996
rect 3858 11936 3922 11940
rect 8952 11996 9016 12000
rect 8952 11940 8956 11996
rect 8956 11940 9012 11996
rect 9012 11940 9016 11996
rect 8952 11936 9016 11940
rect 9032 11996 9096 12000
rect 9032 11940 9036 11996
rect 9036 11940 9092 11996
rect 9092 11940 9096 11996
rect 9032 11936 9096 11940
rect 9112 11996 9176 12000
rect 9112 11940 9116 11996
rect 9116 11940 9172 11996
rect 9172 11940 9176 11996
rect 9112 11936 9176 11940
rect 9192 11996 9256 12000
rect 9192 11940 9196 11996
rect 9196 11940 9252 11996
rect 9252 11940 9256 11996
rect 9192 11936 9256 11940
rect 14285 11996 14349 12000
rect 14285 11940 14289 11996
rect 14289 11940 14345 11996
rect 14345 11940 14349 11996
rect 14285 11936 14349 11940
rect 14365 11996 14429 12000
rect 14365 11940 14369 11996
rect 14369 11940 14425 11996
rect 14425 11940 14429 11996
rect 14365 11936 14429 11940
rect 14445 11996 14509 12000
rect 14445 11940 14449 11996
rect 14449 11940 14505 11996
rect 14505 11940 14509 11996
rect 14445 11936 14509 11940
rect 14525 11996 14589 12000
rect 14525 11940 14529 11996
rect 14529 11940 14585 11996
rect 14585 11940 14589 11996
rect 14525 11936 14589 11940
rect 6285 11452 6349 11456
rect 6285 11396 6289 11452
rect 6289 11396 6345 11452
rect 6345 11396 6349 11452
rect 6285 11392 6349 11396
rect 6365 11452 6429 11456
rect 6365 11396 6369 11452
rect 6369 11396 6425 11452
rect 6425 11396 6429 11452
rect 6365 11392 6429 11396
rect 6445 11452 6509 11456
rect 6445 11396 6449 11452
rect 6449 11396 6505 11452
rect 6505 11396 6509 11452
rect 6445 11392 6509 11396
rect 6525 11452 6589 11456
rect 6525 11396 6529 11452
rect 6529 11396 6585 11452
rect 6585 11396 6589 11452
rect 6525 11392 6589 11396
rect 11618 11452 11682 11456
rect 11618 11396 11622 11452
rect 11622 11396 11678 11452
rect 11678 11396 11682 11452
rect 11618 11392 11682 11396
rect 11698 11452 11762 11456
rect 11698 11396 11702 11452
rect 11702 11396 11758 11452
rect 11758 11396 11762 11452
rect 11698 11392 11762 11396
rect 11778 11452 11842 11456
rect 11778 11396 11782 11452
rect 11782 11396 11838 11452
rect 11838 11396 11842 11452
rect 11778 11392 11842 11396
rect 11858 11452 11922 11456
rect 11858 11396 11862 11452
rect 11862 11396 11918 11452
rect 11918 11396 11922 11452
rect 11858 11392 11922 11396
rect 3618 10908 3682 10912
rect 3618 10852 3622 10908
rect 3622 10852 3678 10908
rect 3678 10852 3682 10908
rect 3618 10848 3682 10852
rect 3698 10908 3762 10912
rect 3698 10852 3702 10908
rect 3702 10852 3758 10908
rect 3758 10852 3762 10908
rect 3698 10848 3762 10852
rect 3778 10908 3842 10912
rect 3778 10852 3782 10908
rect 3782 10852 3838 10908
rect 3838 10852 3842 10908
rect 3778 10848 3842 10852
rect 3858 10908 3922 10912
rect 3858 10852 3862 10908
rect 3862 10852 3918 10908
rect 3918 10852 3922 10908
rect 3858 10848 3922 10852
rect 8952 10908 9016 10912
rect 8952 10852 8956 10908
rect 8956 10852 9012 10908
rect 9012 10852 9016 10908
rect 8952 10848 9016 10852
rect 9032 10908 9096 10912
rect 9032 10852 9036 10908
rect 9036 10852 9092 10908
rect 9092 10852 9096 10908
rect 9032 10848 9096 10852
rect 9112 10908 9176 10912
rect 9112 10852 9116 10908
rect 9116 10852 9172 10908
rect 9172 10852 9176 10908
rect 9112 10848 9176 10852
rect 9192 10908 9256 10912
rect 9192 10852 9196 10908
rect 9196 10852 9252 10908
rect 9252 10852 9256 10908
rect 9192 10848 9256 10852
rect 14285 10908 14349 10912
rect 14285 10852 14289 10908
rect 14289 10852 14345 10908
rect 14345 10852 14349 10908
rect 14285 10848 14349 10852
rect 14365 10908 14429 10912
rect 14365 10852 14369 10908
rect 14369 10852 14425 10908
rect 14425 10852 14429 10908
rect 14365 10848 14429 10852
rect 14445 10908 14509 10912
rect 14445 10852 14449 10908
rect 14449 10852 14505 10908
rect 14505 10852 14509 10908
rect 14445 10848 14509 10852
rect 14525 10908 14589 10912
rect 14525 10852 14529 10908
rect 14529 10852 14585 10908
rect 14585 10852 14589 10908
rect 14525 10848 14589 10852
rect 6285 10364 6349 10368
rect 6285 10308 6289 10364
rect 6289 10308 6345 10364
rect 6345 10308 6349 10364
rect 6285 10304 6349 10308
rect 6365 10364 6429 10368
rect 6365 10308 6369 10364
rect 6369 10308 6425 10364
rect 6425 10308 6429 10364
rect 6365 10304 6429 10308
rect 6445 10364 6509 10368
rect 6445 10308 6449 10364
rect 6449 10308 6505 10364
rect 6505 10308 6509 10364
rect 6445 10304 6509 10308
rect 6525 10364 6589 10368
rect 6525 10308 6529 10364
rect 6529 10308 6585 10364
rect 6585 10308 6589 10364
rect 6525 10304 6589 10308
rect 11618 10364 11682 10368
rect 11618 10308 11622 10364
rect 11622 10308 11678 10364
rect 11678 10308 11682 10364
rect 11618 10304 11682 10308
rect 11698 10364 11762 10368
rect 11698 10308 11702 10364
rect 11702 10308 11758 10364
rect 11758 10308 11762 10364
rect 11698 10304 11762 10308
rect 11778 10364 11842 10368
rect 11778 10308 11782 10364
rect 11782 10308 11838 10364
rect 11838 10308 11842 10364
rect 11778 10304 11842 10308
rect 11858 10364 11922 10368
rect 11858 10308 11862 10364
rect 11862 10308 11918 10364
rect 11918 10308 11922 10364
rect 11858 10304 11922 10308
rect 3618 9820 3682 9824
rect 3618 9764 3622 9820
rect 3622 9764 3678 9820
rect 3678 9764 3682 9820
rect 3618 9760 3682 9764
rect 3698 9820 3762 9824
rect 3698 9764 3702 9820
rect 3702 9764 3758 9820
rect 3758 9764 3762 9820
rect 3698 9760 3762 9764
rect 3778 9820 3842 9824
rect 3778 9764 3782 9820
rect 3782 9764 3838 9820
rect 3838 9764 3842 9820
rect 3778 9760 3842 9764
rect 3858 9820 3922 9824
rect 3858 9764 3862 9820
rect 3862 9764 3918 9820
rect 3918 9764 3922 9820
rect 3858 9760 3922 9764
rect 8952 9820 9016 9824
rect 8952 9764 8956 9820
rect 8956 9764 9012 9820
rect 9012 9764 9016 9820
rect 8952 9760 9016 9764
rect 9032 9820 9096 9824
rect 9032 9764 9036 9820
rect 9036 9764 9092 9820
rect 9092 9764 9096 9820
rect 9032 9760 9096 9764
rect 9112 9820 9176 9824
rect 9112 9764 9116 9820
rect 9116 9764 9172 9820
rect 9172 9764 9176 9820
rect 9112 9760 9176 9764
rect 9192 9820 9256 9824
rect 9192 9764 9196 9820
rect 9196 9764 9252 9820
rect 9252 9764 9256 9820
rect 9192 9760 9256 9764
rect 14285 9820 14349 9824
rect 14285 9764 14289 9820
rect 14289 9764 14345 9820
rect 14345 9764 14349 9820
rect 14285 9760 14349 9764
rect 14365 9820 14429 9824
rect 14365 9764 14369 9820
rect 14369 9764 14425 9820
rect 14425 9764 14429 9820
rect 14365 9760 14429 9764
rect 14445 9820 14509 9824
rect 14445 9764 14449 9820
rect 14449 9764 14505 9820
rect 14505 9764 14509 9820
rect 14445 9760 14509 9764
rect 14525 9820 14589 9824
rect 14525 9764 14529 9820
rect 14529 9764 14585 9820
rect 14585 9764 14589 9820
rect 14525 9760 14589 9764
rect 6285 9276 6349 9280
rect 6285 9220 6289 9276
rect 6289 9220 6345 9276
rect 6345 9220 6349 9276
rect 6285 9216 6349 9220
rect 6365 9276 6429 9280
rect 6365 9220 6369 9276
rect 6369 9220 6425 9276
rect 6425 9220 6429 9276
rect 6365 9216 6429 9220
rect 6445 9276 6509 9280
rect 6445 9220 6449 9276
rect 6449 9220 6505 9276
rect 6505 9220 6509 9276
rect 6445 9216 6509 9220
rect 6525 9276 6589 9280
rect 6525 9220 6529 9276
rect 6529 9220 6585 9276
rect 6585 9220 6589 9276
rect 6525 9216 6589 9220
rect 11618 9276 11682 9280
rect 11618 9220 11622 9276
rect 11622 9220 11678 9276
rect 11678 9220 11682 9276
rect 11618 9216 11682 9220
rect 11698 9276 11762 9280
rect 11698 9220 11702 9276
rect 11702 9220 11758 9276
rect 11758 9220 11762 9276
rect 11698 9216 11762 9220
rect 11778 9276 11842 9280
rect 11778 9220 11782 9276
rect 11782 9220 11838 9276
rect 11838 9220 11842 9276
rect 11778 9216 11842 9220
rect 11858 9276 11922 9280
rect 11858 9220 11862 9276
rect 11862 9220 11918 9276
rect 11918 9220 11922 9276
rect 11858 9216 11922 9220
rect 3618 8732 3682 8736
rect 3618 8676 3622 8732
rect 3622 8676 3678 8732
rect 3678 8676 3682 8732
rect 3618 8672 3682 8676
rect 3698 8732 3762 8736
rect 3698 8676 3702 8732
rect 3702 8676 3758 8732
rect 3758 8676 3762 8732
rect 3698 8672 3762 8676
rect 3778 8732 3842 8736
rect 3778 8676 3782 8732
rect 3782 8676 3838 8732
rect 3838 8676 3842 8732
rect 3778 8672 3842 8676
rect 3858 8732 3922 8736
rect 3858 8676 3862 8732
rect 3862 8676 3918 8732
rect 3918 8676 3922 8732
rect 3858 8672 3922 8676
rect 8952 8732 9016 8736
rect 8952 8676 8956 8732
rect 8956 8676 9012 8732
rect 9012 8676 9016 8732
rect 8952 8672 9016 8676
rect 9032 8732 9096 8736
rect 9032 8676 9036 8732
rect 9036 8676 9092 8732
rect 9092 8676 9096 8732
rect 9032 8672 9096 8676
rect 9112 8732 9176 8736
rect 9112 8676 9116 8732
rect 9116 8676 9172 8732
rect 9172 8676 9176 8732
rect 9112 8672 9176 8676
rect 9192 8732 9256 8736
rect 9192 8676 9196 8732
rect 9196 8676 9252 8732
rect 9252 8676 9256 8732
rect 9192 8672 9256 8676
rect 14285 8732 14349 8736
rect 14285 8676 14289 8732
rect 14289 8676 14345 8732
rect 14345 8676 14349 8732
rect 14285 8672 14349 8676
rect 14365 8732 14429 8736
rect 14365 8676 14369 8732
rect 14369 8676 14425 8732
rect 14425 8676 14429 8732
rect 14365 8672 14429 8676
rect 14445 8732 14509 8736
rect 14445 8676 14449 8732
rect 14449 8676 14505 8732
rect 14505 8676 14509 8732
rect 14445 8672 14509 8676
rect 14525 8732 14589 8736
rect 14525 8676 14529 8732
rect 14529 8676 14585 8732
rect 14585 8676 14589 8732
rect 14525 8672 14589 8676
rect 6285 8188 6349 8192
rect 6285 8132 6289 8188
rect 6289 8132 6345 8188
rect 6345 8132 6349 8188
rect 6285 8128 6349 8132
rect 6365 8188 6429 8192
rect 6365 8132 6369 8188
rect 6369 8132 6425 8188
rect 6425 8132 6429 8188
rect 6365 8128 6429 8132
rect 6445 8188 6509 8192
rect 6445 8132 6449 8188
rect 6449 8132 6505 8188
rect 6505 8132 6509 8188
rect 6445 8128 6509 8132
rect 6525 8188 6589 8192
rect 6525 8132 6529 8188
rect 6529 8132 6585 8188
rect 6585 8132 6589 8188
rect 6525 8128 6589 8132
rect 11618 8188 11682 8192
rect 11618 8132 11622 8188
rect 11622 8132 11678 8188
rect 11678 8132 11682 8188
rect 11618 8128 11682 8132
rect 11698 8188 11762 8192
rect 11698 8132 11702 8188
rect 11702 8132 11758 8188
rect 11758 8132 11762 8188
rect 11698 8128 11762 8132
rect 11778 8188 11842 8192
rect 11778 8132 11782 8188
rect 11782 8132 11838 8188
rect 11838 8132 11842 8188
rect 11778 8128 11842 8132
rect 11858 8188 11922 8192
rect 11858 8132 11862 8188
rect 11862 8132 11918 8188
rect 11918 8132 11922 8188
rect 11858 8128 11922 8132
rect 3618 7644 3682 7648
rect 3618 7588 3622 7644
rect 3622 7588 3678 7644
rect 3678 7588 3682 7644
rect 3618 7584 3682 7588
rect 3698 7644 3762 7648
rect 3698 7588 3702 7644
rect 3702 7588 3758 7644
rect 3758 7588 3762 7644
rect 3698 7584 3762 7588
rect 3778 7644 3842 7648
rect 3778 7588 3782 7644
rect 3782 7588 3838 7644
rect 3838 7588 3842 7644
rect 3778 7584 3842 7588
rect 3858 7644 3922 7648
rect 3858 7588 3862 7644
rect 3862 7588 3918 7644
rect 3918 7588 3922 7644
rect 3858 7584 3922 7588
rect 8952 7644 9016 7648
rect 8952 7588 8956 7644
rect 8956 7588 9012 7644
rect 9012 7588 9016 7644
rect 8952 7584 9016 7588
rect 9032 7644 9096 7648
rect 9032 7588 9036 7644
rect 9036 7588 9092 7644
rect 9092 7588 9096 7644
rect 9032 7584 9096 7588
rect 9112 7644 9176 7648
rect 9112 7588 9116 7644
rect 9116 7588 9172 7644
rect 9172 7588 9176 7644
rect 9112 7584 9176 7588
rect 9192 7644 9256 7648
rect 9192 7588 9196 7644
rect 9196 7588 9252 7644
rect 9252 7588 9256 7644
rect 9192 7584 9256 7588
rect 14285 7644 14349 7648
rect 14285 7588 14289 7644
rect 14289 7588 14345 7644
rect 14345 7588 14349 7644
rect 14285 7584 14349 7588
rect 14365 7644 14429 7648
rect 14365 7588 14369 7644
rect 14369 7588 14425 7644
rect 14425 7588 14429 7644
rect 14365 7584 14429 7588
rect 14445 7644 14509 7648
rect 14445 7588 14449 7644
rect 14449 7588 14505 7644
rect 14505 7588 14509 7644
rect 14445 7584 14509 7588
rect 14525 7644 14589 7648
rect 14525 7588 14529 7644
rect 14529 7588 14585 7644
rect 14585 7588 14589 7644
rect 14525 7584 14589 7588
rect 6285 7100 6349 7104
rect 6285 7044 6289 7100
rect 6289 7044 6345 7100
rect 6345 7044 6349 7100
rect 6285 7040 6349 7044
rect 6365 7100 6429 7104
rect 6365 7044 6369 7100
rect 6369 7044 6425 7100
rect 6425 7044 6429 7100
rect 6365 7040 6429 7044
rect 6445 7100 6509 7104
rect 6445 7044 6449 7100
rect 6449 7044 6505 7100
rect 6505 7044 6509 7100
rect 6445 7040 6509 7044
rect 6525 7100 6589 7104
rect 6525 7044 6529 7100
rect 6529 7044 6585 7100
rect 6585 7044 6589 7100
rect 6525 7040 6589 7044
rect 11618 7100 11682 7104
rect 11618 7044 11622 7100
rect 11622 7044 11678 7100
rect 11678 7044 11682 7100
rect 11618 7040 11682 7044
rect 11698 7100 11762 7104
rect 11698 7044 11702 7100
rect 11702 7044 11758 7100
rect 11758 7044 11762 7100
rect 11698 7040 11762 7044
rect 11778 7100 11842 7104
rect 11778 7044 11782 7100
rect 11782 7044 11838 7100
rect 11838 7044 11842 7100
rect 11778 7040 11842 7044
rect 11858 7100 11922 7104
rect 11858 7044 11862 7100
rect 11862 7044 11918 7100
rect 11918 7044 11922 7100
rect 11858 7040 11922 7044
rect 3618 6556 3682 6560
rect 3618 6500 3622 6556
rect 3622 6500 3678 6556
rect 3678 6500 3682 6556
rect 3618 6496 3682 6500
rect 3698 6556 3762 6560
rect 3698 6500 3702 6556
rect 3702 6500 3758 6556
rect 3758 6500 3762 6556
rect 3698 6496 3762 6500
rect 3778 6556 3842 6560
rect 3778 6500 3782 6556
rect 3782 6500 3838 6556
rect 3838 6500 3842 6556
rect 3778 6496 3842 6500
rect 3858 6556 3922 6560
rect 3858 6500 3862 6556
rect 3862 6500 3918 6556
rect 3918 6500 3922 6556
rect 3858 6496 3922 6500
rect 8952 6556 9016 6560
rect 8952 6500 8956 6556
rect 8956 6500 9012 6556
rect 9012 6500 9016 6556
rect 8952 6496 9016 6500
rect 9032 6556 9096 6560
rect 9032 6500 9036 6556
rect 9036 6500 9092 6556
rect 9092 6500 9096 6556
rect 9032 6496 9096 6500
rect 9112 6556 9176 6560
rect 9112 6500 9116 6556
rect 9116 6500 9172 6556
rect 9172 6500 9176 6556
rect 9112 6496 9176 6500
rect 9192 6556 9256 6560
rect 9192 6500 9196 6556
rect 9196 6500 9252 6556
rect 9252 6500 9256 6556
rect 9192 6496 9256 6500
rect 14285 6556 14349 6560
rect 14285 6500 14289 6556
rect 14289 6500 14345 6556
rect 14345 6500 14349 6556
rect 14285 6496 14349 6500
rect 14365 6556 14429 6560
rect 14365 6500 14369 6556
rect 14369 6500 14425 6556
rect 14425 6500 14429 6556
rect 14365 6496 14429 6500
rect 14445 6556 14509 6560
rect 14445 6500 14449 6556
rect 14449 6500 14505 6556
rect 14505 6500 14509 6556
rect 14445 6496 14509 6500
rect 14525 6556 14589 6560
rect 14525 6500 14529 6556
rect 14529 6500 14585 6556
rect 14585 6500 14589 6556
rect 14525 6496 14589 6500
rect 9444 6352 9508 6356
rect 9444 6296 9458 6352
rect 9458 6296 9508 6352
rect 9444 6292 9508 6296
rect 6285 6012 6349 6016
rect 6285 5956 6289 6012
rect 6289 5956 6345 6012
rect 6345 5956 6349 6012
rect 6285 5952 6349 5956
rect 6365 6012 6429 6016
rect 6365 5956 6369 6012
rect 6369 5956 6425 6012
rect 6425 5956 6429 6012
rect 6365 5952 6429 5956
rect 6445 6012 6509 6016
rect 6445 5956 6449 6012
rect 6449 5956 6505 6012
rect 6505 5956 6509 6012
rect 6445 5952 6509 5956
rect 6525 6012 6589 6016
rect 6525 5956 6529 6012
rect 6529 5956 6585 6012
rect 6585 5956 6589 6012
rect 6525 5952 6589 5956
rect 11618 6012 11682 6016
rect 11618 5956 11622 6012
rect 11622 5956 11678 6012
rect 11678 5956 11682 6012
rect 11618 5952 11682 5956
rect 11698 6012 11762 6016
rect 11698 5956 11702 6012
rect 11702 5956 11758 6012
rect 11758 5956 11762 6012
rect 11698 5952 11762 5956
rect 11778 6012 11842 6016
rect 11778 5956 11782 6012
rect 11782 5956 11838 6012
rect 11838 5956 11842 6012
rect 11778 5952 11842 5956
rect 11858 6012 11922 6016
rect 11858 5956 11862 6012
rect 11862 5956 11918 6012
rect 11918 5956 11922 6012
rect 11858 5952 11922 5956
rect 3618 5468 3682 5472
rect 3618 5412 3622 5468
rect 3622 5412 3678 5468
rect 3678 5412 3682 5468
rect 3618 5408 3682 5412
rect 3698 5468 3762 5472
rect 3698 5412 3702 5468
rect 3702 5412 3758 5468
rect 3758 5412 3762 5468
rect 3698 5408 3762 5412
rect 3778 5468 3842 5472
rect 3778 5412 3782 5468
rect 3782 5412 3838 5468
rect 3838 5412 3842 5468
rect 3778 5408 3842 5412
rect 3858 5468 3922 5472
rect 3858 5412 3862 5468
rect 3862 5412 3918 5468
rect 3918 5412 3922 5468
rect 3858 5408 3922 5412
rect 8952 5468 9016 5472
rect 8952 5412 8956 5468
rect 8956 5412 9012 5468
rect 9012 5412 9016 5468
rect 8952 5408 9016 5412
rect 9032 5468 9096 5472
rect 9032 5412 9036 5468
rect 9036 5412 9092 5468
rect 9092 5412 9096 5468
rect 9032 5408 9096 5412
rect 9112 5468 9176 5472
rect 9112 5412 9116 5468
rect 9116 5412 9172 5468
rect 9172 5412 9176 5468
rect 9112 5408 9176 5412
rect 9192 5468 9256 5472
rect 9192 5412 9196 5468
rect 9196 5412 9252 5468
rect 9252 5412 9256 5468
rect 9192 5408 9256 5412
rect 14285 5468 14349 5472
rect 14285 5412 14289 5468
rect 14289 5412 14345 5468
rect 14345 5412 14349 5468
rect 14285 5408 14349 5412
rect 14365 5468 14429 5472
rect 14365 5412 14369 5468
rect 14369 5412 14425 5468
rect 14425 5412 14429 5468
rect 14365 5408 14429 5412
rect 14445 5468 14509 5472
rect 14445 5412 14449 5468
rect 14449 5412 14505 5468
rect 14505 5412 14509 5468
rect 14445 5408 14509 5412
rect 14525 5468 14589 5472
rect 14525 5412 14529 5468
rect 14529 5412 14585 5468
rect 14585 5412 14589 5468
rect 14525 5408 14589 5412
rect 6285 4924 6349 4928
rect 6285 4868 6289 4924
rect 6289 4868 6345 4924
rect 6345 4868 6349 4924
rect 6285 4864 6349 4868
rect 6365 4924 6429 4928
rect 6365 4868 6369 4924
rect 6369 4868 6425 4924
rect 6425 4868 6429 4924
rect 6365 4864 6429 4868
rect 6445 4924 6509 4928
rect 6445 4868 6449 4924
rect 6449 4868 6505 4924
rect 6505 4868 6509 4924
rect 6445 4864 6509 4868
rect 6525 4924 6589 4928
rect 6525 4868 6529 4924
rect 6529 4868 6585 4924
rect 6585 4868 6589 4924
rect 6525 4864 6589 4868
rect 11618 4924 11682 4928
rect 11618 4868 11622 4924
rect 11622 4868 11678 4924
rect 11678 4868 11682 4924
rect 11618 4864 11682 4868
rect 11698 4924 11762 4928
rect 11698 4868 11702 4924
rect 11702 4868 11758 4924
rect 11758 4868 11762 4924
rect 11698 4864 11762 4868
rect 11778 4924 11842 4928
rect 11778 4868 11782 4924
rect 11782 4868 11838 4924
rect 11838 4868 11842 4924
rect 11778 4864 11842 4868
rect 11858 4924 11922 4928
rect 11858 4868 11862 4924
rect 11862 4868 11918 4924
rect 11918 4868 11922 4924
rect 11858 4864 11922 4868
rect 3618 4380 3682 4384
rect 3618 4324 3622 4380
rect 3622 4324 3678 4380
rect 3678 4324 3682 4380
rect 3618 4320 3682 4324
rect 3698 4380 3762 4384
rect 3698 4324 3702 4380
rect 3702 4324 3758 4380
rect 3758 4324 3762 4380
rect 3698 4320 3762 4324
rect 3778 4380 3842 4384
rect 3778 4324 3782 4380
rect 3782 4324 3838 4380
rect 3838 4324 3842 4380
rect 3778 4320 3842 4324
rect 3858 4380 3922 4384
rect 3858 4324 3862 4380
rect 3862 4324 3918 4380
rect 3918 4324 3922 4380
rect 3858 4320 3922 4324
rect 8952 4380 9016 4384
rect 8952 4324 8956 4380
rect 8956 4324 9012 4380
rect 9012 4324 9016 4380
rect 8952 4320 9016 4324
rect 9032 4380 9096 4384
rect 9032 4324 9036 4380
rect 9036 4324 9092 4380
rect 9092 4324 9096 4380
rect 9032 4320 9096 4324
rect 9112 4380 9176 4384
rect 9112 4324 9116 4380
rect 9116 4324 9172 4380
rect 9172 4324 9176 4380
rect 9112 4320 9176 4324
rect 9192 4380 9256 4384
rect 9192 4324 9196 4380
rect 9196 4324 9252 4380
rect 9252 4324 9256 4380
rect 9192 4320 9256 4324
rect 14285 4380 14349 4384
rect 14285 4324 14289 4380
rect 14289 4324 14345 4380
rect 14345 4324 14349 4380
rect 14285 4320 14349 4324
rect 14365 4380 14429 4384
rect 14365 4324 14369 4380
rect 14369 4324 14425 4380
rect 14425 4324 14429 4380
rect 14365 4320 14429 4324
rect 14445 4380 14509 4384
rect 14445 4324 14449 4380
rect 14449 4324 14505 4380
rect 14505 4324 14509 4380
rect 14445 4320 14509 4324
rect 14525 4380 14589 4384
rect 14525 4324 14529 4380
rect 14529 4324 14585 4380
rect 14585 4324 14589 4380
rect 14525 4320 14589 4324
rect 6285 3836 6349 3840
rect 6285 3780 6289 3836
rect 6289 3780 6345 3836
rect 6345 3780 6349 3836
rect 6285 3776 6349 3780
rect 6365 3836 6429 3840
rect 6365 3780 6369 3836
rect 6369 3780 6425 3836
rect 6425 3780 6429 3836
rect 6365 3776 6429 3780
rect 6445 3836 6509 3840
rect 6445 3780 6449 3836
rect 6449 3780 6505 3836
rect 6505 3780 6509 3836
rect 6445 3776 6509 3780
rect 6525 3836 6589 3840
rect 6525 3780 6529 3836
rect 6529 3780 6585 3836
rect 6585 3780 6589 3836
rect 6525 3776 6589 3780
rect 11618 3836 11682 3840
rect 11618 3780 11622 3836
rect 11622 3780 11678 3836
rect 11678 3780 11682 3836
rect 11618 3776 11682 3780
rect 11698 3836 11762 3840
rect 11698 3780 11702 3836
rect 11702 3780 11758 3836
rect 11758 3780 11762 3836
rect 11698 3776 11762 3780
rect 11778 3836 11842 3840
rect 11778 3780 11782 3836
rect 11782 3780 11838 3836
rect 11838 3780 11842 3836
rect 11778 3776 11842 3780
rect 11858 3836 11922 3840
rect 11858 3780 11862 3836
rect 11862 3780 11918 3836
rect 11918 3780 11922 3836
rect 11858 3776 11922 3780
rect 3618 3292 3682 3296
rect 3618 3236 3622 3292
rect 3622 3236 3678 3292
rect 3678 3236 3682 3292
rect 3618 3232 3682 3236
rect 3698 3292 3762 3296
rect 3698 3236 3702 3292
rect 3702 3236 3758 3292
rect 3758 3236 3762 3292
rect 3698 3232 3762 3236
rect 3778 3292 3842 3296
rect 3778 3236 3782 3292
rect 3782 3236 3838 3292
rect 3838 3236 3842 3292
rect 3778 3232 3842 3236
rect 3858 3292 3922 3296
rect 3858 3236 3862 3292
rect 3862 3236 3918 3292
rect 3918 3236 3922 3292
rect 3858 3232 3922 3236
rect 8952 3292 9016 3296
rect 8952 3236 8956 3292
rect 8956 3236 9012 3292
rect 9012 3236 9016 3292
rect 8952 3232 9016 3236
rect 9032 3292 9096 3296
rect 9032 3236 9036 3292
rect 9036 3236 9092 3292
rect 9092 3236 9096 3292
rect 9032 3232 9096 3236
rect 9112 3292 9176 3296
rect 9112 3236 9116 3292
rect 9116 3236 9172 3292
rect 9172 3236 9176 3292
rect 9112 3232 9176 3236
rect 9192 3292 9256 3296
rect 9192 3236 9196 3292
rect 9196 3236 9252 3292
rect 9252 3236 9256 3292
rect 9192 3232 9256 3236
rect 14285 3292 14349 3296
rect 14285 3236 14289 3292
rect 14289 3236 14345 3292
rect 14345 3236 14349 3292
rect 14285 3232 14349 3236
rect 14365 3292 14429 3296
rect 14365 3236 14369 3292
rect 14369 3236 14425 3292
rect 14425 3236 14429 3292
rect 14365 3232 14429 3236
rect 14445 3292 14509 3296
rect 14445 3236 14449 3292
rect 14449 3236 14505 3292
rect 14505 3236 14509 3292
rect 14445 3232 14509 3236
rect 14525 3292 14589 3296
rect 14525 3236 14529 3292
rect 14529 3236 14585 3292
rect 14585 3236 14589 3292
rect 14525 3232 14589 3236
rect 6285 2748 6349 2752
rect 6285 2692 6289 2748
rect 6289 2692 6345 2748
rect 6345 2692 6349 2748
rect 6285 2688 6349 2692
rect 6365 2748 6429 2752
rect 6365 2692 6369 2748
rect 6369 2692 6425 2748
rect 6425 2692 6429 2748
rect 6365 2688 6429 2692
rect 6445 2748 6509 2752
rect 6445 2692 6449 2748
rect 6449 2692 6505 2748
rect 6505 2692 6509 2748
rect 6445 2688 6509 2692
rect 6525 2748 6589 2752
rect 6525 2692 6529 2748
rect 6529 2692 6585 2748
rect 6585 2692 6589 2748
rect 6525 2688 6589 2692
rect 11618 2748 11682 2752
rect 11618 2692 11622 2748
rect 11622 2692 11678 2748
rect 11678 2692 11682 2748
rect 11618 2688 11682 2692
rect 11698 2748 11762 2752
rect 11698 2692 11702 2748
rect 11702 2692 11758 2748
rect 11758 2692 11762 2748
rect 11698 2688 11762 2692
rect 11778 2748 11842 2752
rect 11778 2692 11782 2748
rect 11782 2692 11838 2748
rect 11838 2692 11842 2748
rect 11778 2688 11842 2692
rect 11858 2748 11922 2752
rect 11858 2692 11862 2748
rect 11862 2692 11918 2748
rect 11918 2692 11922 2748
rect 11858 2688 11922 2692
rect 9444 2680 9508 2684
rect 9444 2624 9494 2680
rect 9494 2624 9508 2680
rect 9444 2620 9508 2624
rect 3618 2204 3682 2208
rect 3618 2148 3622 2204
rect 3622 2148 3678 2204
rect 3678 2148 3682 2204
rect 3618 2144 3682 2148
rect 3698 2204 3762 2208
rect 3698 2148 3702 2204
rect 3702 2148 3758 2204
rect 3758 2148 3762 2204
rect 3698 2144 3762 2148
rect 3778 2204 3842 2208
rect 3778 2148 3782 2204
rect 3782 2148 3838 2204
rect 3838 2148 3842 2204
rect 3778 2144 3842 2148
rect 3858 2204 3922 2208
rect 3858 2148 3862 2204
rect 3862 2148 3918 2204
rect 3918 2148 3922 2204
rect 3858 2144 3922 2148
rect 8952 2204 9016 2208
rect 8952 2148 8956 2204
rect 8956 2148 9012 2204
rect 9012 2148 9016 2204
rect 8952 2144 9016 2148
rect 9032 2204 9096 2208
rect 9032 2148 9036 2204
rect 9036 2148 9092 2204
rect 9092 2148 9096 2204
rect 9032 2144 9096 2148
rect 9112 2204 9176 2208
rect 9112 2148 9116 2204
rect 9116 2148 9172 2204
rect 9172 2148 9176 2204
rect 9112 2144 9176 2148
rect 9192 2204 9256 2208
rect 9192 2148 9196 2204
rect 9196 2148 9252 2204
rect 9252 2148 9256 2204
rect 9192 2144 9256 2148
rect 14285 2204 14349 2208
rect 14285 2148 14289 2204
rect 14289 2148 14345 2204
rect 14345 2148 14349 2204
rect 14285 2144 14349 2148
rect 14365 2204 14429 2208
rect 14365 2148 14369 2204
rect 14369 2148 14425 2204
rect 14425 2148 14429 2204
rect 14365 2144 14429 2148
rect 14445 2204 14509 2208
rect 14445 2148 14449 2204
rect 14449 2148 14505 2204
rect 14505 2148 14509 2204
rect 14445 2144 14509 2148
rect 14525 2204 14589 2208
rect 14525 2148 14529 2204
rect 14529 2148 14585 2204
rect 14585 2148 14589 2204
rect 14525 2144 14589 2148
<< metal4 >>
rect 3610 37024 3931 37584
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3931 37024
rect 3610 35936 3931 36960
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3931 35936
rect 3610 34848 3931 35872
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3931 34848
rect 3610 33760 3931 34784
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3931 33760
rect 3610 32672 3931 33696
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3931 32672
rect 3610 31584 3931 32608
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3931 31584
rect 3610 30496 3931 31520
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3931 30496
rect 3610 29408 3931 30432
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3931 29408
rect 3610 28320 3931 29344
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3931 28320
rect 3610 27232 3931 28256
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3931 27232
rect 3610 26144 3931 27168
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3931 26144
rect 3610 25056 3931 26080
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3931 25056
rect 3610 23968 3931 24992
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3931 23968
rect 3610 22880 3931 23904
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3931 22880
rect 3610 21792 3931 22816
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3931 21792
rect 3610 20704 3931 21728
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3931 20704
rect 3610 19616 3931 20640
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3931 19616
rect 3610 18528 3931 19552
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3931 18528
rect 3610 17440 3931 18464
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3931 17440
rect 3610 16352 3931 17376
rect 6277 37568 6597 37584
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 36480 6597 37504
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 35392 6597 36416
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 34304 6597 35328
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 33216 6597 34240
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 32128 6597 33152
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 31040 6597 32064
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 29952 6597 30976
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 28864 6597 29888
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 27776 6597 28800
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 26688 6597 27712
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 25600 6597 26624
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 24512 6597 25536
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 23424 6597 24448
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 22336 6597 23360
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 21248 6597 22272
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 20160 6597 21184
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 19072 6597 20096
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 17984 6597 19008
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 16896 6597 17920
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 5947 16828 6013 16829
rect 5947 16764 5948 16828
rect 6012 16764 6013 16828
rect 5947 16763 6013 16764
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3931 16352
rect 3610 15264 3931 16288
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3931 15264
rect 3610 14176 3931 15200
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3931 14176
rect 3610 13088 3931 14112
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3931 13088
rect 3610 12000 3931 13024
rect 5950 12205 6010 16763
rect 6277 15808 6597 16832
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 14720 6597 15744
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 13632 6597 14656
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 12544 6597 13568
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 5947 12204 6013 12205
rect 5947 12140 5948 12204
rect 6012 12140 6013 12204
rect 5947 12139 6013 12140
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3931 12000
rect 3610 10912 3931 11936
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3931 10912
rect 3610 9824 3931 10848
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3931 9824
rect 3610 8736 3931 9760
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3931 8736
rect 3610 7648 3931 8672
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3931 7648
rect 3610 6560 3931 7584
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3931 6560
rect 3610 5472 3931 6496
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3931 5472
rect 3610 4384 3931 5408
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3931 4384
rect 3610 3296 3931 4320
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3931 3296
rect 3610 2208 3931 3232
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3931 2208
rect 3610 2128 3931 2144
rect 6277 11456 6597 12480
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 10368 6597 11392
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 9280 6597 10304
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 8192 6597 9216
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 7104 6597 8128
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 6016 6597 7040
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 4928 6597 5952
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 3840 6597 4864
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 2752 6597 3776
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2128 6597 2688
rect 8944 37024 9264 37584
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 35936 9264 36960
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 34848 9264 35872
rect 11610 37568 11930 37584
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 36480 11930 37504
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 35392 11930 36416
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11467 35188 11533 35189
rect 11467 35124 11468 35188
rect 11532 35124 11533 35188
rect 11467 35123 11533 35124
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 33760 9264 34784
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 32672 9264 33696
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 31584 9264 32608
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 30496 9264 31520
rect 9627 31516 9693 31517
rect 9627 31452 9628 31516
rect 9692 31452 9693 31516
rect 9627 31451 9693 31452
rect 9630 31245 9690 31451
rect 9627 31244 9693 31245
rect 9627 31180 9628 31244
rect 9692 31180 9693 31244
rect 9627 31179 9693 31180
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 29408 9264 30432
rect 11470 29613 11530 35123
rect 11610 34304 11930 35328
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 33216 11930 34240
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 32128 11930 33152
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 31040 11930 32064
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 29952 11930 30976
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11467 29612 11533 29613
rect 11467 29548 11468 29612
rect 11532 29548 11533 29612
rect 11467 29547 11533 29548
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 28320 9264 29344
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 27232 9264 28256
rect 11610 28864 11930 29888
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11467 28252 11533 28253
rect 11467 28188 11468 28252
rect 11532 28188 11533 28252
rect 11467 28187 11533 28188
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 26144 9264 27168
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 25056 9264 26080
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 23968 9264 24992
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 22880 9264 23904
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 21792 9264 22816
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 20704 9264 21728
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 19616 9264 20640
rect 11470 19821 11530 28187
rect 11610 27776 11930 28800
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 26688 11930 27712
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 25600 11930 26624
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 24512 11930 25536
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 23424 11930 24448
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 22336 11930 23360
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 21248 11930 22272
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 20160 11930 21184
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11467 19820 11533 19821
rect 11467 19756 11468 19820
rect 11532 19756 11533 19820
rect 11467 19755 11533 19756
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 18528 9264 19552
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 17440 9264 18464
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 16352 9264 17376
rect 11610 19072 11930 20096
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 17984 11930 19008
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 9627 17100 9693 17101
rect 9627 17036 9628 17100
rect 9692 17036 9693 17100
rect 9627 17035 9693 17036
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 15264 9264 16288
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 14176 9264 15200
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 13088 9264 14112
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 12000 9264 13024
rect 9630 12341 9690 17035
rect 11610 16896 11930 17920
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 15808 11930 16832
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 14720 11930 15744
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 13632 11930 14656
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 12544 11930 13568
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 9627 12340 9693 12341
rect 9627 12276 9628 12340
rect 9692 12276 9693 12340
rect 9627 12275 9693 12276
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 10912 9264 11936
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 9824 9264 10848
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 8736 9264 9760
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 7648 9264 8672
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 6560 9264 7584
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 5472 9264 6496
rect 11610 11456 11930 12480
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 10368 11930 11392
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 9280 11930 10304
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 8192 11930 9216
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 7104 11930 8128
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 9443 6356 9509 6357
rect 9443 6292 9444 6356
rect 9508 6292 9509 6356
rect 9443 6291 9509 6292
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 4384 9264 5408
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 3296 9264 4320
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 2208 9264 3232
rect 9446 2685 9506 6291
rect 11610 6016 11930 7040
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 4928 11930 5952
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 3840 11930 4864
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 2752 11930 3776
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 9443 2684 9509 2685
rect 9443 2620 9444 2684
rect 9508 2620 9509 2684
rect 9443 2619 9509 2620
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2128 9264 2144
rect 11610 2128 11930 2688
rect 14277 37024 14597 37584
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 35936 14597 36960
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 34848 14597 35872
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 33760 14597 34784
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 32672 14597 33696
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 31584 14597 32608
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 30496 14597 31520
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 29408 14597 30432
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 28320 14597 29344
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 27232 14597 28256
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 26144 14597 27168
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 25056 14597 26080
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 23968 14597 24992
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 22880 14597 23904
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 21792 14597 22816
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 20704 14597 21728
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 19616 14597 20640
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 18528 14597 19552
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 17440 14597 18464
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 16352 14597 17376
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 15264 14597 16288
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 14176 14597 15200
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 13088 14597 14112
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 12000 14597 13024
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 10912 14597 11936
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 9824 14597 10848
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 8736 14597 9760
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 7648 14597 8672
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 6560 14597 7584
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 5472 14597 6496
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 4384 14597 5408
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 3296 14597 4320
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 2208 14597 3232
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2128 14597 2144
use sky130_fd_sc_hd__decap_4  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6
timestamp 1604681595
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _29_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1932 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_29
timestamp 1604681595
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_25
timestamp 1604681595
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1604681595
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41
timestamp 1604681595
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4140 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45
timestamp 1604681595
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1604681595
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_49
timestamp 1604681595
transform 1 0 5612 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1604681595
transform 1 0 5428 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _42_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5612 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_56
timestamp 1604681595
transform 1 0 6256 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_53 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5980 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53
timestamp 1604681595
transform 1 0 5980 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1604681595
transform 1 0 6072 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60
timestamp 1604681595
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1604681595
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1604681595
transform 1 0 6348 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 6440 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_70
timestamp 1604681595
transform 1 0 7544 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_66
timestamp 1604681595
transform 1 0 7176 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1604681595
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67
timestamp 1604681595
transform 1 0 7268 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_73
timestamp 1604681595
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8188 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_93
timestamp 1604681595
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1604681595
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_97
timestamp 1604681595
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10028 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10396 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_110
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1604681595
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1604681595
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_106
timestamp 1604681595
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11408 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11040 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_118
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_117
timestamp 1604681595
transform 1 0 11868 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 12052 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1604681595
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1604681595
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1604681595
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_129
timestamp 1604681595
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_133 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13340 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145
timestamp 1604681595
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1604681595
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_136
timestamp 1604681595
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_140 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13984 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 1840 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7
timestamp 1604681595
transform 1 0 1748 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_10
timestamp 1604681595
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1604681595
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_41
timestamp 1604681595
transform 1 0 4876 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 6440 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 6256 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5428 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 5796 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_45
timestamp 1604681595
transform 1 0 5244 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_49
timestamp 1604681595
transform 1 0 5612 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_53
timestamp 1604681595
transform 1 0 5980 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_67
timestamp 1604681595
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_71
timestamp 1604681595
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10120 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 9936 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1604681595
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_88
timestamp 1604681595
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 11684 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11132 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 11500 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_107
timestamp 1604681595
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_111
timestamp 1604681595
transform 1 0 11316 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_124
timestamp 1604681595
transform 1 0 12512 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1604681595
transform 1 0 13248 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12696 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13064 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_128
timestamp 1604681595
transform 1 0 12880 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_136 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13616 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_144
timestamp 1604681595
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 14812 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604681595
transform 1 0 2116 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1604681595
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1604681595
transform 1 0 1932 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_7
timestamp 1604681595
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_19
timestamp 1604681595
transform 1 0 2852 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 3864 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 3680 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 3312 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 4876 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_23
timestamp 1604681595
transform 1 0 3220 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_26
timestamp 1604681595
transform 1 0 3496 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_39
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_43
timestamp 1604681595
transform 1 0 5060 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 5244 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_51
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1604681595
transform 1 0 5428 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_55
timestamp 1604681595
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1604681595
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7912 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1604681595
transform 1 0 7360 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_66
timestamp 1604681595
transform 1 0 7176 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_70
timestamp 1604681595
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_83
timestamp 1604681595
transform 1 0 8740 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10028 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1604681595
transform 1 0 8924 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_87
timestamp 1604681595
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_91
timestamp 1604681595
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_95
timestamp 1604681595
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_106
timestamp 1604681595
transform 1 0 10856 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_112
timestamp 1604681595
transform 1 0 11408 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604681595
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1604681595
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_132
timestamp 1604681595
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_136
timestamp 1604681595
transform 1 0 13616 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_144
timestamp 1604681595
transform 1 0 14352 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1604681595
transform 1 0 2668 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_9
timestamp 1604681595
transform 1 0 1932 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_13
timestamp 1604681595
transform 1 0 2300 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_16
timestamp 1604681595
transform 1 0 2576 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4324 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3496 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_21
timestamp 1604681595
transform 1 0 3036 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_25
timestamp 1604681595
transform 1 0 3404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_28
timestamp 1604681595
transform 1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6164 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 5336 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 5704 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_44
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_48
timestamp 1604681595
transform 1 0 5520 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_52
timestamp 1604681595
transform 1 0 5888 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1604681595
transform 1 0 8372 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_71
timestamp 1604681595
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_75
timestamp 1604681595
transform 1 0 8004 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_83
timestamp 1604681595
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 8924 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_87
timestamp 1604681595
transform 1 0 9108 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_102
timestamp 1604681595
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 11224 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11040 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_106
timestamp 1604681595
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_119
timestamp 1604681595
transform 1 0 12052 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_125
timestamp 1604681595
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1604681595
transform 1 0 12788 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_131
timestamp 1604681595
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_143
timestamp 1604681595
transform 1 0 14260 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 14812 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 1932 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_18
timestamp 1604681595
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 3496 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3312 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4508 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_22
timestamp 1604681595
transform 1 0 3128 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_35
timestamp 1604681595
transform 1 0 4324 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_39
timestamp 1604681595
transform 1 0 4692 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 5060 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_52
timestamp 1604681595
transform 1 0 5888 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1604681595
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 8372 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_71
timestamp 1604681595
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_75
timestamp 1604681595
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10580 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_88
timestamp 1604681595
transform 1 0 9200 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_92
timestamp 1604681595
transform 1 0 9568 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_95
timestamp 1604681595
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_99
timestamp 1604681595
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_112
timestamp 1604681595
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_116
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_126
timestamp 1604681595
transform 1 0 12696 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_138
timestamp 1604681595
transform 1 0 13800 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7
timestamp 1604681595
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_9
timestamp 1604681595
transform 1 0 1932 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1604681595
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_13
timestamp 1604681595
transform 1 0 2300 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 2116 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 2116 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_23
timestamp 1604681595
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_41
timestamp 1604681595
transform 1 0 4876 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_33
timestamp 1604681595
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604681595
transform 1 0 4508 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_45
timestamp 1604681595
transform 1 0 5244 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_48
timestamp 1604681595
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5704 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1604681595
transform 1 0 5428 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1604681595
transform 1 0 5060 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1604681595
transform 1 0 5612 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1604681595
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_53
timestamp 1604681595
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_52
timestamp 1604681595
transform 1 0 5888 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 6072 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1604681595
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_71
timestamp 1604681595
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_69
timestamp 1604681595
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_65
timestamp 1604681595
transform 1 0 7084 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7636 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_75
timestamp 1604681595
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1604681595
transform 1 0 8648 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7820 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1604681595
transform 1 0 8372 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_83
timestamp 1604681595
transform 1 0 8740 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_91
timestamp 1604681595
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_87
timestamp 1604681595
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_86
timestamp 1604681595
transform 1 0 9016 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1604681595
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1604681595
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_95
timestamp 1604681595
transform 1 0 9844 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 9936 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_112
timestamp 1604681595
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_109
timestamp 1604681595
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1604681595
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_116
timestamp 1604681595
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_125
timestamp 1604681595
transform 1 0 12604 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_113
timestamp 1604681595
transform 1 0 11500 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_137
timestamp 1604681595
transform 1 0 13708 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_145
timestamp 1604681595
transform 1 0 14444 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_135
timestamp 1604681595
transform 1 0 13524 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_143
timestamp 1604681595
transform 1 0 14260 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 14812 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604681595
transform 1 0 2668 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_9
timestamp 1604681595
transform 1 0 1932 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_13
timestamp 1604681595
transform 1 0 2300 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_16
timestamp 1604681595
transform 1 0 2576 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 4784 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 4232 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_21
timestamp 1604681595
transform 1 0 3036 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_25
timestamp 1604681595
transform 1 0 3404 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_36
timestamp 1604681595
transform 1 0 4416 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1604681595
transform 1 0 6072 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1604681595
transform 1 0 4968 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5612 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_46
timestamp 1604681595
transform 1 0 5336 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_51
timestamp 1604681595
transform 1 0 5796 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_58
timestamp 1604681595
transform 1 0 6440 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7268 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8280 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8648 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_64
timestamp 1604681595
transform 1 0 6992 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_76
timestamp 1604681595
transform 1 0 8096 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_80
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 10212 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1604681595
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_88
timestamp 1604681595
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_97
timestamp 1604681595
transform 1 0 10028 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_101
timestamp 1604681595
transform 1 0 10396 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10948 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1604681595
transform 1 0 12420 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_135
timestamp 1604681595
transform 1 0 13524 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_143
timestamp 1604681595
transform 1 0 14260 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 14812 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604681595
transform 1 0 2668 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_9
timestamp 1604681595
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_13
timestamp 1604681595
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1604681595
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_21
timestamp 1604681595
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_25
timestamp 1604681595
transform 1 0 3404 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_31
timestamp 1604681595
transform 1 0 3956 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_34
timestamp 1604681595
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_38
timestamp 1604681595
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4968 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_51
timestamp 1604681595
transform 1 0 5796 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_55
timestamp 1604681595
transform 1 0 6164 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 7268 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1604681595
transform 1 0 7084 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_83
timestamp 1604681595
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_87
timestamp 1604681595
transform 1 0 9108 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_99
timestamp 1604681595
transform 1 0 10212 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_107
timestamp 1604681595
transform 1 0 10948 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_111
timestamp 1604681595
transform 1 0 11316 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_115
timestamp 1604681595
transform 1 0 11684 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1604681595
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_135
timestamp 1604681595
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_143
timestamp 1604681595
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 14812 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 2116 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_7
timestamp 1604681595
transform 1 0 1748 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_13
timestamp 1604681595
transform 1 0 2300 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_17
timestamp 1604681595
transform 1 0 2668 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_20
timestamp 1604681595
transform 1 0 2944 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1604681595
transform 1 0 4600 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_28
timestamp 1604681595
transform 1 0 3680 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_10_41
timestamp 1604681595
transform 1 0 4876 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 5612 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_46
timestamp 1604681595
transform 1 0 5336 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_58
timestamp 1604681595
transform 1 0 6440 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1604681595
transform 1 0 7176 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 7728 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 8096 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_64
timestamp 1604681595
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_70
timestamp 1604681595
transform 1 0 7544 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_74
timestamp 1604681595
transform 1 0 7912 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_78
timestamp 1604681595
transform 1 0 8280 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_88
timestamp 1604681595
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 11132 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_105
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_125
timestamp 1604681595
transform 1 0 12604 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_137
timestamp 1604681595
transform 1 0 13708 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_145
timestamp 1604681595
transform 1 0 14444 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 2760 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_9
timestamp 1604681595
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_13
timestamp 1604681595
transform 1 0 2300 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_34
timestamp 1604681595
transform 1 0 4232 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_40
timestamp 1604681595
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_53
timestamp 1604681595
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1604681595
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_78
timestamp 1604681595
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_82
timestamp 1604681595
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9016 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 8832 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 10672 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_102
timestamp 1604681595
transform 1 0 10488 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_106
timestamp 1604681595
transform 1 0 10856 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_110
timestamp 1604681595
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_135
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_143
timestamp 1604681595
transform 1 0 14260 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 14812 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2300 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_11
timestamp 1604681595
transform 1 0 2116 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604681595
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_40
timestamp 1604681595
transform 1 0 4784 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 5060 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_59
timestamp 1604681595
transform 1 0 6532 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 7268 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8280 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 8648 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_64
timestamp 1604681595
transform 1 0 6992 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_76
timestamp 1604681595
transform 1 0 8096 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_80
timestamp 1604681595
transform 1 0 8464 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10212 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9844 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_84
timestamp 1604681595
transform 1 0 8832 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_97
timestamp 1604681595
transform 1 0 10028 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_115
timestamp 1604681595
transform 1 0 11684 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_127
timestamp 1604681595
transform 1 0 12788 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_139
timestamp 1604681595
transform 1 0 13892 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_145
timestamp 1604681595
transform 1 0 14444 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 14812 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2300 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 2300 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_11
timestamp 1604681595
transform 1 0 2116 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604681595
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 3864 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 3312 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_22
timestamp 1604681595
transform 1 0 3128 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_26
timestamp 1604681595
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_50
timestamp 1604681595
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_46
timestamp 1604681595
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5336 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_61
timestamp 1604681595
transform 1 0 6716 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_55
timestamp 1604681595
transform 1 0 6164 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_58
timestamp 1604681595
transform 1 0 6440 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_54
timestamp 1604681595
transform 1 0 6072 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_64
timestamp 1604681595
transform 1 0 6992 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_71
timestamp 1604681595
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7452 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_82
timestamp 1604681595
transform 1 0 8648 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_78
timestamp 1604681595
transform 1 0 8280 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_75
timestamp 1604681595
transform 1 0 8004 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8464 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 8280 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8464 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_88
timestamp 1604681595
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_103
timestamp 1604681595
transform 1 0 10580 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_100
timestamp 1604681595
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_96
timestamp 1604681595
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9752 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10672 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_111
timestamp 1604681595
transform 1 0 11316 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_107
timestamp 1604681595
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_113
timestamp 1604681595
transform 1 0 11500 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11500 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11132 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_115
timestamp 1604681595
transform 1 0 11684 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1604681595
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11868 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_119
timestamp 1604681595
transform 1 0 12052 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_135
timestamp 1604681595
transform 1 0 13524 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_143
timestamp 1604681595
transform 1 0 14260 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_131
timestamp 1604681595
transform 1 0 13156 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_143
timestamp 1604681595
transform 1 0 14260 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 14812 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 14812 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_9
timestamp 1604681595
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_13
timestamp 1604681595
transform 1 0 2300 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3772 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3588 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_25
timestamp 1604681595
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_38
timestamp 1604681595
transform 1 0 4600 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_50
timestamp 1604681595
transform 1 0 5704 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_58
timestamp 1604681595
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7912 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_65
timestamp 1604681595
transform 1 0 7084 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_69
timestamp 1604681595
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_73
timestamp 1604681595
transform 1 0 7820 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10120 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_90
timestamp 1604681595
transform 1 0 9384 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_95
timestamp 1604681595
transform 1 0 9844 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_107
timestamp 1604681595
transform 1 0 10948 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_112
timestamp 1604681595
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_116
timestamp 1604681595
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1604681595
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_135
timestamp 1604681595
transform 1 0 13524 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_143
timestamp 1604681595
transform 1 0 14260 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 14812 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_15
timestamp 1604681595
transform 1 0 2484 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3128 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_21
timestamp 1604681595
transform 1 0 3036 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1604681595
transform 1 0 3312 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_28
timestamp 1604681595
transform 1 0 3680 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 6532 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1604681595
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_56
timestamp 1604681595
transform 1 0 6256 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_61
timestamp 1604681595
transform 1 0 6716 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7268 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 8280 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_65
timestamp 1604681595
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_76
timestamp 1604681595
transform 1 0 8096 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_80
timestamp 1604681595
transform 1 0 8464 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_84
timestamp 1604681595
transform 1 0 8832 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_16_102
timestamp 1604681595
transform 1 0 10488 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 11224 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10764 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_107
timestamp 1604681595
transform 1 0 10948 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_119
timestamp 1604681595
transform 1 0 12052 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_131
timestamp 1604681595
transform 1 0 13156 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_143
timestamp 1604681595
transform 1 0 14260 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 14812 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_15
timestamp 1604681595
transform 1 0 2484 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_19
timestamp 1604681595
transform 1 0 2852 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 3128 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_31
timestamp 1604681595
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_35
timestamp 1604681595
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_39
timestamp 1604681595
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_43
timestamp 1604681595
transform 1 0 5060 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1604681595
transform 1 0 5796 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1604681595
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8556 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6900 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7912 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_72
timestamp 1604681595
transform 1 0 7728 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_76
timestamp 1604681595
transform 1 0 8096 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_97
timestamp 1604681595
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_101
timestamp 1604681595
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_114
timestamp 1604681595
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 1604681595
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_135
timestamp 1604681595
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_143
timestamp 1604681595
transform 1 0 14260 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 14812 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_7
timestamp 1604681595
transform 1 0 1748 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_12
timestamp 1604681595
transform 1 0 2208 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_20
timestamp 1604681595
transform 1 0 2944 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3128 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_24
timestamp 1604681595
transform 1 0 3312 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_41
timestamp 1604681595
transform 1 0 4876 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6808 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5612 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_46
timestamp 1604681595
transform 1 0 5336 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_52
timestamp 1604681595
transform 1 0 5888 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_78
timestamp 1604681595
transform 1 0 8280 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_83
timestamp 1604681595
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_87
timestamp 1604681595
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 8924 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1604681595
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 9292 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_97
timestamp 1604681595
transform 1 0 10028 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_101
timestamp 1604681595
transform 1 0 10396 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 10212 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10764 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1604681595
transform 1 0 12236 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_133
timestamp 1604681595
transform 1 0 13340 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_145
timestamp 1604681595
transform 1 0 14444 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 14812 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_9
timestamp 1604681595
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1604681595
transform 1 0 1748 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_17
timestamp 1604681595
transform 1 0 2668 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_13
timestamp 1604681595
transform 1 0 2300 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_19
timestamp 1604681595
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 2760 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 2116 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2024 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1604681595
transform 1 0 2944 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1604681595
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_23
timestamp 1604681595
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 3588 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_40
timestamp 1604681595
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_36
timestamp 1604681595
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4324 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4508 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_20_53
timestamp 1604681595
transform 1 0 5980 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1604681595
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1604681595
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6532 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6716 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 8372 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_71
timestamp 1604681595
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_75
timestamp 1604681595
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_82
timestamp 1604681595
transform 1 0 8648 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_77
timestamp 1604681595
transform 1 0 8188 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_81
timestamp 1604681595
transform 1 0 8556 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 8924 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 8924 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_101
timestamp 1604681595
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_88
timestamp 1604681595
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_102
timestamp 1604681595
transform 1 0 10488 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1604681595
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_105
timestamp 1604681595
transform 1 0 10764 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 11040 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 11224 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1604681595
transform 1 0 11224 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1604681595
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_117
timestamp 1604681595
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 12052 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_119
timestamp 1604681595
transform 1 0 12052 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_135
timestamp 1604681595
transform 1 0 13524 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_143
timestamp 1604681595
transform 1 0 14260 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_131
timestamp 1604681595
transform 1 0 13156 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_143
timestamp 1604681595
transform 1 0 14260 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 14812 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 14812 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2760 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_15
timestamp 1604681595
transform 1 0 2484 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_34
timestamp 1604681595
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_38
timestamp 1604681595
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4968 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_51
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_55
timestamp 1604681595
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 7268 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_66
timestamp 1604681595
transform 1 0 7176 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_69
timestamp 1604681595
transform 1 0 7452 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_73
timestamp 1604681595
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_77
timestamp 1604681595
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_81
timestamp 1604681595
transform 1 0 8556 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 10212 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_91
timestamp 1604681595
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_95
timestamp 1604681595
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_108
timestamp 1604681595
transform 1 0 11040 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_135
timestamp 1604681595
transform 1 0 13524 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_143
timestamp 1604681595
transform 1 0 14260 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 14812 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_15
timestamp 1604681595
transform 1 0 2484 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4508 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 4324 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 3128 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_21
timestamp 1604681595
transform 1 0 3036 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_24
timestamp 1604681595
transform 1 0 3312 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_30
timestamp 1604681595
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 6072 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_46
timestamp 1604681595
transform 1 0 5336 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_50
timestamp 1604681595
transform 1 0 5704 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_57
timestamp 1604681595
transform 1 0 6348 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_61
timestamp 1604681595
transform 1 0 6716 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1604681595
transform 1 0 7636 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 7360 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_67
timestamp 1604681595
transform 1 0 7268 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1604681595
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9936 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10304 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_98
timestamp 1604681595
transform 1 0 10120 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_102
timestamp 1604681595
transform 1 0 10488 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_114
timestamp 1604681595
transform 1 0 11592 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_126
timestamp 1604681595
transform 1 0 12696 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_138
timestamp 1604681595
transform 1 0 13800 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 14812 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_15
timestamp 1604681595
transform 1 0 2484 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_19
timestamp 1604681595
transform 1 0 2852 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 3128 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_23_38
timestamp 1604681595
transform 1 0 4600 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_50
timestamp 1604681595
transform 1 0 5704 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1604681595
transform 1 0 7084 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_74
timestamp 1604681595
transform 1 0 7912 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_78
timestamp 1604681595
transform 1 0 8280 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9936 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9752 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9016 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_88
timestamp 1604681595
transform 1 0 9200 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_92
timestamp 1604681595
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10948 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_105
timestamp 1604681595
transform 1 0 10764 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_109
timestamp 1604681595
transform 1 0 11132 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1604681595
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_135
timestamp 1604681595
transform 1 0 13524 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_143
timestamp 1604681595
transform 1 0 14260 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 14812 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604681595
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_40
timestamp 1604681595
transform 1 0 4784 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1604681595
transform 1 0 6532 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 5336 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 5704 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_44
timestamp 1604681595
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_48
timestamp 1604681595
transform 1 0 5520 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_52
timestamp 1604681595
transform 1 0 5888 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_58
timestamp 1604681595
transform 1 0 6440 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604681595
transform 1 0 8096 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 8556 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_68
timestamp 1604681595
transform 1 0 7360 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_72
timestamp 1604681595
transform 1 0 7728 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_75
timestamp 1604681595
transform 1 0 8004 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_79
timestamp 1604681595
transform 1 0 8372 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_83
timestamp 1604681595
transform 1 0 8740 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9936 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_87
timestamp 1604681595
transform 1 0 9108 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1604681595
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1604681595
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1604681595
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1604681595
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1604681595
transform 1 0 14076 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1604681595
transform 1 0 14444 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 14812 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_9
timestamp 1604681595
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_13
timestamp 1604681595
transform 1 0 2300 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_25
timestamp 1604681595
transform 1 0 3404 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_37
timestamp 1604681595
transform 1 0 4508 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4968 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_51
timestamp 1604681595
transform 1 0 5796 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_55
timestamp 1604681595
transform 1 0 6164 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 6992 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 8648 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_80
timestamp 1604681595
transform 1 0 8464 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9200 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9016 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_84
timestamp 1604681595
transform 1 0 8832 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_104
timestamp 1604681595
transform 1 0 10672 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 10948 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_109
timestamp 1604681595
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_113
timestamp 1604681595
transform 1 0 11500 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1604681595
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_135
timestamp 1604681595
transform 1 0 13524 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_143
timestamp 1604681595
transform 1 0 14260 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 14812 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_20
timestamp 1604681595
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_16
timestamp 1604681595
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_11
timestamp 1604681595
transform 1 0 2116 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604681595
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_24
timestamp 1604681595
transform 1 0 3312 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_30
timestamp 1604681595
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3128 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3680 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 3680 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_37
timestamp 1604681595
transform 1 0 4508 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_40
timestamp 1604681595
transform 1 0 4784 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_41
timestamp 1604681595
transform 1 0 4876 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_44
timestamp 1604681595
transform 1 0 5152 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_48
timestamp 1604681595
transform 1 0 5520 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_44
timestamp 1604681595
transform 1 0 5152 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 5336 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4968 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 5244 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_60
timestamp 1604681595
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_48
timestamp 1604681595
transform 1 0 5520 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5612 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_26_69
timestamp 1604681595
transform 1 0 7452 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_65
timestamp 1604681595
transform 1 0 7084 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 7360 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 7544 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_81
timestamp 1604681595
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_77
timestamp 1604681595
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_73
timestamp 1604681595
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_82
timestamp 1604681595
transform 1 0 8648 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1604681595
transform 1 0 7820 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_93
timestamp 1604681595
transform 1 0 9660 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_85
timestamp 1604681595
transform 1 0 8924 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1604681595
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_103
timestamp 1604681595
transform 1 0 10580 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_98
timestamp 1604681595
transform 1 0 10120 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10396 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9936 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9936 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10948 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10948 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_123
timestamp 1604681595
transform 1 0 12420 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_105
timestamp 1604681595
transform 1 0 10764 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_109
timestamp 1604681595
transform 1 0 11132 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1604681595
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_135
timestamp 1604681595
transform 1 0 13524 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_143
timestamp 1604681595
transform 1 0 14260 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_135
timestamp 1604681595
transform 1 0 13524 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_143
timestamp 1604681595
transform 1 0 14260 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 14812 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 14812 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_11
timestamp 1604681595
transform 1 0 2116 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_23
timestamp 1604681595
transform 1 0 3220 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_30
timestamp 1604681595
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3680 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_40
timestamp 1604681595
transform 1 0 4784 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_36
timestamp 1604681595
transform 1 0 4416 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4968 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 6808 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_58
timestamp 1604681595
transform 1 0 6440 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 7176 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 7728 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_64
timestamp 1604681595
transform 1 0 6992 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_68
timestamp 1604681595
transform 1 0 7360 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_74
timestamp 1604681595
transform 1 0 7912 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10396 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9936 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_84
timestamp 1604681595
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_98
timestamp 1604681595
transform 1 0 10120 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_110
timestamp 1604681595
transform 1 0 11224 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_122
timestamp 1604681595
transform 1 0 12328 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_134
timestamp 1604681595
transform 1 0 13432 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 14812 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_15
timestamp 1604681595
transform 1 0 2484 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_19
timestamp 1604681595
transform 1 0 2852 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 3128 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_38
timestamp 1604681595
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_51
timestamp 1604681595
transform 1 0 5796 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_47
timestamp 1604681595
transform 1 0 5428 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_42
timestamp 1604681595
transform 1 0 4968 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 5244 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 5612 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_55
timestamp 1604681595
transform 1 0 6164 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 8464 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_78
timestamp 1604681595
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_82
timestamp 1604681595
transform 1 0 8648 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10304 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9660 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9292 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_87
timestamp 1604681595
transform 1 0 9108 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_91
timestamp 1604681595
transform 1 0 9476 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_95
timestamp 1604681595
transform 1 0 9844 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 11316 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 11684 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 12052 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_109
timestamp 1604681595
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1604681595
transform 1 0 11500 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_117
timestamp 1604681595
transform 1 0 11868 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_121
timestamp 1604681595
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_135
timestamp 1604681595
transform 1 0 13524 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_143
timestamp 1604681595
transform 1 0 14260 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 14812 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 2392 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_7
timestamp 1604681595
transform 1 0 1748 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_13
timestamp 1604681595
transform 1 0 2300 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_16
timestamp 1604681595
transform 1 0 2576 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 3128 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1604681595
transform 1 0 3312 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_28
timestamp 1604681595
transform 1 0 3680 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_41
timestamp 1604681595
transform 1 0 4876 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1604681595
transform 1 0 5612 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6624 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 5428 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_58
timestamp 1604681595
transform 1 0 6440 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_62
timestamp 1604681595
transform 1 0 6808 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7176 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 6992 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_86
timestamp 1604681595
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1604681595
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_102
timestamp 1604681595
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 11224 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 11040 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_106
timestamp 1604681595
transform 1 0 10856 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_119
timestamp 1604681595
transform 1 0 12052 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 12972 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_127
timestamp 1604681595
transform 1 0 12788 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_131
timestamp 1604681595
transform 1 0 13156 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_143
timestamp 1604681595
transform 1 0 14260 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 14812 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2392 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 2760 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_9
timestamp 1604681595
transform 1 0 1932 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_13
timestamp 1604681595
transform 1 0 2300 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_16
timestamp 1604681595
transform 1 0 2576 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_20
timestamp 1604681595
transform 1 0 2944 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1604681595
transform 1 0 3772 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_25
timestamp 1604681595
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_38
timestamp 1604681595
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_42
timestamp 1604681595
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 5152 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1604681595
transform 1 0 5336 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_49
timestamp 1604681595
transform 1 0 5612 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_56
timestamp 1604681595
transform 1 0 6256 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_53
timestamp 1604681595
transform 1 0 5980 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 6072 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8464 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1604681595
transform 1 0 7360 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 7176 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_77
timestamp 1604681595
transform 1 0 8188 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10028 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9476 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_89
timestamp 1604681595
transform 1 0 9292 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_93
timestamp 1604681595
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_114
timestamp 1604681595
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1604681595
transform 1 0 11224 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_106
timestamp 1604681595
transform 1 0 10856 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 11408 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 11040 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1604681595
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_132
timestamp 1604681595
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_136
timestamp 1604681595
transform 1 0 13616 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_144
timestamp 1604681595
transform 1 0 14352 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 14812 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_11
timestamp 1604681595
transform 1 0 2116 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4508 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_23
timestamp 1604681595
transform 1 0 3220 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_36
timestamp 1604681595
transform 1 0 4416 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1604681595
transform 1 0 6072 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5888 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 5520 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_46
timestamp 1604681595
transform 1 0 5336 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_50
timestamp 1604681595
transform 1 0 5704 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6900 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1604681595
transform 1 0 7728 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8740 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_81
timestamp 1604681595
transform 1 0 8556 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1604681595
transform 1 0 8924 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9108 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_89
timestamp 1604681595
transform 1 0 9292 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 9844 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1604681595
transform 1 0 10028 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_100
timestamp 1604681595
transform 1 0 10304 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 10488 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_104
timestamp 1604681595
transform 1 0 10672 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12604 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1604681595
transform 1 0 11040 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 10856 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 12052 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_117
timestamp 1604681595
transform 1 0 11868 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_121
timestamp 1604681595
transform 1 0 12236 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_134
timestamp 1604681595
transform 1 0 13432 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 14812 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_9
timestamp 1604681595
transform 1 0 1932 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_7
timestamp 1604681595
transform 1 0 1748 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_13
timestamp 1604681595
transform 1 0 2300 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 2576 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 2392 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_18
timestamp 1604681595
transform 1 0 2760 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 2576 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4784 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_32
timestamp 1604681595
transform 1 0 4048 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_30
timestamp 1604681595
transform 1 0 3864 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_42
timestamp 1604681595
transform 1 0 4968 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_50
timestamp 1604681595
transform 1 0 5704 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_44
timestamp 1604681595
transform 1 0 5152 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5152 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_60
timestamp 1604681595
transform 1 0 6624 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1604681595
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_53
timestamp 1604681595
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 6440 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_46
timestamp 1604681595
transform 1 0 5336 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_65
timestamp 1604681595
transform 1 0 7084 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 6900 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_34_82
timestamp 1604681595
transform 1 0 8648 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_77
timestamp 1604681595
transform 1 0 8188 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_83
timestamp 1604681595
transform 1 0 8740 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_79
timestamp 1604681595
transform 1 0 8372 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 8464 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 8556 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6900 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_34_88
timestamp 1604681595
transform 1 0 9200 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_91
timestamp 1604681595
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_87
timestamp 1604681595
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 8924 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9292 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_104
timestamp 1604681595
transform 1 0 10672 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1604681595
transform 1 0 9844 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_34_109
timestamp 1604681595
transform 1 0 11132 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_114
timestamp 1604681595
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1604681595
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_118
timestamp 1604681595
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 11868 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_132
timestamp 1604681595
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_136
timestamp 1604681595
transform 1 0 13616 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_144
timestamp 1604681595
transform 1 0 14352 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_133
timestamp 1604681595
transform 1 0 13340 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1604681595
transform 1 0 14444 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 14812 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 14812 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_9
timestamp 1604681595
transform 1 0 1932 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_13
timestamp 1604681595
transform 1 0 2300 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4784 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 4048 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 3680 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_25
timestamp 1604681595
transform 1 0 3404 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_30
timestamp 1604681595
transform 1 0 3864 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_34
timestamp 1604681595
transform 1 0 4232 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6256 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5888 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_49
timestamp 1604681595
transform 1 0 5612 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1604681595
transform 1 0 6072 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1604681595
transform 1 0 7452 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8464 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6992 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 8280 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_66
timestamp 1604681595
transform 1 0 7176 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_72
timestamp 1604681595
transform 1 0 7728 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 10212 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 10580 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_96
timestamp 1604681595
transform 1 0 9936 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_101
timestamp 1604681595
transform 1 0 10396 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_105
timestamp 1604681595
transform 1 0 10764 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_117
timestamp 1604681595
transform 1 0 11868 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_121
timestamp 1604681595
transform 1 0 12236 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_123
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_135
timestamp 1604681595
transform 1 0 13524 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_143
timestamp 1604681595
transform 1 0 14260 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 14812 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1604681595
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1604681595
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6256 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 5704 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 6072 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_48
timestamp 1604681595
transform 1 0 5520 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_52
timestamp 1604681595
transform 1 0 5888 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7452 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 7820 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_65
timestamp 1604681595
transform 1 0 7084 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_71
timestamp 1604681595
transform 1 0 7636 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_75
timestamp 1604681595
transform 1 0 8004 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 10212 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_87
timestamp 1604681595
transform 1 0 9108 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_91
timestamp 1604681595
transform 1 0 9476 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_93
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_115
timestamp 1604681595
transform 1 0 11684 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_127
timestamp 1604681595
transform 1 0 12788 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_139
timestamp 1604681595
transform 1 0 13892 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_145
timestamp 1604681595
transform 1 0 14444 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 14812 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_15
timestamp 1604681595
transform 1 0 2484 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4232 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 4048 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 3680 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 3312 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_23
timestamp 1604681595
transform 1 0 3220 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_26
timestamp 1604681595
transform 1 0 3496 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_30
timestamp 1604681595
transform 1 0 3864 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_50
timestamp 1604681595
transform 1 0 5704 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_54
timestamp 1604681595
transform 1 0 6072 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1604681595
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 8372 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_71
timestamp 1604681595
transform 1 0 7636 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_75
timestamp 1604681595
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_82
timestamp 1604681595
transform 1 0 8648 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 9752 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 8832 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 10212 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_86
timestamp 1604681595
transform 1 0 9016 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_97
timestamp 1604681595
transform 1 0 10028 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_101
timestamp 1604681595
transform 1 0 10396 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1604681595
transform 1 0 11500 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_121
timestamp 1604681595
transform 1 0 12236 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_123
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_135
timestamp 1604681595
transform 1 0 13524 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_143
timestamp 1604681595
transform 1 0 14260 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 14812 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1604681595
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 4784 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4324 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1604681595
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_32
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_37
timestamp 1604681595
transform 1 0 4508 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 5244 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_38_43
timestamp 1604681595
transform 1 0 5060 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_61
timestamp 1604681595
transform 1 0 6716 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7452 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 6900 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 7268 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 8464 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_65
timestamp 1604681595
transform 1 0 7084 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_78
timestamp 1604681595
transform 1 0 8280 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_82
timestamp 1604681595
transform 1 0 8648 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 9016 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9844 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_88
timestamp 1604681595
transform 1 0 9200 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1604681595
transform 1 0 10028 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1604681595
transform 1 0 11132 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1604681595
transform 1 0 12236 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_133
timestamp 1604681595
transform 1 0 13340 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_145
timestamp 1604681595
transform 1 0 14444 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 14812 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1604681595
transform 1 0 4784 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4324 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4140 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4324 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_27
timestamp 1604681595
transform 1 0 3588 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1604681595
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_32
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_37
timestamp 1604681595
transform 1 0 4508 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_43
timestamp 1604681595
transform 1 0 5060 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_49
timestamp 1604681595
transform 1 0 5612 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_44
timestamp 1604681595
transform 1 0 5152 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 5428 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 5796 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5796 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_60
timestamp 1604681595
transform 1 0 6624 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_57
timestamp 1604681595
transform 1 0 6348 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_53
timestamp 1604681595
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 6808 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7360 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 8464 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7176 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_78
timestamp 1604681595
transform 1 0 8280 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_82
timestamp 1604681595
transform 1 0 8648 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_64
timestamp 1604681595
transform 1 0 6992 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_88
timestamp 1604681595
transform 1 0 9200 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_84
timestamp 1604681595
transform 1 0 8832 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9016 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 8832 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9016 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_40_102
timestamp 1604681595
transform 1 0 10488 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_103
timestamp 1604681595
transform 1 0 10580 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_99
timestamp 1604681595
transform 1 0 10212 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_95
timestamp 1604681595
transform 1 0 9844 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10396 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10028 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_112
timestamp 1604681595
transform 1 0 11408 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_109
timestamp 1604681595
transform 1 0 11132 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 11224 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1604681595
transform 1 0 11224 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_39_120
timestamp 1604681595
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_116
timestamp 1604681595
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_119
timestamp 1604681595
transform 1 0 12052 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_135
timestamp 1604681595
transform 1 0 13524 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_143
timestamp 1604681595
transform 1 0 14260 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_131
timestamp 1604681595
transform 1 0 13156 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_143
timestamp 1604681595
transform 1 0 14260 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 14812 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 14812 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4784 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4600 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 4232 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3864 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_27
timestamp 1604681595
transform 1 0 3588 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_32
timestamp 1604681595
transform 1 0 4048 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_36
timestamp 1604681595
transform 1 0 4416 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 5796 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_49
timestamp 1604681595
transform 1 0 5612 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_53
timestamp 1604681595
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1604681595
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7544 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 7360 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8556 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6992 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_66
timestamp 1604681595
transform 1 0 7176 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_79
timestamp 1604681595
transform 1 0 8372 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_83
timestamp 1604681595
transform 1 0 8740 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9108 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8924 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_103
timestamp 1604681595
transform 1 0 10580 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_111
timestamp 1604681595
transform 1 0 11316 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_107
timestamp 1604681595
transform 1 0 10948 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11500 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11132 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_119
timestamp 1604681595
transform 1 0 12052 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_115
timestamp 1604681595
transform 1 0 11684 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11868 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_135
timestamp 1604681595
transform 1 0 13524 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_143
timestamp 1604681595
transform 1 0 14260 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 14812 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1604681595
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 4784 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604681595
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_38
timestamp 1604681595
transform 1 0 4600 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1604681595
transform 1 0 5704 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_42_42
timestamp 1604681595
transform 1 0 4968 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_59
timestamp 1604681595
transform 1 0 6532 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7820 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7544 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_67
timestamp 1604681595
transform 1 0 7268 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_72
timestamp 1604681595
transform 1 0 7728 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_82
timestamp 1604681595
transform 1 0 8648 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10672 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 9108 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_86
timestamp 1604681595
transform 1 0 9016 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_89
timestamp 1604681595
transform 1 0 9292 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_102
timestamp 1604681595
transform 1 0 10488 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11224 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11040 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_106
timestamp 1604681595
transform 1 0 10856 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_126
timestamp 1604681595
transform 1 0 12696 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_138
timestamp 1604681595
transform 1 0 13800 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 14812 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1604681595
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1604681595
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1604681595
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1604681595
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1604681595
transform 1 0 4692 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 6164 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1604681595
transform 1 0 5796 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_58
timestamp 1604681595
transform 1 0 6440 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_62
timestamp 1604681595
transform 1 0 6808 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 8464 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8280 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 6992 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_66
timestamp 1604681595
transform 1 0 7176 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_72
timestamp 1604681595
transform 1 0 7728 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_75
timestamp 1604681595
transform 1 0 8004 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_43_83
timestamp 1604681595
transform 1 0 8740 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8832 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10396 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10212 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9844 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_93
timestamp 1604681595
transform 1 0 9660 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_97
timestamp 1604681595
transform 1 0 10028 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 11960 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 11408 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 12604 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1604681595
transform 1 0 11224 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_114
timestamp 1604681595
transform 1 0 11592 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_120
timestamp 1604681595
transform 1 0 12144 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_123
timestamp 1604681595
transform 1 0 12420 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12972 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_127
timestamp 1604681595
transform 1 0 12788 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_131
timestamp 1604681595
transform 1 0 13156 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_143
timestamp 1604681595
transform 1 0 14260 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1604681595
transform -1 0 14812 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1604681595
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1604681595
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1604681595
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_27
timestamp 1604681595
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_32
timestamp 1604681595
transform 1 0 4048 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_40
timestamp 1604681595
transform 1 0 4784 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 5428 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4968 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_44
timestamp 1604681595
transform 1 0 5152 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_49
timestamp 1604681595
transform 1 0 5612 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_61
timestamp 1604681595
transform 1 0 6716 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 7176 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 7544 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 8464 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_65
timestamp 1604681595
transform 1 0 7084 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_68
timestamp 1604681595
transform 1 0 7360 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_72
timestamp 1604681595
transform 1 0 7728 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1604681595
transform 1 0 8648 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10396 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8832 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10212 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9200 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_86
timestamp 1604681595
transform 1 0 9016 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_90
timestamp 1604681595
transform 1 0 9384 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_93
timestamp 1604681595
transform 1 0 9660 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1604681595
transform 1 0 11960 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_44_110
timestamp 1604681595
transform 1 0 11224 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_127
timestamp 1604681595
transform 1 0 12788 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_139
timestamp 1604681595
transform 1 0 13892 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_145
timestamp 1604681595
transform 1 0 14444 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1604681595
transform -1 0 14812 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1604681595
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1604681595
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1604681595
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 4784 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4416 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4048 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_27
timestamp 1604681595
transform 1 0 3588 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_31
timestamp 1604681595
transform 1 0 3956 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_34
timestamp 1604681595
transform 1 0 4232 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_38
timestamp 1604681595
transform 1 0 4600 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4968 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 5980 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_51
timestamp 1604681595
transform 1 0 5796 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_55
timestamp 1604681595
transform 1 0 6164 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_62
timestamp 1604681595
transform 1 0 6808 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1604681595
transform 1 0 7176 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 6992 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 8188 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_75
timestamp 1604681595
transform 1 0 8004 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_79
timestamp 1604681595
transform 1 0 8372 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10580 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10396 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10028 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_91
timestamp 1604681595
transform 1 0 9476 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_99
timestamp 1604681595
transform 1 0 10212 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_112
timestamp 1604681595
transform 1 0 11408 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_120
timestamp 1604681595
transform 1 0 12144 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_123
timestamp 1604681595
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_135
timestamp 1604681595
transform 1 0 13524 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_143
timestamp 1604681595
transform 1 0 14260 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1604681595
transform -1 0 14812 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1604681595
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1604681595
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1604681595
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1604681595
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_9
timestamp 1604681595
transform 1 0 1932 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_13
timestamp 1604681595
transform 1 0 2300 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1604681595
transform 1 0 3588 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3404 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3588 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 4600 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1604681595
transform 1 0 3772 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_32
timestamp 1604681595
transform 1 0 4048 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_36
timestamp 1604681595
transform 1 0 4416 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_40
timestamp 1604681595
transform 1 0 4784 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_46
timestamp 1604681595
transform 1 0 5336 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 5152 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4968 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5428 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1604681595
transform 1 0 6348 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_53
timestamp 1604681595
transform 1 0 5980 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_56
timestamp 1604681595
transform 1 0 6256 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 6808 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 6164 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 6992 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 8464 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 8648 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_80
timestamp 1604681595
transform 1 0 8464 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_78
timestamp 1604681595
transform 1 0 8280 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_82
timestamp 1604681595
transform 1 0 8648 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_88
timestamp 1604681595
transform 1 0 9200 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_84
timestamp 1604681595
transform 1 0 8832 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 9016 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 8832 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1604681595
transform 1 0 9016 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1604681595
transform 1 0 9660 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_99
timestamp 1604681595
transform 1 0 10212 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_95
timestamp 1604681595
transform 1 0 9844 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_100
timestamp 1604681595
transform 1 0 10304 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_96
timestamp 1604681595
transform 1 0 9936 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 10120 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10580 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 10028 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_114
timestamp 1604681595
transform 1 0 11592 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_113
timestamp 1604681595
transform 1 0 11500 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_109
timestamp 1604681595
transform 1 0 11132 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_105
timestamp 1604681595
transform 1 0 10764 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11316 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 10948 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_120
timestamp 1604681595
transform 1 0 12144 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_120
timestamp 1604681595
transform 1 0 12144 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_117
timestamp 1604681595
transform 1 0 11868 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 12328 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 11960 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 11960 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1604681595
transform 1 0 12420 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_124
timestamp 1604681595
transform 1 0 12512 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_136
timestamp 1604681595
transform 1 0 13616 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_144
timestamp 1604681595
transform 1 0 14352 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_126
timestamp 1604681595
transform 1 0 12696 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_138
timestamp 1604681595
transform 1 0 13800 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1604681595
transform -1 0 14812 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1604681595
transform -1 0 14812 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1604681595
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1604681595
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1604681595
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4232 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3588 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 4600 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_29
timestamp 1604681595
transform 1 0 3772 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_32
timestamp 1604681595
transform 1 0 4048 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_36
timestamp 1604681595
transform 1 0 4416 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_40
timestamp 1604681595
transform 1 0 4784 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5428 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5152 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_46
timestamp 1604681595
transform 1 0 5336 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1604681595
transform 1 0 8004 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 7820 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_63
timestamp 1604681595
transform 1 0 6900 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_71
timestamp 1604681595
transform 1 0 7636 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 9016 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_84
timestamp 1604681595
transform 1 0 8832 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_88
timestamp 1604681595
transform 1 0 9200 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1604681595
transform 1 0 11960 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_48_109
timestamp 1604681595
transform 1 0 11132 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_117
timestamp 1604681595
transform 1 0 11868 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 12972 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_127
timestamp 1604681595
transform 1 0 12788 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_131
timestamp 1604681595
transform 1 0 13156 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_143
timestamp 1604681595
transform 1 0 14260 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1604681595
transform -1 0 14812 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1604681595
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1604681595
transform 1 0 1380 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_7
timestamp 1604681595
transform 1 0 1748 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_19
timestamp 1604681595
transform 1 0 2852 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 3680 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 3496 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 3128 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_24
timestamp 1604681595
transform 1 0 3312 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 5888 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 6256 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 5520 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_44
timestamp 1604681595
transform 1 0 5152 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_50
timestamp 1604681595
transform 1 0 5704 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1604681595
transform 1 0 6072 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_58
timestamp 1604681595
transform 1 0 6440 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_62
timestamp 1604681595
transform 1 0 6808 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1604681595
transform 1 0 8096 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 7912 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 7544 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_72
timestamp 1604681595
transform 1 0 7728 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10028 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9844 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 9476 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 9108 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_85
timestamp 1604681595
transform 1 0 8924 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_89
timestamp 1604681595
transform 1 0 9292 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_93
timestamp 1604681595
transform 1 0 9660 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 11776 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_113
timestamp 1604681595
transform 1 0 11500 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_118
timestamp 1604681595
transform 1 0 11960 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 13432 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 13800 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_132
timestamp 1604681595
transform 1 0 13248 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_136
timestamp 1604681595
transform 1 0 13616 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_140
timestamp 1604681595
transform 1 0 13984 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1604681595
transform -1 0 14812 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1604681595
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 2116 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_9
timestamp 1604681595
transform 1 0 1932 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_13
timestamp 1604681595
transform 1 0 2300 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4140 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 3312 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_21
timestamp 1604681595
transform 1 0 3036 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_26
timestamp 1604681595
transform 1 0 3496 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_32
timestamp 1604681595
transform 1 0 4048 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5888 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_50_42
timestamp 1604681595
transform 1 0 4968 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_50
timestamp 1604681595
transform 1 0 5704 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_61
timestamp 1604681595
transform 1 0 6716 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 8096 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 6900 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_65
timestamp 1604681595
transform 1 0 7084 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_73
timestamp 1604681595
transform 1 0 7820 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_78
timestamp 1604681595
transform 1 0 8280 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 9660 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_90
timestamp 1604681595
transform 1 0 9384 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 12328 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 11316 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_109
timestamp 1604681595
transform 1 0 11132 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_113
timestamp 1604681595
transform 1 0 11500 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_121
timestamp 1604681595
transform 1 0 12236 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_138
timestamp 1604681595
transform 1 0 13800 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1604681595
transform -1 0 14812 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1604681595
transform 1 0 1748 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1604681595
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 1564 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1604681595
transform 1 0 1380 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_16
timestamp 1604681595
transform 1 0 2576 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 3312 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 3128 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_40
timestamp 1604681595
transform 1 0 4784 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 5060 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 5428 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 5796 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_45
timestamp 1604681595
transform 1 0 5244 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_49
timestamp 1604681595
transform 1 0 5612 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_53
timestamp 1604681595
transform 1 0 5980 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_71
timestamp 1604681595
transform 1 0 7636 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_83
timestamp 1604681595
transform 1 0 8740 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 10580 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 10212 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_95
timestamp 1604681595
transform 1 0 9844 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_101
timestamp 1604681595
transform 1 0 10396 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 11776 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_114
timestamp 1604681595
transform 1 0 11592 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_118
timestamp 1604681595
transform 1 0 11960 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_132
timestamp 1604681595
transform 1 0 13248 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_136
timestamp 1604681595
transform 1 0 13616 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_144
timestamp 1604681595
transform 1 0 14352 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1604681595
transform -1 0 14812 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1604681595
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1604681595
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 1748 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_3
timestamp 1604681595
transform 1 0 1380 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_9
timestamp 1604681595
transform 1 0 1932 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1604681595
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1604681595
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_27
timestamp 1604681595
transform 1 0 3588 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_29
timestamp 1604681595
transform 1 0 3772 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_21
timestamp 1604681595
transform 1 0 3036 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_36
timestamp 1604681595
transform 1 0 4416 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_33
timestamp 1604681595
transform 1 0 4140 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_32
timestamp 1604681595
transform 1 0 4048 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 4232 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4784 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4600 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4784 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_53_49
timestamp 1604681595
transform 1 0 5612 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_42
timestamp 1604681595
transform 1 0 4968 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5060 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_59
timestamp 1604681595
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_55
timestamp 1604681595
transform 1 0 6164 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_60
timestamp 1604681595
transform 1 0 6624 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_52
timestamp 1604681595
transform 1 0 5888 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 5980 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 6348 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_62
timestamp 1604681595
transform 1 0 6808 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 6808 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_67
timestamp 1604681595
transform 1 0 7268 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_70
timestamp 1604681595
transform 1 0 7544 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_64
timestamp 1604681595
transform 1 0 6992 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 7084 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 7636 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 7452 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1604681595
transform 1 0 7636 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_80
timestamp 1604681595
transform 1 0 8464 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8648 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_73
timestamp 1604681595
transform 1 0 7820 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_84
timestamp 1604681595
transform 1 0 8832 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_93
timestamp 1604681595
transform 1 0 9660 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_90
timestamp 1604681595
transform 1 0 9384 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_85
timestamp 1604681595
transform 1 0 8924 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9200 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9016 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9200 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_97
timestamp 1604681595
transform 1 0 10028 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_97
timestamp 1604681595
transform 1 0 10028 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9844 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10212 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_101
timestamp 1604681595
transform 1 0 10396 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 11316 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 10764 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_107
timestamp 1604681595
transform 1 0 10948 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_113
timestamp 1604681595
transform 1 0 11500 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_121
timestamp 1604681595
transform 1 0 12236 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_123
timestamp 1604681595
transform 1 0 12420 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 12972 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_127
timestamp 1604681595
transform 1 0 12788 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_131
timestamp 1604681595
transform 1 0 13156 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_143
timestamp 1604681595
transform 1 0 14260 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_135
timestamp 1604681595
transform 1 0 13524 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_143
timestamp 1604681595
transform 1 0 14260 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1604681595
transform -1 0 14812 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1604681595
transform -1 0 14812 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1604681595
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1604681595
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1604681595
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1604681595
transform 1 0 4876 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_27
timestamp 1604681595
transform 1 0 3588 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_32
timestamp 1604681595
transform 1 0 4048 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_40
timestamp 1604681595
transform 1 0 4784 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6348 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 5336 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_44
timestamp 1604681595
transform 1 0 5152 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_48
timestamp 1604681595
transform 1 0 5520 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_56
timestamp 1604681595
transform 1 0 6256 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1604681595
transform 1 0 8556 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 8004 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_73
timestamp 1604681595
transform 1 0 7820 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_77
timestamp 1604681595
transform 1 0 8188 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10672 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 9016 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_84
timestamp 1604681595
transform 1 0 8832 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_88
timestamp 1604681595
transform 1 0 9200 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_102
timestamp 1604681595
transform 1 0 10488 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 11040 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_106
timestamp 1604681595
transform 1 0 10856 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_110
timestamp 1604681595
transform 1 0 11224 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_122
timestamp 1604681595
transform 1 0 12328 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_134
timestamp 1604681595
transform 1 0 13432 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1604681595
transform -1 0 14812 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1604681595
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1604681595
transform 1 0 1380 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_7
timestamp 1604681595
transform 1 0 1748 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_19
timestamp 1604681595
transform 1 0 2852 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604681595
transform 1 0 4048 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_31
timestamp 1604681595
transform 1 0 3956 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_34
timestamp 1604681595
transform 1 0 4232 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_40
timestamp 1604681595
transform 1 0 4784 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 6164 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4968 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_53
timestamp 1604681595
transform 1 0 5980 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_57
timestamp 1604681595
transform 1 0 6348 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_62
timestamp 1604681595
transform 1 0 6808 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7176 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1604681595
transform 1 0 8740 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6992 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 8188 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 8556 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_75
timestamp 1604681595
transform 1 0 8004 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_79
timestamp 1604681595
transform 1 0 8372 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10304 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10120 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9752 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_92
timestamp 1604681595
transform 1 0 9568 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_96
timestamp 1604681595
transform 1 0 9936 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 11316 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_109
timestamp 1604681595
transform 1 0 11132 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_113
timestamp 1604681595
transform 1 0 11500 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_121
timestamp 1604681595
transform 1 0 12236 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_123
timestamp 1604681595
transform 1 0 12420 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_135
timestamp 1604681595
transform 1 0 13524 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_143
timestamp 1604681595
transform 1 0 14260 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1604681595
transform -1 0 14812 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1604681595
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_9
timestamp 1604681595
transform 1 0 1932 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 4048 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_21
timestamp 1604681595
transform 1 0 3036 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_29
timestamp 1604681595
transform 1 0 3772 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_36
timestamp 1604681595
transform 1 0 4416 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5336 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5152 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_62
timestamp 1604681595
transform 1 0 6808 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1604681595
transform 1 0 7728 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 7176 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 8740 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_68
timestamp 1604681595
transform 1 0 7360 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_81
timestamp 1604681595
transform 1 0 8556 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10212 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 9108 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 10028 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_85
timestamp 1604681595
transform 1 0 8924 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_89
timestamp 1604681595
transform 1 0 9292 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_93
timestamp 1604681595
transform 1 0 9660 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 12420 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 11960 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_115
timestamp 1604681595
transform 1 0 11684 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_120
timestamp 1604681595
transform 1 0 12144 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_125
timestamp 1604681595
transform 1 0 12604 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 12788 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_129
timestamp 1604681595
transform 1 0 12972 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_141
timestamp 1604681595
transform 1 0 14076 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_145
timestamp 1604681595
transform 1 0 14444 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1604681595
transform -1 0 14812 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 1380 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1604681595
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 1932 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604681595
transform 1 0 2668 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2300 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_7
timestamp 1604681595
transform 1 0 1748 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_11
timestamp 1604681595
transform 1 0 2116 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_15
timestamp 1604681595
transform 1 0 2484 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_19
timestamp 1604681595
transform 1 0 2852 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4140 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604681595
transform 1 0 3956 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 3588 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 3220 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_25
timestamp 1604681595
transform 1 0 3404 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_29
timestamp 1604681595
transform 1 0 3772 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 5796 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_49
timestamp 1604681595
transform 1 0 5612 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_53
timestamp 1604681595
transform 1 0 5980 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_57
timestamp 1604681595
transform 1 0 6348 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 7820 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 8740 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 8188 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_71
timestamp 1604681595
transform 1 0 7636 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_75
timestamp 1604681595
transform 1 0 8004 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_79
timestamp 1604681595
transform 1 0 8372 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1604681595
transform 1 0 9292 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 9108 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 10396 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_85
timestamp 1604681595
transform 1 0 8924 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_98
timestamp 1604681595
transform 1 0 10120 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_103
timestamp 1604681595
transform 1 0 10580 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_111
timestamp 1604681595
transform 1 0 11316 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_107
timestamp 1604681595
transform 1 0 10948 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 10764 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1604681595
transform 1 0 11040 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_118
timestamp 1604681595
transform 1 0 11960 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_115
timestamp 1604681595
transform 1 0 11684 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 11776 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 13432 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_132
timestamp 1604681595
transform 1 0 13248 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_136
timestamp 1604681595
transform 1 0 13616 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_144
timestamp 1604681595
transform 1 0 14352 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1604681595
transform -1 0 14812 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 2668 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1604681595
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_9
timestamp 1604681595
transform 1 0 1932 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 4048 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_21
timestamp 1604681595
transform 1 0 3036 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_29
timestamp 1604681595
transform 1 0 3772 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_36
timestamp 1604681595
transform 1 0 4416 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5520 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5336 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6808 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_44
timestamp 1604681595
transform 1 0 5152 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_57
timestamp 1604681595
transform 1 0 6348 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_61
timestamp 1604681595
transform 1 0 6716 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 7360 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7176 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_64
timestamp 1604681595
transform 1 0 6992 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_93
timestamp 1604681595
transform 1 0 9660 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_91
timestamp 1604681595
transform 1 0 9476 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_88
timestamp 1604681595
transform 1 0 9200 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_84
timestamp 1604681595
transform 1 0 8832 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 9292 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_97
timestamp 1604681595
transform 1 0 10028 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 10212 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9844 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1604681595
transform 1 0 10396 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1604681595
transform 1 0 11960 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_58_110
timestamp 1604681595
transform 1 0 11224 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_127
timestamp 1604681595
transform 1 0 12788 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_139
timestamp 1604681595
transform 1 0 13892 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_145
timestamp 1604681595
transform 1 0 14444 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1604681595
transform -1 0 14812 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_7
timestamp 1604681595
transform 1 0 1748 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_9
timestamp 1604681595
transform 1 0 1932 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1932 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1604681595
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1604681595
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 1380 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_11
timestamp 1604681595
transform 1 0 2116 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_17
timestamp 1604681595
transform 1 0 2668 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_13
timestamp 1604681595
transform 1 0 2300 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 2484 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 2116 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 2484 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_19
timestamp 1604681595
transform 1 0 2852 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_29
timestamp 1604681595
transform 1 0 3772 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_25
timestamp 1604681595
transform 1 0 3404 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 3588 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 3036 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_36
timestamp 1604681595
transform 1 0 4416 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_37
timestamp 1604681595
transform 1 0 4508 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604681595
transform 1 0 3956 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 4140 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 4048 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_41
timestamp 1604681595
transform 1 0 4876 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604681595
transform 1 0 4692 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_51
timestamp 1604681595
transform 1 0 5796 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_44
timestamp 1604681595
transform 1 0 5152 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_49
timestamp 1604681595
transform 1 0 5612 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604681595
transform 1 0 5060 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1604681595
transform 1 0 5796 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 5244 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604681595
transform 1 0 5428 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_57
timestamp 1604681595
transform 1 0 6348 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_53
timestamp 1604681595
transform 1 0 5980 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1604681595
transform 1 0 6532 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_59_62
timestamp 1604681595
transform 1 0 6808 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604681595
transform 1 0 8096 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7636 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1604681595
transform 1 0 7452 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 7636 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 6992 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_66
timestamp 1604681595
transform 1 0 7176 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_68
timestamp 1604681595
transform 1 0 7360 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_73
timestamp 1604681595
transform 1 0 7820 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_80
timestamp 1604681595
transform 1 0 8464 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9844 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9660 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9292 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 10672 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_87
timestamp 1604681595
transform 1 0 9108 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_91
timestamp 1604681595
transform 1 0 9476 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_102
timestamp 1604681595
transform 1 0 10488 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_111
timestamp 1604681595
transform 1 0 11316 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_119
timestamp 1604681595
transform 1 0 12052 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_123
timestamp 1604681595
transform 1 0 12420 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_106
timestamp 1604681595
transform 1 0 10856 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_118
timestamp 1604681595
transform 1 0 11960 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_135
timestamp 1604681595
transform 1 0 13524 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_143
timestamp 1604681595
transform 1 0 14260 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_130
timestamp 1604681595
transform 1 0 13064 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_142
timestamp 1604681595
transform 1 0 14168 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1604681595
transform -1 0 14812 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1604681595
transform -1 0 14812 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1604681595
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1604681595
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1604681595
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604681595
transform 1 0 4508 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1604681595
transform 1 0 4324 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_27
timestamp 1604681595
transform 1 0 3588 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_41
timestamp 1604681595
transform 1 0 4876 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604681595
transform 1 0 5612 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1604681595
transform 1 0 5060 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1604681595
transform 1 0 6164 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1604681595
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_45
timestamp 1604681595
transform 1 0 5244 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_53
timestamp 1604681595
transform 1 0 5980 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_57
timestamp 1604681595
transform 1 0 6348 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_62
timestamp 1604681595
transform 1 0 6808 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1604681595
transform 1 0 8188 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604681595
transform 1 0 7084 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1604681595
transform 1 0 7636 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1604681595
transform 1 0 8740 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 8004 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_69
timestamp 1604681595
transform 1 0 7452 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_73
timestamp 1604681595
transform 1 0 7820 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_81
timestamp 1604681595
transform 1 0 8556 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 9660 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 10212 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_85
timestamp 1604681595
transform 1 0 8924 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_97
timestamp 1604681595
transform 1 0 10028 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_101
timestamp 1604681595
transform 1 0 10396 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_113
timestamp 1604681595
transform 1 0 11500 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_121
timestamp 1604681595
transform 1 0 12236 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_123
timestamp 1604681595
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_135
timestamp 1604681595
transform 1 0 13524 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_143
timestamp 1604681595
transform 1 0 14260 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1604681595
transform -1 0 14812 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1604681595
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1604681595
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1604681595
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604681595
transform 1 0 4784 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_27
timestamp 1604681595
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_32
timestamp 1604681595
transform 1 0 4048 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1604681595
transform 1 0 6348 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_44
timestamp 1604681595
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_56
timestamp 1604681595
transform 1 0 6256 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_61
timestamp 1604681595
transform 1 0 6716 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_73
timestamp 1604681595
transform 1 0 7820 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_85
timestamp 1604681595
transform 1 0 8924 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_91
timestamp 1604681595
transform 1 0 9476 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_93
timestamp 1604681595
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_105
timestamp 1604681595
transform 1 0 10764 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_117
timestamp 1604681595
transform 1 0 11868 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_129
timestamp 1604681595
transform 1 0 12972 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_141
timestamp 1604681595
transform 1 0 14076 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_145
timestamp 1604681595
transform 1 0 14444 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1604681595
transform -1 0 14812 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1604681595
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1604681595
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1604681595
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604681595
transform 1 0 4600 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_27
timestamp 1604681595
transform 1 0 3588 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_35
timestamp 1604681595
transform 1 0 4324 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1604681595
transform 1 0 5152 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_42
timestamp 1604681595
transform 1 0 4968 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_46
timestamp 1604681595
transform 1 0 5336 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_58
timestamp 1604681595
transform 1 0 6440 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_62
timestamp 1604681595
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_74
timestamp 1604681595
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_86
timestamp 1604681595
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_98
timestamp 1604681595
transform 1 0 10120 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_110
timestamp 1604681595
transform 1 0 11224 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_123
timestamp 1604681595
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_135
timestamp 1604681595
transform 1 0 13524 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_143
timestamp 1604681595
transform 1 0 14260 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1604681595
transform -1 0 14812 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1604681595
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1604681595
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1604681595
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_27
timestamp 1604681595
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_32
timestamp 1604681595
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_44
timestamp 1604681595
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_56
timestamp 1604681595
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_63
timestamp 1604681595
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_75
timestamp 1604681595
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_87
timestamp 1604681595
transform 1 0 9108 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_94
timestamp 1604681595
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_106
timestamp 1604681595
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_118
timestamp 1604681595
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_125
timestamp 1604681595
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_137
timestamp 1604681595
transform 1 0 13708 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_145
timestamp 1604681595
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1604681595
transform -1 0 14812 0 -1 37536
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 1096 480 1216 6 ccff_head
port 0 nsew default input
rlabel metal3 s 15520 29928 16000 30048 6 ccff_tail
port 1 nsew default tristate
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[0]
port 2 nsew default input
rlabel metal2 s 12162 0 12218 480 6 chany_bottom_in[10]
port 3 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[11]
port 4 nsew default input
rlabel metal2 s 12990 0 13046 480 6 chany_bottom_in[12]
port 5 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[13]
port 6 nsew default input
rlabel metal2 s 13726 0 13782 480 6 chany_bottom_in[14]
port 7 nsew default input
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_in[15]
port 8 nsew default input
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_in[16]
port 9 nsew default input
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_in[17]
port 10 nsew default input
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_in[18]
port 11 nsew default input
rlabel metal2 s 15750 0 15806 480 6 chany_bottom_in[19]
port 12 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[1]
port 13 nsew default input
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_in[2]
port 14 nsew default input
rlabel metal2 s 9402 0 9458 480 6 chany_bottom_in[3]
port 15 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[4]
port 16 nsew default input
rlabel metal2 s 10138 0 10194 480 6 chany_bottom_in[5]
port 17 nsew default input
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_in[6]
port 18 nsew default input
rlabel metal2 s 10966 0 11022 480 6 chany_bottom_in[7]
port 19 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[8]
port 20 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_in[9]
port 21 nsew default input
rlabel metal2 s 202 0 258 480 6 chany_bottom_out[0]
port 22 nsew default tristate
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_out[10]
port 23 nsew default tristate
rlabel metal2 s 4526 0 4582 480 6 chany_bottom_out[11]
port 24 nsew default tristate
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_out[12]
port 25 nsew default tristate
rlabel metal2 s 5354 0 5410 480 6 chany_bottom_out[13]
port 26 nsew default tristate
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_out[14]
port 27 nsew default tristate
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_out[15]
port 28 nsew default tristate
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_out[16]
port 29 nsew default tristate
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_out[17]
port 30 nsew default tristate
rlabel metal2 s 7378 0 7434 480 6 chany_bottom_out[18]
port 31 nsew default tristate
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_out[19]
port 32 nsew default tristate
rlabel metal2 s 570 0 626 480 6 chany_bottom_out[1]
port 33 nsew default tristate
rlabel metal2 s 938 0 994 480 6 chany_bottom_out[2]
port 34 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_out[3]
port 35 nsew default tristate
rlabel metal2 s 1766 0 1822 480 6 chany_bottom_out[4]
port 36 nsew default tristate
rlabel metal2 s 2134 0 2190 480 6 chany_bottom_out[5]
port 37 nsew default tristate
rlabel metal2 s 2594 0 2650 480 6 chany_bottom_out[6]
port 38 nsew default tristate
rlabel metal2 s 2962 0 3018 480 6 chany_bottom_out[7]
port 39 nsew default tristate
rlabel metal2 s 3330 0 3386 480 6 chany_bottom_out[8]
port 40 nsew default tristate
rlabel metal2 s 3790 0 3846 480 6 chany_bottom_out[9]
port 41 nsew default tristate
rlabel metal2 s 8206 39520 8262 40000 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 12162 39520 12218 40000 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 12530 39520 12586 40000 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 12990 39520 13046 40000 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 13358 39520 13414 40000 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 13726 39520 13782 40000 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 14186 39520 14242 40000 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 14554 39520 14610 40000 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 14922 39520 14978 40000 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 15382 39520 15438 40000 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 15750 39520 15806 40000 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 8574 39520 8630 40000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 8942 39520 8998 40000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 9402 39520 9458 40000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 9770 39520 9826 40000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 10138 39520 10194 40000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 10598 39520 10654 40000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 10966 39520 11022 40000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 11334 39520 11390 40000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 11794 39520 11850 40000 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 202 39520 258 40000 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 4158 39520 4214 40000 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 4526 39520 4582 40000 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 4986 39520 5042 40000 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 5354 39520 5410 40000 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 5722 39520 5778 40000 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 6182 39520 6238 40000 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 6550 39520 6606 40000 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 6918 39520 6974 40000 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 7378 39520 7434 40000 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 7746 39520 7802 40000 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 570 39520 626 40000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 938 39520 994 40000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 1398 39520 1454 40000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 1766 39520 1822 40000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 2134 39520 2190 40000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 2594 39520 2650 40000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 2962 39520 3018 40000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 3330 39520 3386 40000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 3790 39520 3846 40000 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 3408 480 3528 6 left_grid_pin_16_
port 82 nsew default tristate
rlabel metal3 s 0 5720 480 5840 6 left_grid_pin_17_
port 83 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 left_grid_pin_18_
port 84 nsew default tristate
rlabel metal3 s 0 10480 480 10600 6 left_grid_pin_19_
port 85 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 left_grid_pin_20_
port 86 nsew default tristate
rlabel metal3 s 0 15104 480 15224 6 left_grid_pin_21_
port 87 nsew default tristate
rlabel metal3 s 0 17552 480 17672 6 left_grid_pin_22_
port 88 nsew default tristate
rlabel metal3 s 0 19864 480 19984 6 left_grid_pin_23_
port 89 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 left_grid_pin_24_
port 90 nsew default tristate
rlabel metal3 s 0 24488 480 24608 6 left_grid_pin_25_
port 91 nsew default tristate
rlabel metal3 s 0 26936 480 27056 6 left_grid_pin_26_
port 92 nsew default tristate
rlabel metal3 s 0 29248 480 29368 6 left_grid_pin_27_
port 93 nsew default tristate
rlabel metal3 s 0 31560 480 31680 6 left_grid_pin_28_
port 94 nsew default tristate
rlabel metal3 s 0 34008 480 34128 6 left_grid_pin_29_
port 95 nsew default tristate
rlabel metal3 s 0 36320 480 36440 6 left_grid_pin_30_
port 96 nsew default tristate
rlabel metal3 s 0 38632 480 38752 6 left_grid_pin_31_
port 97 nsew default tristate
rlabel metal3 s 15520 9936 16000 10056 6 prog_clk
port 98 nsew default input
rlabel metal4 s 3611 2128 3931 37584 6 VPWR
port 99 nsew default input
rlabel metal4 s 6277 2128 6597 37584 6 VGND
port 100 nsew default input
<< properties >>
string FIXED_BBOX 0 0 16000 40000
<< end >>
