* NGSPICE file created from sb_0__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

.subckt sb_0__1_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_left_grid_pin_11_ bottom_left_grid_pin_13_ bottom_left_grid_pin_15_
+ bottom_left_grid_pin_1_ bottom_left_grid_pin_3_ bottom_left_grid_pin_5_ bottom_left_grid_pin_7_
+ bottom_left_grid_pin_9_ bottom_right_grid_pin_11_ chanx_right_in[0] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chany_bottom_in[0] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_out[0] chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3]
+ chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7]
+ chany_bottom_out[8] chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_out[0] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] data_in enable
+ right_bottom_grid_pin_12_ right_top_grid_pin_10_ top_left_grid_pin_11_ top_left_grid_pin_13_
+ top_left_grid_pin_15_ top_left_grid_pin_1_ top_left_grid_pin_3_ top_left_grid_pin_5_
+ top_left_grid_pin_7_ top_left_grid_pin_9_ top_right_grid_pin_11_ vpwr vgnd
XFILLER_39_222 vpwr vgnd scs8hd_fill_2
Xmem_right_track_12.LATCH_1_.latch data_in _181_/A _167_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_100 vpwr vgnd scs8hd_fill_2
XFILLER_7_7 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_115 vgnd vpwr scs8hd_fill_1
XFILLER_9_126 vpwr vgnd scs8hd_fill_2
XFILLER_9_137 vgnd vpwr scs8hd_decap_4
XFILLER_13_155 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__113__B _109_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_3_ mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_129 vpwr vgnd scs8hd_fill_2
XFILLER_6_118 vgnd vpwr scs8hd_decap_8
XFILLER_6_107 vgnd vpwr scs8hd_decap_8
XFILLER_12_32 vpwr vgnd scs8hd_fill_2
XANTENNA__214__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _181_/A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_247 vgnd vpwr scs8hd_decap_12
XANTENNA__108__B _109_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_95 vpwr vgnd scs8hd_fill_2
XFILLER_5_140 vgnd vpwr scs8hd_decap_12
XANTENNA__124__A _101_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _194_/HI _176_/Y mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_184 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _188_/HI mem_bottom_track_17.LATCH_2_.latch/Q
+ mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_200_ _200_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA__209__A _209_/A vgnd vpwr scs8hd_diode_2
X_131_ _110_/A _131_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
XFILLER_2_154 vgnd vpwr scs8hd_decap_12
XFILLER_9_22 vgnd vpwr scs8hd_decap_12
XANTENNA__119__A _108_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_2_.latch data_in mem_bottom_track_17.LATCH_2_.latch/Q _151_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _213_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_242 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_53 vpwr vgnd scs8hd_fill_2
XFILLER_34_96 vgnd vpwr scs8hd_decap_3
XFILLER_34_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB _095_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_257 vgnd vpwr scs8hd_decap_12
X_114_ address[4] _135_/B vgnd vpwr scs8hd_inv_8
XFILLER_38_106 vpwr vgnd scs8hd_fill_2
XANTENNA__121__B _121_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_6_.scs8hd_inv_1 bottom_left_grid_pin_7_ mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_track_0.LATCH_4_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_37_161 vpwr vgnd scs8hd_fill_2
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XFILLER_20_21 vpwr vgnd scs8hd_fill_2
XANTENNA__222__A _222_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[6] mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_56 vgnd vpwr scs8hd_decap_12
XANTENNA__132__A _111_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_109 vpwr vgnd scs8hd_fill_2
XFILLER_34_186 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_1_.latch data_in _183_/A _169_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_208 vgnd vpwr scs8hd_decap_12
XFILLER_25_175 vpwr vgnd scs8hd_fill_2
XFILLER_15_21 vpwr vgnd scs8hd_fill_2
XFILLER_40_178 vgnd vpwr scs8hd_decap_12
XFILLER_40_145 vgnd vpwr scs8hd_decap_8
XFILLER_31_53 vpwr vgnd scs8hd_fill_2
XANTENNA__217__A _217_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_98 vpwr vgnd scs8hd_fill_2
XFILLER_31_75 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ _178_/A mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_0_230 vgnd vpwr scs8hd_decap_4
XFILLER_0_263 vgnd vpwr scs8hd_decap_12
XFILLER_31_123 vgnd vpwr scs8hd_decap_3
XFILLER_16_186 vpwr vgnd scs8hd_fill_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__A _154_/A vgnd vpwr scs8hd_diode_2
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _180_/Y vgnd
+ vpwr scs8hd_diode_2
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _188_/HI vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _191_/HI _182_/Y mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_112 vpwr vgnd scs8hd_fill_2
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_13_178 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _195_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_27_259 vpwr vgnd scs8hd_fill_2
XFILLER_18_259 vgnd vpwr scs8hd_decap_12
XFILLER_26_270 vgnd vpwr scs8hd_decap_4
XFILLER_5_196 vgnd vpwr scs8hd_decap_12
XFILLER_5_152 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__124__B _121_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _109_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_24_218 vgnd vpwr scs8hd_decap_12
X_130_ _109_/A _131_/B _130_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_10 vgnd vpwr scs8hd_decap_4
XANTENNA__225__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_23_65 vgnd vpwr scs8hd_decap_4
XFILLER_2_166 vgnd vpwr scs8hd_decap_12
XANTENNA__119__B _121_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_34 vgnd vpwr scs8hd_decap_3
XFILLER_9_56 vpwr vgnd scs8hd_fill_2
XFILLER_14_251 vgnd vpwr scs8hd_decap_12
XANTENNA__135__A _135_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A top_left_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_113_ _101_/B _109_/B _113_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_86 vgnd vpwr scs8hd_decap_6
XFILLER_34_64 vpwr vgnd scs8hd_fill_2
XFILLER_7_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _182_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _186_/A mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_184 vgnd vpwr scs8hd_decap_4
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XFILLER_20_88 vpwr vgnd scs8hd_fill_2
XFILLER_29_97 vpwr vgnd scs8hd_fill_2
XFILLER_29_53 vpwr vgnd scs8hd_fill_2
XFILLER_6_68 vgnd vpwr scs8hd_decap_12
XANTENNA__132__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_140 vgnd vpwr scs8hd_decap_3
XFILLER_19_162 vpwr vgnd scs8hd_fill_2
XFILLER_34_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_102 vgnd vpwr scs8hd_decap_3
XFILLER_25_198 vpwr vgnd scs8hd_fill_2
XFILLER_25_132 vpwr vgnd scs8hd_fill_2
XFILLER_0_275 vpwr vgnd scs8hd_fill_2
XFILLER_31_179 vpwr vgnd scs8hd_fill_2
XFILLER_31_168 vpwr vgnd scs8hd_fill_2
XFILLER_31_135 vpwr vgnd scs8hd_fill_2
XFILLER_31_113 vgnd vpwr scs8hd_decap_8
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_165 vpwr vgnd scs8hd_fill_2
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__B _168_/B vgnd vpwr scs8hd_diode_2
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A _152_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _173_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _180_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.INVTX1_2_.scs8hd_inv_1_A right_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A bottom_left_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _209_/A vgnd vpwr scs8hd_inv_1
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XANTENNA__138__A _137_/X vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_138 vgnd vpwr scs8hd_decap_4
XFILLER_10_149 vgnd vpwr scs8hd_decap_4
XFILLER_12_12 vpwr vgnd scs8hd_fill_2
XFILLER_12_23 vgnd vpwr scs8hd_decap_4
XFILLER_12_67 vgnd vpwr scs8hd_decap_6
XFILLER_37_75 vgnd vpwr scs8hd_fill_1
XFILLER_37_53 vpwr vgnd scs8hd_fill_2
XFILLER_5_164 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__140__B _141_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_274 vgnd vpwr scs8hd_fill_1
XFILLER_32_230 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_208 vgnd vpwr scs8hd_decap_12
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_99 vgnd vpwr scs8hd_fill_1
XFILLER_2_178 vgnd vpwr scs8hd_decap_12
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_263 vgnd vpwr scs8hd_decap_12
X_189_ _189_/HI _189_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr
+ scs8hd_diode_2
XANTENNA__135__B _135_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_6
XANTENNA__151__A _111_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_88 vpwr vgnd scs8hd_fill_2
X_112_ _152_/A _109_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_119 vgnd vpwr scs8hd_decap_4
XANTENNA__146__A _160_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _175_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _173_/A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_29_10 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_5_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_45 vpwr vgnd scs8hd_fill_2
XFILLER_28_152 vgnd vpwr scs8hd_fill_1
XFILLER_40_114 vgnd vpwr scs8hd_decap_8
XFILLER_15_78 vgnd vpwr scs8hd_decap_3
XFILLER_31_88 vpwr vgnd scs8hd_fill_2
XFILLER_31_22 vpwr vgnd scs8hd_fill_2
XFILLER_31_11 vgnd vpwr scs8hd_decap_3
XFILLER_0_243 vgnd vpwr scs8hd_decap_4
XFILLER_16_122 vpwr vgnd scs8hd_fill_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_199 vpwr vgnd scs8hd_fill_2
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__C _170_/C vgnd vpwr scs8hd_diode_2
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__143__B _141_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_269 vgnd vpwr scs8hd_decap_8
XFILLER_39_214 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_22_136 vgnd vpwr scs8hd_decap_4
XFILLER_22_147 vgnd vpwr scs8hd_decap_6
XFILLER_22_169 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_4.LATCH_1_.latch data_in _175_/A _161_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_26_88 vpwr vgnd scs8hd_fill_2
XFILLER_26_77 vpwr vgnd scs8hd_fill_2
XFILLER_9_107 vpwr vgnd scs8hd_fill_2
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_21_180 vgnd vpwr scs8hd_fill_1
Xmux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _177_/Y mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_3_59 vpwr vgnd scs8hd_fill_2
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_4_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__154__A _154_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_140 vgnd vpwr scs8hd_decap_12
XFILLER_27_206 vpwr vgnd scs8hd_fill_2
Xmux_right_track_14.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_46 vpwr vgnd scs8hd_fill_2
XFILLER_18_206 vgnd vpwr scs8hd_decap_8
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_43 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_121 vgnd vpwr scs8hd_fill_1
Xmem_top_track_0.LATCH_0_.latch data_in mem_top_track_0.LATCH_0_.latch/Q _101_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_176 vgnd vpwr scs8hd_decap_6
XANTENNA__149__A _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_242 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_3_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_34 vpwr vgnd scs8hd_fill_2
XFILLER_2_102 vpwr vgnd scs8hd_fill_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XFILLER_0_38 vpwr vgnd scs8hd_fill_2
XFILLER_0_49 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_9_69 vgnd vpwr scs8hd_decap_4
X_188_ _188_/HI _188_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__135__C _135_/C vgnd vpwr scs8hd_diode_2
XANTENNA__151__B _152_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _179_/A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _193_/HI _174_/Y mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_23 vpwr vgnd scs8hd_fill_2
X_111_ _111_/A _109_/B _111_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__146__B _146_/B vgnd vpwr scs8hd_diode_2
XANTENNA__162__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_131 vpwr vgnd scs8hd_fill_2
XFILLER_37_197 vgnd vpwr scs8hd_decap_12
XFILLER_1_92 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_13 vpwr vgnd scs8hd_fill_2
XFILLER_29_22 vgnd vpwr scs8hd_decap_3
XFILLER_20_68 vgnd vpwr scs8hd_fill_1
XFILLER_29_66 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _196_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XFILLER_34_178 vgnd vpwr scs8hd_fill_1
XFILLER_34_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_175 vpwr vgnd scs8hd_fill_2
XFILLER_19_197 vpwr vgnd scs8hd_fill_2
XANTENNA__157__A _154_/X vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_2_.latch data_in mem_bottom_track_1.LATCH_2_.latch/Q _132_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _192_/HI _185_/Y mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB _110_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_156 vpwr vgnd scs8hd_fill_2
XFILLER_15_13 vpwr vgnd scs8hd_fill_2
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_200 vpwr vgnd scs8hd_fill_2
XFILLER_16_145 vgnd vpwr scs8hd_decap_4
XFILLER_31_148 vgnd vpwr scs8hd_decap_6
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_226 vgnd vpwr scs8hd_decap_12
XFILLER_11_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_115 vpwr vgnd scs8hd_fill_2
XFILLER_30_192 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_23 vpwr vgnd scs8hd_fill_2
XFILLER_26_12 vpwr vgnd scs8hd_fill_2
XFILLER_13_104 vpwr vgnd scs8hd_fill_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_13_159 vpwr vgnd scs8hd_fill_2
XFILLER_21_170 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_27 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ _176_/A mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_8_152 vgnd vpwr scs8hd_fill_1
XANTENNA__170__A _160_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_36 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__080__A enable vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_218 vgnd vpwr scs8hd_decap_12
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
Xmux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _190_/HI _180_/Y mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__149__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XFILLER_32_254 vgnd vpwr scs8hd_decap_12
XANTENNA__165__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_210 vgnd vpwr scs8hd_decap_8
XFILLER_23_221 vpwr vgnd scs8hd_fill_2
XFILLER_23_243 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__075__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.INVTX1_0_.scs8hd_inv_1 chany_top_in[6] mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_210 vgnd vpwr scs8hd_decap_4
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ _187_/HI _187_/LO vgnd vpwr scs8hd_conb_1
Xmux_bottom_track_9.INVTX1_3_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _184_/Y mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_18_57 vgnd vpwr scs8hd_decap_4
X_110_ _110_/A _109_/B _110_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_45 vgnd vpwr scs8hd_decap_8
XFILLER_34_23 vgnd vpwr scs8hd_decap_8
XFILLER_11_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _179_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__146__C _161_/C vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XANTENNA__162__B _161_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_165 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.INVTX1_4_.scs8hd_inv_1 chanx_right_in[3] mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_25 vgnd vpwr scs8hd_decap_4
XFILLER_28_154 vgnd vpwr scs8hd_decap_6
XFILLER_28_121 vpwr vgnd scs8hd_fill_2
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_19_132 vpwr vgnd scs8hd_fill_2
XANTENNA__157__B _161_/B vgnd vpwr scs8hd_diode_2
XANTENNA__173__A _173_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_113 vpwr vgnd scs8hd_fill_2
XFILLER_31_35 vpwr vgnd scs8hd_fill_2
XFILLER_25_179 vpwr vgnd scs8hd_fill_2
XANTENNA__083__A _154_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_25 vpwr vgnd scs8hd_fill_2
XFILLER_15_36 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ _182_/A mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_31_57 vpwr vgnd scs8hd_fill_2
XFILLER_0_234 vgnd vpwr scs8hd_fill_1
XFILLER_31_105 vpwr vgnd scs8hd_fill_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_205 vgnd vpwr scs8hd_fill_1
XFILLER_39_238 vgnd vpwr scs8hd_decap_6
XANTENNA__168__A _154_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_92 vpwr vgnd scs8hd_fill_2
XFILLER_7_70 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_1_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__078__A _077_/X vgnd vpwr scs8hd_diode_2
XFILLER_13_116 vpwr vgnd scs8hd_fill_2
XFILLER_13_138 vpwr vgnd scs8hd_fill_2
XFILLER_13_149 vgnd vpwr scs8hd_decap_4
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_193 vpwr vgnd scs8hd_fill_2
XFILLER_3_39 vgnd vpwr scs8hd_decap_12
XFILLER_12_171 vgnd vpwr scs8hd_decap_3
XANTENNA__170__B _155_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_252 vgnd vpwr scs8hd_decap_12
XFILLER_10_108 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_78 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[4] mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_274 vgnd vpwr scs8hd_fill_1
Xmem_top_track_8.LATCH_1_.latch data_in mem_top_track_8.LATCH_1_.latch/Q _112_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _181_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_266 vgnd vpwr scs8hd_decap_8
XANTENNA__165__B _155_/A vgnd vpwr scs8hd_diode_2
XANTENNA__181__A _181_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vpwr vgnd scs8hd_fill_2
XFILLER_23_14 vgnd vpwr scs8hd_fill_1
XANTENNA__091__A _090_/X vgnd vpwr scs8hd_diode_2
XFILLER_23_69 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
X_186_ _186_/A _186_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _176_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__176__A _176_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_247 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.INVTX1_6_.scs8hd_inv_1 bottom_left_grid_pin_5_ mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_68 vgnd vpwr scs8hd_decap_3
XANTENNA__086__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_11_269 vgnd vpwr scs8hd_decap_8
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_10.INVTX1_0_.scs8hd_inv_1 chany_top_in[5] mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__162__C _161_/C vgnd vpwr scs8hd_diode_2
XFILLER_6_251 vgnd vpwr scs8hd_decap_12
X_169_ _160_/A _155_/A _170_/C _161_/D _169_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_37_188 vgnd vpwr scs8hd_fill_1
XFILLER_37_177 vgnd vpwr scs8hd_decap_6
XFILLER_37_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_199 vpwr vgnd scs8hd_fill_2
XFILLER_28_188 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_210 vpwr vgnd scs8hd_fill_2
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XFILLER_34_158 vgnd vpwr scs8hd_decap_3
XANTENNA__157__C _157_/C vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_9.LATCH_3_.latch data_in mem_bottom_track_9.LATCH_3_.latch/Q _141_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_25_136 vgnd vpwr scs8hd_decap_4
XANTENNA__083__B address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_191 vpwr vgnd scs8hd_fill_2
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_169 vpwr vgnd scs8hd_fill_2
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _174_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_91 vpwr vgnd scs8hd_fill_2
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _168_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_150 vgnd vpwr scs8hd_decap_3
XANTENNA__184__A _184_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__094__A _094_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _178_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_154 vgnd vpwr scs8hd_decap_12
XFILLER_12_150 vgnd vpwr scs8hd_fill_1
XFILLER_12_183 vpwr vgnd scs8hd_fill_2
XFILLER_12_194 vgnd vpwr scs8hd_decap_12
XANTENNA__170__C _170_/C vgnd vpwr scs8hd_diode_2
XANTENNA__179__A _179_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_264 vgnd vpwr scs8hd_decap_12
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
XFILLER_12_16 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB _149_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.tap_buf4_0_.scs8hd_inv_1 mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ _202_/A vgnd vpwr scs8hd_inv_1
XFILLER_37_57 vpwr vgnd scs8hd_fill_2
XFILLER_37_46 vpwr vgnd scs8hd_fill_2
XFILLER_26_253 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_3_.latch data_in mem_top_track_16.LATCH_3_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__089__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_17_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__165__C _157_/C vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ _175_/Y mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_190 vgnd vpwr scs8hd_decap_12
XFILLER_23_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_9_39 vpwr vgnd scs8hd_fill_2
X_185_ _185_/A _185_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_6.INVTX1_1_.scs8hd_inv_1 chany_top_in[8] mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_6 vpwr vgnd scs8hd_fill_2
XFILLER_1_171 vgnd vpwr scs8hd_decap_12
XFILLER_20_259 vgnd vpwr scs8hd_decap_12
XANTENNA__086__B _086_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _176_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_91 vgnd vpwr scs8hd_fill_1
XANTENNA__162__D _162_/D vgnd vpwr scs8hd_diode_2
XFILLER_6_263 vgnd vpwr scs8hd_decap_12
X_168_ _154_/X _168_/B _161_/C _162_/D _168_/Y vgnd vpwr scs8hd_nor4_4
X_099_ address[1] address[2] address[0] _100_/A vgnd vpwr scs8hd_or3_4
XFILLER_37_112 vpwr vgnd scs8hd_fill_2
XFILLER_1_51 vgnd vpwr scs8hd_decap_8
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
XFILLER_1_95 vgnd vpwr scs8hd_decap_12
XFILLER_20_49 vpwr vgnd scs8hd_fill_2
XFILLER_29_36 vpwr vgnd scs8hd_fill_2
XANTENNA__097__A _097_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_93 vgnd vpwr scs8hd_decap_4
XFILLER_34_126 vpwr vgnd scs8hd_fill_2
XFILLER_19_112 vpwr vgnd scs8hd_fill_2
XFILLER_19_145 vpwr vgnd scs8hd_fill_2
XFILLER_35_90 vgnd vpwr scs8hd_decap_3
XANTENNA__157__D _161_/D vgnd vpwr scs8hd_diode_2
XFILLER_40_107 vgnd vpwr scs8hd_decap_3
XANTENNA__083__C _161_/C vgnd vpwr scs8hd_diode_2
XFILLER_0_247 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_17.LATCH_3_.latch data_in mem_bottom_track_17.LATCH_3_.latch/Q _150_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_126 vpwr vgnd scs8hd_fill_2
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_70 vpwr vgnd scs8hd_fill_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XANTENNA__168__C _161_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_251 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.tap_buf4_0_.scs8hd_inv_1 mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ _205_/A vgnd vpwr scs8hd_inv_1
Xmux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _181_/Y mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_8_166 vgnd vpwr scs8hd_decap_12
XANTENNA__170__D _162_/D vgnd vpwr scs8hd_diode_2
XFILLER_35_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_26_221 vgnd vpwr scs8hd_decap_12
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XFILLER_32_213 vgnd vpwr scs8hd_fill_1
XFILLER_17_243 vgnd vpwr scs8hd_fill_1
XANTENNA__165__D _161_/D vgnd vpwr scs8hd_diode_2
XFILLER_4_84 vgnd vpwr scs8hd_decap_8
Xmux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _174_/A mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_257 vgnd vpwr scs8hd_decap_12
XFILLER_2_106 vgnd vpwr scs8hd_decap_12
X_184_ _184_/A _184_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_top_track_0.LATCH_5_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_27 vpwr vgnd scs8hd_fill_2
XFILLER_18_49 vpwr vgnd scs8hd_fill_2
XANTENNA__086__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_11_205 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_80 vgnd vpwr scs8hd_fill_1
X_098_ _085_/B _152_/A _098_/Y vgnd vpwr scs8hd_nor2_4
X_167_ _154_/X _168_/B _161_/C _161_/D _167_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_1_74 vgnd vpwr scs8hd_decap_8
Xmux_right_track_4.INVTX1_1_.scs8hd_inv_1 chany_top_in[7] mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_17 vpwr vgnd scs8hd_fill_2
XFILLER_28_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ _178_/Y mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _113_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_12
XFILLER_10_61 vgnd vpwr scs8hd_fill_1
XFILLER_10_72 vgnd vpwr scs8hd_fill_1
XFILLER_34_105 vpwr vgnd scs8hd_fill_2
XFILLER_19_179 vpwr vgnd scs8hd_fill_2
X_219_ chany_bottom_in[6] chany_top_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_33_193 vpwr vgnd scs8hd_fill_2
XFILLER_15_17 vpwr vgnd scs8hd_fill_2
XFILLER_31_16 vgnd vpwr scs8hd_decap_4
XFILLER_0_259 vpwr vgnd scs8hd_fill_2
XFILLER_0_204 vgnd vpwr scs8hd_decap_12
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_105 vpwr vgnd scs8hd_fill_2
XFILLER_16_149 vgnd vpwr scs8hd_fill_1
XFILLER_24_171 vgnd vpwr scs8hd_decap_8
Xmux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _198_/HI mem_top_track_16.LATCH_2_.latch/Q
+ mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_7 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_193 vpwr vgnd scs8hd_fill_2
XANTENNA__168__D _162_/D vgnd vpwr scs8hd_diode_2
XFILLER_22_119 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_196 vgnd vpwr scs8hd_decap_4
XFILLER_7_73 vpwr vgnd scs8hd_fill_2
XFILLER_7_62 vgnd vpwr scs8hd_decap_8
XFILLER_7_51 vpwr vgnd scs8hd_fill_2
XFILLER_38_263 vgnd vpwr scs8hd_decap_12
XFILLER_26_49 vgnd vpwr scs8hd_decap_12
XFILLER_26_27 vpwr vgnd scs8hd_fill_2
XFILLER_26_16 vpwr vgnd scs8hd_fill_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_108 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _182_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_71 vgnd vpwr scs8hd_decap_4
XFILLER_16_93 vgnd vpwr scs8hd_decap_3
XFILLER_8_101 vpwr vgnd scs8hd_fill_2
XFILLER_8_178 vgnd vpwr scs8hd_decap_12
XFILLER_12_163 vpwr vgnd scs8hd_fill_2
Xmux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ _180_/A mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A top_left_grid_pin_7_ vgnd vpwr scs8hd_diode_2
XFILLER_12_29 vpwr vgnd scs8hd_fill_2
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XFILLER_26_233 vgnd vpwr scs8hd_decap_12
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_92 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_23_225 vgnd vpwr scs8hd_decap_12
XFILLER_23_28 vgnd vpwr scs8hd_decap_4
XFILLER_23_269 vgnd vpwr scs8hd_decap_8
XFILLER_2_118 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_183_ _183_/A _183_/Y vgnd vpwr scs8hd_inv_8
XFILLER_36_9 vgnd vpwr scs8hd_fill_1
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XFILLER_38_80 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _186_/Y mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A bottom_left_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _180_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_217 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 top_left_grid_pin_11_ mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
X_097_ _097_/A _152_/A vgnd vpwr scs8hd_buf_1
X_166_ _161_/A _155_/A _157_/C _162_/D _166_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _186_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_125 vpwr vgnd scs8hd_fill_2
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XFILLER_10_40 vgnd vpwr scs8hd_decap_8
XFILLER_10_84 vpwr vgnd scs8hd_fill_2
XFILLER_19_136 vpwr vgnd scs8hd_fill_2
XFILLER_19_93 vpwr vgnd scs8hd_fill_2
XFILLER_19_158 vpwr vgnd scs8hd_fill_2
X_218_ _218_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
X_149_ _109_/A _152_/B _149_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_3 vgnd vpwr scs8hd_decap_8
XFILLER_25_117 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_150 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_39 vgnd vpwr scs8hd_decap_3
XFILLER_0_249 vgnd vpwr scs8hd_decap_6
XFILLER_0_216 vgnd vpwr scs8hd_fill_1
Xmux_right_track_2.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_109 vpwr vgnd scs8hd_fill_2
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A bottom_left_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_30_175 vgnd vpwr scs8hd_decap_6
XFILLER_7_96 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _189_/HI mem_bottom_track_9.LATCH_2_.latch/Q
+ mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_142 vpwr vgnd scs8hd_fill_2
XFILLER_21_153 vpwr vgnd scs8hd_fill_2
XFILLER_21_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_242 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_142 vpwr vgnd scs8hd_fill_2
XFILLER_32_93 vgnd vpwr scs8hd_fill_1
XFILLER_32_60 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _175_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _182_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_27 vgnd vpwr scs8hd_decap_12
XFILLER_26_212 vpwr vgnd scs8hd_fill_2
XFILLER_26_245 vgnd vpwr scs8hd_decap_8
XFILLER_5_105 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_223 vgnd vpwr scs8hd_decap_12
XFILLER_17_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_237 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_40 vpwr vgnd scs8hd_fill_2
XFILLER_14_215 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_182_ _182_/A _182_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_196 vgnd vpwr scs8hd_decap_12
XANTENNA__100__A _100_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_218 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_2_.scs8hd_inv_1 top_left_grid_pin_15_ mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_229 vgnd vpwr scs8hd_decap_12
Xmux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ _173_/Y mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_83 vpwr vgnd scs8hd_fill_2
XFILLER_10_251 vgnd vpwr scs8hd_decap_12
X_165_ _161_/A _155_/A _157_/C _161_/D _165_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_40_93 vpwr vgnd scs8hd_fill_2
XFILLER_34_7 vgnd vpwr scs8hd_decap_12
X_096_ address[1] address[2] _171_/D _097_/A vgnd vpwr scs8hd_or3_4
XFILLER_37_148 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_1_.latch data_in mem_top_track_0.LATCH_1_.latch/Q _098_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_17 vgnd vpwr scs8hd_decap_3
XFILLER_28_148 vgnd vpwr scs8hd_decap_4
XFILLER_3_269 vgnd vpwr scs8hd_decap_8
XFILLER_3_214 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _177_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_50 vgnd vpwr scs8hd_fill_1
XFILLER_19_72 vpwr vgnd scs8hd_fill_2
XFILLER_34_118 vgnd vpwr scs8hd_decap_8
XFILLER_27_181 vpwr vgnd scs8hd_fill_2
X_148_ _108_/A _152_/B _148_/Y vgnd vpwr scs8hd_nor2_4
X_217_ _217_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_25_3 vpwr vgnd scs8hd_fill_2
X_079_ address[5] _154_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_0_239 vpwr vgnd scs8hd_fill_2
XFILLER_24_195 vgnd vpwr scs8hd_decap_4
XFILLER_24_151 vpwr vgnd scs8hd_fill_2
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_62 vgnd vpwr scs8hd_fill_1
XFILLER_21_95 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB _088_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_154 vgnd vpwr scs8hd_decap_3
XFILLER_30_110 vgnd vpwr scs8hd_fill_1
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_7_31 vgnd vpwr scs8hd_decap_12
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_132 vgnd vpwr scs8hd_decap_4
XFILLER_21_176 vgnd vpwr scs8hd_decap_4
XFILLER_29_210 vgnd vpwr scs8hd_decap_12
XFILLER_12_187 vpwr vgnd scs8hd_fill_2
XFILLER_16_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _152_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_50 vgnd vpwr scs8hd_fill_1
XANTENNA__103__A address[3] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_4_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_39 vgnd vpwr scs8hd_decap_4
XFILLER_5_128 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_3_.latch data_in mem_bottom_track_1.LATCH_3_.latch/Q _131_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_205 vpwr vgnd scs8hd_fill_2
XFILLER_17_235 vgnd vpwr scs8hd_decap_8
Xmux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _179_/Y mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_76 vgnd vpwr scs8hd_decap_3
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_227 vgnd vpwr scs8hd_decap_12
X_181_ _181_/A _181_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_22_271 vgnd vpwr scs8hd_decap_4
XFILLER_13_85 vpwr vgnd scs8hd_fill_2
Xmem_right_track_14.LATCH_0_.latch data_in _186_/A _172_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_208 vgnd vpwr scs8hd_decap_6
XFILLER_9_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
X_095_ _085_/B _111_/A _095_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_263 vgnd vpwr scs8hd_decap_12
X_164_ _161_/A _161_/B _106_/C _162_/D _164_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_24_62 vpwr vgnd scs8hd_fill_2
XFILLER_27_7 vpwr vgnd scs8hd_fill_2
XFILLER_37_127 vpwr vgnd scs8hd_fill_2
XFILLER_37_116 vgnd vpwr scs8hd_decap_6
XANTENNA__111__A _111_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_88 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_28_138 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_12.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_226 vgnd vpwr scs8hd_decap_12
XFILLER_3_204 vgnd vpwr scs8hd_decap_3
XFILLER_10_64 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_116 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_147_ _147_/A _152_/B vgnd vpwr scs8hd_buf_1
X_216_ chany_top_in[0] chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
X_078_ _077_/X _108_/A vgnd vpwr scs8hd_buf_1
XANTENNA__106__A _154_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_160 vgnd vpwr scs8hd_fill_1
XFILLER_18_193 vgnd vpwr scs8hd_decap_4
XFILLER_33_174 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
XFILLER_24_130 vpwr vgnd scs8hd_fill_2
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_top_track_16.LATCH_3_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_30_122 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ _176_/Y mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_7_43 vgnd vpwr scs8hd_decap_6
XFILLER_15_163 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_222 vgnd vpwr scs8hd_decap_12
XFILLER_32_84 vgnd vpwr scs8hd_decap_8
XFILLER_26_258 vgnd vpwr scs8hd_decap_12
XANTENNA__204__A _204_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB _164_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XANTENNA__114__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_239 vgnd vpwr scs8hd_decap_12
X_180_ _180_/A _180_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_20 vpwr vgnd scs8hd_fill_2
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_110 vpwr vgnd scs8hd_fill_2
XANTENNA__109__A _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_232 vgnd vpwr scs8hd_decap_12
XFILLER_34_19 vgnd vpwr scs8hd_fill_1
XFILLER_24_41 vpwr vgnd scs8hd_fill_2
XFILLER_40_84 vgnd vpwr scs8hd_decap_8
XFILLER_6_202 vgnd vpwr scs8hd_decap_12
X_094_ _094_/A _111_/A vgnd vpwr scs8hd_buf_1
X_163_ _161_/A _161_/B _106_/C _161_/D _163_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__111__B _109_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _199_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_2_.latch data_in mem_top_track_8.LATCH_2_.latch/Q _111_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_106 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _181_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ _182_/Y mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_3_238 vgnd vpwr scs8hd_decap_6
XANTENNA__212__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_10_32 vgnd vpwr scs8hd_decap_4
XFILLER_27_194 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_153 vpwr vgnd scs8hd_fill_2
X_215_ chany_top_in[1] chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_35_95 vpwr vgnd scs8hd_fill_2
XFILLER_35_73 vpwr vgnd scs8hd_fill_2
XANTENNA__122__A _111_/A vgnd vpwr scs8hd_diode_2
X_077_ address[1] _086_/B _171_/D _077_/X vgnd vpwr scs8hd_or3_4
XANTENNA__106__B _155_/A vgnd vpwr scs8hd_diode_2
X_146_ _160_/A _146_/B _161_/C _147_/A vgnd vpwr scs8hd_or3_4
XFILLER_33_197 vpwr vgnd scs8hd_fill_2
XFILLER_25_109 vpwr vgnd scs8hd_fill_2
XFILLER_18_172 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_109 vpwr vgnd scs8hd_fill_2
XANTENNA__207__A _207_/A vgnd vpwr scs8hd_diode_2
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_31 vgnd vpwr scs8hd_decap_4
XFILLER_21_42 vpwr vgnd scs8hd_fill_2
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_142 vpwr vgnd scs8hd_fill_2
XFILLER_15_175 vpwr vgnd scs8hd_fill_2
XFILLER_30_145 vgnd vpwr scs8hd_decap_3
XFILLER_7_77 vpwr vgnd scs8hd_fill_2
XFILLER_7_55 vpwr vgnd scs8hd_fill_2
XFILLER_15_197 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _154_/A vgnd vpwr scs8hd_diode_2
X_129_ _108_/A _131_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_3_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_112 vpwr vgnd scs8hd_fill_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_12
XFILLER_29_234 vgnd vpwr scs8hd_decap_8
XFILLER_16_75 vgnd vpwr scs8hd_fill_1
XFILLER_8_105 vgnd vpwr scs8hd_decap_4
XFILLER_12_167 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_204 vpwr vgnd scs8hd_fill_2
XFILLER_35_248 vpwr vgnd scs8hd_fill_2
XFILLER_26_215 vgnd vpwr scs8hd_decap_4
XFILLER_26_204 vgnd vpwr scs8hd_decap_8
Xmem_bottom_track_9.LATCH_4_.latch data_in mem_bottom_track_9.LATCH_4_.latch/Q _140_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__220__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_27_41 vpwr vgnd scs8hd_fill_2
XFILLER_17_204 vpwr vgnd scs8hd_fill_2
XFILLER_17_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _190_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_251 vgnd vpwr scs8hd_decap_12
XFILLER_32_218 vgnd vpwr scs8hd_decap_12
XFILLER_27_96 vpwr vgnd scs8hd_fill_2
XFILLER_17_259 vpwr vgnd scs8hd_fill_2
XFILLER_4_56 vgnd vpwr scs8hd_decap_12
XANTENNA__130__A _109_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _185_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__215__A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_13_65 vpwr vgnd scs8hd_fill_2
XFILLER_38_84 vgnd vpwr scs8hd_decap_8
XANTENNA__109__B _109_/B vgnd vpwr scs8hd_diode_2
XANTENNA__125__A address[6] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_6_.scs8hd_inv_1 bottom_left_grid_pin_9_ mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _178_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
X_162_ _161_/A _161_/B _161_/C _162_/D _162_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_40_30 vgnd vpwr scs8hd_fill_1
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
X_093_ _093_/A address[2] address[0] _094_/A vgnd vpwr scs8hd_or3_4
Xmem_top_track_16.LATCH_4_.latch data_in mem_top_track_16.LATCH_4_.latch/Q _120_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_right_track_10.LATCH_0_.latch data_in _180_/A _166_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_88 vgnd vpwr scs8hd_decap_4
XFILLER_19_53 vpwr vgnd scs8hd_fill_2
XFILLER_35_52 vpwr vgnd scs8hd_fill_2
XFILLER_27_184 vgnd vpwr scs8hd_fill_1
XFILLER_27_140 vgnd vpwr scs8hd_decap_4
XFILLER_19_97 vpwr vgnd scs8hd_fill_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
X_145_ address[5] _160_/A vgnd vpwr scs8hd_inv_8
X_214_ chany_top_in[2] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA__106__C _106_/C vgnd vpwr scs8hd_diode_2
XANTENNA__122__B _121_/B vgnd vpwr scs8hd_diode_2
X_076_ address[0] _171_/D vgnd vpwr scs8hd_inv_8
XFILLER_18_151 vpwr vgnd scs8hd_fill_2
XFILLER_33_154 vgnd vpwr scs8hd_decap_3
XFILLER_33_143 vgnd vpwr scs8hd_decap_4
XFILLER_33_110 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_143 vgnd vpwr scs8hd_decap_8
XFILLER_24_110 vgnd vpwr scs8hd_decap_3
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vgnd vpwr scs8hd_decap_4
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__223__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_30_102 vgnd vpwr scs8hd_decap_8
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_132 vgnd vpwr scs8hd_decap_4
X_128_ _127_/X _131_/B vgnd vpwr scs8hd_buf_1
XANTENNA__133__A _152_/A vgnd vpwr scs8hd_diode_2
XANTENNA__117__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_38_213 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _176_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_157 vpwr vgnd scs8hd_fill_2
XFILLER_29_257 vgnd vpwr scs8hd_decap_12
XANTENNA__218__A _218_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_54 vpwr vgnd scs8hd_fill_2
XFILLER_32_97 vpwr vgnd scs8hd_fill_2
XFILLER_32_64 vpwr vgnd scs8hd_fill_2
XFILLER_32_42 vgnd vpwr scs8hd_decap_8
XFILLER_12_146 vgnd vpwr scs8hd_decap_4
XANTENNA__128__A _127_/X vgnd vpwr scs8hd_diode_2
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _184_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB _108_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_109 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_27_53 vpwr vgnd scs8hd_fill_2
XFILLER_17_249 vgnd vpwr scs8hd_decap_6
XFILLER_40_263 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_17.LATCH_4_.latch data_in mem_bottom_track_17.LATCH_4_.latch/Q _149_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_68 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__130__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_271 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_230 vgnd vpwr scs8hd_decap_12
XFILLER_1_123 vgnd vpwr scs8hd_decap_12
Xmem_right_track_6.LATCH_0_.latch data_in _178_/A _164_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_245 vgnd vpwr scs8hd_decap_12
XANTENNA__141__A _110_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_193 vpwr vgnd scs8hd_fill_2
XANTENNA__226__A _226_/A vgnd vpwr scs8hd_diode_2
X_161_ _161_/A _161_/B _161_/C _161_/D _161_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_24_87 vpwr vgnd scs8hd_fill_2
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
XFILLER_10_200 vgnd vpwr scs8hd_decap_12
XFILLER_40_97 vpwr vgnd scs8hd_fill_2
X_092_ _085_/B _110_/A _092_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_108 vpwr vgnd scs8hd_fill_2
XANTENNA__136__A _135_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _178_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_163 vgnd vpwr scs8hd_decap_3
XFILLER_36_152 vgnd vpwr scs8hd_fill_1
XFILLER_19_65 vgnd vpwr scs8hd_decap_4
Xmux_right_track_12.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[7] mux_right_track_12.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_100 vgnd vpwr scs8hd_fill_1
XFILLER_27_174 vgnd vpwr scs8hd_decap_4
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_213_ _213_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
Xmux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _199_/HI mem_top_track_8.LATCH_2_.latch/Q
+ mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_075_ address[2] _086_/B vgnd vpwr scs8hd_inv_8
X_144_ _101_/B _141_/B _144_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_2.tap_buf4_0_.scs8hd_inv_1 mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _207_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _098_/Y vgnd vpwr scs8hd_diode_2
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_9.INVTX1_5_.scs8hd_inv_1 bottom_left_grid_pin_1_ mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_66 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XANTENNA__117__C _170_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__133__B _131_/B vgnd vpwr scs8hd_diode_2
X_127_ _154_/A _168_/B _170_/C _127_/X vgnd vpwr scs8hd_or3_4
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _217_/A vgnd vpwr scs8hd_inv_1
Xmux_top_track_16.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[2] mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_269 vgnd vpwr scs8hd_decap_8
XFILLER_8_118 vgnd vpwr scs8hd_decap_8
XFILLER_12_125 vpwr vgnd scs8hd_fill_2
XFILLER_16_88 vpwr vgnd scs8hd_fill_2
XFILLER_32_32 vgnd vpwr scs8hd_fill_1
XFILLER_8_129 vgnd vpwr scs8hd_decap_8
XFILLER_11_180 vgnd vpwr scs8hd_fill_1
XANTENNA__144__A _101_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_184 vgnd vpwr scs8hd_decap_12
XFILLER_7_151 vgnd vpwr scs8hd_decap_12
Xmux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _174_/Y mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_32_209 vgnd vpwr scs8hd_decap_4
XFILLER_27_65 vpwr vgnd scs8hd_fill_2
XFILLER_4_154 vgnd vpwr scs8hd_decap_12
XFILLER_4_121 vgnd vpwr scs8hd_decap_12
XANTENNA__139__A _108_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_12 vpwr vgnd scs8hd_fill_2
XFILLER_22_242 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_2_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_89 vpwr vgnd scs8hd_fill_2
XFILLER_38_64 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_135 vgnd vpwr scs8hd_decap_12
XFILLER_13_242 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_257 vgnd vpwr scs8hd_decap_12
XANTENNA__141__B _141_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_161 vpwr vgnd scs8hd_fill_2
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
X_160_ _160_/A _161_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_227 vgnd vpwr scs8hd_decap_12
X_091_ _090_/X _110_/A vgnd vpwr scs8hd_buf_1
XFILLER_10_212 vpwr vgnd scs8hd_fill_2
XFILLER_24_66 vpwr vgnd scs8hd_fill_2
XFILLER_1_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_59 vpwr vgnd scs8hd_fill_2
XANTENNA__152__A _152_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_142 vpwr vgnd scs8hd_fill_2
XFILLER_10_57 vgnd vpwr scs8hd_decap_4
XFILLER_10_68 vgnd vpwr scs8hd_decap_4
XFILLER_19_33 vpwr vgnd scs8hd_fill_2
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_42_145 vgnd vpwr scs8hd_decap_8
XFILLER_42_134 vgnd vpwr scs8hd_decap_8
XFILLER_42_123 vgnd vpwr scs8hd_fill_1
XFILLER_35_43 vpwr vgnd scs8hd_fill_2
X_212_ chany_top_in[4] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
X_143_ _152_/A _141_/B _143_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
XFILLER_33_123 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_131 vgnd vpwr scs8hd_decap_4
XFILLER_33_178 vgnd vpwr scs8hd_decap_3
XANTENNA__147__A _147_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_91 vgnd vpwr scs8hd_fill_1
XFILLER_2_80 vgnd vpwr scs8hd_decap_8
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_9 vgnd vpwr scs8hd_decap_3
Xmux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ _180_/Y mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_30_159 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[5] mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_126_ _146_/B _168_/B vgnd vpwr scs8hd_buf_1
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_6 vgnd vpwr scs8hd_decap_12
Xmux_right_track_10.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[8] mux_right_track_10.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_16_12 vpwr vgnd scs8hd_fill_2
XFILLER_16_23 vpwr vgnd scs8hd_fill_2
XFILLER_32_11 vgnd vpwr scs8hd_decap_3
XFILLER_12_104 vpwr vgnd scs8hd_fill_2
XFILLER_16_78 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _186_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_163 vgnd vpwr scs8hd_decap_12
XANTENNA__144__B _141_/B vgnd vpwr scs8hd_diode_2
X_109_ _109_/A _109_/B _109_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__160__A _160_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_196 vgnd vpwr scs8hd_decap_12
XFILLER_34_251 vgnd vpwr scs8hd_decap_12
XFILLER_27_11 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_22 vpwr vgnd scs8hd_fill_2
XFILLER_25_240 vgnd vpwr scs8hd_decap_4
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_166 vgnd vpwr scs8hd_decap_12
XFILLER_4_133 vgnd vpwr scs8hd_decap_12
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__155__A _155_/A vgnd vpwr scs8hd_diode_2
XANTENNA__139__B _141_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A bottom_left_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_24 vgnd vpwr scs8hd_decap_3
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_22_254 vgnd vpwr scs8hd_fill_1
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_8_6 vgnd vpwr scs8hd_decap_12
XFILLER_1_114 vgnd vpwr scs8hd_decap_8
XFILLER_1_147 vgnd vpwr scs8hd_decap_12
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_210 vgnd vpwr scs8hd_decap_12
XFILLER_9_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_184 vgnd vpwr scs8hd_decap_4
XFILLER_39_173 vpwr vgnd scs8hd_fill_2
XFILLER_24_23 vpwr vgnd scs8hd_fill_2
XFILLER_24_45 vpwr vgnd scs8hd_fill_2
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XFILLER_6_239 vgnd vpwr scs8hd_decap_12
X_090_ _093_/A address[2] _171_/D _090_/X vgnd vpwr scs8hd_or3_4
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _182_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB _172_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__152__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_176 vgnd vpwr scs8hd_decap_3
Xmem_right_track_2.LATCH_0_.latch data_in _174_/A _159_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_36 vgnd vpwr scs8hd_fill_1
XFILLER_19_12 vpwr vgnd scs8hd_fill_2
XFILLER_27_132 vpwr vgnd scs8hd_fill_2
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
XFILLER_35_77 vpwr vgnd scs8hd_fill_2
XFILLER_27_198 vgnd vpwr scs8hd_decap_4
X_211_ chany_top_in[5] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
X_142_ _111_/A _141_/B _142_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A bottom_left_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_110 vpwr vgnd scs8hd_fill_2
XFILLER_18_154 vgnd vpwr scs8hd_decap_6
XFILLER_18_176 vgnd vpwr scs8hd_decap_4
XANTENNA__163__A _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_102 vpwr vgnd scs8hd_fill_2
XFILLER_24_179 vgnd vpwr scs8hd_fill_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_35 vgnd vpwr scs8hd_fill_1
XFILLER_21_46 vpwr vgnd scs8hd_fill_2
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XFILLER_15_102 vgnd vpwr scs8hd_decap_3
XFILLER_15_146 vpwr vgnd scs8hd_fill_2
XFILLER_7_59 vpwr vgnd scs8hd_fill_2
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
X_125_ address[6] _146_/B vgnd vpwr scs8hd_inv_8
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XFILLER_38_205 vgnd vpwr scs8hd_decap_8
XFILLER_23_6 vpwr vgnd scs8hd_fill_2
XANTENNA__158__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_21_116 vgnd vpwr scs8hd_decap_4
XFILLER_21_138 vpwr vgnd scs8hd_fill_2
XFILLER_16_35 vpwr vgnd scs8hd_fill_2
XFILLER_32_23 vgnd vpwr scs8hd_decap_6
Xmem_top_track_0.LATCH_2_.latch data_in mem_top_track_0.LATCH_2_.latch/Q _095_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_138 vpwr vgnd scs8hd_fill_2
XFILLER_20_171 vgnd vpwr scs8hd_decap_3
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
X_108_ _108_/A _109_/B _108_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_175 vgnd vpwr scs8hd_decap_8
XFILLER_11_193 vgnd vpwr scs8hd_decap_12
XFILLER_21_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB _167_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _177_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _222_/A vgnd vpwr scs8hd_inv_1
XFILLER_27_45 vgnd vpwr scs8hd_decap_3
XFILLER_17_208 vgnd vpwr scs8hd_decap_4
XFILLER_17_219 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _191_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_178 vgnd vpwr scs8hd_decap_12
XFILLER_4_145 vgnd vpwr scs8hd_decap_8
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__171__A _154_/X vgnd vpwr scs8hd_diode_2
XFILLER_22_200 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.INVTX1_3_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_36 vpwr vgnd scs8hd_fill_2
XFILLER_13_69 vgnd vpwr scs8hd_decap_3
XFILLER_1_159 vgnd vpwr scs8hd_decap_12
XANTENNA__081__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_222 vgnd vpwr scs8hd_decap_12
XANTENNA__166__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_92 vpwr vgnd scs8hd_fill_2
XFILLER_5_70 vgnd vpwr scs8hd_decap_3
XFILLER_24_79 vpwr vgnd scs8hd_fill_2
XANTENNA__076__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XFILLER_1_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_4_.latch data_in mem_bottom_track_1.LATCH_4_.latch/Q _130_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_4.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_199 vgnd vpwr scs8hd_decap_12
XFILLER_36_188 vgnd vpwr scs8hd_decap_8
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_19_46 vgnd vpwr scs8hd_decap_4
XFILLER_42_125 vgnd vpwr scs8hd_decap_6
XFILLER_35_56 vgnd vpwr scs8hd_decap_3
XFILLER_35_12 vgnd vpwr scs8hd_decap_12
XFILLER_27_155 vpwr vgnd scs8hd_fill_2
XFILLER_27_111 vpwr vgnd scs8hd_fill_2
XFILLER_19_57 vpwr vgnd scs8hd_fill_2
X_141_ _110_/A _141_/B _141_/Y vgnd vpwr scs8hd_nor2_4
X_210_ chany_top_in[6] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_3_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_114 vpwr vgnd scs8hd_fill_2
XFILLER_18_144 vgnd vpwr scs8hd_decap_4
XANTENNA__163__B _161_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _183_/A vgnd vpwr
+ scs8hd_diode_2
Xmem_right_track_14.LATCH_1_.latch data_in _185_/A _171_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_14 vpwr vgnd scs8hd_fill_2
XFILLER_30_128 vgnd vpwr scs8hd_decap_8
XFILLER_15_114 vpwr vgnd scs8hd_fill_2
XFILLER_15_169 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
X_124_ _101_/B _121_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_91 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_5_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__174__A _174_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_58 vpwr vgnd scs8hd_fill_2
XFILLER_32_68 vgnd vpwr scs8hd_decap_3
XANTENNA__084__A _083_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_150 vgnd vpwr scs8hd_fill_1
XFILLER_20_183 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
X_107_ _106_/X _109_/B vgnd vpwr scs8hd_buf_1
XFILLER_7_121 vgnd vpwr scs8hd_fill_1
XFILLER_11_172 vpwr vgnd scs8hd_fill_2
XANTENNA__169__A _160_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_261 vgnd vpwr scs8hd_decap_12
XFILLER_8_70 vgnd vpwr scs8hd_decap_3
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XANTENNA__079__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_25_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_245 vgnd vpwr scs8hd_decap_12
XFILLER_31_212 vgnd vpwr scs8hd_decap_12
XANTENNA__171__B _168_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_212 vpwr vgnd scs8hd_fill_2
XANTENNA__081__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_13_234 vgnd vpwr scs8hd_decap_8
XFILLER_13_245 vgnd vpwr scs8hd_decap_12
XANTENNA__166__B _155_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr
+ scs8hd_diode_2
XANTENNA__182__A _182_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_197 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_215 vgnd vpwr scs8hd_decap_12
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XANTENNA__092__A _085_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__177__A _177_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_10.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XFILLER_19_69 vgnd vpwr scs8hd_fill_1
XFILLER_42_115 vgnd vpwr scs8hd_decap_8
XFILLER_42_104 vgnd vpwr scs8hd_decap_8
XFILLER_35_24 vgnd vpwr scs8hd_decap_8
XFILLER_27_178 vgnd vpwr scs8hd_fill_1
XANTENNA__087__A _087_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_140_ _109_/A _141_/B _140_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_track_16.LATCH_4_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_bottom_track_9.INVTX1_2_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_159 vpwr vgnd scs8hd_fill_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_18_189 vpwr vgnd scs8hd_fill_2
XANTENNA__163__C _106_/C vgnd vpwr scs8hd_diode_2
XFILLER_24_126 vpwr vgnd scs8hd_fill_2
XFILLER_24_115 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_159 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_3_.scs8hd_inv_1 chanx_right_in[0] mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_123_ _152_/A _121_/B _123_/Y vgnd vpwr scs8hd_nor2_4
Xmem_top_track_8.LATCH_3_.latch data_in mem_top_track_8.LATCH_3_.latch/Q _110_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_251 vgnd vpwr scs8hd_decap_12
XFILLER_11_151 vgnd vpwr scs8hd_decap_3
X_106_ _154_/A _155_/A _106_/C _106_/X vgnd vpwr scs8hd_or3_4
XFILLER_22_80 vgnd vpwr scs8hd_fill_1
XANTENNA__169__B _155_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XANTENNA__185__A _185_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_273 vgnd vpwr scs8hd_decap_4
XFILLER_8_93 vgnd vpwr scs8hd_decap_4
XFILLER_27_69 vpwr vgnd scs8hd_fill_2
XFILLER_40_202 vgnd vpwr scs8hd_decap_12
XANTENNA__095__A _085_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_31_224 vgnd vpwr scs8hd_decap_12
XFILLER_16_254 vgnd vpwr scs8hd_fill_1
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_257 vgnd vpwr scs8hd_decap_12
XANTENNA__171__C _106_/C vgnd vpwr scs8hd_diode_2
XFILLER_13_16 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__081__C _135_/C vgnd vpwr scs8hd_diode_2
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_13_257 vgnd vpwr scs8hd_decap_12
XFILLER_28_90 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 chany_top_in[4] mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__166__C _157_/C vgnd vpwr scs8hd_diode_2
XFILLER_39_132 vpwr vgnd scs8hd_fill_2
XFILLER_39_165 vgnd vpwr scs8hd_decap_4
XFILLER_24_15 vpwr vgnd scs8hd_fill_2
XANTENNA__092__B _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_227 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_220 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_9.LATCH_5_.latch data_in mem_bottom_track_9.LATCH_5_.latch/Q _139_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_6 vpwr vgnd scs8hd_fill_2
XFILLER_36_168 vgnd vpwr scs8hd_decap_8
XFILLER_36_146 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
XFILLER_35_47 vgnd vpwr scs8hd_decap_3
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _185_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_5_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_199_ _199_/HI _199_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__163__D _161_/D vgnd vpwr scs8hd_diode_2
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _192_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_4_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_8.INVTX1_4_.scs8hd_inv_1 chanx_right_in[5] mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_38 vgnd vpwr scs8hd_fill_1
XANTENNA__098__A _085_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_138 vpwr vgnd scs8hd_fill_2
XFILLER_23_193 vpwr vgnd scs8hd_fill_2
X_122_ _111_/A _121_/B _122_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_108 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_5_.latch data_in mem_top_track_16.LATCH_5_.latch/Q _119_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_241 vgnd vpwr scs8hd_decap_3
XFILLER_16_16 vpwr vgnd scs8hd_fill_2
XFILLER_12_119 vgnd vpwr scs8hd_decap_4
XFILLER_16_27 vpwr vgnd scs8hd_fill_2
Xmem_right_track_10.LATCH_1_.latch data_in _179_/A _165_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_163 vpwr vgnd scs8hd_fill_2
XFILLER_20_196 vgnd vpwr scs8hd_decap_12
XFILLER_28_263 vgnd vpwr scs8hd_decap_12
XFILLER_7_134 vgnd vpwr scs8hd_decap_3
XFILLER_7_123 vgnd vpwr scs8hd_decap_3
X_105_ _105_/A _106_/C vgnd vpwr scs8hd_buf_1
XFILLER_22_70 vgnd vpwr scs8hd_decap_4
XFILLER_34_200 vpwr vgnd scs8hd_fill_2
XANTENNA__169__C _170_/C vgnd vpwr scs8hd_diode_2
XFILLER_27_26 vpwr vgnd scs8hd_fill_2
XFILLER_27_15 vpwr vgnd scs8hd_fill_2
XFILLER_25_211 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__095__B _111_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_104 vgnd vpwr scs8hd_decap_8
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_236 vgnd vpwr scs8hd_decap_8
XFILLER_16_211 vgnd vpwr scs8hd_decap_3
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_269 vgnd vpwr scs8hd_decap_8
XANTENNA__171__D _171_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_47 vgnd vpwr scs8hd_decap_8
XFILLER_13_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_195 vpwr vgnd scs8hd_fill_2
XANTENNA__166__D _162_/D vgnd vpwr scs8hd_diode_2
XFILLER_5_62 vgnd vpwr scs8hd_decap_8
XFILLER_5_51 vgnd vpwr scs8hd_decap_8
XFILLER_8_251 vgnd vpwr scs8hd_decap_12
XFILLER_39_177 vgnd vpwr scs8hd_decap_6
XFILLER_39_188 vgnd vpwr scs8hd_fill_1
XFILLER_24_27 vpwr vgnd scs8hd_fill_2
XFILLER_24_49 vpwr vgnd scs8hd_fill_2
XFILLER_10_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_81 vpwr vgnd scs8hd_fill_2
XFILLER_5_232 vgnd vpwr scs8hd_decap_12
XFILLER_14_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _184_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_36_125 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_17.LATCH_5_.latch data_in mem_bottom_track_17.LATCH_5_.latch/Q _148_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_136 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_16 vpwr vgnd scs8hd_fill_2
XFILLER_2_202 vgnd vpwr scs8hd_decap_12
XFILLER_33_139 vpwr vgnd scs8hd_fill_2
XFILLER_18_114 vpwr vgnd scs8hd_fill_2
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XFILLER_25_92 vpwr vgnd scs8hd_fill_2
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _187_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_91 vgnd vpwr scs8hd_decap_4
X_198_ _198_/HI _198_/LO vgnd vpwr scs8hd_conb_1
Xmux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_106 vpwr vgnd scs8hd_fill_2
XFILLER_32_194 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[4] mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_right_track_6.LATCH_1_.latch data_in _177_/A _163_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__098__B _152_/A vgnd vpwr scs8hd_diode_2
X_121_ _110_/A _121_/B _121_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_19 vgnd vpwr scs8hd_decap_12
XFILLER_14_172 vgnd vpwr scs8hd_fill_1
XFILLER_16_39 vpwr vgnd scs8hd_fill_2
XFILLER_20_186 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _178_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_113 vpwr vgnd scs8hd_fill_2
X_104_ _135_/A address[4] _135_/C _105_/A vgnd vpwr scs8hd_or3_4
XFILLER_34_212 vpwr vgnd scs8hd_fill_2
XANTENNA__169__D _161_/D vgnd vpwr scs8hd_diode_2
XFILLER_8_40 vgnd vpwr scs8hd_decap_3
XFILLER_8_84 vpwr vgnd scs8hd_fill_2
XFILLER_6_190 vgnd vpwr scs8hd_decap_12
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_25_245 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_93 vpwr vgnd scs8hd_fill_2
XFILLER_3_171 vgnd vpwr scs8hd_decap_12
XFILLER_22_204 vgnd vpwr scs8hd_decap_8
XFILLER_22_259 vgnd vpwr scs8hd_decap_12
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XFILLER_9_208 vgnd vpwr scs8hd_decap_12
XFILLER_0_163 vpwr vgnd scs8hd_fill_2
XFILLER_0_185 vgnd vpwr scs8hd_fill_1
XFILLER_8_263 vgnd vpwr scs8hd_decap_12
XFILLER_39_101 vpwr vgnd scs8hd_fill_2
XFILLER_30_60 vpwr vgnd scs8hd_fill_2
XFILLER_39_91 vpwr vgnd scs8hd_fill_2
XFILLER_27_159 vpwr vgnd scs8hd_fill_2
XFILLER_27_115 vgnd vpwr scs8hd_decap_4
Xmux_right_track_14.tap_buf4_0_.scs8hd_inv_1 mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _201_/A vgnd vpwr scs8hd_inv_1
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XFILLER_33_118 vpwr vgnd scs8hd_fill_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_26_181 vpwr vgnd scs8hd_fill_2
XFILLER_25_71 vpwr vgnd scs8hd_fill_2
XFILLER_18_148 vgnd vpwr scs8hd_fill_1
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XFILLER_41_151 vgnd vpwr scs8hd_decap_12
X_197_ _197_/HI _197_/LO vgnd vpwr scs8hd_conb_1
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _218_/A vgnd vpwr scs8hd_inv_1
XFILLER_32_173 vgnd vpwr scs8hd_decap_12
XFILLER_21_18 vpwr vgnd scs8hd_fill_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
X_120_ _109_/A _121_/B _120_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_173 vgnd vpwr scs8hd_decap_4
Xmux_right_track_4.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_95 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_221 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_121 vpwr vgnd scs8hd_fill_2
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_11_176 vgnd vpwr scs8hd_decap_4
XFILLER_11_187 vgnd vpwr scs8hd_decap_4
X_103_ address[3] _135_/A vgnd vpwr scs8hd_inv_8
XFILLER_19_243 vgnd vpwr scs8hd_fill_1
XFILLER_8_30 vgnd vpwr scs8hd_fill_1
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XFILLER_25_257 vgnd vpwr scs8hd_decap_12
XFILLER_16_224 vgnd vpwr scs8hd_decap_12
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_12.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_120 vgnd vpwr scs8hd_decap_4
XFILLER_0_142 vpwr vgnd scs8hd_fill_2
XFILLER_0_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _204_/A vgnd vpwr scs8hd_inv_1
XFILLER_14_84 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_245 vgnd vpwr scs8hd_decap_12
XANTENNA__101__A _085_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_193 vgnd vpwr scs8hd_decap_3
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_127 vpwr vgnd scs8hd_fill_2
XPHY_83 vgnd vpwr scs8hd_decap_3
XFILLER_41_163 vgnd vpwr scs8hd_decap_12
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
XFILLER_41_82 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
X_196_ _196_/HI _196_/LO vgnd vpwr scs8hd_conb_1
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_5_ mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_17_160 vgnd vpwr scs8hd_fill_1
XFILLER_17_182 vgnd vpwr scs8hd_fill_1
XFILLER_32_141 vgnd vpwr scs8hd_decap_12
XFILLER_17_193 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _187_/HI mem_bottom_track_1.LATCH_2_.latch/Q
+ mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_11_52 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_93 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_179_ _179_/A _179_/Y vgnd vpwr scs8hd_inv_8
XFILLER_37_233 vgnd vpwr scs8hd_decap_8
XFILLER_35_3 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_211 vgnd vpwr scs8hd_decap_3
Xmem_right_track_2.LATCH_1_.latch data_in _173_/A _157_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_111 vpwr vgnd scs8hd_fill_2
X_102_ address[6] _155_/A vgnd vpwr scs8hd_buf_1
XFILLER_22_84 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_97 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_239 vgnd vpwr scs8hd_decap_12
XFILLER_25_269 vgnd vpwr scs8hd_decap_8
XFILLER_16_203 vgnd vpwr scs8hd_decap_8
XFILLER_16_236 vgnd vpwr scs8hd_decap_12
XFILLER_17_73 vgnd vpwr scs8hd_decap_3
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_72 vpwr vgnd scs8hd_fill_2
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_184 vgnd vpwr scs8hd_decap_12
XANTENNA__104__A _135_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_83 vgnd vpwr scs8hd_decap_4
XFILLER_0_132 vgnd vpwr scs8hd_decap_6
XFILLER_0_154 vgnd vpwr scs8hd_fill_1
XFILLER_0_187 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_top_track_0.LATCH_3_.latch data_in mem_top_track_0.LATCH_3_.latch/Q _092_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XFILLER_39_114 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_0_.latch data_in mem_bottom_track_9.LATCH_0_.latch/Q _144_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_136 vpwr vgnd scs8hd_fill_2
XFILLER_40_18 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_19 vpwr vgnd scs8hd_fill_2
XFILLER_14_52 vpwr vgnd scs8hd_fill_2
XFILLER_14_63 vpwr vgnd scs8hd_fill_2
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
XANTENNA__101__B _101_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_2_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 top_left_grid_pin_9_ mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_84 vgnd vpwr scs8hd_decap_3
XFILLER_41_175 vgnd vpwr scs8hd_decap_8
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_26_194 vgnd vpwr scs8hd_decap_8
XFILLER_26_161 vpwr vgnd scs8hd_fill_2
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_62 vpwr vgnd scs8hd_fill_2
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
X_195_ _195_/HI _195_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__112__A _152_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XFILLER_2_88 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_142 vgnd vpwr scs8hd_fill_1
Xmem_top_track_16.LATCH_0_.latch data_in mem_top_track_16.LATCH_0_.latch/Q _124_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_197 vpwr vgnd scs8hd_fill_2
XFILLER_11_75 vgnd vpwr scs8hd_decap_3
XFILLER_36_61 vgnd vpwr scs8hd_fill_1
XANTENNA__107__A _106_/X vgnd vpwr scs8hd_diode_2
XFILLER_14_175 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_178_ _178_/A _178_/Y vgnd vpwr scs8hd_inv_8
XFILLER_37_245 vgnd vpwr scs8hd_decap_12
XFILLER_28_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_5_.latch data_in mem_bottom_track_1.LATCH_5_.latch/Q _129_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_167 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_101_ _085_/B _101_/B _101_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_123 vpwr vgnd scs8hd_fill_2
XFILLER_11_134 vpwr vgnd scs8hd_fill_2
XFILLER_11_156 vgnd vpwr scs8hd_decap_3
XFILLER_22_96 vpwr vgnd scs8hd_fill_2
XFILLER_19_223 vgnd vpwr scs8hd_decap_12
XFILLER_19_245 vpwr vgnd scs8hd_fill_2
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_34_204 vgnd vpwr scs8hd_decap_8
XFILLER_8_32 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB _092_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_7_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__210__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_215 vgnd vpwr scs8hd_decap_4
XFILLER_16_248 vgnd vpwr scs8hd_decap_6
XFILLER_16_259 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _183_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_95 vpwr vgnd scs8hd_fill_2
XFILLER_33_62 vgnd vpwr scs8hd_fill_1
XFILLER_3_196 vgnd vpwr scs8hd_decap_8
XANTENNA__104__B address[4] vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _153_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_262 vpwr vgnd scs8hd_fill_2
XANTENNA__205__A _205_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_40 vgnd vpwr scs8hd_decap_4
XFILLER_12_251 vgnd vpwr scs8hd_decap_12
XANTENNA__115__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_5_88 vpwr vgnd scs8hd_fill_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_181 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_17.LATCH_0_.latch data_in mem_bottom_track_17.LATCH_0_.latch/Q _153_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_4_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_30_41 vgnd vpwr scs8hd_decap_3
XFILLER_5_269 vgnd vpwr scs8hd_decap_8
XFILLER_14_97 vpwr vgnd scs8hd_fill_2
XFILLER_39_83 vpwr vgnd scs8hd_fill_2
XFILLER_39_72 vgnd vpwr scs8hd_decap_8
XFILLER_30_85 vgnd vpwr scs8hd_decap_4
XFILLER_36_129 vpwr vgnd scs8hd_fill_2
XFILLER_29_170 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_3_ vgnd vpwr scs8hd_diode_2
XFILLER_35_162 vpwr vgnd scs8hd_fill_2
XFILLER_35_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_4_.scs8hd_inv_1 chanx_right_in[4] mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_143 vpwr vgnd scs8hd_fill_2
XFILLER_41_132 vpwr vgnd scs8hd_fill_2
XFILLER_41_110 vpwr vgnd scs8hd_fill_2
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr
+ scs8hd_diode_2
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_25_96 vpwr vgnd scs8hd_fill_2
XFILLER_25_52 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
X_194_ _194_/HI _194_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__112__B _109_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XFILLER_32_154 vgnd vpwr scs8hd_decap_8
XFILLER_32_198 vgnd vpwr scs8hd_decap_4
XFILLER_23_132 vpwr vgnd scs8hd_fill_2
XFILLER_23_154 vpwr vgnd scs8hd_fill_2
XANTENNA__213__A _213_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_36_84 vgnd vpwr scs8hd_decap_8
XFILLER_14_110 vpwr vgnd scs8hd_fill_2
XFILLER_14_154 vgnd vpwr scs8hd_decap_3
X_177_ _177_/A _177_/Y vgnd vpwr scs8hd_inv_8
XFILLER_14_187 vgnd vpwr scs8hd_decap_8
XFILLER_14_198 vgnd vpwr scs8hd_decap_12
XANTENNA__123__A _152_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
XFILLER_20_146 vgnd vpwr scs8hd_decap_4
XFILLER_9_180 vgnd vpwr scs8hd_decap_3
XFILLER_20_179 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A bottom_left_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_139 vgnd vpwr scs8hd_decap_12
XFILLER_7_128 vpwr vgnd scs8hd_fill_2
XFILLER_7_117 vgnd vpwr scs8hd_decap_4
XANTENNA__208__A right_top_grid_pin_10_ vgnd vpwr scs8hd_diode_2
XFILLER_11_168 vpwr vgnd scs8hd_fill_2
X_100_ _100_/A _101_/B vgnd vpwr scs8hd_buf_1
XFILLER_22_53 vpwr vgnd scs8hd_fill_2
XFILLER_19_235 vgnd vpwr scs8hd_decap_8
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A _117_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_88 vgnd vpwr scs8hd_decap_4
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_52 vgnd vpwr scs8hd_fill_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XFILLER_17_97 vpwr vgnd scs8hd_fill_2
XANTENNA__104__C _135_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__120__B _121_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_21_274 vgnd vpwr scs8hd_decap_3
Xmux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_3
XFILLER_0_167 vgnd vpwr scs8hd_decap_4
XANTENNA__221__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_4_.latch data_in mem_top_track_8.LATCH_4_.latch/Q _109_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_263 vgnd vpwr scs8hd_decap_12
XANTENNA__115__B _135_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_149 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__131__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_193 vgnd vpwr scs8hd_decap_12
XFILLER_30_64 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_top_track_16.LATCH_5_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA__216__A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_39_62 vpwr vgnd scs8hd_fill_2
XFILLER_36_108 vgnd vpwr scs8hd_decap_8
XFILLER_29_193 vpwr vgnd scs8hd_fill_2
XANTENNA__126__A _146_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_119 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_8
XPHY_75 vgnd vpwr scs8hd_decap_3
X_193_ _193_/HI _193_/LO vgnd vpwr scs8hd_conb_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XFILLER_17_141 vpwr vgnd scs8hd_fill_2
XFILLER_17_163 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_22 vpwr vgnd scs8hd_fill_2
XFILLER_11_99 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_track_1.LATCH_3_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_74 vgnd vpwr scs8hd_decap_8
X_176_ _176_/A _176_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__B _121_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
XFILLER_20_125 vpwr vgnd scs8hd_fill_2
XFILLER_28_203 vgnd vpwr scs8hd_decap_8
XANTENNA__224__A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_32 vpwr vgnd scs8hd_fill_2
XFILLER_22_76 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XFILLER_8_45 vgnd vpwr scs8hd_decap_4
X_159_ _154_/X _161_/B _157_/C _162_/D _159_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__134__A _101_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_3 vpwr vgnd scs8hd_fill_2
XFILLER_25_228 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_10 vgnd vpwr scs8hd_decap_4
XFILLER_17_65 vpwr vgnd scs8hd_fill_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_31 vpwr vgnd scs8hd_fill_2
XANTENNA__219__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__129__A _108_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_146 vgnd vpwr scs8hd_decap_8
XFILLER_0_179 vgnd vpwr scs8hd_decap_6
XFILLER_28_64 vpwr vgnd scs8hd_fill_2
XFILLER_8_202 vgnd vpwr scs8hd_decap_12
XANTENNA__131__B _131_/B vgnd vpwr scs8hd_diode_2
XANTENNA__115__C _135_/C vgnd vpwr scs8hd_diode_2
XFILLER_14_88 vgnd vpwr scs8hd_decap_4
XFILLER_39_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _111_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_5_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_175 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.INVTX1_5_.scs8hd_inv_1 bottom_left_grid_pin_3_ mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
X_192_ _192_/HI _192_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_14.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[3] mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_32_101 vpwr vgnd scs8hd_fill_2
XFILLER_17_175 vgnd vpwr scs8hd_decap_4
XANTENNA__137__A _154_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_56 vgnd vpwr scs8hd_decap_3
XFILLER_36_64 vgnd vpwr scs8hd_fill_1
XFILLER_36_42 vgnd vpwr scs8hd_fill_1
XFILLER_14_145 vpwr vgnd scs8hd_fill_2
X_175_ _175_/A _175_/Y vgnd vpwr scs8hd_inv_8
XFILLER_9_160 vgnd vpwr scs8hd_decap_12
XFILLER_20_104 vpwr vgnd scs8hd_fill_2
XFILLER_28_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_115 vgnd vpwr scs8hd_decap_4
XFILLER_22_88 vpwr vgnd scs8hd_fill_2
XFILLER_19_204 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_2_.scs8hd_inv_1/Y
+ _178_/A mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_19_215 vpwr vgnd scs8hd_fill_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
X_158_ address[0] _162_/D vgnd vpwr scs8hd_buf_1
X_089_ address[1] _093_/A vgnd vpwr scs8hd_inv_8
XANTENNA__134__B _131_/B vgnd vpwr scs8hd_diode_2
XANTENNA__150__A _110_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_262 vgnd vpwr scs8hd_decap_12
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_76 vpwr vgnd scs8hd_fill_2
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__129__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA__145__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_21_243 vgnd vpwr scs8hd_fill_1
XFILLER_28_32 vpwr vgnd scs8hd_fill_2
XFILLER_28_87 vgnd vpwr scs8hd_fill_1
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_12 vpwr vgnd scs8hd_fill_2
XFILLER_14_23 vpwr vgnd scs8hd_fill_2
XFILLER_14_56 vpwr vgnd scs8hd_fill_2
XFILLER_14_67 vgnd vpwr scs8hd_decap_6
XFILLER_30_77 vpwr vgnd scs8hd_fill_2
XFILLER_39_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__142__B _141_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_198 vgnd vpwr scs8hd_decap_3
XFILLER_35_110 vgnd vpwr scs8hd_decap_6
Xmux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _197_/HI mem_top_track_0.LATCH_2_.latch/Q
+ mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_41_102 vpwr vgnd scs8hd_fill_2
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_165 vgnd vpwr scs8hd_fill_1
XFILLER_25_22 vgnd vpwr scs8hd_decap_3
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vpwr vgnd scs8hd_fill_2
XFILLER_41_87 vpwr vgnd scs8hd_fill_2
X_191_ _191_/HI _191_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_220 vgnd vpwr scs8hd_decap_12
XFILLER_17_132 vgnd vpwr scs8hd_decap_3
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
XFILLER_32_124 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__137__B _168_/B vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _101_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_113 vgnd vpwr scs8hd_decap_4
XFILLER_23_179 vpwr vgnd scs8hd_fill_2
XFILLER_11_35 vpwr vgnd scs8hd_fill_2
XFILLER_36_32 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_0_.latch data_in mem_bottom_track_1.LATCH_0_.latch/Q _134_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_135 vgnd vpwr scs8hd_fill_1
XFILLER_14_168 vgnd vpwr scs8hd_decap_4
X_174_ _174_/A _174_/Y vgnd vpwr scs8hd_inv_8
XFILLER_28_7 vpwr vgnd scs8hd_fill_2
XANTENNA__148__A _108_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_172 vgnd vpwr scs8hd_decap_8
Xmux_right_track_12.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[1] mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_138 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_227 vgnd vpwr scs8hd_decap_12
XFILLER_3_80 vgnd vpwr scs8hd_fill_1
XFILLER_7_109 vpwr vgnd scs8hd_fill_2
XFILLER_11_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_4_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_249 vgnd vpwr scs8hd_decap_12
X_226_ _226_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
X_157_ _154_/X _161_/B _157_/C _161_/D _157_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_8_58 vgnd vpwr scs8hd_decap_12
XFILLER_40_6 vgnd vpwr scs8hd_decap_12
X_088_ _085_/B _109_/A _088_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__150__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_274 vgnd vpwr scs8hd_decap_3
XFILLER_18_271 vgnd vpwr scs8hd_decap_4
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_230 vgnd vpwr scs8hd_decap_12
XFILLER_16_219 vgnd vpwr scs8hd_fill_1
XFILLER_17_34 vpwr vgnd scs8hd_fill_2
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_55 vgnd vpwr scs8hd_decap_4
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_274 vgnd vpwr scs8hd_fill_1
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__161__A _161_/A vgnd vpwr scs8hd_diode_2
X_209_ _209_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_90 vpwr vgnd scs8hd_fill_2
XFILLER_21_266 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_104 vpwr vgnd scs8hd_fill_2
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XFILLER_5_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__156__A _171_/D vgnd vpwr scs8hd_diode_2
Xmux_right_track_10.tap_buf4_0_.scs8hd_inv_1 mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ _203_/A vgnd vpwr scs8hd_inv_1
XFILLER_38_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_35 vpwr vgnd scs8hd_fill_2
XFILLER_30_23 vpwr vgnd scs8hd_fill_2
XFILLER_39_32 vgnd vpwr scs8hd_decap_6
XFILLER_39_21 vgnd vpwr scs8hd_decap_4
XFILLER_39_10 vpwr vgnd scs8hd_fill_2
XFILLER_30_89 vgnd vpwr scs8hd_fill_1
XFILLER_39_87 vpwr vgnd scs8hd_fill_2
XFILLER_29_174 vgnd vpwr scs8hd_decap_3
XFILLER_29_163 vgnd vpwr scs8hd_fill_1
XFILLER_4_251 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 top_left_grid_pin_7_ mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_144 vgnd vpwr scs8hd_decap_3
XFILLER_6_91 vgnd vpwr scs8hd_fill_1
XFILLER_26_122 vgnd vpwr scs8hd_decap_8
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vpwr vgnd scs8hd_fill_2
XFILLER_41_136 vgnd vpwr scs8hd_decap_4
XFILLER_41_114 vpwr vgnd scs8hd_fill_2
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_26_177 vpwr vgnd scs8hd_fill_2
XFILLER_25_67 vpwr vgnd scs8hd_fill_2
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
X_190_ _190_/HI _190_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_232 vgnd vpwr scs8hd_decap_12
XFILLER_17_199 vpwr vgnd scs8hd_fill_2
XANTENNA__153__B _152_/B vgnd vpwr scs8hd_diode_2
XANTENNA__137__C _157_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _174_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_136 vgnd vpwr scs8hd_decap_6
XFILLER_23_158 vpwr vgnd scs8hd_fill_2
XFILLER_14_114 vpwr vgnd scs8hd_fill_2
X_173_ _173_/A _173_/Y vgnd vpwr scs8hd_inv_8
XFILLER_35_9 vgnd vpwr scs8hd_fill_1
XANTENNA__148__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__164__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_92 vpwr vgnd scs8hd_fill_2
XFILLER_28_239 vgnd vpwr scs8hd_decap_12
XFILLER_22_24 vgnd vpwr scs8hd_decap_4
XFILLER_22_57 vpwr vgnd scs8hd_fill_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
X_225_ chany_bottom_in[0] chany_top_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_6_154 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.INVTX1_7_.scs8hd_inv_1 bottom_left_grid_pin_11_ mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_156_ _171_/D _161_/D vgnd vpwr scs8hd_buf_1
X_087_ _087_/A _109_/A vgnd vpwr scs8hd_buf_1
XANTENNA__159__A _154_/X vgnd vpwr scs8hd_diode_2
XFILLER_33_253 vpwr vgnd scs8hd_fill_2
XFILLER_33_242 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[1] mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_10.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[2] mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_242 vgnd vpwr scs8hd_decap_12
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_33_89 vgnd vpwr scs8hd_decap_4
XFILLER_3_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_242 vpwr vgnd scs8hd_fill_2
XFILLER_15_253 vpwr vgnd scs8hd_fill_2
XANTENNA__161__B _161_/B vgnd vpwr scs8hd_diode_2
X_208_ right_top_grid_pin_10_ chanx_right_out[0] vgnd vpwr scs8hd_buf_2
X_139_ _108_/A _141_/B _139_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_4.tap_buf4_0_.scs8hd_inv_1 mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ _206_/A vgnd vpwr scs8hd_inv_1
XFILLER_31_3 vgnd vpwr scs8hd_decap_8
XFILLER_2_190 vgnd vpwr scs8hd_decap_12
XFILLER_21_223 vgnd vpwr scs8hd_decap_12
XFILLER_21_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_10.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_23 vpwr vgnd scs8hd_fill_2
XFILLER_28_12 vpwr vgnd scs8hd_fill_2
XFILLER_8_227 vgnd vpwr scs8hd_decap_12
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__172__A _154_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_142 vpwr vgnd scs8hd_fill_2
XFILLER_30_46 vgnd vpwr scs8hd_decap_3
XFILLER_5_208 vgnd vpwr scs8hd_decap_12
XANTENNA__082__A _082_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_197 vpwr vgnd scs8hd_fill_2
XFILLER_29_142 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_4_263 vgnd vpwr scs8hd_decap_12
XFILLER_35_123 vpwr vgnd scs8hd_fill_2
XANTENNA__167__A _154_/X vgnd vpwr scs8hd_diode_2
XFILLER_26_145 vgnd vpwr scs8hd_decap_8
XPHY_13 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A address[1] vgnd vpwr scs8hd_diode_2
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_17_112 vgnd vpwr scs8hd_decap_4
XFILLER_32_137 vpwr vgnd scs8hd_fill_2
XFILLER_17_156 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_0.LATCH_4_.latch data_in mem_top_track_0.LATCH_4_.latch/Q _088_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_26 vgnd vpwr scs8hd_decap_4
Xmem_bottom_track_9.LATCH_1_.latch data_in mem_bottom_track_9.LATCH_1_.latch/Q _143_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _183_/A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_172_ _154_/X _168_/B _106_/C address[0] _172_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _193_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_130 vpwr vgnd scs8hd_fill_2
XFILLER_9_141 vgnd vpwr scs8hd_fill_1
XFILLER_9_152 vpwr vgnd scs8hd_fill_2
XANTENNA__164__B _161_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_196 vgnd vpwr scs8hd_decap_12
XANTENNA__180__A _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[5] mux_right_track_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__090__A _093_/A vgnd vpwr scs8hd_diode_2
X_224_ chany_bottom_in[1] chany_top_out[2] vgnd vpwr scs8hd_buf_2
X_155_ _155_/A _161_/B vgnd vpwr scs8hd_buf_1
XFILLER_6_166 vgnd vpwr scs8hd_decap_12
XFILLER_6_133 vgnd vpwr scs8hd_decap_12
X_086_ address[1] _086_/B address[0] _087_/A vgnd vpwr scs8hd_or3_4
XFILLER_10_173 vgnd vpwr scs8hd_fill_1
XFILLER_33_7 vgnd vpwr scs8hd_decap_8
XFILLER_33_210 vgnd vpwr scs8hd_decap_12
XANTENNA__159__B _161_/B vgnd vpwr scs8hd_diode_2
XANTENNA__175__A _175_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_14 vgnd vpwr scs8hd_fill_1
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__085__A _108_/A vgnd vpwr scs8hd_diode_2
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_35 vpwr vgnd scs8hd_fill_2
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XFILLER_24_254 vgnd vpwr scs8hd_decap_12
XFILLER_17_69 vpwr vgnd scs8hd_fill_2
XFILLER_3_114 vgnd vpwr scs8hd_decap_8
XFILLER_3_147 vgnd vpwr scs8hd_decap_12
Xmem_top_track_16.LATCH_1_.latch data_in mem_top_track_16.LATCH_1_.latch/Q _123_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_207_ _207_/A chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_30_213 vgnd vpwr scs8hd_fill_1
XANTENNA__161__C _161_/C vgnd vpwr scs8hd_diode_2
X_138_ _137_/X _141_/B vgnd vpwr scs8hd_buf_1
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_24_3 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_2_.scs8hd_inv_1/Y
+ _176_/A mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_61 vgnd vpwr scs8hd_fill_1
XFILLER_0_94 vgnd vpwr scs8hd_decap_6
XFILLER_21_235 vgnd vpwr scs8hd_decap_8
XFILLER_0_128 vpwr vgnd scs8hd_fill_2
XFILLER_28_79 vpwr vgnd scs8hd_fill_2
XFILLER_28_46 vpwr vgnd scs8hd_fill_2
XFILLER_8_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_39 vgnd vpwr scs8hd_decap_12
Xmem_right_track_12.LATCH_0_.latch data_in _182_/A _168_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__172__B _168_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_45 vgnd vpwr scs8hd_decap_12
XFILLER_29_132 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_2_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_179 vpwr vgnd scs8hd_fill_2
XANTENNA__183__A _183_/A vgnd vpwr scs8hd_diode_2
XANTENNA__167__B _168_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_6_93 vgnd vpwr scs8hd_decap_3
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _226_/A vgnd vpwr scs8hd_inv_1
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_157 vpwr vgnd scs8hd_fill_2
XFILLER_25_14 vpwr vgnd scs8hd_fill_2
XANTENNA__077__B _086_/B vgnd vpwr scs8hd_diode_2
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XFILLER_34_190 vgnd vpwr scs8hd_fill_1
XANTENNA__093__A _093_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_245 vgnd vpwr scs8hd_decap_12
XFILLER_32_116 vgnd vpwr scs8hd_decap_8
XFILLER_32_105 vpwr vgnd scs8hd_fill_2
XFILLER_17_179 vgnd vpwr scs8hd_fill_1
XANTENNA__178__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_46 vgnd vpwr scs8hd_decap_8
XFILLER_36_13 vgnd vpwr scs8hd_decap_12
XANTENNA__088__A _085_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_57 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_127 vgnd vpwr scs8hd_decap_8
XFILLER_14_149 vgnd vpwr scs8hd_decap_4
X_171_ _154_/X _168_/B _106_/C _171_/D _171_/Y vgnd vpwr scs8hd_nor4_4
Xmem_bottom_track_17.LATCH_1_.latch data_in mem_bottom_track_17.LATCH_1_.latch/Q _152_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB _165_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__164__C _106_/C vgnd vpwr scs8hd_diode_2
XFILLER_20_108 vgnd vpwr scs8hd_decap_4
XFILLER_3_83 vgnd vpwr scs8hd_decap_4
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
XFILLER_11_119 vgnd vpwr scs8hd_fill_1
XFILLER_22_15 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__090__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_27_263 vgnd vpwr scs8hd_decap_12
Xmux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_2_.scs8hd_inv_1/Y
+ _182_/A mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_19_208 vgnd vpwr scs8hd_decap_4
XFILLER_19_219 vpwr vgnd scs8hd_fill_2
X_223_ chany_bottom_in[2] chany_top_out[3] vgnd vpwr scs8hd_buf_2
X_085_ _108_/A _085_/B _085_/Y vgnd vpwr scs8hd_nor2_4
X_154_ _154_/A _154_/X vgnd vpwr scs8hd_buf_1
XFILLER_6_178 vgnd vpwr scs8hd_decap_12
XFILLER_6_145 vgnd vpwr scs8hd_decap_8
XFILLER_10_163 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_222 vgnd vpwr scs8hd_decap_12
XANTENNA__159__C _157_/C vgnd vpwr scs8hd_diode_2
XFILLER_18_230 vgnd vpwr scs8hd_decap_12
XANTENNA__085__B _085_/B vgnd vpwr scs8hd_diode_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_266 vgnd vpwr scs8hd_decap_8
XFILLER_3_159 vgnd vpwr scs8hd_decap_12
XFILLER_30_203 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[6] mux_right_track_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_222 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.LATCH_0_.latch data_in _184_/A _170_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_206_ _206_/A chanx_right_out[2] vgnd vpwr scs8hd_buf_2
X_137_ _154_/A _168_/B _157_/C _137_/X vgnd vpwr scs8hd_or3_4
XFILLER_23_91 vpwr vgnd scs8hd_fill_2
XANTENNA__161__D _161_/D vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_60 vgnd vpwr scs8hd_fill_1
XANTENNA__186__A _186_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_36 vgnd vpwr scs8hd_fill_1
XANTENNA__096__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _180_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_5_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__172__C _106_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A top_left_grid_pin_9_ vgnd vpwr scs8hd_diode_2
XFILLER_14_16 vpwr vgnd scs8hd_fill_2
XFILLER_14_27 vpwr vgnd scs8hd_fill_2
XFILLER_39_68 vpwr vgnd scs8hd_fill_2
XFILLER_39_57 vgnd vpwr scs8hd_decap_4
XFILLER_29_166 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_10.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_158 vpwr vgnd scs8hd_fill_2
XANTENNA__167__C _161_/C vgnd vpwr scs8hd_diode_2
XFILLER_6_83 vpwr vgnd scs8hd_fill_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_25_48 vpwr vgnd scs8hd_fill_2
XPHY_15 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__077__C _171_/D vgnd vpwr scs8hd_diode_2
XPHY_26 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XANTENNA__093__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_257 vgnd vpwr scs8hd_decap_12
Xmem_top_track_8.LATCH_5_.latch data_in mem_top_track_8.LATCH_5_.latch/Q _108_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_31_172 vgnd vpwr scs8hd_decap_4
XFILLER_11_39 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A bottom_left_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_36 vgnd vpwr scs8hd_decap_6
XFILLER_36_25 vgnd vpwr scs8hd_decap_6
XANTENNA__088__B _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_183 vpwr vgnd scs8hd_fill_2
X_170_ _160_/A _155_/A _170_/C _162_/D _170_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_37_209 vgnd vpwr scs8hd_decap_12
XFILLER_13_172 vgnd vpwr scs8hd_decap_4
XFILLER_13_194 vpwr vgnd scs8hd_fill_2
XANTENNA__164__D _162_/D vgnd vpwr scs8hd_diode_2
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
XFILLER_3_51 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__090__C _171_/D vgnd vpwr scs8hd_diode_2
XANTENNA__099__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_27_275 vpwr vgnd scs8hd_fill_2
XFILLER_27_253 vpwr vgnd scs8hd_fill_2
XFILLER_27_242 vpwr vgnd scs8hd_fill_2
X_222_ _222_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
X_153_ _101_/B _152_/B _153_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_8_18 vgnd vpwr scs8hd_decap_12
XFILLER_10_120 vgnd vpwr scs8hd_decap_3
X_084_ _083_/X _085_/B vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__159__D _162_/D vgnd vpwr scs8hd_diode_2
XFILLER_18_242 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_2_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_245 vgnd vpwr scs8hd_decap_8
XFILLER_33_234 vgnd vpwr scs8hd_decap_8
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_6.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_33_48 vgnd vpwr scs8hd_decap_4
XFILLER_33_15 vgnd vpwr scs8hd_fill_1
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB _139_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XFILLER_15_234 vgnd vpwr scs8hd_decap_8
XFILLER_15_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_205_ _205_/A chanx_right_out[3] vgnd vpwr scs8hd_buf_2
X_136_ _135_/X _157_/C vgnd vpwr scs8hd_buf_1
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XFILLER_9_94 vpwr vgnd scs8hd_fill_2
XFILLER_21_204 vpwr vgnd scs8hd_fill_2
XFILLER_21_215 vpwr vgnd scs8hd_fill_2
XFILLER_0_108 vgnd vpwr scs8hd_decap_12
XFILLER_28_59 vgnd vpwr scs8hd_decap_3
XANTENNA__096__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_12_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _197_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _173_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__172__D address[0] vgnd vpwr scs8hd_diode_2
X_119_ _108_/A _121_/B _119_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_38_123 vgnd vpwr scs8hd_fill_1
Xmux_right_track_2.INVTX1_2_.scs8hd_inv_1 right_bottom_grid_pin_12_ mux_right_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_30_27 vpwr vgnd scs8hd_fill_2
XFILLER_14_39 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_101 vpwr vgnd scs8hd_fill_2
XFILLER_29_80 vpwr vgnd scs8hd_fill_2
XFILLER_20_71 vpwr vgnd scs8hd_fill_2
XFILLER_20_93 vpwr vgnd scs8hd_fill_2
XANTENNA__167__D _161_/D vgnd vpwr scs8hd_diode_2
XFILLER_41_118 vpwr vgnd scs8hd_fill_2
XFILLER_34_181 vgnd vpwr scs8hd_decap_3
XFILLER_25_27 vpwr vgnd scs8hd_fill_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XANTENNA__093__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_1_269 vgnd vpwr scs8hd_decap_8
XFILLER_9_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_4_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_137 vpwr vgnd scs8hd_fill_2
XFILLER_15_71 vgnd vpwr scs8hd_decap_4
XFILLER_31_92 vpwr vgnd scs8hd_fill_2
XFILLER_31_195 vpwr vgnd scs8hd_fill_2
XFILLER_31_184 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_173 vgnd vpwr scs8hd_fill_1
XFILLER_7_3 vpwr vgnd scs8hd_fill_2
XFILLER_9_111 vgnd vpwr scs8hd_decap_4
XFILLER_9_144 vgnd vpwr scs8hd_decap_8
XFILLER_13_184 vgnd vpwr scs8hd_fill_1
XFILLER_3_74 vgnd vpwr scs8hd_decap_6
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
XFILLER_3_96 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_4_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_28 vgnd vpwr scs8hd_fill_1
XFILLER_27_210 vgnd vpwr scs8hd_decap_12
XANTENNA__099__B address[2] vgnd vpwr scs8hd_diode_2
X_152_ _152_/A _152_/B _152_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_8.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_083_ _154_/A address[6] _161_/C _083_/X vgnd vpwr scs8hd_or3_4
X_221_ chany_bottom_in[4] chany_top_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_10_176 vgnd vpwr scs8hd_decap_12
XFILLER_12_50 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_37_91 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _177_/A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_202 vgnd vpwr scs8hd_decap_12
XFILLER_17_28 vgnd vpwr scs8hd_decap_4
X_204_ _204_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
XFILLER_15_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_135_ _135_/A _135_/B _135_/C _135_/X vgnd vpwr scs8hd_or3_4
XFILLER_2_150 vgnd vpwr scs8hd_decap_3
XFILLER_0_42 vgnd vpwr scs8hd_decap_4
XFILLER_0_53 vgnd vpwr scs8hd_decap_8
XFILLER_0_75 vgnd vpwr scs8hd_decap_12
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XFILLER_28_16 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__096__C _171_/D vgnd vpwr scs8hd_diode_2
XFILLER_12_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_271 vgnd vpwr scs8hd_decap_4
XFILLER_7_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
X_118_ _117_/X _121_/B vgnd vpwr scs8hd_buf_1
XFILLER_38_157 vgnd vpwr scs8hd_decap_12
XFILLER_38_146 vgnd vpwr scs8hd_decap_6
XFILLER_38_102 vpwr vgnd scs8hd_fill_2
Xmem_right_track_4.LATCH_0_.latch data_in _176_/A _162_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_3 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ _174_/A mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB _085_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_35_127 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_26_105 vpwr vgnd scs8hd_fill_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_25_171 vpwr vgnd scs8hd_fill_2
XFILLER_31_71 vpwr vgnd scs8hd_fill_2
XFILLER_15_83 vpwr vgnd scs8hd_fill_2
XFILLER_15_94 vpwr vgnd scs8hd_fill_2
XFILLER_16_182 vpwr vgnd scs8hd_fill_2
XFILLER_23_119 vgnd vpwr scs8hd_decap_3
XFILLER_11_19 vgnd vpwr scs8hd_fill_1
Xmux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _185_/A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _195_/HI _178_/Y mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_93 vgnd vpwr scs8hd_fill_1
XFILLER_9_156 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_211 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _194_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_222 vgnd vpwr scs8hd_decap_12
XANTENNA__099__C address[0] vgnd vpwr scs8hd_diode_2
X_220_ chany_bottom_in[5] chany_top_out[6] vgnd vpwr scs8hd_buf_2
X_151_ _111_/A _152_/B _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_188 vgnd vpwr scs8hd_decap_12
XFILLER_12_84 vgnd vpwr scs8hd_decap_8
X_082_ _082_/A _161_/C vgnd vpwr scs8hd_buf_1
Xmux_top_track_0.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[0] mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _198_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_258 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_269 vgnd vpwr scs8hd_decap_8
X_203_ _203_/A chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_23_72 vpwr vgnd scs8hd_fill_2
X_134_ _101_/B _131_/B _134_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_2_.scs8hd_inv_1/Y
+ _180_/A mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_1.LATCH_1_.latch data_in mem_bottom_track_1.LATCH_1_.latch/Q _133_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_6 vpwr vgnd scs8hd_fill_2
XFILLER_0_32 vgnd vpwr scs8hd_decap_3
XFILLER_0_87 vgnd vpwr scs8hd_decap_6
XFILLER_9_52 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_206 vgnd vpwr scs8hd_decap_8
XFILLER_12_239 vgnd vpwr scs8hd_decap_12
XFILLER_34_82 vpwr vgnd scs8hd_fill_2
XFILLER_7_232 vgnd vpwr scs8hd_decap_12
X_117_ _154_/A address[6] _170_/C _117_/X vgnd vpwr scs8hd_or3_4
XFILLER_38_169 vgnd vpwr scs8hd_decap_12
XFILLER_38_136 vgnd vpwr scs8hd_decap_4
XFILLER_15_3 vgnd vpwr scs8hd_fill_1
XFILLER_30_18 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _184_/A mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_202 vgnd vpwr scs8hd_decap_12
XFILLER_20_84 vpwr vgnd scs8hd_fill_2
XFILLER_26_139 vgnd vpwr scs8hd_decap_4
XFILLER_25_18 vpwr vgnd scs8hd_fill_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_25_194 vpwr vgnd scs8hd_fill_2
XFILLER_15_40 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__102__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_31_131 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB _163_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_72 vgnd vpwr scs8hd_decap_3
XFILLER_26_61 vpwr vgnd scs8hd_fill_2
XFILLER_13_120 vpwr vgnd scs8hd_fill_2
XFILLER_8_190 vgnd vpwr scs8hd_decap_12
XFILLER_22_19 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _179_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_245 vgnd vpwr scs8hd_decap_8
XFILLER_27_234 vgnd vpwr scs8hd_decap_8
X_150_ _110_/A _152_/B _150_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_112 vgnd vpwr scs8hd_decap_8
XFILLER_10_134 vpwr vgnd scs8hd_fill_2
XFILLER_10_145 vpwr vgnd scs8hd_fill_2
XFILLER_10_167 vgnd vpwr scs8hd_decap_6
XFILLER_12_63 vpwr vgnd scs8hd_fill_2
XFILLER_12_96 vgnd vpwr scs8hd_decap_6
X_081_ address[3] address[4] _135_/C _082_/A vgnd vpwr scs8hd_or3_4
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_71 vgnd vpwr scs8hd_decap_4
XFILLER_5_182 vgnd vpwr scs8hd_fill_1
XFILLER_33_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A top_left_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _174_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_204 vpwr vgnd scs8hd_fill_2
XFILLER_30_207 vgnd vpwr scs8hd_decap_6
X_202_ _202_/A chanx_right_out[6] vgnd vpwr scs8hd_buf_2
X_133_ _152_/A _131_/B _133_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_95 vgnd vpwr scs8hd_decap_4
XFILLER_2_130 vgnd vpwr scs8hd_decap_12
XANTENNA__110__A _110_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_84 vpwr vgnd scs8hd_fill_2
XANTENNA__105__A _105_/A vgnd vpwr scs8hd_diode_2
X_116_ _115_/X _170_/C vgnd vpwr scs8hd_buf_1
XFILLER_38_126 vgnd vpwr scs8hd_fill_1
XFILLER_39_28 vpwr vgnd scs8hd_fill_2
XFILLER_39_17 vpwr vgnd scs8hd_fill_2
XFILLER_29_159 vgnd vpwr scs8hd_decap_4
XFILLER_20_41 vpwr vgnd scs8hd_fill_2
XFILLER_35_118 vpwr vgnd scs8hd_fill_2
XFILLER_28_192 vpwr vgnd scs8hd_fill_2
XFILLER_6_87 vgnd vpwr scs8hd_decap_4
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XFILLER_34_151 vpwr vgnd scs8hd_fill_2
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmem_top_track_8.LATCH_0_.latch data_in mem_top_track_8.LATCH_0_.latch/Q _113_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_184 vgnd vpwr scs8hd_fill_1
XFILLER_25_140 vgnd vpwr scs8hd_fill_1
XFILLER_31_176 vgnd vpwr scs8hd_fill_1
XFILLER_31_154 vgnd vpwr scs8hd_fill_1
XFILLER_31_121 vgnd vpwr scs8hd_fill_1
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_210 vpwr vgnd scs8hd_fill_2
XFILLER_22_132 vpwr vgnd scs8hd_fill_2
XFILLER_22_143 vpwr vgnd scs8hd_fill_2
XFILLER_22_165 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _176_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_187 vpwr vgnd scs8hd_fill_2
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_84 vpwr vgnd scs8hd_fill_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_6
XFILLER_13_132 vgnd vpwr scs8hd_decap_4
XFILLER_13_198 vgnd vpwr scs8hd_decap_12
XANTENNA__113__A _101_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_202 vgnd vpwr scs8hd_fill_1
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
X_080_ enable _135_/C vgnd vpwr scs8hd_inv_8
Xmux_bottom_track_17.INVTX1_7_.scs8hd_inv_1 bottom_left_grid_pin_15_ mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XANTENNA__108__A _108_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_109 vgnd vpwr scs8hd_decap_3
Xmem_top_track_0.LATCH_5_.latch data_in mem_top_track_0.LATCH_5_.latch/Q _085_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_132_ _111_/A _131_/B _132_/Y vgnd vpwr scs8hd_nor2_4
X_201_ _201_/A chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_2_142 vgnd vpwr scs8hd_decap_8
Xmem_bottom_track_9.LATCH_2_.latch data_in mem_bottom_track_9.LATCH_2_.latch/Q _142_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__110__B _109_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_10 vgnd vpwr scs8hd_decap_12
XFILLER_9_65 vpwr vgnd scs8hd_fill_2
XFILLER_21_208 vgnd vpwr scs8hd_decap_4
XFILLER_21_219 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _175_/A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _174_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_230 vgnd vpwr scs8hd_decap_12
XANTENNA__211__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_63 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_11_241 vgnd vpwr scs8hd_decap_3
XFILLER_7_245 vgnd vpwr scs8hd_decap_12
X_115_ address[3] _135_/B _135_/C _115_/X vgnd vpwr scs8hd_or3_4
XANTENNA__121__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_138 vpwr vgnd scs8hd_fill_2
XFILLER_37_193 vpwr vgnd scs8hd_fill_2
XANTENNA__206__A _206_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_29_62 vgnd vpwr scs8hd_decap_4
XFILLER_29_40 vpwr vgnd scs8hd_fill_2
XFILLER_20_53 vpwr vgnd scs8hd_fill_2
XFILLER_20_64 vgnd vpwr scs8hd_decap_4
XFILLER_20_97 vpwr vgnd scs8hd_fill_2
XFILLER_29_84 vpwr vgnd scs8hd_fill_2
XFILLER_28_171 vgnd vpwr scs8hd_decap_6
XANTENNA__116__A _115_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_2_.latch data_in mem_top_track_16.LATCH_2_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_3 vgnd vpwr scs8hd_fill_1
XFILLER_34_174 vgnd vpwr scs8hd_decap_4
XFILLER_34_141 vgnd vpwr scs8hd_decap_8
XFILLER_19_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _196_/HI _183_/Y mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XFILLER_40_133 vgnd vpwr scs8hd_decap_8
XFILLER_25_152 vpwr vgnd scs8hd_fill_2
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
XFILLER_15_75 vgnd vpwr scs8hd_fill_1
XFILLER_16_130 vgnd vpwr scs8hd_decap_6
XFILLER_16_152 vgnd vpwr scs8hd_fill_1
XFILLER_31_199 vpwr vgnd scs8hd_fill_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _189_/HI vgnd vpwr
+ scs8hd_diode_2
.ends

