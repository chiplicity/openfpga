VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__1_
  CLASS BLOCK ;
  FOREIGN sb_0__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 2.400 4.040 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 2.400 10.840 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 2.400 18.320 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.390 137.600 2.670 140.000 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 2.400 25.800 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 137.600 7.270 140.000 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 2.400 ;
    END
  END address[6]
  PIN bottom_left_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 2.400 40.760 ;
    END
  END bottom_left_grid_pin_11_
  PIN bottom_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 137.600 17.390 140.000 ;
    END
  END bottom_left_grid_pin_13_
  PIN bottom_left_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.170 137.600 22.450 140.000 ;
    END
  END bottom_left_grid_pin_15_
  PIN bottom_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 4.800 140.000 5.400 ;
    END
  END bottom_left_grid_pin_1_
  PIN bottom_left_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 2.400 ;
    END
  END bottom_left_grid_pin_3_
  PIN bottom_left_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 2.400 33.280 ;
    END
  END bottom_left_grid_pin_5_
  PIN bottom_left_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 2.400 ;
    END
  END bottom_left_grid_pin_7_
  PIN bottom_left_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.050 137.600 12.330 140.000 ;
    END
  END bottom_left_grid_pin_9_
  PIN bottom_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 27.230 137.600 27.510 140.000 ;
    END
  END bottom_right_grid_pin_11_
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 14.320 140.000 14.920 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 24.520 140.000 25.120 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 2.400 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.290 137.600 32.570 140.000 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.350 137.600 37.630 140.000 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.950 137.600 42.230 140.000 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 34.720 140.000 35.320 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 44.240 140.000 44.840 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 2.400 48.240 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 2.400 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 47.010 137.600 47.290 140.000 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 52.070 137.600 52.350 140.000 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 2.400 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 57.130 137.600 57.410 140.000 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 54.440 140.000 55.040 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 2.400 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 64.640 140.000 65.240 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 62.190 137.600 62.470 140.000 ;
    END
  END chanx_right_out[8]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 2.400 55.040 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 2.400 62.520 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 2.400 70.000 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.250 137.600 67.530 140.000 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.310 137.600 72.590 140.000 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.910 137.600 77.190 140.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 2.400 77.480 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 2.400 84.960 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.970 137.600 82.250 140.000 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.030 137.600 87.310 140.000 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 74.840 140.000 75.440 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 84.360 140.000 84.960 ;
    END
  END chany_bottom_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 94.560 140.000 95.160 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 2.400 92.440 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 2.400 99.240 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 104.760 140.000 105.360 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 2.400 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 2.400 106.720 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 92.090 137.600 92.370 140.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 2.400 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 2.400 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.150 137.600 97.430 140.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.210 137.600 102.490 140.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.270 137.600 107.550 140.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 2.400 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 111.870 137.600 112.150 140.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 2.400 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.930 137.600 117.210 140.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 2.400 114.200 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.990 137.600 122.270 140.000 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 2.400 ;
    END
  END enable
  PIN right_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 2.400 121.680 ;
    END
  END right_bottom_grid_pin_12_
  PIN right_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 114.280 140.000 114.880 ;
    END
  END right_top_grid_pin_10_
  PIN top_left_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 2.400 ;
    END
  END top_left_grid_pin_11_
  PIN top_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 134.680 140.000 135.280 ;
    END
  END top_left_grid_pin_13_
  PIN top_left_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 2.400 129.160 ;
    END
  END top_left_grid_pin_15_
  PIN top_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.050 137.600 127.330 140.000 ;
    END
  END top_left_grid_pin_1_
  PIN top_left_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 132.110 137.600 132.390 140.000 ;
    END
  END top_left_grid_pin_3_
  PIN top_left_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 124.480 140.000 125.080 ;
    END
  END top_left_grid_pin_5_
  PIN top_left_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 2.400 ;
    END
  END top_left_grid_pin_7_
  PIN top_left_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 137.170 137.600 137.450 140.000 ;
    END
  END top_left_grid_pin_9_
  PIN top_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 2.400 136.640 ;
    END
  END top_right_grid_pin_11_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 0.070 0.380 138.390 137.660 ;
      LAYER met2 ;
        RECT 0.090 137.320 2.110 137.770 ;
        RECT 2.950 137.320 6.710 137.770 ;
        RECT 7.550 137.320 11.770 137.770 ;
        RECT 12.610 137.320 16.830 137.770 ;
        RECT 17.670 137.320 21.890 137.770 ;
        RECT 22.730 137.320 26.950 137.770 ;
        RECT 27.790 137.320 32.010 137.770 ;
        RECT 32.850 137.320 37.070 137.770 ;
        RECT 37.910 137.320 41.670 137.770 ;
        RECT 42.510 137.320 46.730 137.770 ;
        RECT 47.570 137.320 51.790 137.770 ;
        RECT 52.630 137.320 56.850 137.770 ;
        RECT 57.690 137.320 61.910 137.770 ;
        RECT 62.750 137.320 66.970 137.770 ;
        RECT 67.810 137.320 72.030 137.770 ;
        RECT 72.870 137.320 76.630 137.770 ;
        RECT 77.470 137.320 81.690 137.770 ;
        RECT 82.530 137.320 86.750 137.770 ;
        RECT 87.590 137.320 91.810 137.770 ;
        RECT 92.650 137.320 96.870 137.770 ;
        RECT 97.710 137.320 101.930 137.770 ;
        RECT 102.770 137.320 106.990 137.770 ;
        RECT 107.830 137.320 111.590 137.770 ;
        RECT 112.430 137.320 116.650 137.770 ;
        RECT 117.490 137.320 121.710 137.770 ;
        RECT 122.550 137.320 126.770 137.770 ;
        RECT 127.610 137.320 131.830 137.770 ;
        RECT 132.670 137.320 136.890 137.770 ;
        RECT 137.730 137.320 138.830 137.770 ;
        RECT 0.090 2.680 138.830 137.320 ;
        RECT 0.090 0.155 2.570 2.680 ;
        RECT 3.410 0.155 8.550 2.680 ;
        RECT 9.390 0.155 14.990 2.680 ;
        RECT 15.830 0.155 21.430 2.680 ;
        RECT 22.270 0.155 27.870 2.680 ;
        RECT 28.710 0.155 34.310 2.680 ;
        RECT 35.150 0.155 40.290 2.680 ;
        RECT 41.130 0.155 46.730 2.680 ;
        RECT 47.570 0.155 53.170 2.680 ;
        RECT 54.010 0.155 59.610 2.680 ;
        RECT 60.450 0.155 66.050 2.680 ;
        RECT 66.890 0.155 72.490 2.680 ;
        RECT 73.330 0.155 78.470 2.680 ;
        RECT 79.310 0.155 84.910 2.680 ;
        RECT 85.750 0.155 91.350 2.680 ;
        RECT 92.190 0.155 97.790 2.680 ;
        RECT 98.630 0.155 104.230 2.680 ;
        RECT 105.070 0.155 110.210 2.680 ;
        RECT 111.050 0.155 116.650 2.680 ;
        RECT 117.490 0.155 123.090 2.680 ;
        RECT 123.930 0.155 129.530 2.680 ;
        RECT 130.370 0.155 135.970 2.680 ;
        RECT 136.810 0.155 138.830 2.680 ;
      LAYER met3 ;
        RECT 2.800 135.680 138.855 136.040 ;
        RECT 2.800 135.640 137.200 135.680 ;
        RECT 0.270 134.280 137.200 135.640 ;
        RECT 0.270 129.560 138.855 134.280 ;
        RECT 2.800 128.160 138.855 129.560 ;
        RECT 0.270 125.480 138.855 128.160 ;
        RECT 0.270 124.080 137.200 125.480 ;
        RECT 0.270 122.080 138.855 124.080 ;
        RECT 2.800 120.680 138.855 122.080 ;
        RECT 0.270 115.280 138.855 120.680 ;
        RECT 0.270 114.600 137.200 115.280 ;
        RECT 2.800 113.880 137.200 114.600 ;
        RECT 2.800 113.200 138.855 113.880 ;
        RECT 0.270 107.120 138.855 113.200 ;
        RECT 2.800 105.760 138.855 107.120 ;
        RECT 2.800 105.720 137.200 105.760 ;
        RECT 0.270 104.360 137.200 105.720 ;
        RECT 0.270 99.640 138.855 104.360 ;
        RECT 2.800 98.240 138.855 99.640 ;
        RECT 0.270 95.560 138.855 98.240 ;
        RECT 0.270 94.160 137.200 95.560 ;
        RECT 0.270 92.840 138.855 94.160 ;
        RECT 2.800 91.440 138.855 92.840 ;
        RECT 0.270 85.360 138.855 91.440 ;
        RECT 2.800 83.960 137.200 85.360 ;
        RECT 0.270 77.880 138.855 83.960 ;
        RECT 2.800 76.480 138.855 77.880 ;
        RECT 0.270 75.840 138.855 76.480 ;
        RECT 0.270 74.440 137.200 75.840 ;
        RECT 0.270 70.400 138.855 74.440 ;
        RECT 2.800 69.000 138.855 70.400 ;
        RECT 0.270 65.640 138.855 69.000 ;
        RECT 0.270 64.240 137.200 65.640 ;
        RECT 0.270 62.920 138.855 64.240 ;
        RECT 2.800 61.520 138.855 62.920 ;
        RECT 0.270 55.440 138.855 61.520 ;
        RECT 2.800 54.040 137.200 55.440 ;
        RECT 0.270 48.640 138.855 54.040 ;
        RECT 2.800 47.240 138.855 48.640 ;
        RECT 0.270 45.240 138.855 47.240 ;
        RECT 0.270 43.840 137.200 45.240 ;
        RECT 0.270 41.160 138.855 43.840 ;
        RECT 2.800 39.760 138.855 41.160 ;
        RECT 0.270 35.720 138.855 39.760 ;
        RECT 0.270 34.320 137.200 35.720 ;
        RECT 0.270 33.680 138.855 34.320 ;
        RECT 2.800 32.280 138.855 33.680 ;
        RECT 0.270 26.200 138.855 32.280 ;
        RECT 2.800 25.520 138.855 26.200 ;
        RECT 2.800 24.800 137.200 25.520 ;
        RECT 0.270 24.120 137.200 24.800 ;
        RECT 0.270 18.720 138.855 24.120 ;
        RECT 2.800 17.320 138.855 18.720 ;
        RECT 0.270 15.320 138.855 17.320 ;
        RECT 0.270 13.920 137.200 15.320 ;
        RECT 0.270 11.240 138.855 13.920 ;
        RECT 2.800 9.840 138.855 11.240 ;
        RECT 0.270 5.800 138.855 9.840 ;
        RECT 0.270 4.440 137.200 5.800 ;
        RECT 2.800 4.400 137.200 4.440 ;
        RECT 2.800 3.040 138.855 4.400 ;
        RECT 0.270 0.175 138.855 3.040 ;
      LAYER met4 ;
        RECT 0.295 10.640 27.655 128.080 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 138.625 128.080 ;
  END
END sb_0__1_
END LIBRARY

