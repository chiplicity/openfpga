VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__0_
  CLASS BLOCK ;
  FOREIGN sb_0__0_ ;
  ORIGIN -0.005 0.000 ;
  SIZE 137.635 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.950 0.000 24.230 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.430 0.000 41.710 2.400 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.910 0.000 59.190 2.400 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.390 0.000 76.670 2.400 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.870 0.000 94.150 2.400 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 111.350 0.000 111.630 2.400 ;
    END
  END address[5]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 89.800 137.640 90.400 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 95.240 137.640 95.840 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 100.000 137.640 100.600 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 105.440 137.640 106.040 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 110.880 137.640 111.480 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 115.640 137.640 116.240 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 121.080 137.640 121.680 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 126.520 137.640 127.120 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 131.280 137.640 131.880 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.240 43.560 137.640 44.160 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.240 48.320 137.640 48.920 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.240 53.760 137.640 54.360 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.240 58.520 137.640 59.120 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.240 63.960 137.640 64.560 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.240 69.400 137.640 70.000 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.240 74.160 137.640 74.760 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.240 79.600 137.640 80.200 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.240 85.040 137.640 85.640 ;
    END
  END chanx_right_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.430 137.600 41.710 140.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.490 137.600 46.770 140.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.550 137.600 51.830 140.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.610 137.600 56.890 140.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.130 137.600 62.410 140.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.190 137.600 67.470 140.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.250 137.600 72.530 140.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.310 137.600 77.590 140.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 82.830 137.600 83.110 140.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.890 137.600 88.170 140.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.950 137.600 93.230 140.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.010 137.600 98.290 140.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.530 137.600 103.810 140.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.590 137.600 108.870 140.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.650 137.600 113.930 140.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 118.710 137.600 118.990 140.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.230 137.600 124.510 140.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.290 137.600 129.570 140.000 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 128.830 0.000 129.110 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.470 0.000 6.750 2.400 ;
    END
  END enable
  PIN right_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 27.920 137.640 28.520 ;
    END
  END right_bottom_grid_pin_11_
  PIN right_bottom_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 32.680 137.640 33.280 ;
    END
  END right_bottom_grid_pin_13_
  PIN right_bottom_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 38.120 137.640 38.720 ;
    END
  END right_bottom_grid_pin_15_
  PIN right_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 2.080 137.640 2.680 ;
    END
  END right_bottom_grid_pin_1_
  PIN right_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 6.840 137.640 7.440 ;
    END
  END right_bottom_grid_pin_3_
  PIN right_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 12.280 137.640 12.880 ;
    END
  END right_bottom_grid_pin_5_
  PIN right_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 17.040 137.640 17.640 ;
    END
  END right_bottom_grid_pin_7_
  PIN right_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 22.480 137.640 23.080 ;
    END
  END right_bottom_grid_pin_9_
  PIN right_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 136.720 137.640 137.320 ;
    END
  END right_top_grid_pin_10_
  PIN top_left_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.790 137.600 26.070 140.000 ;
    END
  END top_left_grid_pin_11_
  PIN top_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.850 137.600 31.130 140.000 ;
    END
  END top_left_grid_pin_13_
  PIN top_left_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.910 137.600 36.190 140.000 ;
    END
  END top_left_grid_pin_15_
  PIN top_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.030 137.600 0.310 140.000 ;
    END
  END top_left_grid_pin_1_
  PIN top_left_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.090 137.600 5.370 140.000 ;
    END
  END top_left_grid_pin_3_
  PIN top_left_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.150 137.600 10.430 140.000 ;
    END
  END top_left_grid_pin_5_
  PIN top_left_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.210 137.600 15.490 140.000 ;
    END
  END top_left_grid_pin_7_
  PIN top_left_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.730 137.600 21.010 140.000 ;
    END
  END top_left_grid_pin_9_
  PIN top_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 134.350 137.600 134.630 140.000 ;
    END
  END top_right_grid_pin_11_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 25.695 10.640 27.295 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 49.025 10.640 50.625 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 3.160 10.795 131.960 127.925 ;
      LAYER met1 ;
        RECT 3.160 10.640 134.650 128.080 ;
      LAYER met2 ;
        RECT 0.590 137.320 4.810 137.600 ;
        RECT 5.650 137.320 9.870 137.600 ;
        RECT 10.710 137.320 14.930 137.600 ;
        RECT 15.770 137.320 20.450 137.600 ;
        RECT 21.290 137.320 25.510 137.600 ;
        RECT 26.350 137.320 30.570 137.600 ;
        RECT 31.410 137.320 35.630 137.600 ;
        RECT 36.470 137.320 41.150 137.600 ;
        RECT 41.990 137.320 46.210 137.600 ;
        RECT 47.050 137.320 51.270 137.600 ;
        RECT 52.110 137.320 56.330 137.600 ;
        RECT 57.170 137.320 61.850 137.600 ;
        RECT 62.690 137.320 66.910 137.600 ;
        RECT 67.750 137.320 71.970 137.600 ;
        RECT 72.810 137.320 77.030 137.600 ;
        RECT 77.870 137.320 82.550 137.600 ;
        RECT 83.390 137.320 87.610 137.600 ;
        RECT 88.450 137.320 92.670 137.600 ;
        RECT 93.510 137.320 97.730 137.600 ;
        RECT 98.570 137.320 103.250 137.600 ;
        RECT 104.090 137.320 108.310 137.600 ;
        RECT 109.150 137.320 113.370 137.600 ;
        RECT 114.210 137.320 118.430 137.600 ;
        RECT 119.270 137.320 123.950 137.600 ;
        RECT 124.790 137.320 129.010 137.600 ;
        RECT 129.850 137.320 134.070 137.600 ;
        RECT 0.030 2.680 134.620 137.320 ;
        RECT 0.030 2.195 6.190 2.680 ;
        RECT 7.030 2.195 23.670 2.680 ;
        RECT 24.510 2.195 41.150 2.680 ;
        RECT 41.990 2.195 58.630 2.680 ;
        RECT 59.470 2.195 76.110 2.680 ;
        RECT 76.950 2.195 93.590 2.680 ;
        RECT 94.430 2.195 111.070 2.680 ;
        RECT 111.910 2.195 128.550 2.680 ;
        RECT 129.390 2.195 134.620 2.680 ;
      LAYER met3 ;
        RECT 0.005 136.320 134.840 137.185 ;
        RECT 0.005 132.280 135.240 136.320 ;
        RECT 0.005 130.880 134.840 132.280 ;
        RECT 0.005 127.520 135.240 130.880 ;
        RECT 0.005 126.120 134.840 127.520 ;
        RECT 0.005 122.080 135.240 126.120 ;
        RECT 0.005 120.680 134.840 122.080 ;
        RECT 0.005 116.640 135.240 120.680 ;
        RECT 0.005 115.240 134.840 116.640 ;
        RECT 0.005 111.880 135.240 115.240 ;
        RECT 0.005 110.480 134.840 111.880 ;
        RECT 0.005 106.440 135.240 110.480 ;
        RECT 0.005 105.040 134.840 106.440 ;
        RECT 0.005 101.000 135.240 105.040 ;
        RECT 0.005 99.600 134.840 101.000 ;
        RECT 0.005 96.240 135.240 99.600 ;
        RECT 0.005 94.840 134.840 96.240 ;
        RECT 0.005 90.800 135.240 94.840 ;
        RECT 0.005 89.400 134.840 90.800 ;
        RECT 0.005 86.040 135.240 89.400 ;
        RECT 0.005 84.640 134.840 86.040 ;
        RECT 0.005 80.600 135.240 84.640 ;
        RECT 0.005 79.200 134.840 80.600 ;
        RECT 0.005 75.160 135.240 79.200 ;
        RECT 0.005 73.760 134.840 75.160 ;
        RECT 0.005 70.400 135.240 73.760 ;
        RECT 0.005 69.000 134.840 70.400 ;
        RECT 0.005 64.960 135.240 69.000 ;
        RECT 0.005 63.560 134.840 64.960 ;
        RECT 0.005 59.520 135.240 63.560 ;
        RECT 0.005 58.120 134.840 59.520 ;
        RECT 0.005 54.760 135.240 58.120 ;
        RECT 0.005 53.360 134.840 54.760 ;
        RECT 0.005 49.320 135.240 53.360 ;
        RECT 0.005 47.920 134.840 49.320 ;
        RECT 0.005 44.560 135.240 47.920 ;
        RECT 0.005 43.160 134.840 44.560 ;
        RECT 0.005 39.120 135.240 43.160 ;
        RECT 0.005 37.720 134.840 39.120 ;
        RECT 0.005 33.680 135.240 37.720 ;
        RECT 0.005 32.280 134.840 33.680 ;
        RECT 0.005 28.920 135.240 32.280 ;
        RECT 0.005 27.520 134.840 28.920 ;
        RECT 0.005 23.480 135.240 27.520 ;
        RECT 0.005 22.080 134.840 23.480 ;
        RECT 0.005 18.040 135.240 22.080 ;
        RECT 0.005 16.640 134.840 18.040 ;
        RECT 0.005 13.280 135.240 16.640 ;
        RECT 0.005 11.880 134.840 13.280 ;
        RECT 0.005 7.840 135.240 11.880 ;
        RECT 0.005 6.440 134.840 7.840 ;
        RECT 0.005 3.080 135.240 6.440 ;
        RECT 0.005 2.215 134.840 3.080 ;
      LAYER met4 ;
        RECT 27.695 10.640 48.625 128.080 ;
        RECT 51.025 10.640 121.545 128.080 ;
  END
END sb_0__0_
END LIBRARY

