//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog netlist for pre-configured FPGA fabric by design: and2
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Wed Oct  7 01:24:55 2020
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

module and2_top_formal_verification (
input [0:0] a_fm,
input [0:0] b_fm,
output [0:0] out_c_fm);

// ----- Local wires for FPGA fabric -----
wire [0:0] set;
wire [0:0] reset;
wire [0:0] clk;
wire [0:95] gfpga_pad_GPIO_PAD;
wire [0:0] enable;
wire [0:15] address;
wire [0:0] data_in;

// ----- FPGA top-level module to be capsulated -----
	fpga_top U0_formal_verification (
		.set(set[0]),
		.reset(reset[0]),
		.clk(clk[0]),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[0:95]),
		.enable(enable[0]),
		.address(address[0:15]),
		.data_in(data_in[0]));

// ----- Begin Connect Global ports of FPGA top module -----
	assign set[0] = 1'b0;
	assign reset[0] = 1'b0;
// ----- End Connect Global ports of FPGA top module -----

// ----- Link BLIF Benchmark I/Os to FPGA I/Os -----
// ----- Blif Benchmark input a is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD[50] -----
	assign gfpga_pad_GPIO_PAD[50] = a_fm[0];
// ----- Blif Benchmark input b is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD[53] -----
	assign gfpga_pad_GPIO_PAD[53] = b_fm[0];
// ----- Blif Benchmark output out_c is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD[54] -----
	assign out_c_fm[0] = gfpga_pad_GPIO_PAD[54];

// ----- Wire unused FPGA I/Os to constants -----
	assign gfpga_pad_GPIO_PAD[0] = 1'b0;
	assign gfpga_pad_GPIO_PAD[1] = 1'b0;
	assign gfpga_pad_GPIO_PAD[2] = 1'b0;
	assign gfpga_pad_GPIO_PAD[3] = 1'b0;
	assign gfpga_pad_GPIO_PAD[4] = 1'b0;
	assign gfpga_pad_GPIO_PAD[5] = 1'b0;
	assign gfpga_pad_GPIO_PAD[6] = 1'b0;
	assign gfpga_pad_GPIO_PAD[7] = 1'b0;
	assign gfpga_pad_GPIO_PAD[8] = 1'b0;
	assign gfpga_pad_GPIO_PAD[9] = 1'b0;
	assign gfpga_pad_GPIO_PAD[10] = 1'b0;
	assign gfpga_pad_GPIO_PAD[11] = 1'b0;
	assign gfpga_pad_GPIO_PAD[12] = 1'b0;
	assign gfpga_pad_GPIO_PAD[13] = 1'b0;
	assign gfpga_pad_GPIO_PAD[14] = 1'b0;
	assign gfpga_pad_GPIO_PAD[15] = 1'b0;
	assign gfpga_pad_GPIO_PAD[16] = 1'b0;
	assign gfpga_pad_GPIO_PAD[17] = 1'b0;
	assign gfpga_pad_GPIO_PAD[18] = 1'b0;
	assign gfpga_pad_GPIO_PAD[19] = 1'b0;
	assign gfpga_pad_GPIO_PAD[20] = 1'b0;
	assign gfpga_pad_GPIO_PAD[21] = 1'b0;
	assign gfpga_pad_GPIO_PAD[22] = 1'b0;
	assign gfpga_pad_GPIO_PAD[23] = 1'b0;
	assign gfpga_pad_GPIO_PAD[24] = 1'b0;
	assign gfpga_pad_GPIO_PAD[25] = 1'b0;
	assign gfpga_pad_GPIO_PAD[26] = 1'b0;
	assign gfpga_pad_GPIO_PAD[27] = 1'b0;
	assign gfpga_pad_GPIO_PAD[28] = 1'b0;
	assign gfpga_pad_GPIO_PAD[29] = 1'b0;
	assign gfpga_pad_GPIO_PAD[30] = 1'b0;
	assign gfpga_pad_GPIO_PAD[31] = 1'b0;
	assign gfpga_pad_GPIO_PAD[32] = 1'b0;
	assign gfpga_pad_GPIO_PAD[33] = 1'b0;
	assign gfpga_pad_GPIO_PAD[34] = 1'b0;
	assign gfpga_pad_GPIO_PAD[35] = 1'b0;
	assign gfpga_pad_GPIO_PAD[36] = 1'b0;
	assign gfpga_pad_GPIO_PAD[37] = 1'b0;
	assign gfpga_pad_GPIO_PAD[38] = 1'b0;
	assign gfpga_pad_GPIO_PAD[39] = 1'b0;
	assign gfpga_pad_GPIO_PAD[40] = 1'b0;
	assign gfpga_pad_GPIO_PAD[41] = 1'b0;
	assign gfpga_pad_GPIO_PAD[42] = 1'b0;
	assign gfpga_pad_GPIO_PAD[43] = 1'b0;
	assign gfpga_pad_GPIO_PAD[44] = 1'b0;
	assign gfpga_pad_GPIO_PAD[45] = 1'b0;
	assign gfpga_pad_GPIO_PAD[46] = 1'b0;
	assign gfpga_pad_GPIO_PAD[47] = 1'b0;
	assign gfpga_pad_GPIO_PAD[48] = 1'b0;
	assign gfpga_pad_GPIO_PAD[49] = 1'b0;
	assign gfpga_pad_GPIO_PAD[51] = 1'b0;
	assign gfpga_pad_GPIO_PAD[52] = 1'b0;
	assign gfpga_pad_GPIO_PAD[55] = 1'b0;
	assign gfpga_pad_GPIO_PAD[56] = 1'b0;
	assign gfpga_pad_GPIO_PAD[57] = 1'b0;
	assign gfpga_pad_GPIO_PAD[58] = 1'b0;
	assign gfpga_pad_GPIO_PAD[59] = 1'b0;
	assign gfpga_pad_GPIO_PAD[60] = 1'b0;
	assign gfpga_pad_GPIO_PAD[61] = 1'b0;
	assign gfpga_pad_GPIO_PAD[62] = 1'b0;
	assign gfpga_pad_GPIO_PAD[63] = 1'b0;
	assign gfpga_pad_GPIO_PAD[64] = 1'b0;
	assign gfpga_pad_GPIO_PAD[65] = 1'b0;
	assign gfpga_pad_GPIO_PAD[66] = 1'b0;
	assign gfpga_pad_GPIO_PAD[67] = 1'b0;
	assign gfpga_pad_GPIO_PAD[68] = 1'b0;
	assign gfpga_pad_GPIO_PAD[69] = 1'b0;
	assign gfpga_pad_GPIO_PAD[70] = 1'b0;
	assign gfpga_pad_GPIO_PAD[71] = 1'b0;
	assign gfpga_pad_GPIO_PAD[72] = 1'b0;
	assign gfpga_pad_GPIO_PAD[73] = 1'b0;
	assign gfpga_pad_GPIO_PAD[74] = 1'b0;
	assign gfpga_pad_GPIO_PAD[75] = 1'b0;
	assign gfpga_pad_GPIO_PAD[76] = 1'b0;
	assign gfpga_pad_GPIO_PAD[77] = 1'b0;
	assign gfpga_pad_GPIO_PAD[78] = 1'b0;
	assign gfpga_pad_GPIO_PAD[79] = 1'b0;
	assign gfpga_pad_GPIO_PAD[80] = 1'b0;
	assign gfpga_pad_GPIO_PAD[81] = 1'b0;
	assign gfpga_pad_GPIO_PAD[82] = 1'b0;
	assign gfpga_pad_GPIO_PAD[83] = 1'b0;
	assign gfpga_pad_GPIO_PAD[84] = 1'b0;
	assign gfpga_pad_GPIO_PAD[85] = 1'b0;
	assign gfpga_pad_GPIO_PAD[86] = 1'b0;
	assign gfpga_pad_GPIO_PAD[87] = 1'b0;
	assign gfpga_pad_GPIO_PAD[88] = 1'b0;
	assign gfpga_pad_GPIO_PAD[89] = 1'b0;
	assign gfpga_pad_GPIO_PAD[90] = 1'b0;
	assign gfpga_pad_GPIO_PAD[91] = 1'b0;
	assign gfpga_pad_GPIO_PAD[92] = 1'b0;
	assign gfpga_pad_GPIO_PAD[93] = 1'b0;
	assign gfpga_pad_GPIO_PAD[94] = 1'b0;
	assign gfpga_pad_GPIO_PAD[95] = 1'b0;

// ----- Begin load bitstream to configuration memories -----
`ifdef ICARUS_SIMULATOR
// ----- Begin assign bitstream to configuration memories -----
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = 16'b1010101000000000;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b010;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7] = 8'b01000010;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7] = 8'b00101000;
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b0;
	assign U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.sb_0__0_.mem_top_track_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_12.mem_out[0:1] = 2'b01;
	assign U0_formal_verification.sb_0__0_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_0__1_.mem_top_track_8.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_0__1_.mem_top_track_16.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_0__1_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_0__2_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_0__2_.mem_top_track_8.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_0__2_.mem_top_track_16.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_0__2_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_17.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_0__3_.mem_right_track_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__3_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.sb_1__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_8.mem_out[0:1] = 2'b01;
	assign U0_formal_verification.sb_1__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_16.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.sb_1__0_.mem_right_track_0.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_1__0_.mem_right_track_8.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_1__0_.mem_right_track_16.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_1__0_.mem_left_track_1.mem_out[0:5] = 6'b100001;
	assign U0_formal_verification.sb_1__0_.mem_left_track_9.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_1__0_.mem_left_track_17.mem_out[0:5] = 6'b010100;
	assign U0_formal_verification.sb_1__1_.mem_top_track_0.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_1__1_.mem_top_track_8.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_1__1_.mem_top_track_16.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_1__1_.mem_right_track_0.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_1__1_.mem_right_track_8.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_1__1_.mem_right_track_16.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_out[0:7] = 8'b01000100;
	assign U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_1__1_.mem_left_track_1.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_1__1_.mem_left_track_9.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_1__1_.mem_left_track_17.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_1__2_.mem_top_track_0.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_1__2_.mem_top_track_8.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_1__2_.mem_top_track_16.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_1__2_.mem_right_track_0.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_1__2_.mem_right_track_8.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_1__2_.mem_right_track_16.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_1__2_.mem_left_track_1.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_1__2_.mem_left_track_9.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_1__2_.mem_left_track_17.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_1__3_.mem_right_track_0.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_1__3_.mem_right_track_8.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_1__3_.mem_right_track_16.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_1__3_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__3_.mem_left_track_1.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_1__3_.mem_left_track_9.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_1__3_.mem_left_track_17.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_2__0_.mem_top_track_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.sb_2__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_16.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.sb_2__0_.mem_right_track_0.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_2__0_.mem_right_track_8.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_2__0_.mem_right_track_16.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_2__0_.mem_left_track_1.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_2__0_.mem_left_track_9.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_2__0_.mem_left_track_17.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_2__1_.mem_top_track_0.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_2__1_.mem_top_track_8.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_2__1_.mem_top_track_16.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_2__1_.mem_right_track_0.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_2__1_.mem_right_track_8.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_2__1_.mem_right_track_16.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_2__1_.mem_left_track_1.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_2__1_.mem_left_track_9.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_2__1_.mem_left_track_17.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_2__2_.mem_top_track_0.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_2__2_.mem_top_track_8.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_2__2_.mem_top_track_16.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_2__2_.mem_right_track_0.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_2__2_.mem_right_track_8.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_2__2_.mem_right_track_16.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_2__2_.mem_left_track_1.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_2__2_.mem_left_track_9.mem_out[0:7] = 8'b00000001;
	assign U0_formal_verification.sb_2__2_.mem_left_track_17.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_2__3_.mem_right_track_0.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_2__3_.mem_right_track_8.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_2__3_.mem_right_track_16.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_2__3_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__3_.mem_left_track_1.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_2__3_.mem_left_track_9.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_2__3_.mem_left_track_17.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_3__0_.mem_top_track_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__0_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_3__1_.mem_top_track_8.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_3__1_.mem_top_track_16.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_3__1_.mem_bottom_track_1.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_3__1_.mem_bottom_track_9.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_3__1_.mem_bottom_track_17.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_3__1_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__1_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_top_track_0.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_3__2_.mem_top_track_8.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_3__2_.mem_top_track_16.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_3__2_.mem_bottom_track_1.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_3__2_.mem_bottom_track_9.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_3__2_.mem_bottom_track_17.mem_out[0:5] = 6'b001001;
	assign U0_formal_verification.sb_3__2_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__2_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_3__3_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_out[0:5] = 6'b010100;
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_out[0:5] = 6'b001010;
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_1__3_.mem_bottom_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__3_.mem_bottom_ipin_1.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__3_.mem_bottom_ipin_2.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__3_.mem_bottom_ipin_3.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__3_.mem_bottom_ipin_4.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__3_.mem_bottom_ipin_5.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__3_.mem_bottom_ipin_6.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__3_.mem_bottom_ipin_7.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__3_.mem_top_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_1__3_.mem_top_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_1__3_.mem_top_ipin_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_2__3_.mem_bottom_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__3_.mem_bottom_ipin_1.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__3_.mem_bottom_ipin_2.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__3_.mem_bottom_ipin_3.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__3_.mem_bottom_ipin_4.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__3_.mem_bottom_ipin_5.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__3_.mem_bottom_ipin_6.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__3_.mem_bottom_ipin_7.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__3_.mem_top_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_2__3_.mem_top_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_2__3_.mem_top_ipin_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_3__0_.mem_bottom_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__0_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_3__0_.mem_bottom_ipin_2.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__0_.mem_top_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__0_.mem_top_ipin_1.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__0_.mem_top_ipin_2.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__0_.mem_top_ipin_3.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__0_.mem_top_ipin_4.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__0_.mem_top_ipin_5.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__0_.mem_top_ipin_6.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__0_.mem_top_ipin_7.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__1_.mem_bottom_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__1_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_3__1_.mem_bottom_ipin_2.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__1_.mem_top_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__1_.mem_top_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_3__1_.mem_top_ipin_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_3__2_.mem_bottom_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__2_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_3__2_.mem_bottom_ipin_2.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__2_.mem_top_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__2_.mem_top_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_3__2_.mem_top_ipin_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_3__3_.mem_bottom_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__3_.mem_bottom_ipin_1.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__3_.mem_bottom_ipin_2.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__3_.mem_bottom_ipin_3.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__3_.mem_bottom_ipin_4.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__3_.mem_bottom_ipin_5.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__3_.mem_bottom_ipin_6.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__3_.mem_bottom_ipin_7.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__3_.mem_top_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cbx_3__3_.mem_top_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_3__3_.mem_top_ipin_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__1_.mem_left_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__1_.mem_right_ipin_1.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__1_.mem_right_ipin_2.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__1_.mem_right_ipin_3.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__1_.mem_right_ipin_4.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__1_.mem_right_ipin_5.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__1_.mem_right_ipin_6.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__1_.mem_right_ipin_7.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__2_.mem_left_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__2_.mem_right_ipin_1.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__2_.mem_right_ipin_2.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__2_.mem_right_ipin_3.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__2_.mem_right_ipin_4.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__2_.mem_right_ipin_5.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__2_.mem_right_ipin_6.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__2_.mem_right_ipin_7.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__3_.mem_left_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__3_.mem_left_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_0__3_.mem_right_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__3_.mem_right_ipin_1.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__3_.mem_right_ipin_2.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__3_.mem_right_ipin_3.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__3_.mem_right_ipin_4.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__3_.mem_right_ipin_5.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__3_.mem_right_ipin_6.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_0__3_.mem_right_ipin_7.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_1__1_.mem_left_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_1__1_.mem_left_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_1__2_.mem_left_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_1__3_.mem_left_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_1__3_.mem_left_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_1__3_.mem_right_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_1__3_.mem_right_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_1__3_.mem_right_ipin_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_2__1_.mem_left_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_2__2_.mem_left_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_2__3_.mem_left_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_2__3_.mem_left_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_2__3_.mem_right_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_2__3_.mem_right_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_2__3_.mem_right_ipin_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_3__1_.mem_left_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__1_.mem_left_ipin_1.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__1_.mem_left_ipin_2.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__1_.mem_left_ipin_3.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__1_.mem_left_ipin_4.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__1_.mem_left_ipin_5.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__1_.mem_left_ipin_6.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__1_.mem_left_ipin_7.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__1_.mem_right_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__1_.mem_right_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_3__1_.mem_right_ipin_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_3__2_.mem_left_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__2_.mem_left_ipin_1.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__2_.mem_left_ipin_2.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__2_.mem_left_ipin_3.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__2_.mem_left_ipin_4.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__2_.mem_left_ipin_5.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__2_.mem_left_ipin_6.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__2_.mem_left_ipin_7.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__2_.mem_right_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__2_.mem_right_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_3__2_.mem_right_ipin_2.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_3__3_.mem_left_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__3_.mem_left_ipin_1.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__3_.mem_left_ipin_2.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__3_.mem_left_ipin_3.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__3_.mem_left_ipin_4.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__3_.mem_left_ipin_5.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__3_.mem_left_ipin_6.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__3_.mem_left_ipin_7.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__3_.mem_right_ipin_0.mem_out[0:5] = 6'b000001;
	assign U0_formal_verification.cby_3__3_.mem_right_ipin_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cby_3__3_.mem_right_ipin_2.mem_out[0:1] = {2{1'b0}};
initial begin
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = 16'b0101010111111111;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7] = 8'b10111101;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.sb_0__0_.mem_top_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_12.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_0__1_.mem_top_track_8.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_0__1_.mem_top_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_0__1_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_0__2_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_0__2_.mem_top_track_8.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_0__2_.mem_top_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_0__2_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_0__3_.mem_right_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_8.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_16.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__0_.mem_right_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__0_.mem_right_track_8.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__0_.mem_right_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__0_.mem_left_track_1.mem_outb[0:5] = 6'b011110;
	force U0_formal_verification.sb_1__0_.mem_left_track_9.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__0_.mem_left_track_17.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_1__1_.mem_top_track_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__1_.mem_top_track_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__1_.mem_top_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__1_.mem_right_track_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__1_.mem_right_track_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__1_.mem_right_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__1_.mem_left_track_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__1_.mem_left_track_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__1_.mem_left_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__2_.mem_top_track_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__2_.mem_top_track_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__2_.mem_top_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__2_.mem_right_track_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__2_.mem_right_track_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__2_.mem_right_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__2_.mem_left_track_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__2_.mem_left_track_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__2_.mem_left_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__3_.mem_right_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__3_.mem_right_track_8.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__3_.mem_right_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_1.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__3_.mem_left_track_9.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_1__3_.mem_left_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__0_.mem_top_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_2__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_16.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_2__0_.mem_right_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__0_.mem_right_track_8.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__0_.mem_right_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__0_.mem_left_track_1.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__0_.mem_left_track_9.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__0_.mem_left_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__1_.mem_top_track_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__1_.mem_top_track_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__1_.mem_top_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__1_.mem_right_track_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__1_.mem_right_track_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__1_.mem_right_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__1_.mem_left_track_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__1_.mem_left_track_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__1_.mem_left_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__2_.mem_top_track_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__2_.mem_top_track_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__2_.mem_top_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__2_.mem_right_track_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__2_.mem_right_track_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__2_.mem_right_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__2_.mem_left_track_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__2_.mem_left_track_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__2_.mem_left_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__3_.mem_right_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__3_.mem_right_track_8.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__3_.mem_right_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_1.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__3_.mem_left_track_9.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_2__3_.mem_left_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__0_.mem_top_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__1_.mem_top_track_8.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__1_.mem_top_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_1.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_9.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__1_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_0.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__2_.mem_top_track_8.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__2_.mem_top_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_1.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_9.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_17.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_3__2_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_outb[0:5] = 6'b110101;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__3_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__3_.mem_bottom_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__3_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__3_.mem_bottom_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__3_.mem_bottom_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__3_.mem_bottom_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__3_.mem_bottom_ipin_6.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__3_.mem_bottom_ipin_7.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_2__3_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__3_.mem_bottom_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__3_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__3_.mem_bottom_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__3_.mem_bottom_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__3_.mem_bottom_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__3_.mem_bottom_ipin_6.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__3_.mem_bottom_ipin_7.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_6.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_7.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__2_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_3__3_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__3_.mem_bottom_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__3_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__3_.mem_bottom_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__3_.mem_bottom_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__3_.mem_bottom_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__3_.mem_bottom_ipin_6.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__3_.mem_bottom_ipin_7.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_6.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_7.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_6.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_7.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__3_.mem_left_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__3_.mem_left_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_6.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__3_.mem_right_ipin_7.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_1__1_.mem_left_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_1__1_.mem_left_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_1__3_.mem_left_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_1__3_.mem_left_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_1__3_.mem_right_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_2__3_.mem_left_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__3_.mem_left_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__3_.mem_right_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_left_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__1_.mem_left_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__1_.mem_left_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__1_.mem_left_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__1_.mem_left_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__1_.mem_left_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__1_.mem_left_ipin_6.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__1_.mem_left_ipin_7.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__1_.mem_right_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__1_.mem_right_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_6.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_7.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__2_.mem_right_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_3__3_.mem_left_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__3_.mem_left_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__3_.mem_left_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__3_.mem_left_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__3_.mem_left_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__3_.mem_left_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__3_.mem_left_ipin_6.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__3_.mem_left_ipin_7.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__3_.mem_right_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_3__3_.mem_right_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_2.mem_outb[0:1] = {2{1'b1}};
end
// ----- End assign bitstream to configuration memories -----
`else
// ----- Begin deposit bitstream to configuration memories -----
initial begin
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], 16'b1010101000000000);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], 16'b0101010111111111);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b010);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b101);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7], 8'b01000010);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7], 8'b10111101);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7], 8'b00101000);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7], 8'b11010111);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_1__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_2__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_3__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_4__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_4.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_4.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_6.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_6.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_8.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_8.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_10.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_10.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_12.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_12.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_14.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_16.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_4.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_4.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_6.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_6.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_8.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_8.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_10.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_10.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_12.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_12.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_14.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_16.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_0.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_0.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_8.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_8.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_16.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_16.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_4.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_4.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_6.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_6.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_8.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_8.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_10.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_10.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_12.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_12.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_14.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_0__2_.mem_top_track_0.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_0__2_.mem_top_track_0.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_0__2_.mem_top_track_8.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_0__2_.mem_top_track_8.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_0__2_.mem_top_track_16.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_0__2_.mem_top_track_16.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_4.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_4.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_6.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_6.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_8.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_8.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_10.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_10.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_12.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_12.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_14.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_17.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_17.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_4.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_4.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_6.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_6.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_8.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_8.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_10.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_10.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_12.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_12.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_14.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_right_track_16.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_3.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_3.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_5.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_5.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_7.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_7.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_9.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_9.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_11.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_11.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_13.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_15.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__3_.mem_bottom_track_17.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_8.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_8.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_14.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_16.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_16.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_0.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_0.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_8.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_8.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_16.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_16.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_1.mem_out[0:5], 6'b100001);
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_1.mem_outb[0:5], 6'b011110);
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_9.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_9.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_17.mem_out[0:5], 6'b010100);
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_17.mem_outb[0:5], 6'b101011);
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_0.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_0.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_8.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_8.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_16.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_16.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_0.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_0.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_8.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_8.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_16.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_16.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_out[0:7], 8'b01000100);
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_outb[0:7], 8'b10111011);
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_1.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_1.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_9.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_9.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_17.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_17.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_1__2_.mem_top_track_0.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_1__2_.mem_top_track_0.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_1__2_.mem_top_track_8.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_1__2_.mem_top_track_8.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_1__2_.mem_top_track_16.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_1__2_.mem_top_track_16.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_0.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_0.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_8.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_8.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_16.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_16.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_1.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_1.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_9.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_9.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_17.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_17.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_1__3_.mem_right_track_0.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_1__3_.mem_right_track_0.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_1__3_.mem_right_track_8.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_1__3_.mem_right_track_8.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_1__3_.mem_right_track_16.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_1__3_.mem_right_track_16.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_3.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_3.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_5.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_5.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_7.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_7.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_9.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_9.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_11.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_11.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_13.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_15.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__3_.mem_bottom_track_17.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__3_.mem_left_track_1.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_1__3_.mem_left_track_1.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_1__3_.mem_left_track_9.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_1__3_.mem_left_track_9.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_1__3_.mem_left_track_17.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_1__3_.mem_left_track_17.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_8.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_8.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_14.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_16.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_16.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.sb_2__0_.mem_right_track_0.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_2__0_.mem_right_track_0.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_2__0_.mem_right_track_8.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_2__0_.mem_right_track_8.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_2__0_.mem_right_track_16.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_2__0_.mem_right_track_16.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_1.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_1.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_9.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_9.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_17.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_17.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_0.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_0.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_8.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_8.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_16.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_16.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_2__1_.mem_right_track_0.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_2__1_.mem_right_track_0.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_2__1_.mem_right_track_8.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_2__1_.mem_right_track_8.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_2__1_.mem_right_track_16.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_2__1_.mem_right_track_16.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_1.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_1.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_9.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_9.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_17.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_17.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_2__2_.mem_top_track_0.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_2__2_.mem_top_track_0.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_2__2_.mem_top_track_8.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_2__2_.mem_top_track_8.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_2__2_.mem_top_track_16.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_2__2_.mem_top_track_16.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_2__2_.mem_right_track_0.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_2__2_.mem_right_track_0.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_2__2_.mem_right_track_8.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_2__2_.mem_right_track_8.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_2__2_.mem_right_track_16.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_2__2_.mem_right_track_16.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_1.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_1.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_9.mem_out[0:7], 8'b00000001);
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_9.mem_outb[0:7], 8'b11111110);
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_17.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_17.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_2__3_.mem_right_track_0.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_2__3_.mem_right_track_0.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_2__3_.mem_right_track_8.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_2__3_.mem_right_track_8.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_2__3_.mem_right_track_16.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_2__3_.mem_right_track_16.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_3.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_3.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_5.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_5.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_7.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_7.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_9.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_9.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_11.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_11.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_13.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_15.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__3_.mem_bottom_track_17.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__3_.mem_left_track_1.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_2__3_.mem_left_track_1.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_2__3_.mem_left_track_9.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_2__3_.mem_left_track_9.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_2__3_.mem_left_track_17.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_2__3_.mem_left_track_17.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_4.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_4.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_6.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_6.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_8.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_8.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_10.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_10.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_12.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_12.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_14.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_top_track_16.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_3.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_3.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_5.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_5.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_7.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_7.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_9.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_9.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_11.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_11.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_13.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_15.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__0_.mem_left_track_17.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__1_.mem_top_track_0.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_3__1_.mem_top_track_0.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_3__1_.mem_top_track_8.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_3__1_.mem_top_track_8.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_3__1_.mem_top_track_16.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_3__1_.mem_top_track_16.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_3__1_.mem_bottom_track_1.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_3__1_.mem_bottom_track_1.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_3__1_.mem_bottom_track_9.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_3__1_.mem_bottom_track_9.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_3__1_.mem_bottom_track_17.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_3__1_.mem_bottom_track_17.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_3.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_3.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_5.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_5.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_7.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_7.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_9.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_9.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_11.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_11.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_13.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_15.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__1_.mem_left_track_17.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__2_.mem_top_track_0.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_3__2_.mem_top_track_0.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_3__2_.mem_top_track_8.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_3__2_.mem_top_track_8.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_3__2_.mem_top_track_16.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_3__2_.mem_top_track_16.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_3__2_.mem_bottom_track_1.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_3__2_.mem_bottom_track_1.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_3__2_.mem_bottom_track_9.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_3__2_.mem_bottom_track_9.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_3__2_.mem_bottom_track_17.mem_out[0:5], 6'b001001);
	$deposit(U0_formal_verification.sb_3__2_.mem_bottom_track_17.mem_outb[0:5], 6'b110110);
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_3.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_3.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_5.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_5.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_7.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_7.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_9.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_9.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_11.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_11.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_13.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_15.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__2_.mem_left_track_17.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_3.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_3.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_5.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_5.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_7.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_7.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_9.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_9.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_11.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_11.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_13.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_15.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_bottom_track_17.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_3.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_3.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_5.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_5.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_7.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_7.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_9.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_9.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_11.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_11.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_13.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_15.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_3__3_.mem_left_track_17.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_out[0:5], 6'b010100);
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_outb[0:5], 6'b101011);
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_out[0:5], 6'b001010);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_outb[0:5], 6'b110101);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_1__3_.mem_bottom_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__3_.mem_bottom_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__3_.mem_bottom_ipin_1.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__3_.mem_bottom_ipin_1.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__3_.mem_bottom_ipin_2.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__3_.mem_bottom_ipin_2.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__3_.mem_bottom_ipin_3.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__3_.mem_bottom_ipin_3.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__3_.mem_bottom_ipin_4.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__3_.mem_bottom_ipin_4.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__3_.mem_bottom_ipin_5.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__3_.mem_bottom_ipin_5.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__3_.mem_bottom_ipin_6.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__3_.mem_bottom_ipin_6.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__3_.mem_bottom_ipin_7.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__3_.mem_bottom_ipin_7.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_1__3_.mem_top_ipin_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_2__3_.mem_bottom_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__3_.mem_bottom_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__3_.mem_bottom_ipin_1.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__3_.mem_bottom_ipin_1.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__3_.mem_bottom_ipin_2.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__3_.mem_bottom_ipin_2.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__3_.mem_bottom_ipin_3.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__3_.mem_bottom_ipin_3.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__3_.mem_bottom_ipin_4.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__3_.mem_bottom_ipin_4.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__3_.mem_bottom_ipin_5.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__3_.mem_bottom_ipin_5.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__3_.mem_bottom_ipin_6.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__3_.mem_bottom_ipin_6.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__3_.mem_bottom_ipin_7.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__3_.mem_bottom_ipin_7.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_2__3_.mem_top_ipin_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_3__0_.mem_bottom_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__0_.mem_bottom_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__0_.mem_bottom_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_3__0_.mem_bottom_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_3__0_.mem_bottom_ipin_2.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__0_.mem_bottom_ipin_2.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_1.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_1.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_2.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_2.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_3.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_3.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_4.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_4.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_5.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_5.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_6.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_6.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_7.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__0_.mem_top_ipin_7.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__1_.mem_bottom_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__1_.mem_bottom_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__1_.mem_bottom_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_3__1_.mem_bottom_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_3__1_.mem_bottom_ipin_2.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__1_.mem_bottom_ipin_2.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_3__1_.mem_top_ipin_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_bottom_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__2_.mem_bottom_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__2_.mem_bottom_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_bottom_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_bottom_ipin_2.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__2_.mem_bottom_ipin_2.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_3__2_.mem_top_ipin_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_3__3_.mem_bottom_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__3_.mem_bottom_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__3_.mem_bottom_ipin_1.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__3_.mem_bottom_ipin_1.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__3_.mem_bottom_ipin_2.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__3_.mem_bottom_ipin_2.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__3_.mem_bottom_ipin_3.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__3_.mem_bottom_ipin_3.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__3_.mem_bottom_ipin_4.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__3_.mem_bottom_ipin_4.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__3_.mem_bottom_ipin_5.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__3_.mem_bottom_ipin_5.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__3_.mem_bottom_ipin_6.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__3_.mem_bottom_ipin_6.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__3_.mem_bottom_ipin_7.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__3_.mem_bottom_ipin_7.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_3__3_.mem_top_ipin_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__1_.mem_left_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_0__1_.mem_left_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_1.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_1.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_2.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_2.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_3.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_3.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_4.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_4.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_5.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_5.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_6.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_6.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_7.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_7.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__2_.mem_left_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_0__2_.mem_left_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_1.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_1.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_2.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_2.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_3.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_3.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_4.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_4.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_5.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_5.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_6.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_6.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_7.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_7.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__3_.mem_left_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__3_.mem_left_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__3_.mem_left_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_0__3_.mem_left_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_0__3_.mem_right_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__3_.mem_right_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__3_.mem_right_ipin_1.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__3_.mem_right_ipin_1.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__3_.mem_right_ipin_2.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__3_.mem_right_ipin_2.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__3_.mem_right_ipin_3.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__3_.mem_right_ipin_3.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__3_.mem_right_ipin_4.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__3_.mem_right_ipin_4.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__3_.mem_right_ipin_5.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__3_.mem_right_ipin_5.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__3_.mem_right_ipin_6.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__3_.mem_right_ipin_6.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_0__3_.mem_right_ipin_7.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_0__3_.mem_right_ipin_7.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_1__1_.mem_left_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_1__1_.mem_left_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_1__1_.mem_left_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_left_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_1__2_.mem_left_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_left_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_1__3_.mem_left_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_1__3_.mem_left_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_1__3_.mem_left_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_1__3_.mem_left_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_1__3_.mem_right_ipin_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_2__3_.mem_left_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_2__3_.mem_left_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_2__3_.mem_left_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_2__3_.mem_left_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_2__3_.mem_right_ipin_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_3__1_.mem_left_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__1_.mem_left_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__1_.mem_left_ipin_1.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__1_.mem_left_ipin_1.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__1_.mem_left_ipin_2.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__1_.mem_left_ipin_2.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__1_.mem_left_ipin_3.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__1_.mem_left_ipin_3.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__1_.mem_left_ipin_4.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__1_.mem_left_ipin_4.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__1_.mem_left_ipin_5.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__1_.mem_left_ipin_5.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__1_.mem_left_ipin_6.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__1_.mem_left_ipin_6.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__1_.mem_left_ipin_7.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__1_.mem_left_ipin_7.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_3__1_.mem_right_ipin_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_3__2_.mem_left_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__2_.mem_left_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__2_.mem_left_ipin_1.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__2_.mem_left_ipin_1.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__2_.mem_left_ipin_2.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__2_.mem_left_ipin_2.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__2_.mem_left_ipin_3.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__2_.mem_left_ipin_3.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__2_.mem_left_ipin_4.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__2_.mem_left_ipin_4.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__2_.mem_left_ipin_5.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__2_.mem_left_ipin_5.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__2_.mem_left_ipin_6.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__2_.mem_left_ipin_6.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__2_.mem_left_ipin_7.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__2_.mem_left_ipin_7.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_3__2_.mem_right_ipin_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_3__3_.mem_left_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__3_.mem_left_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__3_.mem_left_ipin_1.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__3_.mem_left_ipin_1.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__3_.mem_left_ipin_2.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__3_.mem_left_ipin_2.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__3_.mem_left_ipin_3.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__3_.mem_left_ipin_3.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__3_.mem_left_ipin_4.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__3_.mem_left_ipin_4.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__3_.mem_left_ipin_5.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__3_.mem_left_ipin_5.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__3_.mem_left_ipin_6.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__3_.mem_left_ipin_6.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__3_.mem_left_ipin_7.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__3_.mem_left_ipin_7.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_0.mem_out[0:5], 6'b000001);
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_0.mem_outb[0:5], 6'b111110);
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_3__3_.mem_right_ipin_2.mem_outb[0:1], {2{1'b1}});
end
// ----- End deposit bitstream to configuration memories -----
`endif
// ----- End load bitstream to configuration memories -----
endmodule
// ----- END Verilog module for and2_top_formal_verification -----

